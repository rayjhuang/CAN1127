
`timescale 1ns/10ps
`define ATPG // let ANALOG_TOP don't report some dummy messages
`define BENCH bench
`include "../bench/def_bench.v"
module stm_atpg;
`ifdef FSDB
initial begin
	$fsdbDumpfile ("bench_a.fsdb");
	$fsdbDumpvars;
	forever #100_000 $fsdbDumpflush;
end
`endif
initial begin
`ifdef VCD
	$dumpfile ("bench_a.vcd");
	$dumpvars (9,`BENCH);
	$dumpvars (2,stm_atpg);
	forever #100_000 $dumpflush;
`endif
	#200_000_000
	$display ($time,"ns <%m> ERROR: simulation time's up");
	$finish;
end

//pulldown (`DUT.U0_CODE.VSS);
//pulldown (`DUT.U0_CODE.HV_VSS);

reg pd_ena=1;
initial #1000 pd_ena=0;
initial force `DUT_ANA.GATE_A = 'hz; // STIL expects this to be floating, 'cause it is generated by an empty ANALOG_TOP
initial force `DUT_ANA.GATE_B = 'hz;
pulldown (pull0) (pd_gpio2); tranif1 (pd_gpio2,`DUT.GPIO2,pd_ena);
pulldown (pull0) (pd_gpio1); tranif1 (pd_gpio1,`DUT.GPIO1,pd_ena);
pulldown (pull0) (pd_sda);   tranif1 (pd_sda,`  DUT.SDA,  pd_ena); // why STIL floating this?
pulldown (pull0) (pd_scl);   tranif1 (pd_scl,  `DUT.SCL,  pd_ena); // and expected this to be floating?
initial begin
`ifdef MAX $sdf_annotate ("chiptop_ss.sdf",`DUT,,,"MAXIMUM");
`elsif MIN $sdf_annotate ("chiptop_ff.sdf",`DUT,,,"MINIMUM");
`else "ERROR: no SDF case specified"
`endif
	#80 `DUT.U0_ANALOG_TOP.r_rstz = 1;
//	#1000 $finish;
end
`ifdef SF0 // stuck-at-0 fault
initial begin: stuck_0_fault
//	force `REGBNK.csp_regr =0; // atpg_chain failed
//	force `REGBNK.rb_otpwr =0; // pass atpg_chain and atpg_serial2
;
end // stuck_0_fault
`endif

// it's a disaster when a FF sample a X data (no delay in this STD lib)
   pulldown (weak0) (bench.SDA);
   pulldown (weak0) (bench.SCL);
   pulldown (weak0) (bench.GPIO1);
// pulldown (weak0) (bench.GPIO2);

integer idx;
parameter MAX_LENGTH = 1204; // max scan length
parameter N_SIG = 7; // no. of scan signals (in/out/control)
//rameter NP_POS = 8; // position of resetz (negative pulse)
parameter PP_POS = 4; // position of clock (positive pulse)
parameter CK_PERIOD = 50; // ns, defined in STIL (refer to exist.tcl chiptop_11xxa0.spf)
parameter CK_RISE = 4; // x10%, rise at
`define STR_PP "PP 20 40" // positive pulse string, according to CK_RISE
parameter MAX_VEC_WIDTH = 100; // max char per vector
`define SIG_OE 'h60 // output enable for those output signals
`define SIG_BUS \
	bench.GPIO5,\
	bench.GPIO4,\
	bench.GPIO3,\
	bench.GPIO1,\
	bench.SDA,\
	bench.SCL,\
	bench.TST
reg [8*30:0] sig_name [0:N_SIG-1];
initial begin
	sig_name[6]  = "GPIO5";
	sig_name[5]  = "GPIO4";
	sig_name[4]  = {"GPIO3: ",`STR_PP," after POR"};
	sig_name[3]  = "GPIO1";
	sig_name[2]  = "SDA";
	sig_name[1]  = "SCL";
	sig_name[0]  = "TST";
end

`ifdef VEC_VER // verifying vectors
reg [N_SIG-1:0] vec_bus;
wire [N_SIG-1:0] vec_wire = vec_bus;
tran u0 [N_SIG-1:0] ({`SIG_BUS},vec_wire);
initial begin: vector_verify
	reg [8*MAX_VEC_WIDTH-1:0] vec_str;
	reg [7:0] ptr, pos;
	reg flag;
	integer fpr;
	fpr = $fopen(`VEC_VER,"r");
	while (!$feof(fpr)) begin
	   flag = $fgets(vec_str,fpr);
	   if (bench.vector_number<=5
	    || bench.vector_number>=15989 && bench.vector_number<=16000)
	      $display ($time,"ns <%m> vector_number:%0d,vec_str:%0s",bench.vector_number,vec_str);
	   flag = 0;
	   for (idx=0;idx<MAX_VEC_WIDTH;idx=idx+1) begin
	      flag = flag ?vec_str[idx*8+:8]>" " :vec_str[idx*8+:8]==";";
	      if (!flag || vec_str[idx*8+:8]==";") vec_str[idx*8+:8]=0;
	   end
	   ptr =0;
	   for (idx=0;idx<MAX_VEC_WIDTH;idx=idx+1)
	      if (!ptr && vec_str[idx*8+:8]) ptr = idx;
	   if (ptr) begin // a cycle
	      for (idx=0;idx<N_SIG;idx=idx+1) begin
	         pos = N_SIG-1-idx;
	         vec_bus[pos] =
			(pos==PP_POS) ? 'h0 :
//			(pos==NP_POS) ? 'h1 :
				vec_str[(idx+ptr)*8+:8]=="1" ?'h1 :
				vec_str[(idx+ptr)*8+:8]=="0" ?'h0 :
				vec_str[(idx+ptr)*8+:8]=="H" ?'hz :
				vec_str[(idx+ptr)*8+:8]=="L" ?'hz :
				vec_str[(idx+ptr)*8+:8]=="X" ?'hz :'hx;
	      end
#(CK_PERIOD*CK_RISE/10)
	      if (vec_str[(N_SIG-1-PP_POS+ptr)*8+:8]=="1") vec_bus[PP_POS] = 'h1;
//	      if (vec_str[(N_SIG-1-NP_POS+ptr)*8+:8]=="0") vec_bus[NP_POS] = 'h0;
#(CK_PERIOD*4/10)
	      vec_bus[PP_POS] = 'h0;
//	      vec_bus[NP_POS] = 'h1;
#(CK_PERIOD*(10-CK_RISE-4)/10-1)
	      for (idx=0;idx<N_SIG;idx=idx+1) begin
	         pos = N_SIG-1-idx;
	         if (vec_str[(idx+ptr)*8+:8]=="H" && vec_wire[pos]!=='h1 ||
	             vec_str[(idx+ptr)*8+:8]=="L" && vec_wire[pos]!=='h0) begin
	            bench.mismatch_number = bench.mismatch_number +1;
	            $display ($time,"ns <%m> ERROR: %0s mismatch vec:%0d, exp:%c, dat:%x",
			sig_name[pos],bench.vector_number,vec_str[(idx+ptr)*8+:8],vec_wire[pos]);
	         end
	      end
#1	      bench.vector_number = bench.vector_number +1;
	   end
	end
	if (bench.mismatch_number>0)
	   $display ($time,"ns <%m> ERROR: simulation ended at vector: %0d, mismatch: %0d",
							bench.vector_number,bench.mismatch_number);
	else
	   $display ($time,"ns <%m> NOTE: simulation completed at vector: %0d",bench.vector_number);
	$finish;
end

endmodule // stm_atpg
module bench; // a very simple bench for verfying vectors
   integer pattern_number ='hx,
           vector_number =0,
           mismatch_number =0;

   always @(vector_number)
	if (vector_number%1000==0)
	   $display ($time,"ns <%m> vector: %0d, mismatch: %0d",vector_number,mismatch_number);

`ifdef CAN1126A0 chiptop_1126a0
`endif
   U0_DUT (
      .DP(DP),
      .DN(DN),
      .CC1(CC1),
      .CC2(CC2),
      .TST(TST),
      .SCL(SCL),
      .SDA(SDA),
      .GPIO1(GPIO1),
      .GPIO2(GPIO2),
      .GPIO3(GPIO3),
      .GPIO4(GPIO4),
      .GPIO5(GPIO5));
`endif // VEC_VER


`ifdef VEC_GEN // generating vectors
always #1_000_000 begin
	$display ($time,"ns <%m> NOTE: pattern: %0d, vector: %0d",
				bench.pattern_number,bench.vector_number);
end
integer fpw;
initial begin
	fpw = $fopen(`VEC_GEN,"w"); // .txt for auto backup
	$fwrite(fpw,"@@PATTERN DEFINE\n");
	for (idx=0;idx<N_SIG;idx=idx+1) $fwrite(fpw,"\/\/\t%0s\n",sig_name[idx]);
end
reg pp_pulse, np_pulse;
integer pattern_number =-1;
wire pattern_1st = (bench.vector_number <= (MAX_LENGTH+3)); // first MAX_LENGTH+3 vectors are shift-in only
function [7:0] s2char (input sig, oe);
	s2char = sig===0 ?oe ? pattern_1st ?"X" :"L" :"0"
	       : sig===1 ?oe ? pattern_1st ?"X" :"H" :"1" :"X";
endfunction
wire [N_SIG-1:0] sig_bus = { `SIG_BUS },
                 sig_oe = { `SIG_OE };
always @(bench.vector_number) begin
#(CK_PERIOD/2)
	pp_pulse = sig_bus[PP_POS];
//	np_pulse = sig_bus[NP_POS];
	if (pattern_number!=bench.pattern_number && pp_pulse) begin
	   $fwrite(fpw,"P%04d:",bench.pattern_number);
	   pattern_number = bench.pattern_number;
	end
	$fwrite(fpw,"\t");
#(CK_PERIOD/2-1)	
	for (idx=0;idx<N_SIG;idx=idx+1)
	   $fwrite(fpw,"%1c",s2char(
		(idx==PP_POS) ?pp_pulse :
//		(idx==NP_POS) ?np_pulse :
				sig_bus[idx], sig_oe[idx]));
	$fwrite(fpw,";\n");
	if (bench.vector_number%1000==0) $fflush(fpw);
end // before 100ns
`endif // VEC_GEN

endmodule // stm_atpg or the simple bench for verifying

