
module anatop_1127a0 ( CC1, CC2, DP, DN, VFB, CSP, CSN, COMP, SW, BST, VDRV, 
        LG, HG, GATE, BST_SET, DCM_SEL, HGOFF, HGON, LGOFF, LGON, EN_DRV, FSW, 
        EN_OSC, MAXDS, EN_GM, EN_ODLDO, EN_IBUK, EN_CP, EXT_CP, INT_CP, 
        ANTI_INRUSH, PWREN_HOLD, RP_SEL, RP1_EN, RP2_EN, VCONN1_EN, VCONN2_EN, 
        SGP, S20U, S100U, TX_EN, TX_DAT, CC_SEL, TRA, TFA, LSR, RX_DAT, RX_SQL, 
        SEL_RX_TH, DAC1_EN, DPDN_SHORT, DP_2V7_EN, DN_2V7_EN, DP_0P6V_EN, 
        DN_0P6V_EN, DP_DWN_EN, DN_DWN_EN, CC_SLOPE, DAC2, DAC3, DAC1, CV2, 
        LFOSC_ENB, VO_DISCHG, DISCHG_SEL, CMP_SEL_VO10, CMP_SEL_VO20, 
        CMP_SEL_GP1, CMP_SEL_GP2, CMP_SEL_GP3, CMP_SEL_GP4, CMP_SEL_GP5, 
        CMP_SEL_VIN20, CMP_SEL_TS, CMP_SEL_IS, CMP_SEL_CC2, CMP_SEL_CC1, 
        CMP_SEL_CC2_4, CMP_SEL_CC1_4, CMP_SEL_DP, CMP_SEL_DP_3, CMP_SEL_DN, 
        CMP_SEL_DN_3, OCP_EN, COMP_O, CCI2C_EN, UVP_SEL, TM, V5OCP, RSTB, DAC0, 
        SLEEP, OSC_LOW, OSC_STOP, PWRDN, VPP_ZERO, OSC_O, RD_DET, IMP_OSC, 
        DRP_OSC, STB_RP, RD_ENB, OCP, SCP, UVP, LDO3P9V, VPP_SEL, CC1_DOB, 
        CC2_DOB, CC1_DI, CC2_DI, OTPI, OVP_SEL, OVP, DN_COMP, DP_COMP, 
        DPDN_VTH, DPDEN, DPDO, DPIE, DNDEN, DNDO, DNIE, CP_CLKX2, 
        SEL_CONST_OVP, LP_EN, DNCHK_EN, IRP_EN, CCFBEN, REGTRM, AD_RST, 
        AD_HOLD, DN_FAULT, SEL_CCGAIN, VFB_SWB, CPVSEL, CLAMPV_EN, HVNG_CPEN, 
        OCP_SEL, OCP_80M, OCP_160M, DMY_OUT, DMY_IN, VPP_OTP, RSTB_5, V1P1, 
        TS_ANA_R, GP5_ANA_R, GP4_ANA_R, GP3_ANA_R, GP2_ANA_R, GP1_ANA_R, 
        TS_ANA_P, GP5_ANA_P, GP4_ANA_P, GP3_ANA_P, GP2_ANA_P, GP1_ANA_P );
  input [1:0] FSW;
  input [1:0] RP_SEL;
  input [5:1] SGP;
  input [1:0] CC_SLOPE;
  input [7:0] DAC2;
  input [5:0] DAC3;
  input [9:0] DAC1;
  input [3:0] TM;
  input [10:0] DAC0;
  input [1:0] OVP_SEL;
  input [55:0] REGTRM;
  output [3:0] DMY_OUT;
  input [4:0] DMY_IN;
  input BST_SET, DCM_SEL, HGOFF, HGON, LGOFF, LGON, EN_DRV, EN_OSC, MAXDS,
         EN_GM, EN_ODLDO, EN_IBUK, EN_CP, EXT_CP, INT_CP, ANTI_INRUSH,
         PWREN_HOLD, RP1_EN, RP2_EN, VCONN1_EN, VCONN2_EN, S20U, S100U, TX_EN,
         TX_DAT, CC_SEL, TRA, TFA, LSR, SEL_RX_TH, DAC1_EN, DPDN_SHORT,
         DP_2V7_EN, DN_2V7_EN, DP_0P6V_EN, DN_0P6V_EN, DP_DWN_EN, DN_DWN_EN,
         CV2, LFOSC_ENB, VO_DISCHG, DISCHG_SEL, CMP_SEL_VO10, CMP_SEL_VO20,
         CMP_SEL_GP1, CMP_SEL_GP2, CMP_SEL_GP3, CMP_SEL_GP4, CMP_SEL_GP5,
         CMP_SEL_VIN20, CMP_SEL_TS, CMP_SEL_IS, CMP_SEL_CC2, CMP_SEL_CC1,
         CMP_SEL_CC2_4, CMP_SEL_CC1_4, CMP_SEL_DP, CMP_SEL_DP_3, CMP_SEL_DN,
         CMP_SEL_DN_3, OCP_EN, CCI2C_EN, UVP_SEL, SLEEP, OSC_LOW, OSC_STOP,
         PWRDN, VPP_ZERO, STB_RP, RD_ENB, LDO3P9V, VPP_SEL, CC1_DOB, CC2_DOB,
         DPDN_VTH, DPDEN, DPDO, DPIE, DNDEN, DNDO, DNIE, CP_CLKX2,
         SEL_CONST_OVP, LP_EN, DNCHK_EN, IRP_EN, CCFBEN, AD_RST, AD_HOLD,
         SEL_CCGAIN, VFB_SWB, CPVSEL, CLAMPV_EN, HVNG_CPEN, OCP_SEL, TS_ANA_R,
         GP5_ANA_R, GP4_ANA_R, GP3_ANA_R, GP2_ANA_R, GP1_ANA_R;
  output LG, HG, GATE, RX_DAT, RX_SQL, COMP_O, V5OCP, RSTB, OSC_O, RD_DET,
         IMP_OSC, DRP_OSC, OCP, SCP, UVP, CC1_DI, CC2_DI, OTPI, OVP, DN_COMP,
         DP_COMP, DN_FAULT, OCP_80M, OCP_160M, VPP_OTP, RSTB_5, V1P1, TS_ANA_P,
         GP5_ANA_P, GP4_ANA_P, GP3_ANA_P, GP2_ANA_P, GP1_ANA_P;
  inout CC1,  CC2,  DP,  DN,  VFB,  CSP,  CSN,  COMP,  SW,  BST,  VDRV;


endmodule

