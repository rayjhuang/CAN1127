`timescale 1ns/1ns
module mpsse_mst_i2c (
`include "mpsse_mst_bhv.v"
`include "mpsse_i2c_task.v"
endmodule // mpsse_mst_i2c
