#=============================================================================
#Copyright 2022 MACRONIX INTERNATIONAL Co., Ltd.  All Rights Reserved.
#CONFIDENTIAL SOFTWARE/DATA OF MACRONIX INTERNATIONAL Co., Ltd
#=============================================================================
#Program		Single Port SRAM Compiler
#Process		0.18μm CMOS SPDM/SPTM/SPQM BCD(5V/40V)
#Version		1.0
#Date			2022/11/07 14:00:50
#=============================================================================
#Instance Name		MSL18B_1536X8_RW10TM4_16_20221107
#Words			1536
#Bits			8
#Multiplexer Width	16
#=============================================================================
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO MSL18B_1536X8_RW10TM4_16_20221107
  CLASS RING ;
  FOREIGN MSL18B_1536X8_RW10TM4_16_20221107 0 0 ;
  ORIGIN 0 0 ;
  SIZE 317.760 BY 348.410 ;
  SYMMETRY X Y R90 ;
  PIN DO[0]
   DIRECTION OUTPUT ;
   USE SIGNAL ;
   ANTENNADIFFAREA 3.2508 ;
   PORT
     LAYER MET1 ;
     RECT 39.810 22.000 40.710 22.280 ;
     LAYER MET2 ;
     RECT 39.810 22.000 40.710 22.280 ;
     LAYER MET3 ;
     RECT 39.810 22.000 40.710 22.280 ;
   END
  END DO[0]
  PIN DI[0]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3784 ;
   PORT
     LAYER MET1 ;
     RECT 41.725 22.000 42.625 22.280 ;
     LAYER MET2 ;
     RECT 41.725 22.000 42.625 22.280 ;
     LAYER MET3 ;
     RECT 41.725 22.000 42.625 22.280 ;
   END
  END DI[0]
  PIN DO[1]
   DIRECTION OUTPUT ;
   USE SIGNAL ;
   ANTENNADIFFAREA 3.2508 ;
   PORT
     LAYER MET1 ;
     RECT 68.270 22.000 69.170 22.280 ;
     LAYER MET2 ;
     RECT 68.270 22.000 69.170 22.280 ;
     LAYER MET3 ;
     RECT 68.270 22.000 69.170 22.280 ;
   END
  END DO[1]
  PIN DI[1]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3784 ;
   PORT
     LAYER MET1 ;
     RECT 70.185 22.000 71.085 22.280 ;
     LAYER MET2 ;
     RECT 70.185 22.000 71.085 22.280 ;
     LAYER MET3 ;
     RECT 70.185 22.000 71.085 22.280 ;
   END
  END DI[1]
  PIN DO[2]
   DIRECTION OUTPUT ;
   USE SIGNAL ;
   ANTENNADIFFAREA 3.2508 ;
   PORT
     LAYER MET1 ;
     RECT 96.730 22.000 97.630 22.280 ;
     LAYER MET2 ;
     RECT 96.730 22.000 97.630 22.280 ;
     LAYER MET3 ;
     RECT 96.730 22.000 97.630 22.280 ;
   END
  END DO[2]
  PIN DI[2]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3784 ;
   PORT
     LAYER MET1 ;
     RECT 98.645 22.000 99.545 22.280 ;
     LAYER MET2 ;
     RECT 98.645 22.000 99.545 22.280 ;
     LAYER MET3 ;
     RECT 98.645 22.000 99.545 22.280 ;
   END
  END DI[2]
  PIN DO[3]
   DIRECTION OUTPUT ;
   USE SIGNAL ;
   ANTENNADIFFAREA 3.2508 ;
   PORT
     LAYER MET1 ;
     RECT 125.190 22.000 126.090 22.280 ;
     LAYER MET2 ;
     RECT 125.190 22.000 126.090 22.280 ;
     LAYER MET3 ;
     RECT 125.190 22.000 126.090 22.280 ;
   END
  END DO[3]
  PIN DI[3]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3784 ;
   PORT
     LAYER MET1 ;
     RECT 127.105 22.000 128.005 22.280 ;
     LAYER MET2 ;
     RECT 127.105 22.000 128.005 22.280 ;
     LAYER MET3 ;
     RECT 127.105 22.000 128.005 22.280 ;
   END
  END DI[3]
  PIN A[9]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.972 ;
   PORT
     LAYER MET1 ;
     RECT 140.995 22.000 141.895 22.280 ;
     LAYER MET2 ;
     RECT 140.995 22.000 141.895 22.280 ;
     LAYER MET3 ;
     RECT 140.995 22.000 141.895 22.280 ;
   END
  END A[9]
  PIN A[10]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.972 ;
   PORT
     LAYER MET1 ;
     RECT 142.395 22.000 143.295 22.280 ;
     LAYER MET2 ;
     RECT 142.395 22.000 143.295 22.280 ;
     LAYER MET3 ;
     RECT 142.395 22.000 143.295 22.280 ;
   END
  END A[10]
  PIN A[8]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.972 ;
   PORT
     LAYER MET1 ;
     RECT 146.710 22.000 147.610 22.280 ;
     LAYER MET2 ;
     RECT 146.710 22.000 147.610 22.280 ;
     LAYER MET3 ;
     RECT 146.710 22.000 147.610 22.280 ;
   END
  END A[8]
  PIN A[7]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.972 ;
   PORT
     LAYER MET1 ;
     RECT 149.105 22.000 150.005 22.280 ;
     LAYER MET2 ;
     RECT 149.105 22.000 150.005 22.280 ;
     LAYER MET3 ;
     RECT 149.105 22.000 150.005 22.280 ;
   END
  END A[7]
  PIN A[6]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.972 ;
   PORT
     LAYER MET1 ;
     RECT 151.500 22.000 152.400 22.280 ;
     LAYER MET2 ;
     RECT 151.500 22.000 152.400 22.280 ;
     LAYER MET3 ;
     RECT 151.500 22.000 152.400 22.280 ;
   END
  END A[6]
  PIN A[5]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3024 ;
   PORT
     LAYER MET1 ;
     RECT 155.820 22.000 156.720 22.280 ;
     LAYER MET2 ;
     RECT 155.820 22.000 156.720 22.280 ;
     LAYER MET3 ;
     RECT 155.820 22.000 156.720 22.280 ;
   END
  END A[5]
  PIN A[4]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3024 ;
   PORT
     LAYER MET1 ;
     RECT 158.620 22.000 159.520 22.280 ;
     LAYER MET2 ;
     RECT 158.620 22.000 159.520 22.280 ;
     LAYER MET3 ;
     RECT 158.620 22.000 159.520 22.280 ;
   END
  END A[4]
  PIN A[2]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.648 ;
   PORT
     LAYER MET1 ;
     RECT 161.165 22.000 162.065 22.280 ;
     LAYER MET2 ;
     RECT 161.165 22.000 162.065 22.280 ;
     LAYER MET3 ;
     RECT 161.165 22.000 162.065 22.280 ;
   END
  END A[2]
  PIN A[3]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.648 ;
   PORT
     LAYER MET1 ;
     RECT 162.565 22.000 163.465 22.280 ;
     LAYER MET2 ;
     RECT 162.565 22.000 163.465 22.280 ;
     LAYER MET3 ;
     RECT 162.565 22.000 163.465 22.280 ;
   END
  END A[3]
  PIN A[0]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.648 ;
   PORT
     LAYER MET1 ;
     RECT 165.455 22.000 166.355 22.280 ;
     LAYER MET2 ;
     RECT 165.455 22.000 166.355 22.280 ;
     LAYER MET3 ;
     RECT 165.455 22.000 166.355 22.280 ;
   END
  END A[0]
  PIN A[1]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.648 ;
   PORT
     LAYER MET1 ;
     RECT 169.085 22.000 169.985 22.280 ;
     LAYER MET2 ;
     RECT 169.085 22.000 169.985 22.280 ;
     LAYER MET3 ;
     RECT 169.085 22.000 169.985 22.280 ;
   END
  END A[1]
  PIN OEB
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.27 ;
   PORT
     LAYER MET1 ;
     RECT 170.690 22.000 171.590 22.280 ;
     LAYER MET2 ;
     RECT 170.690 22.000 171.590 22.280 ;
     LAYER MET3 ;
     RECT 170.690 22.000 171.590 22.280 ;
   END
  END OEB
  PIN WEB
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.0792 ;
   PORT
     LAYER MET1 ;
     RECT 172.190 22.000 173.090 22.280 ;
     LAYER MET2 ;
     RECT 172.190 22.000 173.090 22.280 ;
     LAYER MET3 ;
     RECT 172.190 22.000 173.090 22.280 ;
   END
  END WEB
  PIN CK
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.252 ;
   PORT
     LAYER MET1 ;
     RECT 173.690 22.000 174.590 22.280 ;
     LAYER MET2 ;
     RECT 173.690 22.000 174.590 22.280 ;
     LAYER MET3 ;
     RECT 173.690 22.000 174.590 22.280 ;
   END
  END CK
  PIN CSB
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 3.06 ;
   PORT
     LAYER MET1 ;
     RECT 175.295 22.000 176.195 22.280 ;
     LAYER MET2 ;
     RECT 175.295 22.000 176.195 22.280 ;
     LAYER MET3 ;
     RECT 175.295 22.000 176.195 22.280 ;
   END
  END CSB
  PIN DO[4]
   DIRECTION OUTPUT ;
   USE SIGNAL ;
   ANTENNADIFFAREA 3.2508 ;
   PORT
     LAYER MET1 ;
     RECT 196.205 22.000 197.105 22.280 ;
     LAYER MET2 ;
     RECT 196.205 22.000 197.105 22.280 ;
     LAYER MET3 ;
     RECT 196.205 22.000 197.105 22.280 ;
   END
  END DO[4]
  PIN DI[4]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3784 ;
   PORT
     LAYER MET1 ;
     RECT 198.120 22.000 199.020 22.280 ;
     LAYER MET2 ;
     RECT 198.120 22.000 199.020 22.280 ;
     LAYER MET3 ;
     RECT 198.120 22.000 199.020 22.280 ;
   END
  END DI[4]
  PIN DO[5]
   DIRECTION OUTPUT ;
   USE SIGNAL ;
   ANTENNADIFFAREA 3.2508 ;
   PORT
     LAYER MET1 ;
     RECT 224.665 22.000 225.565 22.280 ;
     LAYER MET2 ;
     RECT 224.665 22.000 225.565 22.280 ;
     LAYER MET3 ;
     RECT 224.665 22.000 225.565 22.280 ;
   END
  END DO[5]
  PIN DI[5]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3784 ;
   PORT
     LAYER MET1 ;
     RECT 226.580 22.000 227.480 22.280 ;
     LAYER MET2 ;
     RECT 226.580 22.000 227.480 22.280 ;
     LAYER MET3 ;
     RECT 226.580 22.000 227.480 22.280 ;
   END
  END DI[5]
  PIN DO[6]
   DIRECTION OUTPUT ;
   USE SIGNAL ;
   ANTENNADIFFAREA 3.2508 ;
   PORT
     LAYER MET1 ;
     RECT 253.125 22.000 254.025 22.280 ;
     LAYER MET2 ;
     RECT 253.125 22.000 254.025 22.280 ;
     LAYER MET3 ;
     RECT 253.125 22.000 254.025 22.280 ;
   END
  END DO[6]
  PIN DI[6]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3784 ;
   PORT
     LAYER MET1 ;
     RECT 255.040 22.000 255.940 22.280 ;
     LAYER MET2 ;
     RECT 255.040 22.000 255.940 22.280 ;
     LAYER MET3 ;
     RECT 255.040 22.000 255.940 22.280 ;
   END
  END DI[6]
  PIN DO[7]
   DIRECTION OUTPUT ;
   USE SIGNAL ;
   ANTENNADIFFAREA 3.2508 ;
   PORT
     LAYER MET1 ;
     RECT 281.585 22.000 282.485 22.280 ;
     LAYER MET2 ;
     RECT 281.585 22.000 282.485 22.280 ;
     LAYER MET3 ;
     RECT 281.585 22.000 282.485 22.280 ;
   END
  END DO[7]
  PIN DI[7]
   DIRECTION INPUT ;
   USE SIGNAL ;
   ANTENNAGATEAREA 0.3784 ;
   PORT
     LAYER MET1 ;
     RECT 283.500 22.000 284.400 22.280 ;
     LAYER MET2 ;
     RECT 283.500 22.000 284.400 22.280 ;
     LAYER MET3 ;
     RECT 283.500 22.000 284.400 22.280 ;
   END
  END DI[7]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER MET3 ;
      RECT 0.0 0.0 10.000 348.410 ;
      LAYER MET3 ;
      RECT 307.760 0.0 317.760 348.410 ;
      LAYER MET2 ;
      RECT 0.0 0.0 317.760 10.000 ;
      LAYER MET2 ;
      RECT 0.0 338.410 317.760 348.410 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER MET3 ;
      RECT 11.000 11.000 21.000 337.410 ;
      LAYER MET3 ;
      RECT 296.760 11.000 306.760 337.410 ;
      LAYER MET2 ;
      RECT 11.000 11.000 306.760 21.000 ;
      LAYER MET2 ;
      RECT 11.000 327.410 306.760 337.410 ;
    END
  END GND
  OBS
    LAYER VIA1 ;
     RECT 22.000 22.510 295.760 325.900 ;
    LAYER VIA2 ;
     RECT 22.000 22.560 295.760 325.850 ;
    LAYER VIA1 ;
     RECT 22.000 325.900 295.760 326.410 ;
    LAYER VIA2 ;
     RECT 22.000 325.850 295.760 326.410 ;
    LAYER VIA1 ;
     RECT 22.000 22.000 295.760 22.510 ;
    LAYER VIA2 ;
     RECT 22.000 22.000 295.760 22.560 ;
    LAYER MET1 ;
     RECT 22.000 22.510 295.760 325.900 ;
    LAYER MET1 ;
     RECT 22.000 325.900 295.760 326.410 ;
    LAYER MET1 ;
     RECT 22.000 22.000 39.580 22.510 ;
    LAYER MET1 ;
     RECT 40.940 22.000 41.495 22.510 ;
    LAYER MET1 ;
     RECT 42.855 22.000 68.040 22.510 ;
    LAYER MET1 ;
     RECT 69.400 22.000 69.955 22.510 ;
    LAYER MET1 ;
     RECT 71.315 22.000 96.500 22.510 ;
    LAYER MET1 ;
     RECT 97.860 22.000 98.415 22.510 ;
    LAYER MET1 ;
     RECT 99.775 22.000 124.960 22.510 ;
    LAYER MET1 ;
     RECT 126.320 22.000 126.875 22.510 ;
    LAYER MET1 ;
     RECT 128.235 22.000 140.765 22.510 ;
    LAYER MET1 ;
     RECT 142.125 22.000 142.165 22.510 ;
    LAYER MET1 ;
     RECT 143.525 22.000 146.480 22.510 ;
    LAYER MET1 ;
     RECT 147.840 22.000 148.875 22.510 ;
    LAYER MET1 ;
     RECT 150.235 22.000 151.270 22.510 ;
    LAYER MET1 ;
     RECT 152.630 22.000 155.590 22.510 ;
    LAYER MET1 ;
     RECT 156.950 22.000 158.390 22.510 ;
    LAYER MET1 ;
     RECT 159.750 22.000 160.935 22.510 ;
    LAYER MET1 ;
     RECT 162.295 22.000 162.335 22.510 ;
    LAYER MET1 ;
     RECT 163.695 22.000 165.225 22.510 ;
    LAYER MET1 ;
     RECT 166.585 22.000 168.855 22.510 ;
    LAYER MET1 ;
     RECT 170.215 22.000 170.460 22.510 ;
    LAYER MET1 ;
     RECT 171.820 22.000 171.960 22.510 ;
    LAYER MET1 ;
     RECT 173.320 22.000 173.460 22.510 ;
    LAYER MET1 ;
     RECT 174.820 22.000 175.065 22.510 ;
    LAYER MET1 ;
     RECT 176.425 22.000 195.975 22.510 ;
    LAYER MET1 ;
     RECT 197.335 22.000 197.890 22.510 ;
    LAYER MET1 ;
     RECT 199.250 22.000 224.435 22.510 ;
    LAYER MET1 ;
     RECT 225.795 22.000 226.350 22.510 ;
    LAYER MET1 ;
     RECT 227.710 22.000 252.895 22.510 ;
    LAYER MET1 ;
     RECT 254.255 22.000 254.810 22.510 ;
    LAYER MET1 ;
     RECT 256.170 22.000 281.355 22.510 ;
    LAYER MET1 ;
     RECT 282.715 22.000 283.270 22.510 ;
    LAYER MET1 ;
     RECT 284.630 22.000 295.760 22.510 ;
    LAYER MET2 ;
     RECT 22.000 22.560 295.760 325.850 ;
    LAYER MET2 ;
     RECT 22.000 325.850 295.760 326.410 ;
    LAYER MET2 ;
     RECT 22.000 22.000 39.530 22.560 ;
    LAYER MET2 ;
     RECT 40.990 22.000 41.445 22.560 ;
    LAYER MET2 ;
     RECT 42.905 22.000 67.990 22.560 ;
    LAYER MET2 ;
     RECT 69.450 22.000 69.905 22.560 ;
    LAYER MET2 ;
     RECT 71.365 22.000 96.450 22.560 ;
    LAYER MET2 ;
     RECT 97.910 22.000 98.365 22.560 ;
    LAYER MET2 ;
     RECT 99.825 22.000 124.910 22.560 ;
    LAYER MET2 ;
     RECT 126.370 22.000 126.825 22.560 ;
    LAYER MET2 ;
     RECT 128.285 22.000 140.715 22.560 ;
    LAYER MET2 ;
     RECT 143.575 22.000 146.430 22.560 ;
    LAYER MET2 ;
     RECT 147.890 22.000 148.825 22.560 ;
    LAYER MET2 ;
     RECT 150.285 22.000 151.220 22.560 ;
    LAYER MET2 ;
     RECT 152.680 22.000 155.540 22.560 ;
    LAYER MET2 ;
     RECT 157.000 22.000 158.340 22.560 ;
    LAYER MET2 ;
     RECT 159.800 22.000 160.885 22.560 ;
    LAYER MET2 ;
     RECT 163.745 22.000 165.175 22.560 ;
    LAYER MET2 ;
     RECT 166.635 22.000 168.805 22.560 ;
    LAYER MET2 ;
     RECT 170.265 22.000 170.410 22.560 ;
    LAYER MET2 ;
     RECT 171.870 22.000 171.910 22.560 ;
    LAYER MET2 ;
     RECT 173.370 22.000 173.410 22.560 ;
    LAYER MET2 ;
     RECT 174.870 22.000 175.015 22.560 ;
    LAYER MET2 ;
     RECT 176.475 22.000 195.925 22.560 ;
    LAYER MET2 ;
     RECT 197.385 22.000 197.840 22.560 ;
    LAYER MET2 ;
     RECT 199.300 22.000 224.385 22.560 ;
    LAYER MET2 ;
     RECT 225.845 22.000 226.300 22.560 ;
    LAYER MET2 ;
     RECT 227.760 22.000 252.845 22.560 ;
    LAYER MET2 ;
     RECT 254.305 22.000 254.760 22.560 ;
    LAYER MET2 ;
     RECT 256.220 22.000 281.305 22.560 ;
    LAYER MET2 ;
     RECT 282.765 22.000 283.220 22.560 ;
    LAYER MET2 ;
     RECT 284.680 22.000 295.760 22.560 ;
    LAYER MET3 ;
     RECT 22.000 22.560 295.760 325.850 ;
    LAYER MET3 ;
     RECT 22.000 325.850 295.760 326.410 ;
    LAYER MET3 ;
     RECT 22.000 22.000 39.530 22.560 ;
    LAYER MET3 ;
     RECT 40.990 22.000 41.445 22.560 ;
    LAYER MET3 ;
     RECT 42.905 22.000 67.990 22.560 ;
    LAYER MET3 ;
     RECT 69.450 22.000 69.905 22.560 ;
    LAYER MET3 ;
     RECT 71.365 22.000 96.450 22.560 ;
    LAYER MET3 ;
     RECT 97.910 22.000 98.365 22.560 ;
    LAYER MET3 ;
     RECT 99.825 22.000 124.910 22.560 ;
    LAYER MET3 ;
     RECT 126.370 22.000 126.825 22.560 ;
    LAYER MET3 ;
     RECT 128.285 22.000 140.715 22.560 ;
    LAYER MET3 ;
     RECT 143.575 22.000 146.430 22.560 ;
    LAYER MET3 ;
     RECT 147.890 22.000 148.825 22.560 ;
    LAYER MET3 ;
     RECT 150.285 22.000 151.220 22.560 ;
    LAYER MET3 ;
     RECT 152.680 22.000 155.540 22.560 ;
    LAYER MET3 ;
     RECT 157.000 22.000 158.340 22.560 ;
    LAYER MET3 ;
     RECT 159.800 22.000 160.885 22.560 ;
    LAYER MET3 ;
     RECT 163.745 22.000 165.175 22.560 ;
    LAYER MET3 ;
     RECT 166.635 22.000 168.805 22.560 ;
    LAYER MET3 ;
     RECT 170.265 22.000 170.410 22.560 ;
    LAYER MET3 ;
     RECT 171.870 22.000 171.910 22.560 ;
    LAYER MET3 ;
     RECT 173.370 22.000 173.410 22.560 ;
    LAYER MET3 ;
     RECT 174.870 22.000 175.015 22.560 ;
    LAYER MET3 ;
     RECT 176.475 22.000 195.925 22.560 ;
    LAYER MET3 ;
     RECT 197.385 22.000 197.840 22.560 ;
    LAYER MET3 ;
     RECT 199.300 22.000 224.385 22.560 ;
    LAYER MET3 ;
     RECT 225.845 22.000 226.300 22.560 ;
    LAYER MET3 ;
     RECT 227.760 22.000 252.845 22.560 ;
    LAYER MET3 ;
     RECT 254.305 22.000 254.760 22.560 ;
    LAYER MET3 ;
     RECT 256.220 22.000 281.305 22.560 ;
    LAYER MET3 ;
     RECT 282.765 22.000 283.220 22.560 ;
    LAYER MET3 ;
     RECT 284.680 22.000 295.760 22.560 ;
    LAYER MET2 ;
    RECT 0.000 47.985 22.000 48.885 ;
    LAYER VIA2 ;
    RECT 0.140 48.305 9.760 48.565 ;
    LAYER MET2 ;
    RECT 0.000 63.700 22.000 65.130 ;
    LAYER VIA2 ;
    RECT 0.140 64.025 9.760 64.805 ;
    LAYER MET2 ;
    RECT 0.000 72.430 22.000 73.330 ;
    LAYER VIA2 ;
    RECT 0.140 72.750 9.760 73.010 ;
    LAYER MET2 ;
    RECT 0.000 79.895 22.000 81.495 ;
    LAYER VIA2 ;
    RECT 0.140 80.045 9.760 81.345 ;
    LAYER MET2 ;
    RECT 0.000 84.965 22.000 86.315 ;
    LAYER VIA2 ;
    RECT 0.140 85.250 9.760 86.030 ;
    LAYER MET2 ;
    RECT 0.000 56.850 22.000 57.750 ;
    LAYER VIA2 ;
    RECT 0.140 57.170 9.760 57.430 ;
    LAYER MET2 ;
    RECT 0.000 45.940 22.000 46.480 ;
    LAYER VIA2 ;
    RECT 0.140 46.080 9.760 46.340 ;
    LAYER MET2 ;
    RECT 0.000 41.680 22.000 43.640 ;
    LAYER VIA2 ;
    RECT 0.140 42.010 9.760 43.310 ;
    LAYER MET2 ;
    RECT 0.000 35.140 22.000 37.340 ;
    LAYER VIA2 ;
    RECT 0.140 35.330 9.760 37.150 ;
    LAYER MET2 ;
    RECT 0.000 26.020 22.000 28.470 ;
    LAYER VIA2 ;
    RECT 0.140 26.335 9.760 28.155 ;
    LAYER MET3 ;
    RECT 21.000 88.405 22.000 89.405 ;
    LAYER MET3 ;
    RECT 21.000 70.955 22.000 71.855 ;
    LAYER MET3 ;
    RECT 21.000 60.000 22.000 61.400 ;
    LAYER MET3 ;
    RECT 21.000 51.950 22.000 52.850 ;
    LAYER MET3 ;
    RECT 21.000 44.900 22.000 45.440 ;
    LAYER MET3 ;
    RECT 21.000 37.840 22.000 39.140 ;
    LAYER MET3 ;
    RECT 21.000 31.540 22.000 32.840 ;
    LAYER MET3 ;
    RECT 21.000 22.740 22.000 23.840 ;
    LAYER MET3 ;
    RECT 46.325 0.000 47.745 22.000 ;
    LAYER MET3 ;
    RECT 103.245 0.000 104.665 22.000 ;
    LAYER VIA2 ;
    RECT 46.645 0.190 47.425 9.810 ;
    LAYER VIA2 ;
    RECT 103.565 0.190 104.345 9.810 ;
    LAYER MET3 ;
    RECT 37.735 0.000 38.635 22.000 ;
    LAYER MET3 ;
    RECT 94.655 0.000 95.555 22.000 ;
    LAYER VIA2 ;
    RECT 38.055 0.190 38.315 9.810 ;
    LAYER VIA2 ;
    RECT 94.975 0.190 95.235 9.810 ;
    LAYER MET3 ;
    RECT 28.280 0.000 29.700 22.000 ;
    LAYER MET3 ;
    RECT 85.200 0.000 86.620 22.000 ;
    LAYER VIA2 ;
    RECT 28.600 0.190 29.380 9.810 ;
    LAYER VIA2 ;
    RECT 85.520 0.190 86.300 9.810 ;
    LAYER MET2 ;
    RECT 50.755 21.000 51.655 22.000 ;
    LAYER MET2 ;
    RECT 107.675 21.000 108.575 22.000 ;
    LAYER MET2 ;
    RECT 33.840 21.000 35.260 22.000 ;
    LAYER MET2 ;
    RECT 90.760 21.000 92.180 22.000 ;
    LAYER MET2 ;
    RECT 31.670 21.000 32.570 22.000 ;
    LAYER MET2 ;
    RECT 88.590 21.000 89.490 22.000 ;
    LAYER MET2 ;
    RECT 24.850 21.000 26.270 22.000 ;
    LAYER MET2 ;
    RECT 81.770 21.000 83.190 22.000 ;
    LAYER MET3 ;
    RECT 74.785 0.000 76.205 22.000 ;
    LAYER MET3 ;
    RECT 131.705 0.000 133.125 22.000 ;
    LAYER VIA2 ;
    RECT 75.105 0.190 75.885 9.810 ;
    LAYER VIA2 ;
    RECT 132.025 0.190 132.805 9.810 ;
    LAYER MET3 ;
    RECT 66.195 0.000 67.095 22.000 ;
    LAYER MET3 ;
    RECT 123.115 0.000 124.015 22.000 ;
    LAYER VIA2 ;
    RECT 66.515 0.190 66.775 9.810 ;
    LAYER VIA2 ;
    RECT 123.435 0.190 123.695 9.810 ;
    LAYER MET3 ;
    RECT 56.740 0.000 58.160 22.000 ;
    LAYER MET3 ;
    RECT 113.660 0.000 115.080 22.000 ;
    LAYER VIA2 ;
    RECT 57.060 0.190 57.840 9.810 ;
    LAYER VIA2 ;
    RECT 113.980 0.190 114.760 9.810 ;
    LAYER MET2 ;
    RECT 79.215 21.000 80.115 22.000 ;
    LAYER MET2 ;
    RECT 136.135 21.000 137.035 22.000 ;
    LAYER MET2 ;
    RECT 62.300 21.000 63.720 22.000 ;
    LAYER MET2 ;
    RECT 119.220 21.000 120.640 22.000 ;
    LAYER MET2 ;
    RECT 60.130 21.000 61.030 22.000 ;
    LAYER MET2 ;
    RECT 117.050 21.000 117.950 22.000 ;
    LAYER MET2 ;
    RECT 53.310 21.000 54.730 22.000 ;
    LAYER MET2 ;
    RECT 110.230 21.000 111.650 22.000 ;
    LAYER MET3 ;
    RECT 139.595 0.000 140.495 22.000 ;
    LAYER VIA2 ;
    RECT 139.915 0.190 140.175 9.810 ;
    LAYER MET3 ;
    RECT 157.220 0.000 158.120 22.000 ;
    LAYER VIA2 ;
    RECT 157.540 0.190 157.800 9.810 ;
    LAYER MET3 ;
    RECT 145.310 0.000 146.210 22.000 ;
    LAYER VIA2 ;
    RECT 145.630 0.190 145.890 9.810 ;
    LAYER MET3 ;
    RECT 163.965 0.000 164.865 22.000 ;
    LAYER VIA2 ;
    RECT 164.285 0.190 164.545 9.810 ;
    LAYER MET3 ;
    RECT 167.685 0.000 168.585 22.000 ;
    LAYER VIA2 ;
    RECT 168.005 0.190 168.265 9.810 ;
    LAYER MET2 ;
    RECT 154.420 21.000 155.320 22.000 ;
    LAYER MET2 ;
    RECT 152.900 21.000 153.800 22.000 ;
    LAYER MET2 ;
    RECT 143.795 21.000 144.695 22.000 ;
    LAYER MET3 ;
    RECT 176.710 0.000 177.610 22.000 ;
    LAYER VIA2 ;
    RECT 177.030 0.190 177.290 9.810 ;
    LAYER MET2 ;
    RECT 178.110 21.000 179.010 22.000 ;
    LAYER MET3 ;
    RECT 202.720 0.000 204.140 22.000 ;
    LAYER MET3 ;
    RECT 259.640 0.000 261.060 22.000 ;
    LAYER VIA2 ;
    RECT 203.040 0.190 203.820 9.810 ;
    LAYER VIA2 ;
    RECT 259.960 0.190 260.740 9.810 ;
    LAYER MET3 ;
    RECT 194.130 0.000 195.030 22.000 ;
    LAYER MET3 ;
    RECT 251.050 0.000 251.950 22.000 ;
    LAYER VIA2 ;
    RECT 194.450 0.190 194.710 9.810 ;
    LAYER VIA2 ;
    RECT 251.370 0.190 251.630 9.810 ;
    LAYER MET3 ;
    RECT 184.675 0.000 186.095 22.000 ;
    LAYER MET3 ;
    RECT 241.595 0.000 243.015 22.000 ;
    LAYER VIA2 ;
    RECT 184.995 0.190 185.775 9.810 ;
    LAYER VIA2 ;
    RECT 241.915 0.190 242.695 9.810 ;
    LAYER MET2 ;
    RECT 207.150 21.000 208.050 22.000 ;
    LAYER MET2 ;
    RECT 264.070 21.000 264.970 22.000 ;
    LAYER MET2 ;
    RECT 190.235 21.000 191.655 22.000 ;
    LAYER MET2 ;
    RECT 247.155 21.000 248.575 22.000 ;
    LAYER MET2 ;
    RECT 188.065 21.000 188.965 22.000 ;
    LAYER MET2 ;
    RECT 244.985 21.000 245.885 22.000 ;
    LAYER MET2 ;
    RECT 181.245 21.000 182.665 22.000 ;
    LAYER MET2 ;
    RECT 238.165 21.000 239.585 22.000 ;
    LAYER MET3 ;
    RECT 231.180 0.000 232.600 22.000 ;
    LAYER MET3 ;
    RECT 288.100 0.000 289.520 22.000 ;
    LAYER VIA2 ;
    RECT 231.500 0.190 232.280 9.810 ;
    LAYER VIA2 ;
    RECT 288.420 0.190 289.200 9.810 ;
    LAYER MET3 ;
    RECT 222.590 0.000 223.490 22.000 ;
    LAYER MET3 ;
    RECT 279.510 0.000 280.410 22.000 ;
    LAYER VIA2 ;
    RECT 222.910 0.190 223.170 9.810 ;
    LAYER VIA2 ;
    RECT 279.830 0.190 280.090 9.810 ;
    LAYER MET3 ;
    RECT 213.135 0.000 214.555 22.000 ;
    LAYER MET3 ;
    RECT 270.055 0.000 271.475 22.000 ;
    LAYER VIA2 ;
    RECT 213.455 0.190 214.235 9.810 ;
    LAYER VIA2 ;
    RECT 270.375 0.190 271.155 9.810 ;
    LAYER MET2 ;
    RECT 235.610 21.000 236.510 22.000 ;
    LAYER MET2 ;
    RECT 292.530 21.000 293.430 22.000 ;
    LAYER MET2 ;
    RECT 218.695 21.000 220.115 22.000 ;
    LAYER MET2 ;
    RECT 275.615 21.000 277.035 22.000 ;
    LAYER MET2 ;
    RECT 216.525 21.000 217.425 22.000 ;
    LAYER MET2 ;
    RECT 273.445 21.000 274.345 22.000 ;
    LAYER MET2 ;
    RECT 209.705 21.000 211.125 22.000 ;
    LAYER MET2 ;
    RECT 266.625 21.000 268.045 22.000 ;
    LAYER MET2 ;
    RECT 295.760 47.985 317.760 48.885 ;
    LAYER VIA2 ;
    RECT 307.900 48.305 317.520 48.565 ;
    LAYER MET2 ;
    RECT 295.760 26.020 317.760 28.470 ;
    LAYER VIA2 ;
    RECT 307.900 26.335 317.520 28.155 ;
    LAYER MET2 ;
    RECT 295.760 35.140 317.760 37.340 ;
    LAYER VIA2 ;
    RECT 307.900 35.330 317.520 37.150 ;
    LAYER MET2 ;
    RECT 295.760 41.680 317.760 43.640 ;
    LAYER VIA2 ;
    RECT 307.900 42.010 317.520 43.310 ;
    LAYER MET2 ;
    RECT 295.760 45.940 317.760 46.480 ;
    LAYER VIA2 ;
    RECT 307.900 46.080 317.520 46.340 ;
    LAYER MET2 ;
    RECT 295.760 56.850 317.760 57.750 ;
    LAYER VIA2 ;
    RECT 307.900 57.170 317.520 57.430 ;
    LAYER MET2 ;
    RECT 295.760 84.965 317.760 86.315 ;
    LAYER VIA2 ;
    RECT 307.900 85.250 317.520 86.030 ;
    LAYER MET2 ;
    RECT 295.760 79.895 317.760 81.495 ;
    LAYER VIA2 ;
    RECT 307.900 80.045 317.520 81.345 ;
    LAYER MET2 ;
    RECT 295.760 72.430 317.760 73.330 ;
    LAYER VIA2 ;
    RECT 307.900 72.750 317.520 73.010 ;
    LAYER MET2 ;
    RECT 295.760 63.700 317.760 65.130 ;
    LAYER VIA2 ;
    RECT 307.900 64.025 317.520 64.805 ;
    LAYER MET3 ;
    RECT 295.760 22.740 296.760 23.840 ;
    LAYER MET3 ;
    RECT 295.760 31.540 296.760 32.840 ;
    LAYER MET3 ;
    RECT 295.760 37.840 296.760 39.140 ;
    LAYER MET3 ;
    RECT 295.760 44.900 296.760 45.440 ;
    LAYER MET3 ;
    RECT 295.760 51.950 296.760 52.850 ;
    LAYER MET3 ;
    RECT 295.760 60.000 296.760 61.400 ;
    LAYER MET3 ;
    RECT 295.760 70.955 296.760 71.855 ;
    LAYER MET3 ;
    RECT 295.760 88.405 296.760 89.405 ;
    LAYER MET2 ;
    RECT 0.000 90.810 22.000 91.350 ;
    LAYER VIA2 ;
    RECT 0.140 90.950 9.760 91.210 ;
    LAYER MET2 ;
    RECT 0.000 95.570 22.000 96.110 ;
    LAYER VIA2 ;
    RECT 0.140 95.710 9.760 95.970 ;
    LAYER MET2 ;
    RECT 0.000 90.810 22.000 91.350 ;
    LAYER VIA2 ;
    RECT 0.140 90.950 9.760 91.210 ;
    LAYER MET3 ;
    RECT 21.000 94.130 22.000 95.110 ;
    LAYER MET3 ;
    RECT 21.000 91.810 22.000 92.790 ;
    LAYER MET2 ;
    RECT 0.000 100.330 22.000 100.870 ;
    LAYER MET2 ;
    RECT 0.000 105.090 22.000 105.630 ;
    LAYER MET2 ;
    RECT 0.000 109.850 22.000 110.390 ;
    LAYER MET2 ;
    RECT 0.000 114.610 22.000 115.150 ;
    LAYER MET2 ;
    RECT 0.000 119.370 22.000 119.910 ;
    LAYER MET2 ;
    RECT 0.000 124.130 22.000 124.670 ;
    LAYER MET2 ;
    RECT 0.000 128.890 22.000 129.430 ;
    LAYER MET2 ;
    RECT 0.000 133.650 22.000 134.190 ;
    LAYER MET2 ;
    RECT 0.000 138.410 22.000 138.950 ;
    LAYER MET2 ;
    RECT 0.000 143.170 22.000 143.710 ;
    LAYER MET2 ;
    RECT 0.000 147.930 22.000 148.470 ;
    LAYER MET2 ;
    RECT 0.000 152.690 22.000 153.230 ;
    LAYER MET2 ;
    RECT 0.000 157.450 22.000 157.990 ;
    LAYER MET2 ;
    RECT 0.000 162.210 22.000 162.750 ;
    LAYER MET2 ;
    RECT 0.000 166.970 22.000 167.510 ;
    LAYER MET2 ;
    RECT 0.000 171.730 22.000 172.270 ;
    LAYER MET2 ;
    RECT 0.000 176.490 22.000 177.030 ;
    LAYER MET2 ;
    RECT 0.000 181.250 22.000 181.790 ;
    LAYER MET2 ;
    RECT 0.000 186.010 22.000 186.550 ;
    LAYER MET2 ;
    RECT 0.000 190.770 22.000 191.310 ;
    LAYER MET2 ;
    RECT 0.000 195.530 22.000 196.070 ;
    LAYER MET2 ;
    RECT 0.000 200.290 22.000 200.830 ;
    LAYER MET2 ;
    RECT 0.000 205.050 22.000 205.590 ;
    LAYER MET2 ;
    RECT 0.000 209.810 22.000 210.350 ;
    LAYER MET2 ;
    RECT 0.000 214.570 22.000 215.110 ;
    LAYER MET2 ;
    RECT 0.000 219.330 22.000 219.870 ;
    LAYER MET2 ;
    RECT 0.000 224.090 22.000 224.630 ;
    LAYER MET2 ;
    RECT 0.000 228.850 22.000 229.390 ;
    LAYER MET2 ;
    RECT 0.000 233.610 22.000 234.150 ;
    LAYER MET2 ;
    RECT 0.000 238.370 22.000 238.910 ;
    LAYER MET2 ;
    RECT 0.000 243.130 22.000 243.670 ;
    LAYER MET2 ;
    RECT 0.000 247.890 22.000 248.430 ;
    LAYER MET2 ;
    RECT 0.000 252.650 22.000 253.190 ;
    LAYER MET2 ;
    RECT 0.000 257.410 22.000 257.950 ;
    LAYER MET2 ;
    RECT 0.000 262.170 22.000 262.710 ;
    LAYER MET2 ;
    RECT 0.000 266.930 22.000 267.470 ;
    LAYER MET2 ;
    RECT 0.000 271.690 22.000 272.230 ;
    LAYER MET2 ;
    RECT 0.000 276.450 22.000 276.990 ;
    LAYER MET2 ;
    RECT 0.000 281.210 22.000 281.750 ;
    LAYER MET2 ;
    RECT 0.000 285.970 22.000 286.510 ;
    LAYER MET2 ;
    RECT 0.000 290.730 22.000 291.270 ;
    LAYER MET2 ;
    RECT 0.000 295.490 22.000 296.030 ;
    LAYER MET2 ;
    RECT 0.000 300.250 22.000 300.790 ;
    LAYER MET2 ;
    RECT 0.000 305.010 22.000 305.550 ;
    LAYER MET2 ;
    RECT 0.000 309.770 22.000 310.310 ;
    LAYER MET2 ;
    RECT 0.000 314.530 22.000 315.070 ;
    LAYER MET2 ;
    RECT 0.000 319.290 22.000 319.830 ;
    LAYER VIA2 ;
    RECT 0.140 100.470 9.760 100.730 ;
    LAYER VIA2 ;
    RECT 0.140 105.230 9.760 105.490 ;
    LAYER VIA2 ;
    RECT 0.140 109.990 9.760 110.250 ;
    LAYER VIA2 ;
    RECT 0.140 114.750 9.760 115.010 ;
    LAYER VIA2 ;
    RECT 0.140 119.510 9.760 119.770 ;
    LAYER VIA2 ;
    RECT 0.140 124.270 9.760 124.530 ;
    LAYER VIA2 ;
    RECT 0.140 129.030 9.760 129.290 ;
    LAYER VIA2 ;
    RECT 0.140 133.790 9.760 134.050 ;
    LAYER VIA2 ;
    RECT 0.140 138.550 9.760 138.810 ;
    LAYER VIA2 ;
    RECT 0.140 143.310 9.760 143.570 ;
    LAYER VIA2 ;
    RECT 0.140 148.070 9.760 148.330 ;
    LAYER VIA2 ;
    RECT 0.140 152.830 9.760 153.090 ;
    LAYER VIA2 ;
    RECT 0.140 157.590 9.760 157.850 ;
    LAYER VIA2 ;
    RECT 0.140 162.350 9.760 162.610 ;
    LAYER VIA2 ;
    RECT 0.140 167.110 9.760 167.370 ;
    LAYER VIA2 ;
    RECT 0.140 171.870 9.760 172.130 ;
    LAYER VIA2 ;
    RECT 0.140 176.630 9.760 176.890 ;
    LAYER VIA2 ;
    RECT 0.140 181.390 9.760 181.650 ;
    LAYER VIA2 ;
    RECT 0.140 186.150 9.760 186.410 ;
    LAYER VIA2 ;
    RECT 0.140 190.910 9.760 191.170 ;
    LAYER VIA2 ;
    RECT 0.140 195.670 9.760 195.930 ;
    LAYER VIA2 ;
    RECT 0.140 200.430 9.760 200.690 ;
    LAYER VIA2 ;
    RECT 0.140 205.190 9.760 205.450 ;
    LAYER VIA2 ;
    RECT 0.140 209.950 9.760 210.210 ;
    LAYER VIA2 ;
    RECT 0.140 214.710 9.760 214.970 ;
    LAYER VIA2 ;
    RECT 0.140 219.470 9.760 219.730 ;
    LAYER VIA2 ;
    RECT 0.140 224.230 9.760 224.490 ;
    LAYER VIA2 ;
    RECT 0.140 228.990 9.760 229.250 ;
    LAYER VIA2 ;
    RECT 0.140 233.750 9.760 234.010 ;
    LAYER VIA2 ;
    RECT 0.140 238.510 9.760 238.770 ;
    LAYER VIA2 ;
    RECT 0.140 243.270 9.760 243.530 ;
    LAYER VIA2 ;
    RECT 0.140 248.030 9.760 248.290 ;
    LAYER VIA2 ;
    RECT 0.140 252.790 9.760 253.050 ;
    LAYER VIA2 ;
    RECT 0.140 257.550 9.760 257.810 ;
    LAYER VIA2 ;
    RECT 0.140 262.310 9.760 262.570 ;
    LAYER VIA2 ;
    RECT 0.140 267.070 9.760 267.330 ;
    LAYER VIA2 ;
    RECT 0.140 271.830 9.760 272.090 ;
    LAYER VIA2 ;
    RECT 0.140 276.590 9.760 276.850 ;
    LAYER VIA2 ;
    RECT 0.140 281.350 9.760 281.610 ;
    LAYER VIA2 ;
    RECT 0.140 286.110 9.760 286.370 ;
    LAYER VIA2 ;
    RECT 0.140 290.870 9.760 291.130 ;
    LAYER VIA2 ;
    RECT 0.140 295.630 9.760 295.890 ;
    LAYER VIA2 ;
    RECT 0.140 300.390 9.760 300.650 ;
    LAYER VIA2 ;
    RECT 0.140 305.150 9.760 305.410 ;
    LAYER VIA2 ;
    RECT 0.140 309.910 9.760 310.170 ;
    LAYER VIA2 ;
    RECT 0.140 314.670 9.760 314.930 ;
    LAYER VIA2 ;
    RECT 0.140 319.430 9.760 319.690 ;
    LAYER MET2 ;
    RECT 0.000 95.570 22.000 96.110 ;
    LAYER MET2 ;
    RECT 0.000 100.330 22.000 100.870 ;
    LAYER MET2 ;
    RECT 0.000 105.090 22.000 105.630 ;
    LAYER MET2 ;
    RECT 0.000 109.850 22.000 110.390 ;
    LAYER MET2 ;
    RECT 0.000 114.610 22.000 115.150 ;
    LAYER MET2 ;
    RECT 0.000 119.370 22.000 119.910 ;
    LAYER MET2 ;
    RECT 0.000 124.130 22.000 124.670 ;
    LAYER MET2 ;
    RECT 0.000 128.890 22.000 129.430 ;
    LAYER MET2 ;
    RECT 0.000 133.650 22.000 134.190 ;
    LAYER MET2 ;
    RECT 0.000 138.410 22.000 138.950 ;
    LAYER MET2 ;
    RECT 0.000 143.170 22.000 143.710 ;
    LAYER MET2 ;
    RECT 0.000 147.930 22.000 148.470 ;
    LAYER MET2 ;
    RECT 0.000 152.690 22.000 153.230 ;
    LAYER MET2 ;
    RECT 0.000 157.450 22.000 157.990 ;
    LAYER MET2 ;
    RECT 0.000 162.210 22.000 162.750 ;
    LAYER MET2 ;
    RECT 0.000 166.970 22.000 167.510 ;
    LAYER MET2 ;
    RECT 0.000 171.730 22.000 172.270 ;
    LAYER MET2 ;
    RECT 0.000 176.490 22.000 177.030 ;
    LAYER MET2 ;
    RECT 0.000 181.250 22.000 181.790 ;
    LAYER MET2 ;
    RECT 0.000 186.010 22.000 186.550 ;
    LAYER MET2 ;
    RECT 0.000 190.770 22.000 191.310 ;
    LAYER MET2 ;
    RECT 0.000 195.530 22.000 196.070 ;
    LAYER MET2 ;
    RECT 0.000 200.290 22.000 200.830 ;
    LAYER MET2 ;
    RECT 0.000 205.050 22.000 205.590 ;
    LAYER MET2 ;
    RECT 0.000 209.810 22.000 210.350 ;
    LAYER MET2 ;
    RECT 0.000 214.570 22.000 215.110 ;
    LAYER MET2 ;
    RECT 0.000 219.330 22.000 219.870 ;
    LAYER MET2 ;
    RECT 0.000 224.090 22.000 224.630 ;
    LAYER MET2 ;
    RECT 0.000 228.850 22.000 229.390 ;
    LAYER MET2 ;
    RECT 0.000 233.610 22.000 234.150 ;
    LAYER MET2 ;
    RECT 0.000 238.370 22.000 238.910 ;
    LAYER MET2 ;
    RECT 0.000 243.130 22.000 243.670 ;
    LAYER MET2 ;
    RECT 0.000 247.890 22.000 248.430 ;
    LAYER MET2 ;
    RECT 0.000 252.650 22.000 253.190 ;
    LAYER MET2 ;
    RECT 0.000 257.410 22.000 257.950 ;
    LAYER MET2 ;
    RECT 0.000 262.170 22.000 262.710 ;
    LAYER MET2 ;
    RECT 0.000 266.930 22.000 267.470 ;
    LAYER MET2 ;
    RECT 0.000 271.690 22.000 272.230 ;
    LAYER MET2 ;
    RECT 0.000 276.450 22.000 276.990 ;
    LAYER MET2 ;
    RECT 0.000 281.210 22.000 281.750 ;
    LAYER MET2 ;
    RECT 0.000 285.970 22.000 286.510 ;
    LAYER MET2 ;
    RECT 0.000 290.730 22.000 291.270 ;
    LAYER MET2 ;
    RECT 0.000 295.490 22.000 296.030 ;
    LAYER MET2 ;
    RECT 0.000 300.250 22.000 300.790 ;
    LAYER MET2 ;
    RECT 0.000 305.010 22.000 305.550 ;
    LAYER MET2 ;
    RECT 0.000 309.770 22.000 310.310 ;
    LAYER MET2 ;
    RECT 0.000 314.530 22.000 315.070 ;
    LAYER VIA2 ;
    RECT 0.140 95.710 9.760 95.970 ;
    LAYER VIA2 ;
    RECT 0.140 100.470 9.760 100.730 ;
    LAYER VIA2 ;
    RECT 0.140 105.230 9.760 105.490 ;
    LAYER VIA2 ;
    RECT 0.140 109.990 9.760 110.250 ;
    LAYER VIA2 ;
    RECT 0.140 114.750 9.760 115.010 ;
    LAYER VIA2 ;
    RECT 0.140 119.510 9.760 119.770 ;
    LAYER VIA2 ;
    RECT 0.140 124.270 9.760 124.530 ;
    LAYER VIA2 ;
    RECT 0.140 129.030 9.760 129.290 ;
    LAYER VIA2 ;
    RECT 0.140 133.790 9.760 134.050 ;
    LAYER VIA2 ;
    RECT 0.140 138.550 9.760 138.810 ;
    LAYER VIA2 ;
    RECT 0.140 143.310 9.760 143.570 ;
    LAYER VIA2 ;
    RECT 0.140 148.070 9.760 148.330 ;
    LAYER VIA2 ;
    RECT 0.140 152.830 9.760 153.090 ;
    LAYER VIA2 ;
    RECT 0.140 157.590 9.760 157.850 ;
    LAYER VIA2 ;
    RECT 0.140 162.350 9.760 162.610 ;
    LAYER VIA2 ;
    RECT 0.140 167.110 9.760 167.370 ;
    LAYER VIA2 ;
    RECT 0.140 171.870 9.760 172.130 ;
    LAYER VIA2 ;
    RECT 0.140 176.630 9.760 176.890 ;
    LAYER VIA2 ;
    RECT 0.140 181.390 9.760 181.650 ;
    LAYER VIA2 ;
    RECT 0.140 186.150 9.760 186.410 ;
    LAYER VIA2 ;
    RECT 0.140 190.910 9.760 191.170 ;
    LAYER VIA2 ;
    RECT 0.140 195.670 9.760 195.930 ;
    LAYER VIA2 ;
    RECT 0.140 200.430 9.760 200.690 ;
    LAYER VIA2 ;
    RECT 0.140 205.190 9.760 205.450 ;
    LAYER VIA2 ;
    RECT 0.140 209.950 9.760 210.210 ;
    LAYER VIA2 ;
    RECT 0.140 214.710 9.760 214.970 ;
    LAYER VIA2 ;
    RECT 0.140 219.470 9.760 219.730 ;
    LAYER VIA2 ;
    RECT 0.140 224.230 9.760 224.490 ;
    LAYER VIA2 ;
    RECT 0.140 228.990 9.760 229.250 ;
    LAYER VIA2 ;
    RECT 0.140 233.750 9.760 234.010 ;
    LAYER VIA2 ;
    RECT 0.140 238.510 9.760 238.770 ;
    LAYER VIA2 ;
    RECT 0.140 243.270 9.760 243.530 ;
    LAYER VIA2 ;
    RECT 0.140 248.030 9.760 248.290 ;
    LAYER VIA2 ;
    RECT 0.140 252.790 9.760 253.050 ;
    LAYER VIA2 ;
    RECT 0.140 257.550 9.760 257.810 ;
    LAYER VIA2 ;
    RECT 0.140 262.310 9.760 262.570 ;
    LAYER VIA2 ;
    RECT 0.140 267.070 9.760 267.330 ;
    LAYER VIA2 ;
    RECT 0.140 271.830 9.760 272.090 ;
    LAYER VIA2 ;
    RECT 0.140 276.590 9.760 276.850 ;
    LAYER VIA2 ;
    RECT 0.140 281.350 9.760 281.610 ;
    LAYER VIA2 ;
    RECT 0.140 286.110 9.760 286.370 ;
    LAYER VIA2 ;
    RECT 0.140 290.870 9.760 291.130 ;
    LAYER VIA2 ;
    RECT 0.140 295.630 9.760 295.890 ;
    LAYER VIA2 ;
    RECT 0.140 300.390 9.760 300.650 ;
    LAYER VIA2 ;
    RECT 0.140 305.150 9.760 305.410 ;
    LAYER VIA2 ;
    RECT 0.140 309.910 9.760 310.170 ;
    LAYER VIA2 ;
    RECT 0.140 314.670 9.760 314.930 ;
    LAYER MET3 ;
    RECT 21.000 98.890 22.000 99.870 ;
    LAYER MET3 ;
    RECT 21.000 103.650 22.000 104.630 ;
    LAYER MET3 ;
    RECT 21.000 108.410 22.000 109.390 ;
    LAYER MET3 ;
    RECT 21.000 113.170 22.000 114.150 ;
    LAYER MET3 ;
    RECT 21.000 117.930 22.000 118.910 ;
    LAYER MET3 ;
    RECT 21.000 122.690 22.000 123.670 ;
    LAYER MET3 ;
    RECT 21.000 127.450 22.000 128.430 ;
    LAYER MET3 ;
    RECT 21.000 132.210 22.000 133.190 ;
    LAYER MET3 ;
    RECT 21.000 136.970 22.000 137.950 ;
    LAYER MET3 ;
    RECT 21.000 141.730 22.000 142.710 ;
    LAYER MET3 ;
    RECT 21.000 146.490 22.000 147.470 ;
    LAYER MET3 ;
    RECT 21.000 151.250 22.000 152.230 ;
    LAYER MET3 ;
    RECT 21.000 156.010 22.000 156.990 ;
    LAYER MET3 ;
    RECT 21.000 160.770 22.000 161.750 ;
    LAYER MET3 ;
    RECT 21.000 165.530 22.000 166.510 ;
    LAYER MET3 ;
    RECT 21.000 170.290 22.000 171.270 ;
    LAYER MET3 ;
    RECT 21.000 175.050 22.000 176.030 ;
    LAYER MET3 ;
    RECT 21.000 179.810 22.000 180.790 ;
    LAYER MET3 ;
    RECT 21.000 184.570 22.000 185.550 ;
    LAYER MET3 ;
    RECT 21.000 189.330 22.000 190.310 ;
    LAYER MET3 ;
    RECT 21.000 194.090 22.000 195.070 ;
    LAYER MET3 ;
    RECT 21.000 198.850 22.000 199.830 ;
    LAYER MET3 ;
    RECT 21.000 203.610 22.000 204.590 ;
    LAYER MET3 ;
    RECT 21.000 208.370 22.000 209.350 ;
    LAYER MET3 ;
    RECT 21.000 213.130 22.000 214.110 ;
    LAYER MET3 ;
    RECT 21.000 217.890 22.000 218.870 ;
    LAYER MET3 ;
    RECT 21.000 222.650 22.000 223.630 ;
    LAYER MET3 ;
    RECT 21.000 227.410 22.000 228.390 ;
    LAYER MET3 ;
    RECT 21.000 232.170 22.000 233.150 ;
    LAYER MET3 ;
    RECT 21.000 236.930 22.000 237.910 ;
    LAYER MET3 ;
    RECT 21.000 241.690 22.000 242.670 ;
    LAYER MET3 ;
    RECT 21.000 246.450 22.000 247.430 ;
    LAYER MET3 ;
    RECT 21.000 251.210 22.000 252.190 ;
    LAYER MET3 ;
    RECT 21.000 255.970 22.000 256.950 ;
    LAYER MET3 ;
    RECT 21.000 260.730 22.000 261.710 ;
    LAYER MET3 ;
    RECT 21.000 265.490 22.000 266.470 ;
    LAYER MET3 ;
    RECT 21.000 270.250 22.000 271.230 ;
    LAYER MET3 ;
    RECT 21.000 275.010 22.000 275.990 ;
    LAYER MET3 ;
    RECT 21.000 279.770 22.000 280.750 ;
    LAYER MET3 ;
    RECT 21.000 284.530 22.000 285.510 ;
    LAYER MET3 ;
    RECT 21.000 289.290 22.000 290.270 ;
    LAYER MET3 ;
    RECT 21.000 294.050 22.000 295.030 ;
    LAYER MET3 ;
    RECT 21.000 298.810 22.000 299.790 ;
    LAYER MET3 ;
    RECT 21.000 303.570 22.000 304.550 ;
    LAYER MET3 ;
    RECT 21.000 308.330 22.000 309.310 ;
    LAYER MET3 ;
    RECT 21.000 313.090 22.000 314.070 ;
    LAYER MET3 ;
    RECT 21.000 317.850 22.000 318.830 ;
    LAYER MET3 ;
    RECT 21.000 96.570 22.000 97.550 ;
    LAYER MET3 ;
    RECT 21.000 101.330 22.000 102.310 ;
    LAYER MET3 ;
    RECT 21.000 106.090 22.000 107.070 ;
    LAYER MET3 ;
    RECT 21.000 110.850 22.000 111.830 ;
    LAYER MET3 ;
    RECT 21.000 115.610 22.000 116.590 ;
    LAYER MET3 ;
    RECT 21.000 120.370 22.000 121.350 ;
    LAYER MET3 ;
    RECT 21.000 125.130 22.000 126.110 ;
    LAYER MET3 ;
    RECT 21.000 129.890 22.000 130.870 ;
    LAYER MET3 ;
    RECT 21.000 134.650 22.000 135.630 ;
    LAYER MET3 ;
    RECT 21.000 139.410 22.000 140.390 ;
    LAYER MET3 ;
    RECT 21.000 144.170 22.000 145.150 ;
    LAYER MET3 ;
    RECT 21.000 148.930 22.000 149.910 ;
    LAYER MET3 ;
    RECT 21.000 153.690 22.000 154.670 ;
    LAYER MET3 ;
    RECT 21.000 158.450 22.000 159.430 ;
    LAYER MET3 ;
    RECT 21.000 163.210 22.000 164.190 ;
    LAYER MET3 ;
    RECT 21.000 167.970 22.000 168.950 ;
    LAYER MET3 ;
    RECT 21.000 172.730 22.000 173.710 ;
    LAYER MET3 ;
    RECT 21.000 177.490 22.000 178.470 ;
    LAYER MET3 ;
    RECT 21.000 182.250 22.000 183.230 ;
    LAYER MET3 ;
    RECT 21.000 187.010 22.000 187.990 ;
    LAYER MET3 ;
    RECT 21.000 191.770 22.000 192.750 ;
    LAYER MET3 ;
    RECT 21.000 196.530 22.000 197.510 ;
    LAYER MET3 ;
    RECT 21.000 201.290 22.000 202.270 ;
    LAYER MET3 ;
    RECT 21.000 206.050 22.000 207.030 ;
    LAYER MET3 ;
    RECT 21.000 210.810 22.000 211.790 ;
    LAYER MET3 ;
    RECT 21.000 215.570 22.000 216.550 ;
    LAYER MET3 ;
    RECT 21.000 220.330 22.000 221.310 ;
    LAYER MET3 ;
    RECT 21.000 225.090 22.000 226.070 ;
    LAYER MET3 ;
    RECT 21.000 229.850 22.000 230.830 ;
    LAYER MET3 ;
    RECT 21.000 234.610 22.000 235.590 ;
    LAYER MET3 ;
    RECT 21.000 239.370 22.000 240.350 ;
    LAYER MET3 ;
    RECT 21.000 244.130 22.000 245.110 ;
    LAYER MET3 ;
    RECT 21.000 248.890 22.000 249.870 ;
    LAYER MET3 ;
    RECT 21.000 253.650 22.000 254.630 ;
    LAYER MET3 ;
    RECT 21.000 258.410 22.000 259.390 ;
    LAYER MET3 ;
    RECT 21.000 263.170 22.000 264.150 ;
    LAYER MET3 ;
    RECT 21.000 267.930 22.000 268.910 ;
    LAYER MET3 ;
    RECT 21.000 272.690 22.000 273.670 ;
    LAYER MET3 ;
    RECT 21.000 277.450 22.000 278.430 ;
    LAYER MET3 ;
    RECT 21.000 282.210 22.000 283.190 ;
    LAYER MET3 ;
    RECT 21.000 286.970 22.000 287.950 ;
    LAYER MET3 ;
    RECT 21.000 291.730 22.000 292.710 ;
    LAYER MET3 ;
    RECT 21.000 296.490 22.000 297.470 ;
    LAYER MET3 ;
    RECT 21.000 301.250 22.000 302.230 ;
    LAYER MET3 ;
    RECT 21.000 306.010 22.000 306.990 ;
    LAYER MET3 ;
    RECT 21.000 310.770 22.000 311.750 ;
    LAYER MET3 ;
    RECT 21.000 315.530 22.000 316.510 ;
    LAYER MET2 ;
    RECT 0.000 319.290 22.000 319.830 ;
    LAYER VIA2 ;
    RECT 0.140 319.430 9.760 319.690 ;
    LAYER MET2 ;
    RECT 0.000 324.050 22.000 324.590 ;
    LAYER VIA2 ;
    RECT 0.140 324.190 9.760 324.450 ;
    LAYER MET3 ;
    RECT 21.000 320.290 22.000 321.270 ;
    LAYER MET3 ;
    RECT 21.000 322.610 22.000 323.590 ;
    LAYER MET2 ;
    RECT 0.000 324.050 22.000 324.590 ;
    LAYER VIA2 ;
    RECT 0.140 324.190 9.760 324.450 ;
    LAYER MET3 ;
    RECT 37.575 326.410 38.405 348.410 ;
    LAYER MET3 ;
    RECT 94.495 326.410 95.325 348.410 ;
    LAYER VIA2 ;
    RECT 37.860 338.600 38.120 348.220 ;
    LAYER VIA2 ;
    RECT 94.780 338.600 95.040 348.220 ;
    LAYER MET2 ;
    RECT 66.035 326.410 66.865 327.410 ;
    LAYER MET2 ;
    RECT 122.955 326.410 123.785 327.410 ;
    LAYER MET3 ;
    RECT 136.970 326.410 138.220 348.410 ;
    LAYER VIA2 ;
    RECT 137.205 338.600 137.985 348.220 ;
    LAYER MET2 ;
    RECT 138.680 326.410 139.930 327.410 ;
    LAYER MET3 ;
    RECT 144.660 326.410 145.260 348.410 ;
    LAYER VIA2 ;
    RECT 144.830 338.600 145.090 348.220 ;
    LAYER MET2 ;
    RECT 143.600 326.410 144.200 327.410 ;
    LAYER MET3 ;
    RECT 165.830 326.410 169.040 348.410 ;
    LAYER VIA2 ;
    RECT 166.005 338.600 168.865 348.220 ;
    LAYER MET3 ;
    RECT 162.430 326.410 163.850 348.410 ;
    LAYER VIA2 ;
    RECT 162.750 338.600 163.530 348.220 ;
    LAYER MET3 ;
    RECT 154.430 326.410 155.030 348.410 ;
    LAYER VIA2 ;
    RECT 154.600 338.600 154.860 348.220 ;
    LAYER MET2 ;
    RECT 174.200 326.410 175.100 327.410 ;
    LAYER MET2 ;
    RECT 169.840 326.410 170.740 327.410 ;
    LAYER MET2 ;
    RECT 171.380 326.410 173.340 327.410 ;
    LAYER MET2 ;
    RECT 159.830 326.410 161.630 327.410 ;
    LAYER MET2 ;
    RECT 153.370 326.410 153.970 327.410 ;
    LAYER MET2 ;
    RECT 295.760 90.810 317.760 91.350 ;
    LAYER VIA2 ;
    RECT 307.900 90.950 317.520 91.210 ;
    LAYER MET2 ;
    RECT 295.760 90.810 317.760 91.350 ;
    LAYER VIA2 ;
    RECT 307.900 90.950 317.520 91.210 ;
    LAYER MET2 ;
    RECT 295.760 95.570 317.760 96.110 ;
    LAYER VIA2 ;
    RECT 307.900 95.710 317.520 95.970 ;
    LAYER MET3 ;
    RECT 295.760 91.810 296.760 92.790 ;
    LAYER MET3 ;
    RECT 295.760 94.130 296.760 95.110 ;
    LAYER MET2 ;
    RECT 295.760 95.570 317.760 96.110 ;
    LAYER MET2 ;
    RECT 295.760 100.330 317.760 100.870 ;
    LAYER MET2 ;
    RECT 295.760 105.090 317.760 105.630 ;
    LAYER MET2 ;
    RECT 295.760 109.850 317.760 110.390 ;
    LAYER MET2 ;
    RECT 295.760 114.610 317.760 115.150 ;
    LAYER MET2 ;
    RECT 295.760 119.370 317.760 119.910 ;
    LAYER MET2 ;
    RECT 295.760 124.130 317.760 124.670 ;
    LAYER MET2 ;
    RECT 295.760 128.890 317.760 129.430 ;
    LAYER MET2 ;
    RECT 295.760 133.650 317.760 134.190 ;
    LAYER MET2 ;
    RECT 295.760 138.410 317.760 138.950 ;
    LAYER MET2 ;
    RECT 295.760 143.170 317.760 143.710 ;
    LAYER MET2 ;
    RECT 295.760 147.930 317.760 148.470 ;
    LAYER MET2 ;
    RECT 295.760 152.690 317.760 153.230 ;
    LAYER MET2 ;
    RECT 295.760 157.450 317.760 157.990 ;
    LAYER MET2 ;
    RECT 295.760 162.210 317.760 162.750 ;
    LAYER MET2 ;
    RECT 295.760 166.970 317.760 167.510 ;
    LAYER MET2 ;
    RECT 295.760 171.730 317.760 172.270 ;
    LAYER MET2 ;
    RECT 295.760 176.490 317.760 177.030 ;
    LAYER MET2 ;
    RECT 295.760 181.250 317.760 181.790 ;
    LAYER MET2 ;
    RECT 295.760 186.010 317.760 186.550 ;
    LAYER MET2 ;
    RECT 295.760 190.770 317.760 191.310 ;
    LAYER MET2 ;
    RECT 295.760 195.530 317.760 196.070 ;
    LAYER MET2 ;
    RECT 295.760 200.290 317.760 200.830 ;
    LAYER MET2 ;
    RECT 295.760 205.050 317.760 205.590 ;
    LAYER MET2 ;
    RECT 295.760 209.810 317.760 210.350 ;
    LAYER MET2 ;
    RECT 295.760 214.570 317.760 215.110 ;
    LAYER MET2 ;
    RECT 295.760 219.330 317.760 219.870 ;
    LAYER MET2 ;
    RECT 295.760 224.090 317.760 224.630 ;
    LAYER MET2 ;
    RECT 295.760 228.850 317.760 229.390 ;
    LAYER MET2 ;
    RECT 295.760 233.610 317.760 234.150 ;
    LAYER MET2 ;
    RECT 295.760 238.370 317.760 238.910 ;
    LAYER MET2 ;
    RECT 295.760 243.130 317.760 243.670 ;
    LAYER MET2 ;
    RECT 295.760 247.890 317.760 248.430 ;
    LAYER MET2 ;
    RECT 295.760 252.650 317.760 253.190 ;
    LAYER MET2 ;
    RECT 295.760 257.410 317.760 257.950 ;
    LAYER MET2 ;
    RECT 295.760 262.170 317.760 262.710 ;
    LAYER MET2 ;
    RECT 295.760 266.930 317.760 267.470 ;
    LAYER MET2 ;
    RECT 295.760 271.690 317.760 272.230 ;
    LAYER MET2 ;
    RECT 295.760 276.450 317.760 276.990 ;
    LAYER VIA2 ;
    RECT 307.900 95.710 317.520 95.970 ;
    LAYER VIA2 ;
    RECT 307.900 100.470 317.520 100.730 ;
    LAYER VIA2 ;
    RECT 307.900 105.230 317.520 105.490 ;
    LAYER VIA2 ;
    RECT 307.900 109.990 317.520 110.250 ;
    LAYER VIA2 ;
    RECT 307.900 114.750 317.520 115.010 ;
    LAYER VIA2 ;
    RECT 307.900 119.510 317.520 119.770 ;
    LAYER VIA2 ;
    RECT 307.900 124.270 317.520 124.530 ;
    LAYER VIA2 ;
    RECT 307.900 129.030 317.520 129.290 ;
    LAYER VIA2 ;
    RECT 307.900 133.790 317.520 134.050 ;
    LAYER VIA2 ;
    RECT 307.900 138.550 317.520 138.810 ;
    LAYER VIA2 ;
    RECT 307.900 143.310 317.520 143.570 ;
    LAYER VIA2 ;
    RECT 307.900 148.070 317.520 148.330 ;
    LAYER VIA2 ;
    RECT 307.900 152.830 317.520 153.090 ;
    LAYER VIA2 ;
    RECT 307.900 157.590 317.520 157.850 ;
    LAYER VIA2 ;
    RECT 307.900 162.350 317.520 162.610 ;
    LAYER VIA2 ;
    RECT 307.900 167.110 317.520 167.370 ;
    LAYER VIA2 ;
    RECT 307.900 171.870 317.520 172.130 ;
    LAYER VIA2 ;
    RECT 307.900 176.630 317.520 176.890 ;
    LAYER VIA2 ;
    RECT 307.900 181.390 317.520 181.650 ;
    LAYER VIA2 ;
    RECT 307.900 186.150 317.520 186.410 ;
    LAYER VIA2 ;
    RECT 307.900 190.910 317.520 191.170 ;
    LAYER VIA2 ;
    RECT 307.900 195.670 317.520 195.930 ;
    LAYER VIA2 ;
    RECT 307.900 200.430 317.520 200.690 ;
    LAYER VIA2 ;
    RECT 307.900 205.190 317.520 205.450 ;
    LAYER VIA2 ;
    RECT 307.900 209.950 317.520 210.210 ;
    LAYER VIA2 ;
    RECT 307.900 214.710 317.520 214.970 ;
    LAYER VIA2 ;
    RECT 307.900 219.470 317.520 219.730 ;
    LAYER VIA2 ;
    RECT 307.900 224.230 317.520 224.490 ;
    LAYER VIA2 ;
    RECT 307.900 228.990 317.520 229.250 ;
    LAYER VIA2 ;
    RECT 307.900 233.750 317.520 234.010 ;
    LAYER VIA2 ;
    RECT 307.900 238.510 317.520 238.770 ;
    LAYER VIA2 ;
    RECT 307.900 243.270 317.520 243.530 ;
    LAYER VIA2 ;
    RECT 307.900 248.030 317.520 248.290 ;
    LAYER VIA2 ;
    RECT 307.900 252.790 317.520 253.050 ;
    LAYER VIA2 ;
    RECT 307.900 257.550 317.520 257.810 ;
    LAYER VIA2 ;
    RECT 307.900 262.310 317.520 262.570 ;
    LAYER VIA2 ;
    RECT 307.900 267.070 317.520 267.330 ;
    LAYER VIA2 ;
    RECT 307.900 271.830 317.520 272.090 ;
    LAYER VIA2 ;
    RECT 307.900 276.590 317.520 276.850 ;
    LAYER MET2 ;
    RECT 295.760 100.330 317.760 100.870 ;
    LAYER MET2 ;
    RECT 295.760 105.090 317.760 105.630 ;
    LAYER MET2 ;
    RECT 295.760 109.850 317.760 110.390 ;
    LAYER MET2 ;
    RECT 295.760 114.610 317.760 115.150 ;
    LAYER MET2 ;
    RECT 295.760 119.370 317.760 119.910 ;
    LAYER MET2 ;
    RECT 295.760 124.130 317.760 124.670 ;
    LAYER MET2 ;
    RECT 295.760 128.890 317.760 129.430 ;
    LAYER MET2 ;
    RECT 295.760 133.650 317.760 134.190 ;
    LAYER MET2 ;
    RECT 295.760 138.410 317.760 138.950 ;
    LAYER MET2 ;
    RECT 295.760 143.170 317.760 143.710 ;
    LAYER MET2 ;
    RECT 295.760 147.930 317.760 148.470 ;
    LAYER MET2 ;
    RECT 295.760 152.690 317.760 153.230 ;
    LAYER MET2 ;
    RECT 295.760 157.450 317.760 157.990 ;
    LAYER MET2 ;
    RECT 295.760 162.210 317.760 162.750 ;
    LAYER MET2 ;
    RECT 295.760 166.970 317.760 167.510 ;
    LAYER MET2 ;
    RECT 295.760 171.730 317.760 172.270 ;
    LAYER MET2 ;
    RECT 295.760 176.490 317.760 177.030 ;
    LAYER MET2 ;
    RECT 295.760 181.250 317.760 181.790 ;
    LAYER MET2 ;
    RECT 295.760 186.010 317.760 186.550 ;
    LAYER MET2 ;
    RECT 295.760 190.770 317.760 191.310 ;
    LAYER MET2 ;
    RECT 295.760 195.530 317.760 196.070 ;
    LAYER MET2 ;
    RECT 295.760 200.290 317.760 200.830 ;
    LAYER MET2 ;
    RECT 295.760 205.050 317.760 205.590 ;
    LAYER MET2 ;
    RECT 295.760 209.810 317.760 210.350 ;
    LAYER MET2 ;
    RECT 295.760 214.570 317.760 215.110 ;
    LAYER MET2 ;
    RECT 295.760 219.330 317.760 219.870 ;
    LAYER MET2 ;
    RECT 295.760 224.090 317.760 224.630 ;
    LAYER MET2 ;
    RECT 295.760 228.850 317.760 229.390 ;
    LAYER MET2 ;
    RECT 295.760 233.610 317.760 234.150 ;
    LAYER MET2 ;
    RECT 295.760 238.370 317.760 238.910 ;
    LAYER MET2 ;
    RECT 295.760 243.130 317.760 243.670 ;
    LAYER MET2 ;
    RECT 295.760 247.890 317.760 248.430 ;
    LAYER MET2 ;
    RECT 295.760 252.650 317.760 253.190 ;
    LAYER MET2 ;
    RECT 295.760 257.410 317.760 257.950 ;
    LAYER MET2 ;
    RECT 295.760 262.170 317.760 262.710 ;
    LAYER MET2 ;
    RECT 295.760 266.930 317.760 267.470 ;
    LAYER MET2 ;
    RECT 295.760 271.690 317.760 272.230 ;
    LAYER MET2 ;
    RECT 295.760 276.450 317.760 276.990 ;
    LAYER MET2 ;
    RECT 295.760 281.210 317.760 281.750 ;
    LAYER VIA2 ;
    RECT 307.900 100.470 317.520 100.730 ;
    LAYER VIA2 ;
    RECT 307.900 105.230 317.520 105.490 ;
    LAYER VIA2 ;
    RECT 307.900 109.990 317.520 110.250 ;
    LAYER VIA2 ;
    RECT 307.900 114.750 317.520 115.010 ;
    LAYER VIA2 ;
    RECT 307.900 119.510 317.520 119.770 ;
    LAYER VIA2 ;
    RECT 307.900 124.270 317.520 124.530 ;
    LAYER VIA2 ;
    RECT 307.900 129.030 317.520 129.290 ;
    LAYER VIA2 ;
    RECT 307.900 133.790 317.520 134.050 ;
    LAYER VIA2 ;
    RECT 307.900 138.550 317.520 138.810 ;
    LAYER VIA2 ;
    RECT 307.900 143.310 317.520 143.570 ;
    LAYER VIA2 ;
    RECT 307.900 148.070 317.520 148.330 ;
    LAYER VIA2 ;
    RECT 307.900 152.830 317.520 153.090 ;
    LAYER VIA2 ;
    RECT 307.900 157.590 317.520 157.850 ;
    LAYER VIA2 ;
    RECT 307.900 162.350 317.520 162.610 ;
    LAYER VIA2 ;
    RECT 307.900 167.110 317.520 167.370 ;
    LAYER VIA2 ;
    RECT 307.900 171.870 317.520 172.130 ;
    LAYER VIA2 ;
    RECT 307.900 176.630 317.520 176.890 ;
    LAYER VIA2 ;
    RECT 307.900 181.390 317.520 181.650 ;
    LAYER VIA2 ;
    RECT 307.900 186.150 317.520 186.410 ;
    LAYER VIA2 ;
    RECT 307.900 190.910 317.520 191.170 ;
    LAYER VIA2 ;
    RECT 307.900 195.670 317.520 195.930 ;
    LAYER VIA2 ;
    RECT 307.900 200.430 317.520 200.690 ;
    LAYER VIA2 ;
    RECT 307.900 205.190 317.520 205.450 ;
    LAYER VIA2 ;
    RECT 307.900 209.950 317.520 210.210 ;
    LAYER VIA2 ;
    RECT 307.900 214.710 317.520 214.970 ;
    LAYER VIA2 ;
    RECT 307.900 219.470 317.520 219.730 ;
    LAYER VIA2 ;
    RECT 307.900 224.230 317.520 224.490 ;
    LAYER VIA2 ;
    RECT 307.900 228.990 317.520 229.250 ;
    LAYER VIA2 ;
    RECT 307.900 233.750 317.520 234.010 ;
    LAYER VIA2 ;
    RECT 307.900 238.510 317.520 238.770 ;
    LAYER VIA2 ;
    RECT 307.900 243.270 317.520 243.530 ;
    LAYER VIA2 ;
    RECT 307.900 248.030 317.520 248.290 ;
    LAYER VIA2 ;
    RECT 307.900 252.790 317.520 253.050 ;
    LAYER VIA2 ;
    RECT 307.900 257.550 317.520 257.810 ;
    LAYER VIA2 ;
    RECT 307.900 262.310 317.520 262.570 ;
    LAYER VIA2 ;
    RECT 307.900 267.070 317.520 267.330 ;
    LAYER VIA2 ;
    RECT 307.900 271.830 317.520 272.090 ;
    LAYER VIA2 ;
    RECT 307.900 276.590 317.520 276.850 ;
    LAYER VIA2 ;
    RECT 307.900 281.350 317.520 281.610 ;
    LAYER MET3 ;
    RECT 295.760 96.570 296.760 97.550 ;
    LAYER MET3 ;
    RECT 295.760 101.330 296.760 102.310 ;
    LAYER MET3 ;
    RECT 295.760 106.090 296.760 107.070 ;
    LAYER MET3 ;
    RECT 295.760 110.850 296.760 111.830 ;
    LAYER MET3 ;
    RECT 295.760 115.610 296.760 116.590 ;
    LAYER MET3 ;
    RECT 295.760 120.370 296.760 121.350 ;
    LAYER MET3 ;
    RECT 295.760 125.130 296.760 126.110 ;
    LAYER MET3 ;
    RECT 295.760 129.890 296.760 130.870 ;
    LAYER MET3 ;
    RECT 295.760 134.650 296.760 135.630 ;
    LAYER MET3 ;
    RECT 295.760 139.410 296.760 140.390 ;
    LAYER MET3 ;
    RECT 295.760 144.170 296.760 145.150 ;
    LAYER MET3 ;
    RECT 295.760 148.930 296.760 149.910 ;
    LAYER MET3 ;
    RECT 295.760 153.690 296.760 154.670 ;
    LAYER MET3 ;
    RECT 295.760 158.450 296.760 159.430 ;
    LAYER MET3 ;
    RECT 295.760 163.210 296.760 164.190 ;
    LAYER MET3 ;
    RECT 295.760 167.970 296.760 168.950 ;
    LAYER MET3 ;
    RECT 295.760 172.730 296.760 173.710 ;
    LAYER MET3 ;
    RECT 295.760 177.490 296.760 178.470 ;
    LAYER MET3 ;
    RECT 295.760 182.250 296.760 183.230 ;
    LAYER MET3 ;
    RECT 295.760 187.010 296.760 187.990 ;
    LAYER MET3 ;
    RECT 295.760 191.770 296.760 192.750 ;
    LAYER MET3 ;
    RECT 295.760 196.530 296.760 197.510 ;
    LAYER MET3 ;
    RECT 295.760 201.290 296.760 202.270 ;
    LAYER MET3 ;
    RECT 295.760 206.050 296.760 207.030 ;
    LAYER MET3 ;
    RECT 295.760 210.810 296.760 211.790 ;
    LAYER MET3 ;
    RECT 295.760 215.570 296.760 216.550 ;
    LAYER MET3 ;
    RECT 295.760 220.330 296.760 221.310 ;
    LAYER MET3 ;
    RECT 295.760 225.090 296.760 226.070 ;
    LAYER MET3 ;
    RECT 295.760 229.850 296.760 230.830 ;
    LAYER MET3 ;
    RECT 295.760 234.610 296.760 235.590 ;
    LAYER MET3 ;
    RECT 295.760 239.370 296.760 240.350 ;
    LAYER MET3 ;
    RECT 295.760 244.130 296.760 245.110 ;
    LAYER MET3 ;
    RECT 295.760 248.890 296.760 249.870 ;
    LAYER MET3 ;
    RECT 295.760 253.650 296.760 254.630 ;
    LAYER MET3 ;
    RECT 295.760 258.410 296.760 259.390 ;
    LAYER MET3 ;
    RECT 295.760 263.170 296.760 264.150 ;
    LAYER MET3 ;
    RECT 295.760 267.930 296.760 268.910 ;
    LAYER MET3 ;
    RECT 295.760 272.690 296.760 273.670 ;
    LAYER MET3 ;
    RECT 295.760 277.450 296.760 278.430 ;
    LAYER MET3 ;
    RECT 295.760 98.890 296.760 99.870 ;
    LAYER MET3 ;
    RECT 295.760 103.650 296.760 104.630 ;
    LAYER MET3 ;
    RECT 295.760 108.410 296.760 109.390 ;
    LAYER MET3 ;
    RECT 295.760 113.170 296.760 114.150 ;
    LAYER MET3 ;
    RECT 295.760 117.930 296.760 118.910 ;
    LAYER MET3 ;
    RECT 295.760 122.690 296.760 123.670 ;
    LAYER MET3 ;
    RECT 295.760 127.450 296.760 128.430 ;
    LAYER MET3 ;
    RECT 295.760 132.210 296.760 133.190 ;
    LAYER MET3 ;
    RECT 295.760 136.970 296.760 137.950 ;
    LAYER MET3 ;
    RECT 295.760 141.730 296.760 142.710 ;
    LAYER MET3 ;
    RECT 295.760 146.490 296.760 147.470 ;
    LAYER MET3 ;
    RECT 295.760 151.250 296.760 152.230 ;
    LAYER MET3 ;
    RECT 295.760 156.010 296.760 156.990 ;
    LAYER MET3 ;
    RECT 295.760 160.770 296.760 161.750 ;
    LAYER MET3 ;
    RECT 295.760 165.530 296.760 166.510 ;
    LAYER MET3 ;
    RECT 295.760 170.290 296.760 171.270 ;
    LAYER MET3 ;
    RECT 295.760 175.050 296.760 176.030 ;
    LAYER MET3 ;
    RECT 295.760 179.810 296.760 180.790 ;
    LAYER MET3 ;
    RECT 295.760 184.570 296.760 185.550 ;
    LAYER MET3 ;
    RECT 295.760 189.330 296.760 190.310 ;
    LAYER MET3 ;
    RECT 295.760 194.090 296.760 195.070 ;
    LAYER MET3 ;
    RECT 295.760 198.850 296.760 199.830 ;
    LAYER MET3 ;
    RECT 295.760 203.610 296.760 204.590 ;
    LAYER MET3 ;
    RECT 295.760 208.370 296.760 209.350 ;
    LAYER MET3 ;
    RECT 295.760 213.130 296.760 214.110 ;
    LAYER MET3 ;
    RECT 295.760 217.890 296.760 218.870 ;
    LAYER MET3 ;
    RECT 295.760 222.650 296.760 223.630 ;
    LAYER MET3 ;
    RECT 295.760 227.410 296.760 228.390 ;
    LAYER MET3 ;
    RECT 295.760 232.170 296.760 233.150 ;
    LAYER MET3 ;
    RECT 295.760 236.930 296.760 237.910 ;
    LAYER MET3 ;
    RECT 295.760 241.690 296.760 242.670 ;
    LAYER MET3 ;
    RECT 295.760 246.450 296.760 247.430 ;
    LAYER MET3 ;
    RECT 295.760 251.210 296.760 252.190 ;
    LAYER MET3 ;
    RECT 295.760 255.970 296.760 256.950 ;
    LAYER MET3 ;
    RECT 295.760 260.730 296.760 261.710 ;
    LAYER MET3 ;
    RECT 295.760 265.490 296.760 266.470 ;
    LAYER MET3 ;
    RECT 295.760 270.250 296.760 271.230 ;
    LAYER MET3 ;
    RECT 295.760 275.010 296.760 275.990 ;
    LAYER MET3 ;
    RECT 295.760 279.770 296.760 280.750 ;
    LAYER MET2 ;
    RECT 295.760 281.210 317.760 281.750 ;
    LAYER VIA2 ;
    RECT 307.900 281.350 317.520 281.610 ;
    LAYER MET3 ;
    RECT 295.760 282.210 296.760 283.190 ;
    LAYER MET2 ;
    RECT 295.760 285.970 317.760 286.510 ;
    LAYER VIA2 ;
    RECT 307.900 286.110 317.520 286.370 ;
    LAYER MET3 ;
    RECT 295.760 284.530 296.760 285.510 ;
    LAYER MET2 ;
    RECT 295.760 285.970 317.760 286.510 ;
    LAYER MET2 ;
    RECT 295.760 290.730 317.760 291.270 ;
    LAYER MET2 ;
    RECT 295.760 295.490 317.760 296.030 ;
    LAYER MET2 ;
    RECT 295.760 300.250 317.760 300.790 ;
    LAYER MET2 ;
    RECT 295.760 305.010 317.760 305.550 ;
    LAYER MET2 ;
    RECT 295.760 309.770 317.760 310.310 ;
    LAYER MET2 ;
    RECT 295.760 314.530 317.760 315.070 ;
    LAYER VIA2 ;
    RECT 307.900 286.110 317.520 286.370 ;
    LAYER VIA2 ;
    RECT 307.900 290.870 317.520 291.130 ;
    LAYER VIA2 ;
    RECT 307.900 295.630 317.520 295.890 ;
    LAYER VIA2 ;
    RECT 307.900 300.390 317.520 300.650 ;
    LAYER VIA2 ;
    RECT 307.900 305.150 317.520 305.410 ;
    LAYER VIA2 ;
    RECT 307.900 309.910 317.520 310.170 ;
    LAYER VIA2 ;
    RECT 307.900 314.670 317.520 314.930 ;
    LAYER MET2 ;
    RECT 295.760 290.730 317.760 291.270 ;
    LAYER MET2 ;
    RECT 295.760 295.490 317.760 296.030 ;
    LAYER MET2 ;
    RECT 295.760 300.250 317.760 300.790 ;
    LAYER MET2 ;
    RECT 295.760 305.010 317.760 305.550 ;
    LAYER MET2 ;
    RECT 295.760 309.770 317.760 310.310 ;
    LAYER MET2 ;
    RECT 295.760 314.530 317.760 315.070 ;
    LAYER MET2 ;
    RECT 295.760 319.290 317.760 319.830 ;
    LAYER VIA2 ;
    RECT 307.900 290.870 317.520 291.130 ;
    LAYER VIA2 ;
    RECT 307.900 295.630 317.520 295.890 ;
    LAYER VIA2 ;
    RECT 307.900 300.390 317.520 300.650 ;
    LAYER VIA2 ;
    RECT 307.900 305.150 317.520 305.410 ;
    LAYER VIA2 ;
    RECT 307.900 309.910 317.520 310.170 ;
    LAYER VIA2 ;
    RECT 307.900 314.670 317.520 314.930 ;
    LAYER VIA2 ;
    RECT 307.900 319.430 317.520 319.690 ;
    LAYER MET3 ;
    RECT 295.760 286.970 296.760 287.950 ;
    LAYER MET3 ;
    RECT 295.760 291.730 296.760 292.710 ;
    LAYER MET3 ;
    RECT 295.760 296.490 296.760 297.470 ;
    LAYER MET3 ;
    RECT 295.760 301.250 296.760 302.230 ;
    LAYER MET3 ;
    RECT 295.760 306.010 296.760 306.990 ;
    LAYER MET3 ;
    RECT 295.760 310.770 296.760 311.750 ;
    LAYER MET3 ;
    RECT 295.760 315.530 296.760 316.510 ;
    LAYER MET3 ;
    RECT 295.760 289.290 296.760 290.270 ;
    LAYER MET3 ;
    RECT 295.760 294.050 296.760 295.030 ;
    LAYER MET3 ;
    RECT 295.760 298.810 296.760 299.790 ;
    LAYER MET3 ;
    RECT 295.760 303.570 296.760 304.550 ;
    LAYER MET3 ;
    RECT 295.760 308.330 296.760 309.310 ;
    LAYER MET3 ;
    RECT 295.760 313.090 296.760 314.070 ;
    LAYER MET3 ;
    RECT 295.760 317.850 296.760 318.830 ;
    LAYER MET2 ;
    RECT 295.760 319.290 317.760 319.830 ;
    LAYER VIA2 ;
    RECT 307.900 319.430 317.520 319.690 ;
    LAYER MET2 ;
    RECT 295.760 324.050 317.760 324.590 ;
    LAYER VIA2 ;
    RECT 307.900 324.190 317.520 324.450 ;
    LAYER MET3 ;
    RECT 295.760 320.290 296.760 321.270 ;
    LAYER MET3 ;
    RECT 295.760 322.610 296.760 323.590 ;
    LAYER MET3 ;
    RECT 177.825 326.410 179.075 348.410 ;
    LAYER VIA2 ;
    RECT 178.060 338.600 178.840 348.220 ;
    LAYER MET2 ;
    RECT 179.535 326.410 180.785 327.410 ;
    LAYER MET3 ;
    RECT 193.970 326.410 194.800 348.410 ;
    LAYER MET3 ;
    RECT 250.890 326.410 251.720 348.410 ;
    LAYER VIA2 ;
    RECT 194.255 338.600 194.515 348.220 ;
    LAYER VIA2 ;
    RECT 251.175 338.600 251.435 348.220 ;
    LAYER MET2 ;
    RECT 222.430 326.410 223.260 327.410 ;
    LAYER MET2 ;
    RECT 279.350 326.410 280.180 327.410 ;
    LAYER MET2 ;
    RECT 295.760 324.050 317.760 324.590 ;
    LAYER VIA2 ;
    RECT 307.900 324.190 317.520 324.450 ;
    LAYER VIA2 ;
    RECT 0.190 0.190 9.810 9.810 ;
    LAYER VIA2 ;
    RECT 11.190 11.190 20.810 20.810 ;
    LAYER VIA2 ;
    RECT 307.950 0.190 317.570 9.810 ;
    LAYER VIA2 ;
    RECT 296.950 11.190 306.570 20.810 ;
    LAYER VIA2 ;
    RECT 296.950 327.600 306.570 337.220 ;
    LAYER VIA2 ;
    RECT 307.950 338.600 317.570 348.220 ;
    LAYER VIA2 ;
    RECT 11.190 327.600 20.810 337.220 ;
    LAYER VIA2 ;
    RECT 0.190 338.600 9.810 348.220 ;
    END 
  END MSL18B_1536X8_RW10TM4_16_20221107
END LIBRARY
