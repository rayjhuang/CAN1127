
module chiptop_1127a0 ( CSP, CSN, VFB, COM, SW, BST, VDRV, LG, HG, GATE, DP, 
        DN, CC1, CC2, TST, GPIO_TS, SCL, SDA, GPIO1, GPIO2, GPIO3, GPIO4, 
        GPIO5 );
  input TST;
  output LG, HG, GATE;
  inout CSP,  CSN,  VFB,  COM,  SW,  BST,  VDRV,  DP,  DN,  CC1,  CC2, 
     GPIO_TS,  SCL,  SDA,  GPIO1,  GPIO2,  GPIO3,  GPIO4,  GPIO5;
  wire   SRAM_WEB, SRAM_CEB, SRAM_OEB, PWREN_HOLD, RD_ENB, STB_RP, DRP_OSC,
         IMP_OSC, TX_EN, TX_DAT, RX_DAT, RX_SQL, DAC1_EN, AD_RST, AD_HOLD,
         COMP_O, CCI2C_EN, RSTB, SLEEP, OSC_LOW, OSC_STOP, PWRDN, VPP_0V,
         VPP_SEL, LDO3P9V, OSC_O, RD_DET, OCP_SEL, CC1_DOB, CC2_DOB, CC1_DI,
         CC2_DI, DP_COMP, DN_COMP, DN_FAULT, LFOSC_ENB, VPP_OTP, IO_RSTB5,
         V1P1, ANAP_TS, TS_ANA_R, ANAP_GP1, GP1_ANA_R, ANAP_GP2, GP2_ANA_R,
         ANAP_GP3, GP3_ANA_R, ANAP_GP4, GP4_ANA_R, ANAP_GP5, GP5_ANA_R, DI_TST,
         DI_TS, SRAM_CLK, PMEM_RE, PMEM_PGM, PMEM_CSB, do_ccctl_0_,
         do_srcctl_0, tm_atpg, n1, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, net1, net2, net3, net4;
  wire   [10:0] SRAM_A;
  wire   [7:0] SRAM_D;
  wire   [7:0] xdat_o;
  wire   [7:0] ANAOPT;
  wire   [1:0] FSW;
  wire   [1:0] RP_EN;
  wire   [1:0] VCONN_EN;
  wire   [17:0] SAMPL_SEL;
  wire   [7:0] DUMMY_IN;
  wire   [55:0] REGTRM;
  wire   [7:0] PWR_I;
  wire   [1:0] OVP_SEL;
  wire   [5:0] DAC3_V;
  wire   [10:0] DAC0;
  wire   [3:0] ANA_TM;
  wire   [9:0] DAC1;
  wire   [1:0] RP_SEL;
  wire   [1:0] IE_GPIO;
  wire   [6:0] DI_GPIO;
  wire   [6:0] OE_GPIO;
  wire   [6:0] DO_GPIO;
  wire   [6:0] PU_GPIO;
  wire   [6:0] PD_GPIO;
  wire   [3:0] DO_TS;
  wire   [1:0] PMEM_CLK;
  wire   [7:0] PMEM_Q1;
  wire   [7:0] PMEM_Q0;
  wire   [1:0] PMEM_SAP;
  wire   [1:0] PMEM_TWLB;
  wire   [15:0] PMEM_A;
  wire   [7:0] bck_regx0;
  wire   [7:2] bck_regx1;
  wire   [7:2] do_xana1;
  wire   [7:0] do_xana0;
  wire   [3:0] do_regx_xtm;
  wire   [5:2] do_cvctl;
  wire   [3:0] do_vooc;
  wire   [5:0] do_dpdm;
  wire   [5:4] do_srcctl;
  wire   [7:0] do_cctrx;
  wire   [3:0] di_xanav;
  wire   [5:0] srci;
  tri   CSP;
  tri   CSN;
  tri   VFB;
  tri   COM;
  tri   SW;
  tri   BST;
  tri   VDRV;
  tri   DP;
  tri   DN;
  tri   CC1;
  tri   CC2;
  tri   TST;
  tri   GPIO_TS;
  tri   SCL;
  tri   SDA;
  tri   GPIO1;
  tri   GPIO2;
  tri   GPIO3;
  tri   GPIO4;
  tri   GPIO5;

  anatop_1127a0 U0_ANALOG_TOP ( .CC1(CC1), .CC2(CC2), .DP(DP), .DN(DN), .VFB(
        VFB), .CSP(CSP), .CSN(CSN), .COM(COM), .SW(SW), .BST(BST), .VDRV(VDRV), 
        .LG(LG), .HG(HG), .GATE(GATE), .BST_SET(bck_regx0[0]), .DCM_SEL(
        bck_regx0[1]), .HGOFF(bck_regx0[2]), .HGON(bck_regx0[4]), .LGOFF(
        bck_regx0[3]), .LGON(bck_regx0[5]), .EN_DRV(bck_regx0[6]), .FSW(FSW), 
        .EN_OSC(bck_regx1[2]), .MAXDS(bck_regx1[3]), .EN_GM(bck_regx1[4]), 
        .EN_ODLDO(bck_regx1[5]), .EN_IBUK(bck_regx1[6]), .CP_EN(do_srcctl_0), 
        .EXT_CP(bck_regx1[7]), .INT_CP(bck_regx0[7]), .ANTI_INRUSH(do_cvctl[5]), .PWREN_HOLD(PWREN_HOLD), .RP_SEL(RP_SEL), .RP1_EN(RP_EN[0]), .RP2_EN(
        RP_EN[1]), .VCONN1_EN(VCONN_EN[0]), .VCONN2_EN(VCONN_EN[1]), .SGP({
        do_cctrx[0], do_regx_xtm}), .S20U(do_cctrx[1]), .S100U(do_cctrx[2]), 
        .TX_EN(TX_EN), .TX_DAT(TX_DAT), .CC_SEL(do_ccctl_0_), .TRA(do_cctrx[4]), .TFA(do_cctrx[5]), .LSR(do_cctrx[6]), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), 
        .SEL_RX_TH(do_cctrx[7]), .DAC1_EN(DAC1_EN), .DPDN_SHORT(do_dpdm[0]), 
        .DP_2V7_EN(do_dpdm[4]), .DN_2V7_EN(do_dpdm[3]), .DP_0P6V_EN(
        do_xana1[3]), .DN_0P6V_EN(do_xana1[2]), .DP_DWN_EN(do_dpdm[2]), 
        .DN_DWN_EN(do_dpdm[1]), .PWR_I(PWR_I), .DAC3(DAC3_V), .DAC1(DAC1), 
        .CV2(do_xana0[0]), .LFOSC_ENB(LFOSC_ENB), .VO_DISCHG(do_srcctl[4]), 
        .DISCHG_SEL(do_srcctl[5]), .CMP_SEL_VO10(SAMPL_SEL[1]), .CMP_SEL_VO20(
        SAMPL_SEL[10]), .CMP_SEL_GP1(SAMPL_SEL[17]), .CMP_SEL_GP2(
        SAMPL_SEL[16]), .CMP_SEL_GP3(SAMPL_SEL[15]), .CMP_SEL_GP4(
        SAMPL_SEL[14]), .CMP_SEL_GP5(SAMPL_SEL[13]), .CMP_SEL_VIN20(
        SAMPL_SEL[0]), .CMP_SEL_TS(SAMPL_SEL[3]), .CMP_SEL_IS(SAMPL_SEL[2]), 
        .CMP_SEL_CC2(SAMPL_SEL[7]), .CMP_SEL_CC1(SAMPL_SEL[6]), 
        .CMP_SEL_CC2_4(SAMPL_SEL[12]), .CMP_SEL_CC1_4(SAMPL_SEL[11]), 
        .CMP_SEL_DP(SAMPL_SEL[4]), .CMP_SEL_DP_3(SAMPL_SEL[8]), .CMP_SEL_DN(
        SAMPL_SEL[5]), .CMP_SEL_DN_3(SAMPL_SEL[9]), .OCP_EN(do_cvctl[2]), 
        .CS_EN(do_cctrx[3]), .COMP_O(COMP_O), .CCI2C_EN(CCI2C_EN), .UVP_SEL(
        do_xana0[7]), .TM(ANA_TM), .V5OCP(srci[4]), .RSTB(RSTB), .DAC0(DAC0), 
        .SLEEP(SLEEP), .OSC_LOW(OSC_LOW), .OSC_STOP(OSC_STOP), .PWRDN(PWRDN), 
        .VPP_ZERO(VPP_0V), .OSC_O(OSC_O), .RD_DET(RD_DET), .IMP_OSC(IMP_OSC), 
        .DRP_OSC(DRP_OSC), .STB_RP(STB_RP), .RD_ENB(RD_ENB), .OCP(srci[1]), 
        .SCP(srci[3]), .UVP(srci[0]), .LDO3P9V(LDO3P9V), .VPP_SEL(VPP_SEL), 
        .CC1_DOB(CC1_DOB), .CC2_DOB(CC2_DOB), .CC1_DI(CC1_DI), .CC2_DI(CC2_DI), 
        .OTPI(srci[5]), .OVP_SEL(OVP_SEL), .OVP(srci[2]), .DN_COMP(DN_COMP), 
        .DP_COMP(DP_COMP), .DPDN_VTH(do_xana0[5]), .DPDEN(do_vooc[3]), .DPDO(
        do_vooc[2]), .DPIE(do_dpdm[5]), .DNDEN(do_vooc[1]), .DNDO(do_vooc[0]), 
        .DNIE(do_dpdm[5]), .DUMMY_IN(DUMMY_IN), .CP_CLKX2(ANAOPT[7]), 
        .SEL_CONST_OVP(ANAOPT[6]), .LP_EN(ANAOPT[5]), .DNCHK_EN(ANAOPT[3]), 
        .IRP_EN(ANAOPT[2]), .CCBFEN(ANAOPT[0]), .REGTRM(REGTRM), .AD_RST(
        AD_RST), .AD_HOLD(AD_HOLD), .DN_FAULT(DN_FAULT), .SEL_CCGAIN(
        do_xana0[3]), .VFB_SW(do_xana0[1]), .CPVSEL(do_xana1[6]), .CLAMPV_EN(
        do_xana1[5]), .HVNG_CPEN(do_xana1[7]), .OCP_SEL(OCP_SEL), .OCP_80M(
        di_xanav[1]), .OCP_160M(di_xanav[0]), .OPTO1(di_xanav[2]), .OPTO2(
        di_xanav[3]), .VPP_OTP(VPP_OTP), .RSTB_5(IO_RSTB5), .V1P1(V1P1), 
        .TS_ANA_R(TS_ANA_R), .GP5_ANA_R(GP5_ANA_R), .GP4_ANA_R(GP4_ANA_R), 
        .GP3_ANA_R(GP3_ANA_R), .GP2_ANA_R(GP2_ANA_R), .GP1_ANA_R(GP1_ANA_R), 
        .TS_ANA_P(ANAP_TS), .GP5_ANA_P(ANAP_GP5), .GP4_ANA_P(ANAP_GP4), 
        .GP3_ANA_P(ANAP_GP3), .GP2_ANA_P(ANAP_GP2), .GP1_ANA_P(ANAP_GP1) );
  IODMURUDA_A0 PAD_SCL ( .PAD(SCL), .IE(IE_GPIO[1]), .DI(DI_GPIO[0]), .OE(
        OE_GPIO[0]), .DO(DO_GPIO[0]), .PU(PU_GPIO[0]), .PD(PD_GPIO[0]), 
        .ANA_R(), .RSTB_5(IO_RSTB5), .VB(V1P1) );
  IODMURUDA_A0 PAD_SDA ( .PAD(SDA), .IE(IE_GPIO[1]), .DI(DI_GPIO[1]), .OE(
        OE_GPIO[1]), .DO(DO_GPIO[1]), .PU(PU_GPIO[1]), .PD(PD_GPIO[1]), 
        .ANA_R(), .RSTB_5(IO_RSTB5), .VB(V1P1) );
  IOBMURUDA_A0 PAD_TST ( .PAD(TST), .IE(1'b1), .DI(DI_TST), .OE(1'b0), .DO(
        1'b0), .PU(1'b0), .PD(1'b1), .ANA_R(), .RSTB_5(IO_RSTB5), .VB(V1P1) );
  IOBMURUDA_A1 PAD_GPIO1 ( .PAD(GPIO1), .IE(IE_GPIO[0]), .DI(DI_GPIO[2]), .OE(
        OE_GPIO[2]), .DO(DO_GPIO[2]), .PU(PU_GPIO[2]), .PD(PD_GPIO[2]), 
        .ANA_R(GP1_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP1) );
  IOBMURUDA_A1 PAD_GPIO2 ( .PAD(GPIO2), .IE(IE_GPIO[0]), .DI(DI_GPIO[3]), .OE(
        OE_GPIO[3]), .DO(DO_GPIO[3]), .PU(PU_GPIO[3]), .PD(PD_GPIO[3]), 
        .ANA_R(GP2_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP2) );
  IOBMURUDA_A1 PAD_GPIO3 ( .PAD(GPIO3), .IE(IE_GPIO[0]), .DI(DI_GPIO[4]), .OE(
        OE_GPIO[4]), .DO(DO_GPIO[4]), .PU(PU_GPIO[4]), .PD(PD_GPIO[4]), 
        .ANA_R(GP3_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP3) );
  IOBMURUDA_A1 PAD_GPIO4 ( .PAD(GPIO4), .IE(IE_GPIO[0]), .DI(DI_GPIO[5]), .OE(
        OE_GPIO[5]), .DO(DO_GPIO[5]), .PU(PU_GPIO[5]), .PD(PD_GPIO[5]), 
        .ANA_R(GP4_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP4) );
  IOBMURUDA_A1 PAD_GPIO5 ( .PAD(GPIO5), .IE(IE_GPIO[0]), .DI(DI_GPIO[6]), .OE(
        OE_GPIO[6]), .DO(DO_GPIO[6]), .PU(PU_GPIO[6]), .PD(PD_GPIO[6]), 
        .ANA_R(GP5_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP5) );
  IOBMURUDA_A1 PAD_GPIO_TS ( .PAD(GPIO_TS), .IE(IE_GPIO[0]), .DI(DI_TS), .OE(
        DO_TS[2]), .DO(DO_TS[3]), .PU(DO_TS[1]), .PD(DO_TS[0]), .ANA_R(
        TS_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_TS) );
  MSL18B_1536X8_RW10TM4_16_20221107 U0_SRAM ( .DO(xdat_o), .CK(SRAM_CLK), 
        .CSB(SRAM_CEB), .OEB(SRAM_OEB), .WEB(SRAM_WEB), .A(SRAM_A), .DI(SRAM_D) );
  ATO0008KX8MX180LBX4DA U0_CODE_0_ ( .A(PMEM_A), .CSB(PMEM_CSB), .CLK(
        PMEM_CLK[0]), .PGM(n1), .RE(PMEM_RE), .TWLB(PMEM_TWLB), .VSS(), 
        .VDD(), .VDDP(VPP_OTP), .SAP(PMEM_SAP), .Q(PMEM_Q0) );
  ATO0008KX8MX180LBX4DA U0_CODE_1_ ( .A(PMEM_A), .CSB(PMEM_CSB), .CLK(
        PMEM_CLK[1]), .PGM(PMEM_PGM), .RE(PMEM_RE), .TWLB(PMEM_TWLB), .VSS(
        ), .VDD(), .VDDP(VPP_OTP), .SAP(PMEM_SAP), .Q(PMEM_Q1) );
  core_a0 U0_CORE ( .SRCI(srci), .XANAV({1'b0, di_xanav}), .BCK_REGX({
        bck_regx1, FSW, bck_regx0}), .ANA_REGX({do_xana1[7:5], 
        SYNOPSYS_UNCONNECTED_1, do_xana1[3:2], SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, do_xana0[7], SYNOPSYS_UNCONNECTED_4, 
        do_xana0[5], SYNOPSYS_UNCONNECTED_5, do_xana0[3], 
        SYNOPSYS_UNCONNECTED_6, do_xana0[1:0]}), .LFOSC_ENB(LFOSC_ENB), 
        .STB_RP(STB_RP), .RD_ENB(RD_ENB), .OCP_SEL(OCP_SEL), .PWREN_HOLD(
        PWREN_HOLD), .CC1_DI(CC1_DI), .CC2_DI(CC2_DI), .DRP_OSC(DRP_OSC), 
        .IMP_OSC(IMP_OSC), .CC1_DOB(CC1_DOB), .CC2_DOB(CC2_DOB), .DAC1_EN(
        DAC1_EN), .SH_RST(AD_RST), .SH_HOLD(AD_HOLD), .LDO3P9V(LDO3P9V), .XTM(
        do_regx_xtm), .DO_CVCTL({OVP_SEL, do_cvctl[5], SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, do_cvctl[2], SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10}), .DO_CCTRX(do_cctrx), .DO_SRCCTL({
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, do_srcctl, VCONN_EN, 
        SYNOPSYS_UNCONNECTED_13, do_srcctl_0}), .DO_CCCTL({RP_EN, RP_SEL, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, do_ccctl_0_}), .DO_DAC0(DAC0), .DO_DPDN(
        do_dpdm), .DO_VOOC(do_vooc), .DO_PWR_I(PWR_I), .PMEM_A(PMEM_A), 
        .PMEM_Q0(PMEM_Q0), .PMEM_Q1(PMEM_Q1), .PMEM_TWLB(PMEM_TWLB), 
        .PMEM_SAP(PMEM_SAP), .PMEM_CLK(PMEM_CLK), .PMEM_CSB(PMEM_CSB), 
        .PMEM_RE(PMEM_RE), .PMEM_PGM(PMEM_PGM), .VPP_SEL(VPP_SEL), .VPP_0V(
        VPP_0V), .SRAM_WEB(SRAM_WEB), .SRAM_CEB(SRAM_CEB), .SRAM_OEB(SRAM_OEB), 
        .SRAM_CLK(SRAM_CLK), .SRAM_A(SRAM_A), .SRAM_D(SRAM_D), .SRAM_RDAT(
        xdat_o), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .RD_DET(RD_DET), .TX_DAT(
        TX_DAT), .TX_EN(TX_EN), .OSC_STOP(OSC_STOP), .OSC_LOW(OSC_LOW), 
        .SLEEP(SLEEP), .PWRDN(PWRDN), .OCDRV_ENZ(), .DAC1_V(DAC1), .SAMPL_SEL(
        SAMPL_SEL), .DAC1_COMP(COMP_O), .CCI2C_EN(CCI2C_EN), .ANA_TM(ANA_TM), 
        .DM_FAULT(DN_FAULT), .DM_COMP(DN_COMP), .DP_COMP(DP_COMP), .DI_GPIO(
        DI_GPIO), .DO_GPIO(DO_GPIO), .OE_GPIO(OE_GPIO), .GPIO_PU(PU_GPIO), 
        .GPIO_PD(PD_GPIO), .GPIO_IE(IE_GPIO), .DO_TS(DO_TS), .DI_TS(DI_TS), 
        .REGTRM(REGTRM), .ANAOPT({ANAOPT[7:5], SYNOPSYS_UNCONNECTED_17, 
        ANAOPT[3:2], SYNOPSYS_UNCONNECTED_18, ANAOPT[0]}), .DUMMY_IN(DUMMY_IN), 
        .DAC3_V(DAC3_V), .i_clk(OSC_O), .i_rstz(RSTB), .atpg_en(tm_atpg), 
        .di_tst(DI_TST), .tm_atpg(tm_atpg) );
  BUFX12 U3 ( .A(PMEM_PGM), .Y(n1) );
endmodule


module core_a0 ( SRCI, XANAV, BCK_REGX, ANA_REGX, LFOSC_ENB, STB_RP, RD_ENB, 
        OCP_SEL, PWREN_HOLD, CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, CC1_DOB, 
        CC2_DOB, DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, XTM, DO_CVCTL, DO_CCTRX, 
        DO_SRCCTL, DO_CCCTL, DO_DAC0, DO_DPDN, DO_VOOC, DO_PWR_I, PMEM_A, 
        PMEM_Q0, PMEM_Q1, PMEM_TWLB, PMEM_SAP, PMEM_CLK, PMEM_CSB, PMEM_RE, 
        PMEM_PGM, VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, 
        SRAM_A, SRAM_D, SRAM_RDAT, RX_DAT, RX_SQL, RD_DET, TX_DAT, TX_EN, 
        OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, DAC1_V, SAMPL_SEL, 
        DAC1_COMP, CCI2C_EN, ANA_TM, DM_FAULT, DM_COMP, DP_COMP, DI_GPIO, 
        DO_GPIO, OE_GPIO, GPIO_PU, GPIO_PD, GPIO_IE, DO_TS, DI_TS, REGTRM, 
        ANAOPT, DUMMY_IN, DAC3_V, i_clk, i_rstz, atpg_en, di_tst, tm_atpg );
  input [5:0] SRCI;
  input [4:0] XANAV;
  output [15:0] BCK_REGX;
  output [15:0] ANA_REGX;
  output [3:0] XTM;
  output [7:0] DO_CVCTL;
  output [7:0] DO_CCTRX;
  output [7:0] DO_SRCCTL;
  output [7:0] DO_CCCTL;
  output [10:0] DO_DAC0;
  output [5:0] DO_DPDN;
  output [3:0] DO_VOOC;
  output [7:0] DO_PWR_I;
  output [15:0] PMEM_A;
  input [7:0] PMEM_Q0;
  input [7:0] PMEM_Q1;
  output [1:0] PMEM_TWLB;
  output [1:0] PMEM_SAP;
  output [1:0] PMEM_CLK;
  output [10:0] SRAM_A;
  output [7:0] SRAM_D;
  input [7:0] SRAM_RDAT;
  output [9:0] DAC1_V;
  output [17:0] SAMPL_SEL;
  output [3:0] ANA_TM;
  input [6:0] DI_GPIO;
  output [6:0] DO_GPIO;
  output [6:0] OE_GPIO;
  output [6:0] GPIO_PU;
  output [6:0] GPIO_PD;
  output [1:0] GPIO_IE;
  output [3:0] DO_TS;
  output [55:0] REGTRM;
  output [7:0] ANAOPT;
  output [7:0] DUMMY_IN;
  output [5:0] DAC3_V;
  input CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, RX_DAT, RX_SQL, RD_DET, DAC1_COMP,
         DM_FAULT, DM_COMP, DP_COMP, DI_TS, i_clk, i_rstz, atpg_en, di_tst;
  output LFOSC_ENB, STB_RP, RD_ENB, OCP_SEL, PWREN_HOLD, CC1_DOB, CC2_DOB,
         DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, PMEM_CSB, PMEM_RE, PMEM_PGM,
         VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, TX_DAT,
         TX_EN, OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, CCI2C_EN, tm_atpg;
  wire   N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N268, n653, n654, aswclk, detclk, tclk_sel, s_clk, aswkup, x_clk,
         t_di_gpio4, t_pmem_clk, pmem_csb, t_pmem_csb, r_osc_gate, t_osc_gate,
         g_clk, xram_ce, iram_ce, sram_en, r_i2c_attr, esfrm_oe, esfrm_we,
         sfrack, ictlr_psrack, esfrm_rrdy, memwr, memrd, memrd_c, memack,
         o_cpurst, hit_xd, hit_xr, hit_ps, hit_ps_c, mcu_ram_r, mcu_ram_w,
         regx_re, iram_we, xram_we, regx_we, bist_en, bist_wr, srstz,
         prl_cany0w, prl_cany0r, mempsrd, r_bclk_sel, r_hold_mcu, t0_intr,
         fcp_intr, dpdm_urx, s0_rxdoe, mcuo_scl, mcuo_sda, mempsack, mempswr,
         mempsrd_c, sfr_w, sfr_r, ictlr_psack, ictlr_inc, set_hold, bkpt_hold,
         bkpt_ena, r_psrd, r_pswr, prl_cany0, prl_c0set, pmem_pgm, pmem_re,
         we_twlb, r_otp_wpls, pwrdn_rst, r_otp_pwdn_en, ramacc, frc_lg_on,
         frc_hg_off, cc1_di, cc2_di, r_sleep, ps_pwrdn, r_pwrdn, r_ocdrv_enz,
         r_osc_stop, r_pwrv_upd, r_otpi_gate, r_fcpre, r_fortxdat, r_fortxrdy,
         r_fortxen, r_gpio_tm, pid_goidle, pid_gobusy, bus_idle, sse_idle,
         r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, r_unlock, r_first, r_last,
         r_fiforst, r_set_cpmsgid, r_txendk, r_txshrt, r_auto_discard,
         r_dat_portrole, r_dat_datarole, r_pshords, r_discard, r_strtch,
         r_i2c_ninc, r_i2c_fwnak, r_i2c_fwack, hwi2c_stretch, i2c_ev_6_,
         i2c_ev_3, i2c_ev_2, prl_discard, prl_GCTxDone, pff_obsd, pff_empty,
         pff_full, ptx_ack, clk_1p0m, clk_500, prstz, sse_rdrdy, upd_rdrdy,
         sse_prefetch, slvo_sda, slvo_re, slvo_early, dm_comp, dp_comp,
         di_sqlch, ptx_cc, ptx_oe, sh_rst, sh_hold, fcp_oe, fcp_do,
         sdischg_duty, clk_100k, r_imp_osc, clk_500k, r_vpp_en, r_vpp0v_en,
         di_ts, di_aswk_0, r_xana_23, r_xana_19, r_xana_18, divff_o1, clk_50k,
         N448, o_dodat0_15_, o_dodat5_2_, N568, N569, N570, N571, N572, N575,
         N576, N577, N578, N579, N580, N581, N582, N583, N584, N1477, N1482,
         net8852, n123, n126, n128, n507, n508, n509, n510, n348, n345, n344,
         n347, n346, n27, n56, n57, n58, n500, n502, n503, n511, n514, n515,
         n516, n517, n6, n11, n19, n20, n534, n644, n646, n647, n648, n649,
         n650, n651, n652, n686, n687, n688, n724, n774, n775, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n868, n869, n870, n871, n872, n873, n874, n884, n889, n895,
         n916, n922, n942, n949, n957, n958, n959, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n981,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1099, n1108, n1109, n1110, n1117, n1120,
         n1130, n1131, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1145, n1, n2, n3, n4, n5, n7, n8, n10, n12, n13, n14, n15,
         n16, n17, n18, n22, n24, n25, n26, n30, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n124, n125, n127, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106;
  wire   [9:0] aswclk_ps;
  wire   [9:0] detclk_ps;
  wire   [1:0] pmem_clk;
  wire   [7:0] sse_wdat;
  wire   [7:0] prx_fifowdat;
  wire   [7:0] sse_adr;
  wire   [7:0] prl_cany0adr;
  wire   [7:0] esfrm_wdat;
  wire   [6:0] esfrm_adr;
  wire   [7:0] mcu_esfrrdat;
  wire   [7:0] delay_inst;
  wire   [7:0] esfrm_rdat;
  wire   [3:0] r_pg0_sel;
  wire   [15:0] memaddr;
  wire   [15:0] memaddr_c;
  wire   [7:0] memdatao;
  wire   [7:0] idat_adr;
  wire   [7:0] idat_wdat;
  wire   [10:0] iram_a;
  wire   [10:0] xram_a;
  wire   [7:0] iram_d;
  wire   [7:0] xram_d;
  wire   [1:0] sram_rdat;
  wire   [7:0] regx_rdat;
  wire   [10:0] bist_adr;
  wire   [7:0] bist_wdat;
  wire   [7:0] memdatai;
  wire   [7:0] ictlr_inst;
  wire   [15:0] mcu_pc;
  wire   [22:16] mcu_dbgpo;
  wire   [3:2] sfr_intr;
  wire   [7:0] exint;
  wire   [7:0] ff_p0;
  wire   [6:0] do_p0;
  wire   [7:0] sfr_rdat;
  wire   [7:0] sfr_wdat;
  wire   [6:0] sfr_adr;
  wire   [14:0] bkpt_pc;
  wire   [14:0] r_inst_ofs;
  wire   [7:0] pmem_q0;
  wire   [7:0] pmem_q1;
  wire   [1:0] pmem_twlb;
  wire   [1:0] wd_twlb;
  wire   [1:0] r_sqlch;
  wire   [3:2] r_ccrx;
  wire   [1:0] r_rxdb_opt;
  wire   [7:4] r_pwrctl;
  wire   [5:2] di_pro;
  wire   [1:0] lg_pulse_len;
  wire   [7:0] r_srcctl;
  wire   [7:0] r_dpdmctl;
  wire   [11:0] r_fw_pwrv;
  wire   [5:0] r_cvcwr;
  wire   [15:0] r_cvofs;
  wire   [7:0] r_cctrx;
  wire   [7:0] r_ccctl;
  wire   [6:0] r_fcpwr;
  wire   [7:0] fcp_r_dat;
  wire   [7:0] fcp_r_sta;
  wire   [7:0] fcp_r_msk;
  wire   [7:0] fcp_r_ctl;
  wire   [7:0] fcp_r_crc;
  wire   [7:0] fcp_r_acc;
  wire   [7:0] fcp_r_tui;
  wire   [7:0] r_accctl;
  wire   [7:5] r_comp_opt;
  wire   [14:0] sfr_dacwr;
  wire   [17:0] r_dac_en;
  wire   [17:0] r_sar_en;
  wire   [7:0] r_isofs;
  wire   [7:0] r_adofs;
  wire   [7:0] dac_r_ctl;
  wire   [7:0] dac_r_cmpsta;
  wire   [17:0] dac_r_comp;
  wire   [143:0] dac_r_vs;
  wire   [5:0] x_daclsb;
  wire   [6:0] REVID;
  wire   [6:0] r_pu_gpio;
  wire   [6:0] r_pd_gpio;
  wire   [6:0] r_gpio_oe;
  wire   [1:0] r_gpio_ie;
  wire   [55:0] r_regtrm;
  wire   [3:0] r_ana_tm;
  wire   [7:0] i2c_ltbuf;
  wire   [7:0] i2c_lt_ofs;
  wire   [4:0] r_txnumk;
  wire   [1:0] r_auto_gdcrc;
  wire   [1:0] r_spec;
  wire   [1:0] r_dat_spec;
  wire   [6:0] r_txauto;
  wire   [6:0] r_rxords_ena;
  wire   [7:1] r_i2c_deva;
  wire   [2:0] prl_cpmsgid;
  wire   [1:0] pff_ack;
  wire   [7:0] pff_rdat;
  wire   [15:0] pff_rxpart;
  wire   [5:0] pff_ptr;
  wire   [6:0] prx_setsta;
  wire   [1:0] prx_rst;
  wire   [4:0] prx_rcvinf;
  wire   [5:0] prx_adpn;
  wire   [3:0] prx_fsm;
  wire   [2:0] ptx_fsm;
  wire   [3:0] prl_fsm;
  wire   [3:0] slvo_ev;
  wire   [1:0] r_i2cslv_route;
  wire   [5:4] r_i2crout;
  wire   [1:0] r_i2cmcu_route;
  wire   [18:17] upd_dbgpo;
  wire   [7:0] r_dacwdat;
  wire   [17:8] wr_dacv;
  wire   [10:7] r_dacwr;
  wire   [17:0] dacmux_sel;
  wire   [3:0] comp_smpl;
  wire   [7:0] r_cvcwdat;
  wire   [7:0] r_sdischg;
  wire   [7:0] r_vcomp;
  wire   [7:0] r_idacsh;
  wire   [7:0] r_cvofsx;
  wire   [7:0] r_xtm;
  wire   [6:0] bist_r_ctl;
  wire   [1:0] regx_hitbst;
  wire   [7:0] bist_r_dat;
  wire   [1:0] regx_wrpwm;
  wire   [15:0] r_pwm;
  wire   [1:0] r_sap;
  wire   [3:0] lt_gpi;
  wire   [6:0] r_do_ts;
  wire   [3:0] r_dpdo_sel;
  wire   [3:0] r_dndo_sel;
  wire   [4:2] di_aswk;
  wire   [7:0] r_bck0;
  wire   [7:0] r_bck1;
  wire   [15:0] r_xana;
  wire   [4:0] di_xanav;
  wire   [7:0] r_aopt;
  wire   [6:0] di_gpio;
  wire   [7:6] do_opt;
  wire   [1:0] pwm_o;
  wire   [15:0] d_dodat;
  wire   [3:0] r_lt_gpi;

  CKBUFX1 U0_ASWCLK_BUF_0_ ( .A(aswclk_ps[0]), .Y(aswclk_ps[1]) );
  CKBUFX1 U0_ASWCLK_BUF_1_ ( .A(aswclk_ps[1]), .Y(aswclk_ps[2]) );
  CKBUFX1 U0_ASWCLK_BUF_2_ ( .A(aswclk_ps[2]), .Y(aswclk_ps[3]) );
  CKBUFX1 U0_ASWCLK_BUF_3_ ( .A(aswclk_ps[3]), .Y(aswclk_ps[4]) );
  CKBUFX1 U0_ASWCLK_BUF_4_ ( .A(aswclk_ps[4]), .Y(aswclk_ps[5]) );
  CKBUFX1 U0_ASWCLK_BUF_5_ ( .A(aswclk_ps[5]), .Y(aswclk_ps[6]) );
  CKBUFX1 U0_ASWCLK_BUF_6_ ( .A(aswclk_ps[6]), .Y(aswclk_ps[7]) );
  CKBUFX1 U0_ASWCLK_BUF_7_ ( .A(aswclk_ps[7]), .Y(aswclk_ps[8]) );
  CKBUFX1 U0_ASWCLK_BUF_8_ ( .A(aswclk_ps[8]), .Y(aswclk_ps[9]) );
  CKBUFX1 U0_ASWCLK_BUF_9_ ( .A(aswclk_ps[9]), .Y(aswclk) );
  CKBUFX1 U0_DETCLK_BUF_0_ ( .A(detclk_ps[0]), .Y(detclk_ps[1]) );
  CKBUFX1 U0_DETCLK_BUF_1_ ( .A(detclk_ps[1]), .Y(detclk_ps[2]) );
  CKBUFX1 U0_DETCLK_BUF_2_ ( .A(detclk_ps[2]), .Y(detclk_ps[3]) );
  CKBUFX1 U0_DETCLK_BUF_3_ ( .A(detclk_ps[3]), .Y(detclk_ps[4]) );
  CKBUFX1 U0_DETCLK_BUF_4_ ( .A(detclk_ps[4]), .Y(detclk_ps[5]) );
  CKBUFX1 U0_DETCLK_BUF_5_ ( .A(detclk_ps[5]), .Y(detclk_ps[6]) );
  CKBUFX1 U0_DETCLK_BUF_6_ ( .A(detclk_ps[6]), .Y(detclk_ps[7]) );
  CKBUFX1 U0_DETCLK_BUF_7_ ( .A(detclk_ps[7]), .Y(detclk_ps[8]) );
  CKBUFX1 U0_DETCLK_BUF_8_ ( .A(detclk_ps[8]), .Y(detclk_ps[9]) );
  CKBUFX1 U0_DETCLK_BUF_9_ ( .A(detclk_ps[9]), .Y(detclk) );
  AND2X1 U0_SCAN_EN ( .A(DI_GPIO[2]), .B(n90), .Y(n6) );
  CKMUX2X1 U0_CLK_MUX ( .D0(i_clk), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(s_clk)
         );
  CKMUX2X1 U0_DCLKMUX ( .D0(RD_DET), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        detclk_ps[0]) );
  CKMUX2X1 U0_ACLKMUX ( .D0(aswkup), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        aswclk_ps[0]) );
  CKBUFX1 U0_MCK_BUF ( .A(i_clk), .Y(x_clk) );
  CKBUFX1 U0_TCK_BUF ( .A(DI_GPIO[4]), .Y(t_di_gpio4) );
  CKBUFX1 U0_BUF_NEG0 ( .A(pmem_clk[0]), .Y(t_pmem_clk) );
  CKBUFX1 U0_BUF_NEG1 ( .A(pmem_csb), .Y(t_pmem_csb) );
  CKBUFX1 U0_BUF_NEG2 ( .A(r_osc_gate), .Y(t_osc_gate) );
  CLKDLX1 U0_MCLK_ICG ( .CK(s_clk), .E(n339), .SE(n91), .ECK(g_clk) );
  CLKDLX1 U0_SRAM_ICG ( .CK(g_clk), .E(sram_en), .SE(n91), .ECK(SRAM_CLK) );
  INVX1 U0_REVIDZ_0_ ( .A(1'b0), .Y(REVID[0]) );
  INVX1 U0_REVIDZ_1_ ( .A(1'b1), .Y(REVID[1]) );
  INVX1 U0_REVIDZ_2_ ( .A(1'b1), .Y(REVID[2]) );
  INVX1 U0_REVIDZ_3_ ( .A(1'b1), .Y(REVID[3]) );
  INVX1 U0_REVIDZ_4_ ( .A(1'b0), .Y(REVID[4]) );
  INVX1 U0_REVIDZ_5_ ( .A(1'b0), .Y(REVID[5]) );
  INVX1 U0_REVIDZ_6_ ( .A(1'b1), .Y(REVID[6]) );
  INVX1 U108 ( .A(n58), .Y(n56) );
  INVX1 U120 ( .A(n58), .Y(n57) );
  INVX1 U175 ( .A(srstz), .Y(n58) );
  MUX2X1 U1009 ( .D0(n653), .D1(DUMMY_IN[7]), .S(n6), .Y(DO_GPIO[6]) );
  MUX2X1 U1010 ( .D0(n654), .D1(PMEM_A[15]), .S(n6), .Y(DO_GPIO[5]) );
  mpb_a0 u0_mpb ( .i_rd({prl_cany0r, n724}), .i_wr({prl_cany0w, i2c_ev_3}), 
        .wdat0(sse_wdat), .wdat1(prx_fifowdat), .addr0(sse_adr), .addr1(
        prl_cany0adr), .r_i2c_attr(r_i2c_attr), .esfrm_oe(esfrm_oe), 
        .esfrm_we(esfrm_we), .sfrack(sfrack), .esfrm_wdat(esfrm_wdat), 
        .esfrm_adr(esfrm_adr), .mcu_esfr_rdat(mcu_esfrrdat), .delay_rdat(
        delay_inst), .delay_rrdy(ictlr_psrack), .esfrm_rrdy(esfrm_rrdy), 
        .esfrm_rdat(esfrm_rdat), .channel_sel(1'b0), .r_pg0_sel(r_pg0_sel), 
        .dma_w(1'b0), .dma_r(1'b0), .dma_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_wdat({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_ack(), .memaddr(memaddr), 
        .memaddr_c({memaddr_c[15:7], n2, n49, memaddr_c[4], n4, memaddr_c[2:0]}), .memwr(memwr), .memrd(memrd), .memrd_c(memrd_c), .cpurst(o_cpurst), 
        .memdatao(memdatao), .memack(memack), .hit_xd(hit_xd), .hit_xr(hit_xr), 
        .hit_ps(hit_ps), .hit_ps_c(hit_ps_c), .idat_r(mcu_ram_r), .idat_w(
        mcu_ram_w), .idat_adr(idat_adr), .idat_wdat(idat_wdat), .iram_ce(
        iram_ce), .xram_ce(xram_ce), .regx_re(regx_re), .iram_we(iram_we), 
        .xram_we(xram_we), .regx_we(regx_we), .iram_a(iram_a), .xram_a(xram_a), 
        .iram_d(iram_d), .xram_d(xram_d), .iram_rdat({n15, n1136, n1135, n1139, 
        n1140, n1145, sram_rdat}), .xram_rdat({n16, n1136, n1135, n1139, n1140, 
        n1145, sram_rdat}), .regx_rdat(regx_rdat), .bist_en(n22), .bist_wr(
        bist_wr), .bist_adr(bist_adr), .bist_wdat(bist_wdat), .bist_xram(1'b0), 
        .mclk(g_clk), .srstz(n57), .test_si(n644), .test_so(n534), .test_se(n6) );
  mcu51_a0 u0_mcu ( .bclki2c(r_bclk_sel), .pc_ini({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .slp2wakeup(1'b0), .r_hold_mcu(r_hold_mcu), .wdt_slow(1'b0), .wdtov({n644, 
        SYNOPSYS_UNCONNECTED_1}), .mdubsy(), .cs_run(), .t0_intr(t0_intr), 
        .clki2c(g_clk), .clkmdu(g_clk), .clkur0(g_clk), .clktm0(g_clk), 
        .clktm1(g_clk), .clkwdt(g_clk), .i2c_autoack(1'b0), .i2c_con_ens1(), 
        .clkcpu(g_clk), .clkper(g_clk), .reset(n58), .ro(o_cpurst), .port0i({
        n1142, di_gpio[6:4], n1141, di_gpio[2:0]}), .exint_9(fcp_intr), 
        .exint({exint[7:4], n688, n687, exint[1:0]}), .clkcpuen(), .clkperen(), 
        .port0o({SYNOPSYS_UNCONNECTED_2, do_p0}), .port0ff(ff_p0), .rxd0o(
        do_opt[7]), .txd0(do_opt[6]), .rxd0i(dpdm_urx), .rxd0oe(s0_rxdoe), 
        .scli(n508), .sdai(n510), .sclo(mcuo_scl), .sdao(mcuo_sda), 
        .waitstaten(), .mempsack(mempsack), .memack(memack), .memdatai(
        memdatai), .memdatao(memdatao), .memaddr(memaddr), .mempswr(mempswr), 
        .mempsrd(mempsrd), .memwr(memwr), .memrd(memrd), .memdatao_comb({
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10}), .memaddr_comb(
        memaddr_c), .mempswr_comb(), .mempsrd_comb(mempsrd_c), .memwr_comb(), 
        .memrd_comb(memrd_c), .ramdatai({n15, n1136, n1135, n1139, n1140, 
        n1145, sram_rdat}), .ramdatao(idat_wdat), .ramaddr(idat_adr), .ramwe(
        mcu_ram_w), .ramoe(mcu_ram_r), .dbgpo({SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, mcu_dbgpo, mcu_pc}), 
        .sfrack(sfrack), .sfrdatai(sfr_rdat), .sfrdatao(sfr_wdat), .sfraddr(
        sfr_adr), .sfrwe(sfr_w), .sfroe(sfr_r), .esfrm_wrdata(esfrm_wdat), 
        .esfrm_addr(esfrm_adr), .esfrm_we(esfrm_we), .esfrm_oe(esfrm_oe), 
        .esfrm_rddata(mcu_esfrrdat), .test_si2(DI_GPIO[1]), .test_si1(n647), 
        .test_so1(n646), .test_se(n6) );
  ictlr_a0 u0_ictlr ( .bkpt_ena(bkpt_ena), .bkpt_pc(bkpt_pc), .memaddr_c({
        memaddr_c[14:7], n2, n49, memaddr_c[4], n4, memaddr_c[2:0]}), 
        .memaddr(memaddr[14:0]), .mcu_psr_c(mempsrd_c), .mcu_psw(mempswr), 
        .hit_ps_c(hit_ps_c), .hit_ps(hit_ps), .mempsack(ictlr_psack), 
        .memdatao(memdatao), .o_set_hold(set_hold), .o_bkp_hold(bkpt_hold), 
        .o_ofs_inc(ictlr_inc), .o_inst(ictlr_inst), .d_inst(delay_inst), 
        .sfr_psrack(ictlr_psrack), .sfr_psofs(r_inst_ofs), .sfr_psr(r_psrd), 
        .sfr_psw(r_pswr), .dw_rst(prl_c0set), .dw_ena(n26), .sfr_wdat({n69, 
        n67, sfr_wdat[5], n65, n62, n60, n55, n52}), .pmem_pgm(pmem_pgm), 
        .pmem_re(pmem_re), .pmem_csb(pmem_csb), .pmem_clk(pmem_clk), .pmem_a(
        PMEM_A), .pmem_q0(pmem_q0), .pmem_q1(pmem_q1), .pmem_twlb(pmem_twlb), 
        .wd_twlb(wd_twlb), .we_twlb(we_twlb), .pwrdn_rst(pwrdn_rst), 
        .r_pwdn_en(r_otp_pwdn_en), .r_multi(r_otp_wpls), .r_hold_mcu(
        r_hold_mcu), .clk(g_clk), .srst(o_cpurst), .test_si3(n646), .test_si2(
        slvo_sda), .test_si1(n652), .test_so2(n647), .test_so1(n651), 
        .test_se(n6) );
  regbank_a0 u0_regbank ( .srci({di_pro[5], n1137, n1143, di_pro[2], n126, 
        n128}), .lg_pulse_len(lg_pulse_len), .dm_fault(n1138), .cc1_di(cc1_di), 
        .cc2_di(cc2_di), .di_rd_det(di_aswk[2]), .i_tmrf(t0_intr), .i_vcbyval(
        r_xtm[4]), .dnchk_en(o_dodat5_2_), .r_pwrv_upd(r_pwrv_upd), .aswkup(
        aswkup), .lg_dischg(frc_lg_on), .frc_hg_off(frc_hg_off), .ps_pwrdn(
        ps_pwrdn), .r_sleep(r_sleep), .r_pwrdn(r_pwrdn), .r_ocdrv_enz(
        r_ocdrv_enz), .r_osc_stop(r_osc_stop), .r_osc_lo(o_dodat0_15_), 
        .r_osc_gate(r_osc_gate), .r_fw_pwrv(r_fw_pwrv), .r_cvcwr(r_cvcwr[1:0]), 
        .r_cvofs(r_cvofs), .r_otpi_gate(r_otpi_gate), .r_pwrctl(r_pwrctl), 
        .r_pwr_i(DO_PWR_I), .r_cvctl(DO_CVCTL), .r_srcctl(r_srcctl), 
        .r_dpdmctl(r_dpdmctl), .r_ccrx({r_sqlch, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, r_ccrx, r_rxdb_opt}), .r_cctrx(r_cctrx), 
        .r_ccctl(r_ccctl), .r_fcpwr(r_fcpwr), .r_fcpre(r_fcpre), .fcp_r_dat(
        fcp_r_dat), .fcp_r_sta(fcp_r_sta), .fcp_r_msk(fcp_r_msk), .fcp_r_ctl(
        fcp_r_ctl), .fcp_r_crc(fcp_r_crc), .fcp_r_acc(fcp_r_acc), .fcp_r_tui(
        fcp_r_tui), .r_accctl(r_accctl), .r_bclk_sel(r_bclk_sel), .r_dacwr(
        sfr_dacwr), .r_dac_en(r_dac_en[7:0]), .r_sar_en(r_sar_en[7:0]), 
        .r_adofs(r_adofs), .r_isofs(r_isofs), .x_daclsb(x_daclsb), 
        .r_comp_opt({r_comp_opt, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26}), .dac_r_ctl(
        dac_r_ctl), .dac_r_comp(dac_r_comp[7:0]), .dac_r_cmpsta(dac_r_cmpsta), 
        .dac_r_vs(dac_r_vs[63:0]), .REVID(REVID), .atpg_en(n90), .sfr_r(sfr_r), 
        .sfr_w(sfr_w), .set_hold(set_hold), .bkpt_hold(bkpt_hold), .cpurst(
        o_cpurst), .sfr_addr({1'b1, sfr_adr}), .sfr_wdat({n69, n67, 
        sfr_wdat[5], n64, n62, n60, n55, n52}), .sfr_rdat(sfr_rdat), .ff_p0(
        ff_p0), .di_p0({n1142, di_gpio[6:4], n1141, di_gpio[2:0]}), 
        .ictlr_idle(pmem_csb), .ictlr_inc(ictlr_inc), .r_inst_ofs(r_inst_ofs), 
        .r_psrd(r_psrd), .r_pswr(r_pswr), .r_fortxdat(r_fortxdat), 
        .r_fortxrdy(r_fortxrdy), .r_fortxen(r_fortxen), .r_ana_tm(r_ana_tm), 
        .r_gpio_tm(r_gpio_tm), .r_gpio_ie(r_gpio_ie), .r_gpio_oe(r_gpio_oe), 
        .r_gpio_pu(r_pu_gpio), .r_gpio_pd(r_pd_gpio), .r_gpio_s0({N268, N267, 
        N266}), .r_gpio_s1({N265, N264, N263}), .r_gpio_s2({N262, N261, N260}), 
        .r_gpio_s3({N259, N258, N257}), .r_regtrm(r_regtrm), .i_pc(mcu_pc), 
        .i_goidle(pid_goidle), .i_gobusy(pid_gobusy), .i_i2c_idle(sse_idle), 
        .bus_idle(bus_idle), .i2c_stretch(hwi2c_stretch), .i_i2c_rwbuf(
        sse_wdat), .i_i2c_ltbuf(i2c_ltbuf), .i_i2c_ofs(i2c_lt_ofs), .o_intr({
        exint[6], sfr_intr, exint[5:4]}), .r_auto_gdcrc(r_auto_gdcrc), 
        .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), .r_fifopsh(r_fifopsh), 
        .r_fifopop(r_fifopop), .r_unlock(r_unlock), .r_first(r_first), 
        .r_last(r_last), .r_fiforst(r_fiforst), .r_set_cpmsgid(r_set_cpmsgid), 
        .r_txendk(r_txendk), .r_txnumk(r_txnumk), .r_txshrt(r_txshrt), 
        .r_auto_discard(r_auto_discard), .r_hold_mcu(r_hold_mcu), .r_txauto(
        r_txauto), .r_rxords_ena(r_rxords_ena), .r_spec(r_spec), .r_dat_spec(
        r_dat_spec), .r_dat_portrole(r_dat_portrole), .r_dat_datarole(
        r_dat_datarole), .r_discard(r_discard), .r_pshords(r_pshords), 
        .r_pg0_sel(r_pg0_sel), .r_strtch(r_strtch), .r_i2c_attr(r_i2c_attr), 
        .r_i2c_ninc(r_i2c_ninc), .r_hwi2c_en(), .r_i2c_fwnak(r_i2c_fwnak), 
        .r_i2c_fwack(r_i2c_fwack), .r_i2c_deva(r_i2c_deva), .i2c_ev({n724, 
        i2c_ev_6_, slvo_ev[3:2], i2c_ev_3, i2c_ev_2, slvo_ev[1:0]}), 
        .prl_c0set(prl_c0set), .prl_cany0(n25), .prl_discard(prl_discard), 
        .prl_GCTxDone(prl_GCTxDone), .prl_cpmsgid(prl_cpmsgid), .pff_ack(
        pff_ack), .prx_rst(prx_rst), .pff_obsd(pff_obsd), .pff_full(pff_full), 
        .pff_empty(pff_empty), .ptx_ack(ptx_ack), .pff_ptr(pff_ptr), 
        .prx_adpn(prx_adpn), .pff_rdat(pff_rdat), .pff_rxpart(pff_rxpart), 
        .prx_rcvinf(prx_rcvinf), .ptx_fsm(ptx_fsm), .prx_fsm(prx_fsm), 
        .prl_fsm(prl_fsm), .prx_setsta(prx_setsta), .clk_1p0m(clk_1p0m), 
        .clk_500(clk_500), .clk(g_clk), .xrstz(i_rstz), .xclk(s_clk), .dbgpo({
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58}), .srstz(srstz), 
        .prstz(prstz), .test_si2(r_pwm[15]), .test_si1(n651), .test_so2(n20), 
        .test_so1(n650), .test_se(n6) );
  i2cslv_a0 u0_i2cslv ( .i_sda(n509), .i_scl(n507), .o_sda(slvo_sda), .i_deva(
        r_i2c_deva), .i_inc(n686), .i_fwnak(r_i2c_fwnak), .i_fwack(r_i2c_fwack), .o_we(i2c_ev_3), .o_re(slvo_re), .o_r_early(slvo_early), .o_idle(sse_idle), 
        .o_dec(), .o_busev(slvo_ev), .o_ofs(sse_adr), .o_lt_ofs(i2c_lt_ofs), 
        .o_wdat(sse_wdat), .o_lt_buf(i2c_ltbuf), .o_dbgpo({
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66}), .i_rdat(esfrm_rdat), .i_rd_mem(sse_rdrdy), .i_clk(g_clk), .i_rstz(srstz), .i_prefetch(
        sse_prefetch), .test_si(n648), .test_se(n6) );
  updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 u0_updphy ( .i_cc(n27), .i_cc_49(n123), 
        .i_sqlch(di_sqlch), .r_sqlch(r_sqlch), .r_adprx_en(r_ccrx[3]), 
        .r_adp2nd(r_ccrx[2]), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), 
        .r_fifopsh(r_fifopsh), .r_fifopop(r_fifopop), .r_fiforst(r_fiforst), 
        .r_unlock(r_unlock), .r_first(r_first), .r_last(r_last), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_rdy(upd_rdrdy), .r_wdat({n69, n67, 
        sfr_wdat[5], n64, n62, n60, n54, n52}), .r_rdat(esfrm_rdat), 
        .r_txnumk(r_txnumk), .r_txendk(r_txendk), .r_txshrt(r_txshrt), 
        .r_auto_discard(r_auto_discard), .r_txauto(r_txauto), .r_rxords_ena(
        r_rxords_ena), .r_spec(r_spec), .r_dat_spec(r_dat_spec), 
        .r_auto_gdcrc(r_auto_gdcrc), .r_rxdb_opt(r_rxdb_opt), .r_pshords(
        r_pshords), .r_dat_portrole(r_dat_portrole), .r_dat_datarole(
        r_dat_datarole), .r_discard(r_discard), .pid_goidle(pid_goidle), 
        .pid_gobusy(pid_gobusy), .pff_ack(pff_ack), .pff_rdat(pff_rdat), 
        .pff_rxpart(pff_rxpart), .prx_rcvinf(prx_rcvinf), .pff_obsd(pff_obsd), 
        .pff_ptr(pff_ptr), .pff_empty(pff_empty), .pff_full(pff_full), 
        .ptx_ack(ptx_ack), .ptx_cc(ptx_cc), .ptx_oe(ptx_oe), .prx_setsta(
        prx_setsta), .prx_rst(prx_rst), .prl_c0set(prl_c0set), .prl_cany0(
        prl_cany0), .prl_cany0r(prl_cany0r), .prl_cany0w(prl_cany0w), 
        .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_cany0adr(
        prl_cany0adr), .prl_cpmsgid(prl_cpmsgid), .prx_fifowdat(prx_fifowdat), 
        .ptx_fsm(ptx_fsm), .prl_fsm(prl_fsm), .prx_fsm(prx_fsm), .prx_adpn(
        prx_adpn), .dbgpo({SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, upd_dbgpo, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .clk(g_clk), 
        .srstz(prstz), .test_si(bist_r_ctl[3]), .test_so(n11), .test_se(n6) );
  dacmux_a0 u0_dacmux ( .clk(g_clk), .srstz(n56), .i_comp(n1142), .r_comp_opt(
        r_comp_opt), .r_wdat(r_dacwdat), .r_adofs(r_adofs), .r_isofs(r_isofs), 
        .r_wr({r_dacwr, sfr_dacwr[14:8]}), .dacv_wr({wr_dacv, sfr_dacwr[7:0]}), 
        .o_dacv(dac_r_vs), .o_shrst(sh_rst), .o_hold(sh_hold), .o_dac1(DAC1_V), 
        .o_daci_sel(dacmux_sel), .o_dat(dac_r_comp), .r_dac_en(r_dac_en), 
        .r_sar_en(r_sar_en), .o_dactl(dac_r_ctl), .o_cmpsta(dac_r_cmpsta), 
        .x_daclsb(x_daclsb), .o_intr(exint[7]), .o_smpl({
        SYNOPSYS_UNCONNECTED_97, comp_smpl}), .test_si2(r_vcomp[7]), 
        .test_si1(DI_GPIO[0]), .test_so1(n652), .test_se(n6) );
  fcp_a0 u0_fcp ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(1'b0), .intr(
        fcp_intr), .tx_en(fcp_oe), .tx_dat(fcp_do), .r_dat(fcp_r_dat), .r_sta(
        fcp_r_sta), .r_ctl(fcp_r_ctl), .r_msk(fcp_r_msk), .r_crc(fcp_r_crc), 
        .r_acc(fcp_r_acc), .r_dpdmsta(r_accctl), .r_wdat({n69, n67, 
        sfr_wdat[5], n64, n62, n60, n54, n51}), .r_wr(r_fcpwr), .r_re(r_fcpre), 
        .clk(g_clk), .srstz(srstz), .r_tui(fcp_r_tui), .test_si(n649), 
        .test_so(n648), .test_se(n6) );
  cvctl_a0 u0_cvctl ( .r_cvcwr(r_cvcwr), .wdat(r_cvcwdat), .r_sdischg(
        r_sdischg), .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), .r_cvofsx(r_cvofsx), .r_cvofs(r_cvofs), .sdischg_duty(sdischg_duty), .r_hlsb_en(r_pwrctl[4]), 
        .r_hlsb_sel(r_pwrctl[5]), .r_hlsb_freq(r_xtm[5]), .r_hlsb_duty(
        r_xtm[6]), .r_fw_pwrv(r_fw_pwrv), .r_dac0(DO_DAC0), .r_dac3(DAC3_V), 
        .clk_100k(clk_100k), .clk(g_clk), .srstz(srstz), .test_si(d_dodat[15]), 
        .test_se(n6) );
  regx_a0 u0_regx ( .regx_r(regx_re), .regx_w(regx_we), .di_drposc(di_aswk_0), 
        .di_imposc(di_aswk[4]), .di_rd_det(di_aswk[2]), .clk_500k(clk_500k), 
        .r_imp_osc(r_imp_osc), .regx_addr({xram_a[6:4], n7, xram_a[2:0]}), 
        .regx_wdat(xram_d), .regx_rdat(regx_rdat), .regx_hitbst(regx_hitbst), 
        .regx_wrpwm(regx_wrpwm), .regx_wrcvc({r_cvcwr[2], r_cvcwr[5:3]}), 
        .r_sdischg(r_sdischg), .r_bistctl(bist_r_ctl), .r_bistdat(bist_r_dat), 
        .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), .r_cvofsx(r_cvofsx), .r_pwm(
        r_pwm), .regx_wrdac({wr_dacv[17:16], r_dacwr[10:9], wr_dacv[15:8], 
        r_dacwr[8:7]}), .dac_r_vs(dac_r_vs[143:64]), .dac_comp(
        dac_r_comp[17:8]), .r_dac_en(r_dac_en[17:8]), .r_sar_en(r_sar_en[17:8]), .r_aopt(r_aopt), .r_xtm(r_xtm), .r_adummyi(DUMMY_IN), .r_bck0(r_bck0), 
        .r_bck1(r_bck1), .r_bck2({SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, lg_pulse_len}), .r_i2crout({r_i2crout, 
        r_i2cmcu_route, r_i2cslv_route}), .r_xana({r_xana_23, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, r_xana_19, r_xana_18, OCP_SEL, PWREN_HOLD, 
        r_xana}), .di_xana(di_xanav), .lt_gpi(lt_gpi), .di_tst(di_tst), 
        .bkpt_pc(bkpt_pc), .bkpt_ena(bkpt_ena), .we_twlb(we_twlb), .r_vpp_en(
        r_vpp_en), .r_vpp0v_en(r_vpp0v_en), .r_otp_pwdn_en(r_otp_pwdn_en), 
        .r_otp_wpls(r_otp_wpls), .wd_twlb(wd_twlb), .r_sap(r_sap), .r_twlb(
        pmem_twlb), .upd_pwrv(r_pwrv_upd), .ramacc(ramacc), .sse_idle(sse_idle), .bus_idle(bus_idle), .r_do_ts(r_do_ts), .r_dpdo_sel(r_dpdo_sel), 
        .r_dndo_sel(r_dndo_sel), .di_ts(di_ts), .detclk(detclk), .aswclk(
        aswclk), .atpg_en(n91), .di_aswk({di_aswk[4], n1138, di_aswk[2], 1'b0, 
        di_aswk_0}), .clk(g_clk), .rrstz(n57), .test_si2(n11), .test_si1(n20), 
        .test_so1(n19), .test_se(n6) );
  srambist_a0 u0_srambist ( .clk(g_clk), .srstz(srstz), .reg_hit(regx_hitbst), 
        .reg_w(regx_we), .reg_r(regx_re), .reg_wdat(xram_d), .iram_rdat({n15, 
        n1136, n1135, n1139, n1140, n1145, sram_rdat}), .xram_rdat({n16, n1136, 
        n1135, n1139, n1140, n1145, sram_rdat}), .bist_en(bist_en), 
        .bist_xram(), .bist_wr(bist_wr), .bist_adr(bist_adr), .bist_wdat(
        bist_wdat), .o_bistctl(bist_r_ctl), .o_bistdat(bist_r_dat), .test_si(
        n19), .test_se(n6) );
  divclk_a0 u0_divclk ( .mclk(g_clk), .srstz(n56), .atpg_en(n71), .clk_1p0m(
        clk_1p0m), .clk_500k(clk_500k), .clk_100k(clk_100k), .clk_50k(clk_50k), 
        .clk_500(clk_500), .divff_o1(divff_o1), .divff_o2(), .test_si(
        r_sar_en[17]), .test_so(n649), .test_se(n6) );
  glpwm_a0_0 u0_pwm_0_ ( .clk(g_clk), .rstz(n57), .clk_base(clk_50k), .we(
        regx_wrpwm[0]), .wdat(xram_d), .r_pwm(r_pwm[7:0]), .pwm_o(pwm_o[0]), 
        .test_si(n534), .test_se(n6) );
  glpwm_a0_1 u0_pwm_1_ ( .clk(g_clk), .rstz(n57), .clk_base(clk_50k), .we(
        regx_wrpwm[1]), .wdat(xram_d), .r_pwm(r_pwm[15:8]), .pwm_o(pwm_o[1]), 
        .test_si(r_pwm[7]), .test_se(n6) );
  SNPS_CLOCK_GATE_HIGH_core_a0 clk_gate_d_dodat_reg ( .CLK(g_clk), .EN(N568), 
        .ENCLK(net8852), .TE(n6) );
  DLNQX1 r_lt_gpi_reg_0_ ( .D(DI_GPIO[3]), .XG(i_rstz), .Q(r_lt_gpi[0]) );
  DLNQX1 r_lt_gpi_reg_2_ ( .D(DI_GPIO[1]), .XG(i_rstz), .Q(r_lt_gpi[2]) );
  DLNQX1 r_lt_gpi_reg_1_ ( .D(DI_GPIO[2]), .XG(i_rstz), .Q(r_lt_gpi[1]) );
  DLNQX1 r_lt_gpi_reg_3_ ( .D(DI_GPIO[0]), .XG(i_rstz), .Q(r_lt_gpi[3]) );
  SDFFQX1 d_dodat_reg_1_ ( .D(N583), .SIN(d_dodat[0]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[1]) );
  SDFFQX1 d_dodat_reg_0_ ( .D(N584), .SIN(n650), .SMC(n6), .C(net8852), .Q(
        d_dodat[0]) );
  SDFFQX1 d_dodat_reg_5_ ( .D(N579), .SIN(d_dodat[4]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[5]) );
  SDFFQX1 d_dodat_reg_11_ ( .D(N1477), .SIN(d_dodat[10]), .SMC(n6), .C(net8852), .Q(d_dodat[11]) );
  SDFFQX1 d_dodat_reg_12_ ( .D(N572), .SIN(d_dodat[11]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[12]) );
  SDFFQX1 d_dodat_reg_4_ ( .D(N580), .SIN(d_dodat[3]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[4]) );
  SDFFQX1 d_dodat_reg_13_ ( .D(N571), .SIN(d_dodat[12]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[13]) );
  SDFFQX1 d_dodat_reg_15_ ( .D(N569), .SIN(d_dodat[14]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[15]) );
  SDFFQX1 d_dodat_reg_14_ ( .D(N570), .SIN(d_dodat[13]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[14]) );
  SDFFQX1 d_dodat_reg_6_ ( .D(N578), .SIN(d_dodat[5]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[6]) );
  SDFFQX1 d_dodat_reg_9_ ( .D(N575), .SIN(d_dodat[8]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[9]) );
  SDFFQX1 d_dodat_reg_3_ ( .D(N581), .SIN(d_dodat[2]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[3]) );
  SDFFQX1 d_dodat_reg_8_ ( .D(N576), .SIN(d_dodat[7]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[8]) );
  SDFFQX1 d_dodat_reg_10_ ( .D(N1482), .SIN(d_dodat[9]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[10]) );
  SDFFQX1 d_dodat_reg_7_ ( .D(N577), .SIN(d_dodat[6]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[7]) );
  SDFFQX1 d_dodat_reg_2_ ( .D(N582), .SIN(d_dodat[1]), .SMC(n6), .C(net8852), 
        .Q(d_dodat[2]) );
  MUX4X1 U667 ( .D0(n284), .D1(n300), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N266), 
        .S1(N267), .Y(n517) );
  MUX4X1 U666 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N266), .S1(N267), .Y(n516) );
  MUX4X1 U654 ( .D0(n284), .D1(n300), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N260), 
        .S1(N261), .Y(n511) );
  MUX4X1 U653 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N260), .S1(N261), .Y(n503) );
  MUX2X1 U652 ( .D0(n511), .D1(n503), .S(N262), .Y(N448) );
  MUX4X1 U670 ( .D0(n284), .D1(n300), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N263), 
        .S1(N264), .Y(n515) );
  MUX4X1 U669 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N263), .S1(N264), .Y(n514) );
  MUX2X1 U668 ( .D0(n515), .D1(n514), .S(N265), .Y(DO_GPIO[1]) );
  MUX4X1 U650 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N257), .S1(N258), .Y(n500) );
  MUX4X1 U651 ( .D0(n284), .D1(n300), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N257), 
        .S1(N258), .Y(n502) );
  INVX1 U3 ( .A(memaddr_c[6]), .Y(n1) );
  INVX3 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(memaddr_c[3]), .Y(n3) );
  INVX3 U6 ( .A(n3), .Y(n4) );
  INVX1 U7 ( .A(xram_a[3]), .Y(n5) );
  INVX3 U8 ( .A(n5), .Y(n7) );
  AO2222XL U9 ( .A(n1137), .B(n197), .C(mcu_dbgpo[16]), .D(n234), .E(pmem_pgm), 
        .F(n233), .G(comp_smpl[3]), .H(n232), .Y(n198) );
  OR2X1 U10 ( .A(wr_dacv[10]), .B(wr_dacv[9]), .Y(n254) );
  AND2X1 U11 ( .A(r_vpp0v_en), .B(ps_pwrdn), .Y(pwrdn_rst) );
  AND2X1 U12 ( .A(n261), .B(n262), .Y(sse_prefetch) );
  BUFX3 U13 ( .A(memaddr_c[5]), .Y(n49) );
  AO2222XL U14 ( .A(n237), .B(r_accctl[4]), .C(n236), .D(fcp_oe), .E(n213), 
        .F(r_ccctl[0]), .G(n228), .H(n1142), .Y(n203) );
  NOR43XL U15 ( .B(n201), .C(n200), .D(n199), .A(n198), .Y(n202) );
  OAI22X1 U16 ( .A(n243), .B(n341), .C(n245), .D(n212), .Y(n221) );
  AOI211X1 U17 ( .C(n1099), .D(n230), .A(n218), .B(n217), .Y(n219) );
  AOI22X1 U18 ( .A(n216), .B(n123), .C(n27), .D(n214), .Y(n8) );
  MUX2X1 U19 ( .D0(xram_d[0]), .D1(n52), .S(n260), .Y(r_dacwdat[0]) );
  MUX2X1 U20 ( .D0(n517), .D1(n516), .S(N268), .Y(DO_GPIO[0]) );
  AOI21AX1 U21 ( .B(SRAM_RDAT[7]), .C(n98), .A(n783), .Y(n10) );
  OA21X1 U22 ( .B(hit_xr), .C(hit_xd), .A(memrd), .Y(n12) );
  INVX8 U23 ( .A(n30), .Y(PMEM_PGM) );
  INVXL U24 ( .A(n12), .Y(n13) );
  INVXL U25 ( .A(n12), .Y(n14) );
  INVXL U26 ( .A(n10), .Y(n15) );
  INVXL U27 ( .A(n10), .Y(n16) );
  BUFX3 U28 ( .A(iram_ce), .Y(n17) );
  BUFX3 U29 ( .A(xram_ce), .Y(n18) );
  BUFX3 U30 ( .A(n345), .Y(PMEM_TWLB[0]) );
  NOR21XL U31 ( .B(pmem_twlb[0]), .A(atpg_en), .Y(n345) );
  BUFX3 U32 ( .A(bist_en), .Y(n22) );
  BUFX3 U33 ( .A(n344), .Y(PMEM_TWLB[1]) );
  NOR21XL U34 ( .B(pmem_twlb[1]), .A(atpg_en), .Y(n344) );
  NOR8X1 U35 ( .A(n259), .B(wr_dacv[13]), .C(n258), .D(n257), .E(n256), .F(
        r_dacwr[7]), .G(n255), .H(n254), .Y(n260) );
  INVX1 U36 ( .A(prl_cany0), .Y(n24) );
  INVX1 U37 ( .A(n24), .Y(n25) );
  INVX1 U38 ( .A(n24), .Y(n26) );
  BUFX4 U39 ( .A(n347), .Y(PMEM_SAP[0]) );
  NOR21XL U40 ( .B(r_sap[0]), .A(n102), .Y(n347) );
  BUFX4 U41 ( .A(n346), .Y(PMEM_SAP[1]) );
  NOR21XL U42 ( .B(r_sap[1]), .A(atpg_en), .Y(n346) );
  INVX1 U43 ( .A(n348), .Y(n30) );
  NOR21XL U44 ( .B(pmem_pgm), .A(n102), .Y(n348) );
  MUX2X1 U45 ( .D0(xram_d[1]), .D1(n55), .S(n50), .Y(r_dacwdat[1]) );
  OR2X2 U46 ( .A(wr_dacv[12]), .B(wr_dacv[11]), .Y(n255) );
  OR2X2 U47 ( .A(wr_dacv[17]), .B(wr_dacv[16]), .Y(n258) );
  MUX2XL U48 ( .D0(xram_d[7]), .D1(n69), .S(n50), .Y(r_dacwdat[7]) );
  MUX2XL U49 ( .D0(xram_d[5]), .D1(sfr_wdat[5]), .S(n50), .Y(r_dacwdat[5]) );
  MUX2XL U50 ( .D0(xram_d[2]), .D1(sfr_wdat[2]), .S(n50), .Y(r_dacwdat[2]) );
  MUX2XL U51 ( .D0(xram_d[3]), .D1(n62), .S(n50), .Y(r_dacwdat[3]) );
  XNOR2XL U52 ( .A(n32), .B(n224), .Y(N580) );
  XOR3X1 U53 ( .A(n223), .B(dacmux_sel[4]), .C(n222), .Y(n32) );
  AO22XL U54 ( .A(iram_a[6]), .B(iram_ce), .C(xram_a[6]), .D(xram_ce), .Y(
        SRAM_A[6]) );
  AO22XL U55 ( .A(iram_a[5]), .B(iram_ce), .C(xram_a[5]), .D(xram_ce), .Y(
        SRAM_A[5]) );
  XNOR2XL U56 ( .A(n33), .B(n205), .Y(N578) );
  XNOR3X1 U57 ( .A(n653), .B(SRAM_D[2]), .C(SRAM_A[6]), .Y(n33) );
  XOR3X1 U58 ( .A(n204), .B(dacmux_sel[6]), .C(DAC1_V[0]), .Y(n205) );
  XNOR2XL U59 ( .A(n34), .B(n250), .Y(N579) );
  XNOR3X1 U60 ( .A(n654), .B(SRAM_A[5]), .C(SRAM_D[1]), .Y(n34) );
  XOR3X1 U61 ( .A(n249), .B(dacmux_sel[5]), .C(DO_PWR_I[5]), .Y(n250) );
  OR4X1 U62 ( .A(n248), .B(n247), .C(n35), .D(n36), .Y(n654) );
  OAI222XL U63 ( .A(n995), .B(n242), .C(n241), .D(n240), .E(n239), .F(n238), 
        .Y(n35) );
  OAI222XL U64 ( .A(n775), .B(n246), .C(n916), .D(n245), .E(n244), .F(n243), 
        .Y(n36) );
  INVX1 U65 ( .A(fcp_oe), .Y(n320) );
  NOR21XL U66 ( .B(r_srcctl[7]), .A(n85), .Y(DO_SRCCTL[7]) );
  NOR21XL U67 ( .B(r_srcctl[6]), .A(n87), .Y(DO_SRCCTL[6]) );
  NOR21XL U68 ( .B(r_ccctl[1]), .A(n84), .Y(DO_CCCTL[1]) );
  NOR21XL U69 ( .B(r_aopt[1]), .A(n80), .Y(ANAOPT[1]) );
  NOR21XL U70 ( .B(r_aopt[4]), .A(n80), .Y(ANAOPT[4]) );
  NOR21XL U71 ( .B(r_xana[12]), .A(n80), .Y(ANA_REGX[12]) );
  NOR21XL U72 ( .B(r_xana[2]), .A(n81), .Y(ANA_REGX[2]) );
  NOR21XL U73 ( .B(r_xana[4]), .A(n81), .Y(ANA_REGX[4]) );
  NOR21XL U74 ( .B(r_xana[6]), .A(n81), .Y(ANA_REGX[6]) );
  NOR21XL U75 ( .B(r_xana[8]), .A(n82), .Y(ANA_REGX[8]) );
  NOR21XL U76 ( .B(r_xana[9]), .A(n82), .Y(ANA_REGX[9]) );
  NOR21XL U77 ( .B(r_ccctl[2]), .A(n84), .Y(DO_CCCTL[2]) );
  NOR21XL U78 ( .B(r_ccctl[3]), .A(n84), .Y(DO_CCCTL[3]) );
  INVX1 U79 ( .A(n103), .Y(n78) );
  INVX1 U80 ( .A(n103), .Y(n77) );
  INVX1 U81 ( .A(n92), .Y(n76) );
  INVX1 U82 ( .A(n92), .Y(n75) );
  INVX1 U83 ( .A(n96), .Y(n74) );
  INVX1 U84 ( .A(n97), .Y(n72) );
  INVX1 U85 ( .A(n101), .Y(n73) );
  INVX1 U86 ( .A(n99), .Y(n79) );
  INVX1 U87 ( .A(n100), .Y(n83) );
  INVX1 U88 ( .A(n92), .Y(n80) );
  INVX1 U89 ( .A(n103), .Y(n81) );
  INVX1 U90 ( .A(n98), .Y(n82) );
  INVX1 U91 ( .A(n93), .Y(n84) );
  INVX1 U92 ( .A(n93), .Y(n86) );
  INVX1 U93 ( .A(n103), .Y(n85) );
  INVX1 U94 ( .A(n93), .Y(n87) );
  INVX1 U95 ( .A(n94), .Y(n71) );
  INVX1 U96 ( .A(n95), .Y(n88) );
  INVX1 U97 ( .A(n97), .Y(n90) );
  INVX1 U98 ( .A(n94), .Y(n91) );
  INVX1 U99 ( .A(n63), .Y(n62) );
  INVX1 U100 ( .A(r_dacwr[8]), .Y(n253) );
  OR4X1 U101 ( .A(n1117), .B(n1108), .C(n942), .D(n922), .Y(n37) );
  INVX1 U102 ( .A(n215), .Y(n230) );
  NAND21X1 U103 ( .B(n266), .A(n103), .Y(SRAM_CEB) );
  INVX1 U104 ( .A(n264), .Y(n265) );
  NAND43X1 U105 ( .B(r_cvcwr[2]), .C(r_cvcwr[5]), .D(r_cvcwr[4]), .A(n263), 
        .Y(n264) );
  INVX1 U106 ( .A(r_cvcwr[3]), .Y(n263) );
  INVX1 U107 ( .A(n1108), .Y(n176) );
  INVX1 U109 ( .A(n922), .Y(n243) );
  INVX1 U110 ( .A(n1117), .Y(n183) );
  INVX1 U111 ( .A(n53), .Y(n52) );
  INVX1 U112 ( .A(n61), .Y(n60) );
  INVX1 U113 ( .A(n66), .Y(n64) );
  INVX1 U114 ( .A(n70), .Y(n69) );
  INVX1 U115 ( .A(n68), .Y(n67) );
  INVX1 U116 ( .A(n59), .Y(n55) );
  INVX1 U117 ( .A(n66), .Y(n65) );
  INVX1 U118 ( .A(n59), .Y(n54) );
  INVX1 U119 ( .A(n53), .Y(n51) );
  INVX1 U121 ( .A(n103), .Y(n89) );
  INVX1 U122 ( .A(n102), .Y(n94) );
  INVX1 U123 ( .A(n91), .Y(n98) );
  INVX1 U124 ( .A(atpg_en), .Y(n96) );
  INVX1 U125 ( .A(n102), .Y(n97) );
  INVX1 U126 ( .A(atpg_en), .Y(n99) );
  INVX1 U127 ( .A(n102), .Y(n100) );
  INVX1 U128 ( .A(n102), .Y(n101) );
  INVX1 U129 ( .A(atpg_en), .Y(n95) );
  INVX1 U130 ( .A(n102), .Y(n92) );
  INVX1 U131 ( .A(atpg_en), .Y(n93) );
  NAND21X1 U132 ( .B(r_dacwr[10]), .A(n252), .Y(n257) );
  NAND21X1 U133 ( .B(wr_dacv[8]), .A(n253), .Y(n256) );
  INVX1 U134 ( .A(r_dacwr[9]), .Y(n252) );
  INVX1 U135 ( .A(sfr_wdat[3]), .Y(n63) );
  NAND43X1 U136 ( .B(n237), .C(n236), .D(n234), .A(n242), .Y(n1108) );
  OR4X1 U137 ( .A(n37), .B(n193), .C(n196), .D(n192), .Y(n215) );
  OR2X1 U138 ( .A(n191), .B(n197), .Y(n922) );
  OAI31XL U139 ( .A(n192), .B(n196), .C(n37), .D(n269), .Y(n267) );
  INVX1 U140 ( .A(n213), .Y(n242) );
  INVX1 U141 ( .A(sram_en), .Y(n266) );
  INVX1 U142 ( .A(n958), .Y(n284) );
  INVX1 U143 ( .A(n863), .Y(SRAM_D[7]) );
  OR2X1 U144 ( .A(n214), .B(n216), .Y(n227) );
  OR2X1 U145 ( .A(n228), .B(n227), .Y(n1117) );
  NAND21X1 U146 ( .B(n232), .A(n179), .Y(n192) );
  OR2X1 U147 ( .A(n235), .B(n231), .Y(n942) );
  INVX1 U148 ( .A(n233), .Y(n179) );
  INVX1 U149 ( .A(n196), .Y(n245) );
  INVX1 U150 ( .A(n237), .Y(n239) );
  INVX1 U151 ( .A(n236), .Y(n241) );
  INVX1 U152 ( .A(n232), .Y(n181) );
  INVX1 U153 ( .A(s0_rxdoe), .Y(n338) );
  XOR2X1 U154 ( .A(DAC3_V[4]), .B(n864), .Y(n223) );
  INVX1 U155 ( .A(n864), .Y(SRAM_D[0]) );
  INVX1 U156 ( .A(sfr_wdat[0]), .Y(n53) );
  NOR2X1 U157 ( .A(n298), .B(n304), .Y(n1015) );
  INVX1 U158 ( .A(sfr_wdat[4]), .Y(n66) );
  INVX1 U159 ( .A(sfr_wdat[6]), .Y(n68) );
  INVX1 U160 ( .A(sfr_wdat[7]), .Y(n70) );
  INVX1 U161 ( .A(sfr_wdat[2]), .Y(n61) );
  INVX1 U162 ( .A(sfr_wdat[1]), .Y(n59) );
  NOR2X1 U163 ( .A(n89), .B(n287), .Y(STB_RP) );
  OAI21X1 U164 ( .B(xram_we), .C(iram_we), .A(n93), .Y(SRAM_WEB) );
  AOI21X1 U165 ( .B(n297), .C(n303), .A(n91), .Y(CCI2C_EN) );
  OR2X1 U166 ( .A(iram_we), .B(xram_we), .Y(n993) );
  NOR2X1 U167 ( .A(n88), .B(n277), .Y(OSC_STOP) );
  NOR2X1 U168 ( .A(n88), .B(n281), .Y(DO_SRCCTL[0]) );
  NOR2X1 U169 ( .A(n88), .B(n279), .Y(DO_SRCCTL[3]) );
  NOR2X1 U170 ( .A(n89), .B(n278), .Y(DO_SRCCTL[2]) );
  NOR2X1 U171 ( .A(n89), .B(n274), .Y(OSC_LOW) );
  XOR2X1 U172 ( .A(DO_DAC0[0]), .B(DAC3_V[5]), .Y(n249) );
  INVX1 U173 ( .A(n193), .Y(n269) );
  INVX1 U174 ( .A(n103), .Y(n102) );
  INVX1 U176 ( .A(n1120), .Y(n167) );
  XOR2X1 U177 ( .A(n210), .B(n209), .Y(N570) );
  XOR3X1 U178 ( .A(dacmux_sel[14]), .B(DAC1_V[8]), .C(n206), .Y(n210) );
  XOR3X1 U179 ( .A(n266), .B(n208), .C(n868), .Y(n209) );
  XOR2X1 U180 ( .A(DO_DAC0[9]), .B(TX_EN), .Y(n206) );
  INVX1 U181 ( .A(n987), .Y(n208) );
  OAI22X1 U182 ( .A(n895), .B(n315), .C(n287), .D(n314), .Y(n1034) );
  INVX1 U183 ( .A(r_xana_19), .Y(n287) );
  MUX2X1 U184 ( .D0(xram_d[4]), .D1(n65), .S(n50), .Y(r_dacwdat[4]) );
  NOR21XL U185 ( .B(dacmux_sel[9]), .A(n72), .Y(SAMPL_SEL[9]) );
  NOR21XL U186 ( .B(dacmux_sel[8]), .A(n72), .Y(SAMPL_SEL[8]) );
  NOR21XL U187 ( .B(dacmux_sel[7]), .A(n72), .Y(SAMPL_SEL[7]) );
  NOR21XL U188 ( .B(dacmux_sel[5]), .A(n72), .Y(SAMPL_SEL[5]) );
  NOR21XL U189 ( .B(dacmux_sel[4]), .A(n72), .Y(SAMPL_SEL[4]) );
  NOR21XL U190 ( .B(dacmux_sel[12]), .A(n73), .Y(SAMPL_SEL[12]) );
  NOR21XL U191 ( .B(dacmux_sel[6]), .A(n72), .Y(SAMPL_SEL[6]) );
  NOR21XL U192 ( .B(dacmux_sel[2]), .A(n72), .Y(SAMPL_SEL[2]) );
  NOR21XL U193 ( .B(dacmux_sel[3]), .A(n72), .Y(SAMPL_SEL[3]) );
  NOR21XL U194 ( .B(dacmux_sel[0]), .A(n73), .Y(SAMPL_SEL[0]) );
  NOR21XL U195 ( .B(dacmux_sel[13]), .A(n73), .Y(SAMPL_SEL[13]) );
  NOR21XL U196 ( .B(dacmux_sel[14]), .A(n73), .Y(SAMPL_SEL[14]) );
  NOR21XL U197 ( .B(dacmux_sel[15]), .A(n73), .Y(SAMPL_SEL[15]) );
  NOR21XL U198 ( .B(dacmux_sel[16]), .A(n73), .Y(SAMPL_SEL[16]) );
  NOR21XL U199 ( .B(dacmux_sel[17]), .A(n73), .Y(SAMPL_SEL[17]) );
  NOR21XL U200 ( .B(dacmux_sel[1]), .A(n73), .Y(SAMPL_SEL[1]) );
  XNOR2XL U201 ( .A(n968), .B(n969), .Y(N572) );
  XNOR2XL U202 ( .A(n970), .B(n971), .Y(n969) );
  XNOR2XL U203 ( .A(n275), .B(n972), .Y(n968) );
  XNOR2XL U204 ( .A(dacmux_sel[12]), .B(DO_DAC0[7]), .Y(n970) );
  XOR2X1 U205 ( .A(n152), .B(n151), .Y(N577) );
  XNOR3X1 U206 ( .A(n150), .B(n149), .C(n148), .Y(n152) );
  XOR3X1 U207 ( .A(SRAM_D[3]), .B(SRAM_A[7]), .C(n949), .Y(n151) );
  INVX1 U208 ( .A(DAC1_V[1]), .Y(n149) );
  INVX1 U209 ( .A(n126), .Y(n341) );
  INVX1 U210 ( .A(n289), .Y(o_dodat5_2_) );
  AOI222XL U211 ( .A(n310), .B(di_sqlch), .C(n1063), .D(n272), .E(n312), .F(
        cc1_di), .Y(n1074) );
  AOI222XL U212 ( .A(n310), .B(n123), .C(n1063), .D(TX_DAT), .E(n312), .F(
        cc2_di), .Y(n1062) );
  AOI221XL U213 ( .A(n1026), .B(n1137), .C(n1027), .D(di_pro[5]), .E(n1044), 
        .Y(n1041) );
  OAI22X1 U214 ( .A(n286), .B(n1029), .C(n340), .D(n1030), .Y(n1044) );
  AOI221XL U215 ( .A(n1063), .B(di_pro[5]), .C(n312), .D(n1142), .E(n1064), 
        .Y(n1061) );
  OAI22X1 U216 ( .A(n341), .B(n313), .C(n278), .D(n1065), .Y(n1064) );
  AOI221XL U217 ( .A(n317), .B(n1143), .C(n316), .D(di_pro[2]), .E(n1043), .Y(
        n1042) );
  ENOX1 U218 ( .A(n341), .B(n315), .C(n128), .D(n1026), .Y(n1043) );
  AND2X1 U219 ( .A(dacmux_sel[11]), .B(n94), .Y(SAMPL_SEL[11]) );
  INVX1 U220 ( .A(di_gpio[2]), .Y(n276) );
  INVX1 U221 ( .A(n1138), .Y(n340) );
  NOR2X1 U222 ( .A(n88), .B(n321), .Y(SAMPL_SEL[10]) );
  INVX1 U223 ( .A(dacmux_sel[10]), .Y(n321) );
  MUX2BXL U224 ( .D0(xram_d[6]), .D1(n68), .S(n50), .Y(r_dacwdat[6]) );
  INVX1 U225 ( .A(DO_PWR_I[4]), .Y(n222) );
  OA21X1 U226 ( .B(n216), .C(n228), .A(n123), .Y(n217) );
  AOI222XL U227 ( .A(n800), .B(n817), .C(n802), .D(n818), .E(n304), .F(n819), 
        .Y(n508) );
  AOI222XL U228 ( .A(n800), .B(n801), .C(n802), .D(n803), .E(n304), .F(n804), 
        .Y(n510) );
  OAI22AX1 U229 ( .D(n820), .C(n821), .A(di_gpio[0]), .B(n820), .Y(n817) );
  NAND2X1 U230 ( .A(n816), .B(n334), .Y(n820) );
  EORX1 U231 ( .A(n822), .B(n823), .C(n823), .D(di_gpio[1]), .Y(n821) );
  NAND2X1 U232 ( .A(n811), .B(n333), .Y(n823) );
  INVX1 U233 ( .A(di_pro[5]), .Y(n140) );
  AOI222XL U234 ( .A(n805), .B(n801), .C(n806), .D(n803), .E(n298), .F(n804), 
        .Y(n509) );
  AOI222XL U235 ( .A(n805), .B(n817), .C(n806), .D(n818), .E(n298), .F(n819), 
        .Y(n507) );
  AOI221XL U236 ( .A(n310), .B(di_pro[2]), .C(n1054), .D(n128), .E(n1075), .Y(
        n1073) );
  OAI22X1 U237 ( .A(n1069), .B(n286), .C(n279), .D(n309), .Y(n1075) );
  NOR2X1 U238 ( .A(n89), .B(n322), .Y(SH_RST) );
  NAND21X1 U239 ( .B(n186), .A(n185), .Y(DO_GPIO[2]) );
  AO2222XL U240 ( .A(di_pro[5]), .B(n191), .C(mcu_dbgpo[20]), .D(n177), .E(
        N448), .F(n267), .G(r_osc_stop), .H(n231), .Y(n186) );
  OA2222XL U241 ( .A(n245), .B(n184), .C(n183), .D(n182), .E(n181), .F(n180), 
        .G(n179), .H(n178), .Y(n185) );
  NAND32X1 U242 ( .B(n197), .C(n235), .A(n176), .Y(n177) );
  XNOR2XL U243 ( .A(n288), .B(dacmux_sel[11]), .Y(n1004) );
  XNOR2XL U244 ( .A(r_xana_19), .B(r_srcctl[0]), .Y(n971) );
  XNOR2XL U245 ( .A(n1002), .B(n1003), .Y(N1477) );
  XNOR2XL U246 ( .A(n1005), .B(n871), .Y(n1002) );
  XNOR2XL U247 ( .A(DO_DAC0[6]), .B(n1004), .Y(n1003) );
  XNOR2XL U248 ( .A(DAC1_V[5]), .B(n863), .Y(n1005) );
  XOR2X1 U249 ( .A(n190), .B(n189), .Y(N582) );
  XOR3X1 U250 ( .A(dacmux_sel[2]), .B(DO_PWR_I[2]), .C(n188), .Y(n189) );
  XOR3X1 U251 ( .A(o_dodat5_2_), .B(n187), .C(DO_GPIO[2]), .Y(n190) );
  XOR2X1 U252 ( .A(DAC3_V[2]), .B(n889), .Y(n188) );
  XOR2X1 U253 ( .A(n175), .B(n174), .Y(N581) );
  XNOR3X1 U254 ( .A(n173), .B(dacmux_sel[3]), .C(n172), .Y(n175) );
  XOR3X1 U255 ( .A(n46), .B(DO_GPIO[3]), .C(SRAM_A[3]), .Y(n174) );
  INVX1 U256 ( .A(DO_PWR_I[3]), .Y(n172) );
  INVX1 U257 ( .A(n1142), .Y(n180) );
  INVX1 U258 ( .A(di_pro[2]), .Y(n244) );
  INVX1 U259 ( .A(n1137), .Y(n142) );
  INVX1 U260 ( .A(di_sqlch), .Y(n182) );
  NOR3XL U261 ( .A(n802), .B(n806), .C(n342), .Y(n27) );
  INVX1 U262 ( .A(n123), .Y(n342) );
  INVX1 U263 ( .A(cc2_di), .Y(n165) );
  INVX1 U264 ( .A(cc1_di), .Y(n184) );
  NAND2X1 U265 ( .A(n1143), .B(n191), .Y(n195) );
  OAI2B11X1 U266 ( .D(regx_rdat[7]), .C(n828), .A(n829), .B(n830), .Y(
        memdatai[7]) );
  AOI22X1 U267 ( .A(n831), .B(n16), .C(ictlr_inst[7]), .D(n14), .Y(n830) );
  AOI22X1 U268 ( .A(xram_d[7]), .B(xram_we), .C(iram_we), .D(iram_d[7]), .Y(
        n863) );
  AO22XL U269 ( .A(iram_a[4]), .B(iram_ce), .C(xram_a[4]), .D(xram_ce), .Y(
        SRAM_A[4]) );
  AO21X1 U270 ( .B(n170), .C(n162), .A(n226), .Y(n237) );
  OAI21BBX1 U271 ( .A(n170), .B(n160), .C(n793), .Y(n236) );
  AO21X1 U272 ( .B(n162), .C(n154), .A(n211), .Y(n213) );
  OR2X1 U273 ( .A(n18), .B(n17), .Y(sram_en) );
  OAI22X1 U274 ( .A(n301), .B(n1010), .C(mcuo_scl), .D(n305), .Y(n958) );
  XNOR3X1 U275 ( .A(n38), .B(n39), .C(SRAM_D[6]), .Y(N1482) );
  XNOR3X1 U276 ( .A(DO_DAC0[5]), .B(dacmux_sel[10]), .C(DAC1_V[4]), .Y(n38) );
  XNOR2XL U277 ( .A(n872), .B(SRAM_A[10]), .Y(n39) );
  AO21X1 U278 ( .B(n168), .C(n48), .A(n163), .Y(n191) );
  OAI21BBX1 U279 ( .A(n168), .B(n160), .C(n791), .Y(n234) );
  AO22XL U280 ( .A(iram_a[3]), .B(iram_ce), .C(n7), .D(xram_ce), .Y(SRAM_A[3])
         );
  XOR2X1 U281 ( .A(n129), .B(n127), .Y(N576) );
  XNOR3X1 U282 ( .A(n125), .B(n124), .C(n122), .Y(n129) );
  XOR3X1 U283 ( .A(SRAM_D[4]), .B(SRAM_A[8]), .C(n874), .Y(n127) );
  INVX1 U284 ( .A(DAC1_V[2]), .Y(n124) );
  XOR2X1 U285 ( .A(n118), .B(n117), .Y(N575) );
  XNOR3X1 U286 ( .A(n116), .B(n115), .C(n114), .Y(n118) );
  XOR3X1 U287 ( .A(SRAM_D[5]), .B(SRAM_A[9]), .C(n873), .Y(n117) );
  INVX1 U288 ( .A(DAC1_V[3]), .Y(n115) );
  XOR2X1 U289 ( .A(n137), .B(n136), .Y(N584) );
  XOR3X1 U290 ( .A(DO_PWR_I[0]), .B(DAC3_V[0]), .C(dacmux_sel[16]), .Y(n136)
         );
  XOR3X1 U291 ( .A(dacmux_sel[0]), .B(DO_GPIO[0]), .C(SRAM_A[0]), .Y(n137) );
  XOR2X1 U292 ( .A(n135), .B(n134), .Y(N583) );
  XOR3X1 U293 ( .A(dacmux_sel[17]), .B(DO_PWR_I[1]), .C(n133), .Y(n134) );
  XOR3X1 U294 ( .A(dacmux_sel[1]), .B(n132), .C(SRAM_A[1]), .Y(n135) );
  XOR2X1 U295 ( .A(DAC3_V[1]), .B(DO_GPIO[1]), .Y(n133) );
  OR2X1 U296 ( .A(slvo_early), .B(slvo_re), .Y(n724) );
  INVX1 U297 ( .A(n981), .Y(n337) );
  INVX1 U298 ( .A(n1131), .Y(n157) );
  INVX1 U299 ( .A(n107), .Y(n168) );
  NAND32X1 U300 ( .B(n270), .C(n158), .A(n157), .Y(n107) );
  INVX1 U301 ( .A(SRAM_A[2]), .Y(n187) );
  NOR2X1 U302 ( .A(n89), .B(n949), .Y(DO_TS[3]) );
  NOR2X1 U303 ( .A(n89), .B(n870), .Y(OE_GPIO[4]) );
  NOR2X1 U304 ( .A(n88), .B(n871), .Y(OE_GPIO[3]) );
  NOR2X1 U305 ( .A(n89), .B(n872), .Y(OE_GPIO[2]) );
  INVX1 U306 ( .A(n153), .Y(n170) );
  NAND21X1 U307 ( .B(n270), .A(n1130), .Y(n153) );
  NAND2X1 U308 ( .A(n868), .B(n93), .Y(OE_GPIO[6]) );
  NAND2X1 U309 ( .A(n869), .B(n92), .Y(OE_GPIO[5]) );
  INVX1 U310 ( .A(pwm_o[0]), .Y(n285) );
  OAI2B11X1 U311 ( .D(regx_rdat[5]), .C(n828), .A(n829), .B(n834), .Y(
        memdatai[5]) );
  AOI22X1 U312 ( .A(n831), .B(n1135), .C(ictlr_inst[5]), .D(n14), .Y(n834) );
  OAI2B11X1 U313 ( .D(regx_rdat[3]), .C(n828), .A(n829), .B(n836), .Y(
        memdatai[3]) );
  AOI22X1 U314 ( .A(n831), .B(n1140), .C(ictlr_inst[3]), .D(n14), .Y(n836) );
  OAI2B11X1 U315 ( .D(regx_rdat[4]), .C(n828), .A(n829), .B(n835), .Y(
        memdatai[4]) );
  AOI22X1 U316 ( .A(n831), .B(n1139), .C(ictlr_inst[4]), .D(n13), .Y(n835) );
  OAI2B11X1 U317 ( .D(regx_rdat[6]), .C(n828), .A(n829), .B(n833), .Y(
        memdatai[6]) );
  AOI22X1 U318 ( .A(n831), .B(n1136), .C(ictlr_inst[6]), .D(n14), .Y(n833) );
  OAI21BBX1 U319 ( .A(n154), .B(n48), .C(n786), .Y(n196) );
  AO21X1 U320 ( .B(n162), .C(n168), .A(n225), .Y(n232) );
  AO21X1 U321 ( .B(n160), .C(n154), .A(n138), .Y(n233) );
  OAI2B11X1 U322 ( .D(regx_rdat[2]), .C(n828), .A(n829), .B(n837), .Y(
        memdatai[2]) );
  AOI22X1 U323 ( .A(n831), .B(n1145), .C(ictlr_inst[2]), .D(n13), .Y(n837) );
  OAI21BBX1 U324 ( .A(n168), .B(n167), .C(n787), .Y(n216) );
  OAI21BBX1 U325 ( .A(n166), .B(n48), .C(n784), .Y(n197) );
  AO21X1 U326 ( .B(n166), .C(n162), .A(n161), .Y(n231) );
  OAI2B11X1 U327 ( .D(regx_rdat[1]), .C(n828), .A(n829), .B(n838), .Y(
        memdatai[1]) );
  AOI22X1 U328 ( .A(n831), .B(sram_rdat[1]), .C(ictlr_inst[1]), .D(n13), .Y(
        n838) );
  AO22X1 U329 ( .A(iram_d[5]), .B(iram_we), .C(xram_d[5]), .D(xram_we), .Y(
        SRAM_D[5]) );
  OAI2B11X1 U330 ( .D(regx_rdat[0]), .C(n828), .A(n829), .B(n839), .Y(
        memdatai[0]) );
  AOI22X1 U331 ( .A(n831), .B(sram_rdat[0]), .C(ictlr_inst[0]), .D(n13), .Y(
        n839) );
  AO22X1 U332 ( .A(iram_d[6]), .B(iram_we), .C(xram_d[6]), .D(xram_we), .Y(
        SRAM_D[6]) );
  MUX2X1 U333 ( .D0(xram_d[0]), .D1(n52), .S(n265), .Y(r_cvcwdat[0]) );
  MUX2X1 U334 ( .D0(xram_d[2]), .D1(sfr_wdat[2]), .S(n265), .Y(r_cvcwdat[2])
         );
  MUX2X1 U335 ( .D0(xram_d[1]), .D1(n55), .S(n265), .Y(r_cvcwdat[1]) );
  MUX2X1 U336 ( .D0(xram_d[5]), .D1(sfr_wdat[5]), .S(n265), .Y(r_cvcwdat[5])
         );
  MUX2X1 U337 ( .D0(xram_d[4]), .D1(n65), .S(n265), .Y(r_cvcwdat[4]) );
  MUX2X1 U338 ( .D0(xram_d[6]), .D1(n67), .S(n265), .Y(r_cvcwdat[6]) );
  MUX2BXL U339 ( .D0(xram_d[3]), .D1(n63), .S(n265), .Y(r_cvcwdat[3]) );
  MUX2BXL U340 ( .D0(xram_d[7]), .D1(n70), .S(n265), .Y(r_cvcwdat[7]) );
  AO21X1 U341 ( .B(n170), .C(n48), .A(n169), .Y(n228) );
  OAI21BBX1 U342 ( .A(n166), .B(n160), .C(n792), .Y(n235) );
  OAI21BBX1 U343 ( .A(n166), .B(n167), .C(n788), .Y(n214) );
  NOR2X1 U344 ( .A(n89), .B(n873), .Y(OE_GPIO[1]) );
  NOR2X1 U345 ( .A(n89), .B(n874), .Y(OE_GPIO[0]) );
  INVX1 U346 ( .A(n798), .Y(n211) );
  INVX1 U347 ( .A(n797), .Y(n226) );
  INVX1 U348 ( .A(n796), .Y(n161) );
  INVX1 U349 ( .A(n783), .Y(n163) );
  INVX1 U350 ( .A(n959), .Y(n300) );
  INVX1 U351 ( .A(n805), .Y(n301) );
  INVX1 U352 ( .A(n800), .Y(n305) );
  AO22X1 U353 ( .A(iram_d[4]), .B(iram_we), .C(xram_d[4]), .D(xram_we), .Y(
        SRAM_D[4]) );
  NAND21X1 U354 ( .B(n995), .A(n196), .Y(n201) );
  INVX1 U355 ( .A(n785), .Y(n169) );
  INVX1 U356 ( .A(n795), .Y(n225) );
  INVX1 U357 ( .A(n794), .Y(n138) );
  AO22X1 U358 ( .A(iram_d[3]), .B(iram_we), .C(xram_d[3]), .D(xram_we), .Y(
        SRAM_D[3]) );
  AO22X1 U359 ( .A(iram_d[2]), .B(iram_we), .C(xram_d[2]), .D(xram_we), .Y(
        SRAM_D[2]) );
  INVX1 U360 ( .A(n916), .Y(n272) );
  INVX1 U361 ( .A(n1088), .Y(n141) );
  INVX1 U362 ( .A(n1087), .Y(n139) );
  AOI22X1 U363 ( .A(xram_d[0]), .B(xram_we), .C(iram_d[0]), .D(iram_we), .Y(
        n864) );
  AO22X1 U364 ( .A(iram_d[1]), .B(iram_we), .C(xram_d[1]), .D(xram_we), .Y(
        SRAM_D[1]) );
  NOR2X1 U365 ( .A(n88), .B(n275), .Y(DO_VOOC[0]) );
  NAND21X1 U366 ( .B(n13), .A(hit_xr), .Y(n828) );
  NOR21XL U367 ( .B(n987), .A(n86), .Y(DO_VOOC[2]) );
  NOR2X1 U368 ( .A(n13), .B(hit_xr), .Y(n831) );
  OAI22X1 U369 ( .A(n1010), .B(n297), .C(mcuo_scl), .D(n303), .Y(n155) );
  AOI221XL U370 ( .A(n1026), .B(pwm_o[0]), .C(n1027), .D(pwm_o[1]), .E(n1028), 
        .Y(n1025) );
  OAI22X1 U371 ( .A(n277), .B(n1029), .C(n274), .D(n1030), .Y(n1028) );
  INVX1 U372 ( .A(n46), .Y(CC1_DOB) );
  OAI22X1 U373 ( .A(n281), .B(n1069), .C(n309), .D(n326), .Y(n1068) );
  INVX1 U374 ( .A(r_srcctl[0]), .Y(n281) );
  INVX1 U375 ( .A(r_srcctl[2]), .Y(n278) );
  INVX1 U376 ( .A(r_srcctl[3]), .Y(n279) );
  INVX1 U377 ( .A(n802), .Y(n303) );
  INVX1 U378 ( .A(n806), .Y(n297) );
  NOR21XL U379 ( .B(n978), .A(n86), .Y(DO_VOOC[1]) );
  INVX1 U380 ( .A(n995), .Y(TX_DAT) );
  OAI32X1 U381 ( .A(n313), .B(n318), .C(n336), .D(n309), .E(n319), .Y(n1079)
         );
  OAI22X1 U382 ( .A(n1010), .B(n1048), .C(mcuo_scl), .D(n1049), .Y(n1014) );
  INVX1 U383 ( .A(r_osc_stop), .Y(n277) );
  AND2X1 U384 ( .A(n994), .B(n94), .Y(DO_VOOC[3]) );
  INVX1 U385 ( .A(n1065), .Y(n310) );
  INVX1 U386 ( .A(n1069), .Y(n312) );
  INVX1 U387 ( .A(n979), .Y(n293) );
  INVX1 U388 ( .A(n1029), .Y(n316) );
  INVX1 U389 ( .A(n1063), .Y(n309) );
  INVX1 U390 ( .A(n1027), .Y(n315) );
  INVX1 U391 ( .A(n1049), .Y(n304) );
  INVX1 U392 ( .A(o_dodat0_15_), .Y(n274) );
  INVX1 U393 ( .A(n1048), .Y(n298) );
  INVX1 U394 ( .A(n1054), .Y(n313) );
  INVX1 U395 ( .A(n1026), .Y(n314) );
  XNOR2XL U396 ( .A(n973), .B(n974), .Y(N571) );
  XNOR2XL U397 ( .A(n977), .B(n978), .Y(n973) );
  XNOR2XL U398 ( .A(n975), .B(n976), .Y(n974) );
  XNOR2XL U399 ( .A(n979), .B(n869), .Y(n977) );
  XNOR2XL U400 ( .A(r_srcctl[1]), .B(dacmux_sel[13]), .Y(n976) );
  XNOR2XL U401 ( .A(o_dodat0_15_), .B(dacmux_sel[15]), .Y(n991) );
  XNOR2XL U402 ( .A(n988), .B(n989), .Y(N569) );
  XNOR2XL U403 ( .A(n992), .B(n993), .Y(n988) );
  XNOR2XL U404 ( .A(n990), .B(n991), .Y(n989) );
  XNOR2XL U405 ( .A(n994), .B(n995), .Y(n992) );
  INVX1 U406 ( .A(dacmux_sel[7]), .Y(n148) );
  INVX1 U407 ( .A(dacmux_sel[8]), .Y(n122) );
  INVX1 U408 ( .A(dacmux_sel[9]), .Y(n114) );
  INVX1 U409 ( .A(n1030), .Y(n317) );
  INVX1 U410 ( .A(n47), .Y(CC2_DOB) );
  NOR2X1 U411 ( .A(n916), .B(n87), .Y(TX_EN) );
  NAND2X1 U412 ( .A(n288), .B(n92), .Y(RD_ENB) );
  NOR2X1 U413 ( .A(n88), .B(n889), .Y(BCK_REGX[2]) );
  NOR2X1 U414 ( .A(n90), .B(n289), .Y(ANAOPT[3]) );
  NOR21XL U415 ( .B(PWRDN), .A(n318), .Y(VPP_0V) );
  INVX1 U416 ( .A(r_osc_gate), .Y(n339) );
  NOR2X1 U417 ( .A(n336), .B(n87), .Y(PWRDN) );
  NOR2X1 U418 ( .A(sh_hold), .B(n322), .Y(N568) );
  NOR2X1 U419 ( .A(n88), .B(n895), .Y(BCK_REGX[5]) );
  NOR2X1 U420 ( .A(n88), .B(n884), .Y(DO_SRCCTL[4]) );
  NOR2X1 U421 ( .A(n89), .B(n979), .Y(ANAOPT[5]) );
  OR2X1 U422 ( .A(sh_hold), .B(n91), .Y(SH_HOLD) );
  INVX1 U423 ( .A(di_gpio[0]), .Y(n283) );
  NAND2X1 U424 ( .A(n326), .B(n92), .Y(SLEEP) );
  NOR2X1 U425 ( .A(n88), .B(n319), .Y(BCK_REGX[4]) );
  XOR2X1 U426 ( .A(DAC3_V[3]), .B(n895), .Y(n173) );
  XOR2X1 U427 ( .A(r_srcctl[3]), .B(DO_DAC0[3]), .Y(n125) );
  XOR2X1 U428 ( .A(r_srcctl[2]), .B(DO_DAC0[4]), .Y(n116) );
  XOR2X1 U429 ( .A(DO_PWR_I[7]), .B(DO_DAC0[2]), .Y(n150) );
  XOR2X1 U430 ( .A(DO_PWR_I[6]), .B(DO_DAC0[1]), .Y(n204) );
  XNOR2XL U431 ( .A(DO_DAC0[8]), .B(DAC1_V[7]), .Y(n975) );
  XNOR2XL U432 ( .A(DO_DAC0[10]), .B(DAC1_V[9]), .Y(n990) );
  XNOR2XL U433 ( .A(DAC1_V[6]), .B(n870), .Y(n972) );
  AND2X1 U434 ( .A(n724), .B(n262), .Y(i2c_ev_6_) );
  INVX1 U435 ( .A(n862), .Y(n327) );
  INVX1 U436 ( .A(n884), .Y(n132) );
  OAI21BX1 U437 ( .C(n110), .B(n774), .A(n775), .Y(n193) );
  NOR21XL U438 ( .B(r_srcctl[1]), .A(n86), .Y(DO_SRCCTL[1]) );
  OR2X2 U439 ( .A(pmem_csb), .B(n90), .Y(PMEM_CSB) );
  NAND2X1 U440 ( .A(n271), .B(n343), .Y(n1120) );
  NAND2X1 U441 ( .A(n93), .B(n775), .Y(tclk_sel) );
  INVX1 U442 ( .A(n967), .Y(n121) );
  INVX1 U443 ( .A(atpg_en), .Y(n103) );
  NOR2X1 U444 ( .A(n90), .B(n270), .Y(lt_gpi[0]) );
  NOR2X1 U445 ( .A(n90), .B(n271), .Y(lt_gpi[2]) );
  NOR2X1 U446 ( .A(n90), .B(n343), .Y(lt_gpi[3]) );
  NAND2X1 U447 ( .A(n335), .B(n92), .Y(OCDRV_ENZ) );
  NAND42X1 U448 ( .C(n221), .D(n220), .A(n40), .B(n219), .Y(DO_GPIO[4]) );
  AOI222XL U449 ( .A(dm_comp), .B(n236), .C(upd_dbgpo[18]), .D(n214), .E(
        r_dpdmctl[4]), .F(n237), .Y(n40) );
  AO2222XL U450 ( .A(o_dodat0_15_), .B(n231), .C(n230), .D(n229), .E(n228), 
        .F(dp_comp), .G(upd_dbgpo[17]), .H(n227), .Y(n248) );
  NAND32X1 U451 ( .B(n203), .C(n41), .A(n202), .Y(n653) );
  NAND3X1 U452 ( .A(n195), .B(n194), .C(n8), .Y(n41) );
  AO2222XL U453 ( .A(mcu_dbgpo[19]), .B(n235), .C(mcu_dbgpo[22]), .D(n234), 
        .E(pmem_re), .F(n233), .G(comp_smpl[2]), .H(n232), .Y(n247) );
  MUX4X1 U454 ( .D0(n105), .D1(n1023), .D2(n1036), .D3(n1022), .S0(
        r_dpdo_sel[3]), .S1(r_dpdo_sel[2]), .Y(n987) );
  AO21X1 U455 ( .B(n1019), .C(n273), .A(n1037), .Y(n105) );
  OAI22X1 U456 ( .A(n1041), .B(n273), .C(r_dpdo_sel[1]), .D(n1042), .Y(n1036)
         );
  OAI22X1 U457 ( .A(n1024), .B(n273), .C(r_dpdo_sel[1]), .D(n1025), .Y(n1023)
         );
  NAND4X1 U458 ( .A(n42), .B(n43), .C(n44), .D(n171), .Y(DO_GPIO[3]) );
  AOI21X1 U459 ( .B(n128), .C(n922), .A(n1109), .Y(n42) );
  AOI22X1 U460 ( .A(mcu_dbgpo[16]), .B(n942), .C(mcu_dbgpo[21]), .D(n1108), 
        .Y(n43) );
  OA22X1 U461 ( .A(n245), .B(n165), .C(n179), .D(n164), .Y(n44) );
  OAI21BBX1 U462 ( .A(DRP_OSC), .B(n100), .C(n791), .Y(di_aswk_0) );
  AOI222XL U463 ( .A(comp_smpl[0]), .B(n232), .C(prx_rcvinf[4]), .D(n227), .E(
        n228), .F(n123), .Y(n171) );
  INVX1 U464 ( .A(r_xana_18), .Y(n288) );
  OAI22X1 U465 ( .A(n1032), .B(n273), .C(r_dpdo_sel[1]), .D(n1033), .Y(n1022)
         );
  AOI221XL U466 ( .A(n317), .B(o_dodat5_2_), .C(r_srcctl[5]), .D(n316), .E(
        n1035), .Y(n1032) );
  AOI221XL U467 ( .A(n317), .B(di_aswk[4]), .C(n316), .D(di_aswk_0), .E(n1034), 
        .Y(n1033) );
  OAI22X1 U468 ( .A(n884), .B(n315), .C(n319), .D(n314), .Y(n1035) );
  AOI221XL U469 ( .A(n1026), .B(di_aswk[2]), .C(r_bck0[3]), .D(n1027), .E(
        n1031), .Y(n1024) );
  OAI22X1 U470 ( .A(n889), .B(n1029), .C(n1030), .D(n288), .Y(n1031) );
  AO21X1 U471 ( .B(SRCI[1]), .C(n93), .A(n211), .Y(n126) );
  GEN2XL U472 ( .D(n147), .E(n146), .C(n145), .B(r_do_ts[6]), .A(n144), .Y(
        n949) );
  OA22X1 U473 ( .A(n142), .B(n141), .C(n140), .D(n139), .Y(n146) );
  OA21X1 U474 ( .B(n1084), .C(n291), .A(n143), .Y(n144) );
  AOI21X1 U475 ( .B(n1093), .C(r_do_ts[4]), .A(n290), .Y(n147) );
  AO21X1 U476 ( .B(RX_DAT), .C(n97), .A(n226), .Y(n123) );
  AO21X1 U477 ( .B(SRCI[5]), .C(n101), .A(n138), .Y(di_pro[5]) );
  AO21X1 U478 ( .B(SRCI[2]), .C(n93), .A(n226), .Y(di_pro[2]) );
  AO21X1 U479 ( .B(RX_SQL), .C(n92), .A(n161), .Y(di_sqlch) );
  OAI21BBX1 U480 ( .A(CC2_DI), .B(n101), .C(n792), .Y(cc2_di) );
  OAI21BBX1 U481 ( .A(CC1_DI), .B(n101), .C(n793), .Y(cc1_di) );
  OAI21BBX1 U482 ( .A(DI_GPIO[2]), .B(n100), .C(n788), .Y(di_gpio[2]) );
  OAI21BBX1 U483 ( .A(DM_FAULT), .B(n101), .C(n794), .Y(n1138) );
  AO21X1 U484 ( .B(IMP_OSC), .C(n103), .A(n169), .Y(di_aswk[4]) );
  AO21X1 U485 ( .B(SRCI[0]), .C(n98), .A(n163), .Y(n128) );
  OAI21BBX1 U486 ( .A(DI_GPIO[3]), .B(n99), .C(n787), .Y(n1141) );
  OAI22X1 U487 ( .A(n854), .B(n295), .C(r_i2crout[5]), .D(n855), .Y(dpdm_urx)
         );
  AOI22AXL U488 ( .A(r_pwrctl[7]), .B(n294), .D(r_pwrctl[7]), .C(n856), .Y(
        n854) );
  AOI22X1 U489 ( .A(r_pwrctl[6]), .B(n294), .C(n856), .D(n323), .Y(n855) );
  INVX1 U490 ( .A(n819), .Y(n294) );
  OAI22AX1 U491 ( .D(n840), .C(n841), .A(n283), .B(n840), .Y(exint[1]) );
  NAND2X1 U492 ( .A(n847), .B(N266), .Y(n840) );
  OAI22AX1 U493 ( .D(n842), .C(n843), .A(di_gpio[1]), .B(n842), .Y(n841) );
  NAND3X1 U494 ( .A(N263), .B(n332), .C(N265), .Y(n842) );
  OAI22AX1 U495 ( .D(n848), .C(n849), .A(n283), .B(n848), .Y(exint[0]) );
  NAND2X1 U496 ( .A(n847), .B(n334), .Y(n848) );
  OAI22AX1 U497 ( .D(n850), .C(n851), .A(di_gpio[1]), .B(n850), .Y(n849) );
  NAND3X1 U498 ( .A(n333), .B(n332), .C(N265), .Y(n850) );
  AOI22AXL U499 ( .A(n857), .B(n858), .D(n858), .C(n283), .Y(n856) );
  OAI22AX1 U500 ( .D(n859), .C(n860), .A(di_gpio[1]), .B(n859), .Y(n857) );
  AOI32X1 U501 ( .A(N258), .B(N259), .C(n861), .D(n327), .E(n276), .Y(n860) );
  NOR3XL U502 ( .A(n331), .B(n1141), .C(n327), .Y(n861) );
  XOR2X1 U503 ( .A(r_aopt[3]), .B(n45), .Y(n289) );
  NAND2X1 U504 ( .A(di_aswk[4]), .B(r_imp_osc), .Y(n45) );
  NOR2X1 U505 ( .A(n1141), .B(N258), .Y(n814) );
  AOI32X1 U506 ( .A(n814), .B(n844), .C(n845), .D(n328), .E(n276), .Y(n843) );
  NOR2X1 U507 ( .A(n331), .B(n329), .Y(n845) );
  INVX1 U508 ( .A(n844), .Y(n328) );
  NAND2X1 U509 ( .A(n846), .B(N260), .Y(n844) );
  AOI32X1 U510 ( .A(N259), .B(n814), .C(n852), .D(n853), .E(n276), .Y(n851) );
  NOR2X1 U511 ( .A(N257), .B(n853), .Y(n852) );
  NOR21XL U512 ( .B(n846), .A(N260), .Y(n853) );
  AOI221XL U513 ( .A(n1087), .B(di_xanav[1]), .C(n1088), .D(di_xanav[0]), .E(
        n1091), .Y(n145) );
  OAI21X1 U514 ( .B(n1092), .C(n291), .A(n290), .Y(n1091) );
  AOI22X1 U515 ( .A(r_do_ts[3]), .B(n1143), .C(n126), .D(n292), .Y(n1092) );
  AOI22X1 U516 ( .A(r_dndo_sel[3]), .B(n1059), .C(n1060), .D(n307), .Y(n1052)
         );
  OAI22X1 U517 ( .A(n1066), .B(n308), .C(r_dndo_sel[2]), .D(n1067), .Y(n1059)
         );
  OAI22X1 U518 ( .A(n1061), .B(n308), .C(r_dndo_sel[2]), .D(n1062), .Y(n1060)
         );
  AOI221XL U519 ( .A(n310), .B(o_dodat0_15_), .C(n1054), .D(pwm_o[1]), .E(
        n1068), .Y(n1067) );
  OAI22X1 U520 ( .A(n1038), .B(n273), .C(r_dpdo_sel[1]), .D(n1039), .Y(n1037)
         );
  AOI221XL U521 ( .A(n317), .B(cc2_di), .C(n316), .D(cc1_di), .E(n1040), .Y(
        n1038) );
  AOI22X1 U522 ( .A(n317), .B(n123), .C(n316), .D(di_sqlch), .Y(n1039) );
  OAI22X1 U523 ( .A(n995), .B(n315), .C(n916), .D(n314), .Y(n1040) );
  AOI22X1 U524 ( .A(r_dndo_sel[3]), .B(n1071), .C(n1072), .D(n307), .Y(n1051)
         );
  OAI22X1 U525 ( .A(n1076), .B(n308), .C(r_dndo_sel[2]), .D(n1077), .Y(n1071)
         );
  OAI22X1 U526 ( .A(n1073), .B(n308), .C(r_dndo_sel[2]), .D(n1074), .Y(n1072)
         );
  AOI221XL U527 ( .A(n312), .B(CC1_DOB), .C(n293), .D(n310), .E(n1079), .Y(
        n1076) );
  INVX1 U528 ( .A(n1050), .Y(n275) );
  OAI221X1 U529 ( .A(r_dpdmctl[0]), .B(n1051), .C(n1052), .D(n324), .E(n1053), 
        .Y(n1050) );
  INVX1 U530 ( .A(r_dpdmctl[0]), .Y(n324) );
  OAI211X1 U531 ( .C(fcp_do), .D(n320), .A(n1054), .B(n1055), .Y(n1053) );
  AO21X1 U532 ( .B(DAC1_COMP), .C(n96), .A(n211), .Y(n1142) );
  AO21X1 U533 ( .B(SRCI[4]), .C(n93), .A(n225), .Y(n1137) );
  AO21X1 U534 ( .B(SRCI[3]), .C(n100), .A(n161), .Y(n1143) );
  AO21X1 U535 ( .B(DP_COMP), .C(n99), .A(n225), .Y(dp_comp) );
  OAI21BBX1 U536 ( .A(DM_COMP), .B(n101), .C(n791), .Y(dm_comp) );
  OAI21BBX1 U537 ( .A(RD_DET), .B(n101), .C(n792), .Y(di_aswk[2]) );
  OAI22AX1 U538 ( .D(n807), .C(n808), .A(di_gpio[0]), .B(n807), .Y(n801) );
  NAND2X1 U539 ( .A(N266), .B(n816), .Y(n807) );
  EORX1 U540 ( .A(n809), .B(n810), .C(n810), .D(di_gpio[1]), .Y(n808) );
  NAND2X1 U541 ( .A(N263), .B(n811), .Y(n810) );
  AOI221XL U542 ( .A(n310), .B(di_aswk[4]), .C(n1054), .D(r_vpp_en), .E(n1070), 
        .Y(n1066) );
  OAI22X1 U543 ( .A(n47), .B(n1069), .C(n884), .D(n309), .Y(n1070) );
  AND2X1 U544 ( .A(n1085), .B(n1086), .Y(n143) );
  AOI31X1 U545 ( .A(r_do_ts[5]), .B(dp_comp), .C(n1088), .D(r_do_ts[6]), .Y(
        n1085) );
  OAI21X1 U546 ( .B(n290), .C(dm_comp), .A(n1087), .Y(n1086) );
  AOI21X1 U547 ( .B(n824), .C(di_gpio[2]), .A(n825), .Y(n822) );
  AOI31X1 U548 ( .A(n331), .B(n329), .C(n814), .D(n824), .Y(n825) );
  NOR2X1 U549 ( .A(n815), .B(N260), .Y(n824) );
  AOI21X1 U550 ( .B(n812), .C(di_gpio[2]), .A(n813), .Y(n809) );
  AOI31X1 U551 ( .A(n814), .B(n329), .C(N257), .D(n812), .Y(n813) );
  NOR2X1 U552 ( .A(n330), .B(n815), .Y(n812) );
  ENOX1 U553 ( .A(n340), .B(n292), .C(n292), .D(t_pmem_clk), .Y(n1093) );
  INVX1 U554 ( .A(sh_rst), .Y(n322) );
  OAI21BBX1 U555 ( .A(XANAV[0]), .B(n101), .C(n790), .Y(di_xanav[0]) );
  OAI21BBX1 U556 ( .A(XANAV[1]), .B(n101), .C(n789), .Y(di_xanav[1]) );
  OAI22X1 U557 ( .A(dp_comp), .B(n295), .C(r_i2crout[5]), .D(dm_comp), .Y(n819) );
  OAI22X1 U558 ( .A(r_i2crout[5]), .B(dp_comp), .C(dm_comp), .D(n295), .Y(n804) );
  OAI22X1 U559 ( .A(r_i2crout[4]), .B(cc2_di), .C(cc1_di), .D(n296), .Y(n818)
         );
  OAI22X1 U560 ( .A(cc2_di), .B(n296), .C(r_i2crout[4]), .D(cc1_di), .Y(n803)
         );
  OAI21BBX1 U561 ( .A(DI_GPIO[5]), .B(n100), .C(n785), .Y(di_gpio[5]) );
  OAI21BBX1 U562 ( .A(DI_GPIO[6]), .B(n100), .C(n784), .Y(di_gpio[6]) );
  OAI21BBX1 U563 ( .A(DI_TS), .B(n99), .C(n793), .Y(di_ts) );
  NAND21X1 U564 ( .B(n267), .A(i_rstz), .Y(n981) );
  NOR32XL U565 ( .B(n269), .C(n981), .A(r_gpio_oe[5]), .Y(n869) );
  AO22XL U566 ( .A(iram_a[2]), .B(iram_ce), .C(xram_a[2]), .D(xram_ce), .Y(
        SRAM_A[2]) );
  OAI211X1 U567 ( .C(r_gpio_tm), .D(di_tst), .A(n103), .B(i_rstz), .Y(n1131)
         );
  AO21X1 U568 ( .B(n111), .C(n981), .A(n121), .Y(n872) );
  OAI221X1 U569 ( .A(n862), .B(s0_rxdoe), .C(n815), .D(n1001), .E(r_gpio_oe[2]), .Y(n111) );
  AOI22X1 U570 ( .A(n300), .B(N260), .C(n284), .D(n330), .Y(n1001) );
  AO22XL U571 ( .A(iram_a[1]), .B(iram_ce), .C(xram_a[1]), .D(xram_ce), .Y(
        SRAM_A[1]) );
  AO22XL U572 ( .A(iram_a[0]), .B(iram_ce), .C(xram_a[0]), .D(xram_ce), .Y(
        SRAM_A[0]) );
  AO22X1 U573 ( .A(iram_a[9]), .B(iram_ce), .C(xram_a[9]), .D(xram_ce), .Y(
        SRAM_A[9]) );
  AO22X1 U574 ( .A(iram_a[8]), .B(n17), .C(xram_a[8]), .D(n18), .Y(SRAM_A[8])
         );
  AO22X1 U575 ( .A(iram_a[7]), .B(n17), .C(xram_a[7]), .D(n18), .Y(SRAM_A[7])
         );
  AO22X1 U576 ( .A(iram_a[10]), .B(iram_ce), .C(xram_a[10]), .D(xram_ce), .Y(
        SRAM_A[10]) );
  XNOR2XL U577 ( .A(do_p0[4]), .B(n285), .Y(n1099) );
  XOR2X1 U578 ( .A(do_p0[5]), .B(pwm_o[1]), .Y(n229) );
  OAI21X1 U579 ( .B(n337), .C(n1006), .A(n967), .Y(n871) );
  AND3X1 U580 ( .A(n1007), .B(n1008), .C(r_gpio_oe[3]), .Y(n1006) );
  NAND4X1 U581 ( .A(N258), .B(N259), .C(N257), .D(n338), .Y(n1008) );
  NAND32X1 U582 ( .B(N258), .C(N259), .A(n1009), .Y(n1007) );
  NOR2X1 U583 ( .A(n1131), .B(r_lt_gpi[1]), .Y(n1130) );
  NOR2X1 U584 ( .A(n268), .B(n1110), .Y(n1109) );
  INVX1 U585 ( .A(n267), .Y(n268) );
  AOI22X1 U586 ( .A(n502), .B(n329), .C(n500), .D(N259), .Y(n1110) );
  INVX1 U587 ( .A(n207), .Y(n868) );
  NAND32X1 U588 ( .B(n337), .C(r_gpio_oe[6]), .A(n269), .Y(n207) );
  NOR2X1 U589 ( .A(n337), .B(r_gpio_oe[4]), .Y(n870) );
  OA22X1 U590 ( .A(n1089), .B(n290), .C(n1090), .D(r_do_ts[5]), .Y(n1084) );
  AOI22X1 U591 ( .A(divff_o1), .B(n292), .C(r_do_ts[3]), .D(x_clk), .Y(n1090)
         );
  AOI22X1 U592 ( .A(pwm_o[0]), .B(n292), .C(r_do_ts[3]), .D(pwm_o[1]), .Y(
        n1089) );
  INVX1 U593 ( .A(n109), .Y(n154) );
  NAND21X1 U594 ( .B(r_lt_gpi[0]), .A(n1130), .Y(n109) );
  OAI21BBX1 U595 ( .A(XANAV[2]), .B(n99), .C(n788), .Y(di_xanav[2]) );
  OAI21BBX1 U596 ( .A(XANAV[3]), .B(n99), .C(n787), .Y(di_xanav[3]) );
  OAI21X1 U597 ( .B(pmem_pgm), .C(hwi2c_stretch), .A(r_strtch), .Y(n1010) );
  NAND21X1 U598 ( .B(n94), .A(d_dodat[3]), .Y(n787) );
  NAND21X1 U599 ( .B(n94), .A(d_dodat[2]), .Y(n788) );
  NAND21X1 U600 ( .B(n95), .A(d_dodat[15]), .Y(n791) );
  NAND21X1 U601 ( .B(n95), .A(d_dodat[6]), .Y(n784) );
  NAND21X1 U602 ( .B(n94), .A(d_dodat[14]), .Y(n792) );
  NAND21X1 U603 ( .B(n95), .A(d_dodat[7]), .Y(n783) );
  NAND21X1 U604 ( .B(n95), .A(d_dodat[9]), .Y(n797) );
  NAND21X1 U605 ( .B(n95), .A(d_dodat[10]), .Y(n796) );
  NAND21X1 U606 ( .B(n95), .A(d_dodat[8]), .Y(n798) );
  OAI22X1 U607 ( .A(slvo_sda), .B(n301), .C(mcuo_sda), .D(n305), .Y(n959) );
  NAND32X1 U608 ( .B(n121), .C(n120), .A(r_gpio_oe[0]), .Y(n874) );
  AO22X1 U609 ( .A(n816), .B(n957), .C(n119), .D(n338), .Y(n120) );
  INVX1 U610 ( .A(n858), .Y(n119) );
  OAI22X1 U611 ( .A(N266), .B(n958), .C(n334), .D(n959), .Y(n957) );
  NAND42X1 U612 ( .C(r_pg0_sel[1]), .D(r_pg0_sel[0]), .A(r_pg0_sel[3]), .B(
        r_pg0_sel[2]), .Y(n261) );
  NAND32X1 U613 ( .B(n121), .C(n113), .A(r_gpio_oe[1]), .Y(n873) );
  AO22X1 U614 ( .A(n811), .B(n966), .C(n112), .D(n338), .Y(n113) );
  INVX1 U615 ( .A(n859), .Y(n112) );
  OAI22X1 U616 ( .A(N263), .B(n958), .C(n333), .D(n959), .Y(n966) );
  NAND21X1 U617 ( .B(n215), .A(do_p0[6]), .Y(n194) );
  NOR2X1 U618 ( .A(r_i2cmcu_route[0]), .B(r_i2cmcu_route[1]), .Y(n800) );
  NOR2X1 U619 ( .A(r_i2cslv_route[0]), .B(r_i2cslv_route[1]), .Y(n805) );
  OAI22X1 U620 ( .A(N257), .B(n958), .C(n331), .D(n959), .Y(n1009) );
  NAND2X1 U621 ( .A(d_dodat[13]), .B(n87), .Y(n793) );
  INVX1 U622 ( .A(n159), .Y(n166) );
  NAND32X1 U623 ( .B(r_lt_gpi[0]), .C(n158), .A(n157), .Y(n159) );
  NAND21X1 U624 ( .B(n94), .A(d_dodat[4]), .Y(n786) );
  NAND21X1 U625 ( .B(n95), .A(d_dodat[5]), .Y(n785) );
  NAND21X1 U626 ( .B(n95), .A(d_dodat[12]), .Y(n794) );
  NAND21X1 U627 ( .B(n94), .A(d_dodat[11]), .Y(n795) );
  OA21X1 U628 ( .B(n942), .C(n234), .A(mcu_dbgpo[18]), .Y(n218) );
  INVX1 U629 ( .A(sse_adr[7]), .Y(n262) );
  NAND2X1 U630 ( .A(mcu_dbgpo[17]), .B(n942), .Y(n199) );
  MUX2IX1 U631 ( .D0(ptx_cc), .D1(r_fortxdat), .S(r_fortxrdy), .Y(n995) );
  NAND21X1 U632 ( .B(n92), .A(d_dodat[1]), .Y(n789) );
  NAND21X1 U633 ( .B(n98), .A(d_dodat[0]), .Y(n790) );
  NAND3X1 U634 ( .A(N268), .B(N267), .C(N266), .Y(n858) );
  NOR2X1 U635 ( .A(ptx_oe), .B(r_fortxen), .Y(n916) );
  NOR2X1 U636 ( .A(n306), .B(r_i2cmcu_route[1]), .Y(n802) );
  NOR2X1 U637 ( .A(n302), .B(r_i2cslv_route[1]), .Y(n806) );
  NOR2X1 U638 ( .A(r_do_ts[3]), .B(r_do_ts[4]), .Y(n1088) );
  NOR2X1 U639 ( .A(n292), .B(r_do_ts[4]), .Y(n1087) );
  NAND3X1 U640 ( .A(N262), .B(N260), .C(N261), .Y(n862) );
  OAI31XL U641 ( .A(n826), .B(o_cpurst), .C(hit_ps), .D(n827), .Y(mempsack) );
  NOR2X1 U642 ( .A(mempsrd), .B(mempswr), .Y(n826) );
  NAND2X1 U643 ( .A(ictlr_psack), .B(hit_ps), .Y(n827) );
  INVX1 U644 ( .A(N260), .Y(n330) );
  INVX1 U645 ( .A(N259), .Y(n329) );
  INVX1 U646 ( .A(r_do_ts[3]), .Y(n292) );
  NAND3X1 U647 ( .A(N265), .B(N264), .C(N263), .Y(n859) );
  INVX1 U648 ( .A(r_i2cslv_route[0]), .Y(n302) );
  INVX1 U649 ( .A(r_i2cmcu_route[0]), .Y(n306) );
  INVX1 U655 ( .A(r_do_ts[5]), .Y(n290) );
  INVX1 U656 ( .A(r_do_ts[4]), .Y(n291) );
  INVX1 U657 ( .A(N266), .Y(n334) );
  INVX1 U658 ( .A(N257), .Y(n331) );
  INVX1 U659 ( .A(N263), .Y(n333) );
  NOR2X1 U660 ( .A(N265), .B(N264), .Y(n811) );
  NOR2X1 U661 ( .A(N268), .B(N267), .Y(n816) );
  AOI221XL U662 ( .A(t_osc_gate), .B(n1063), .C(n312), .D(n280), .E(n1078), 
        .Y(n1077) );
  INVX1 U663 ( .A(n889), .Y(n280) );
  OAI22X1 U664 ( .A(n285), .B(n313), .C(n277), .D(n1065), .Y(n1078) );
  OR2X1 U665 ( .A(N262), .B(N261), .Y(n815) );
  INVX1 U671 ( .A(slvo_sda), .Y(n212) );
  INVX1 U672 ( .A(r_vpp_en), .Y(n164) );
  INVX1 U673 ( .A(r_dpdmctl[6]), .Y(n238) );
  INVX1 U674 ( .A(fcp_do), .Y(n240) );
  OAI21BBX1 U675 ( .A(SRAM_RDAT[4]), .B(n98), .C(n786), .Y(n1139) );
  OAI21BBX1 U676 ( .A(SRAM_RDAT[5]), .B(n98), .C(n785), .Y(n1135) );
  OAI21BBX1 U677 ( .A(SRAM_RDAT[6]), .B(n98), .C(n784), .Y(n1136) );
  OAI21BBX1 U678 ( .A(SRAM_RDAT[3]), .B(n98), .C(n787), .Y(n1140) );
  OAI21BBX1 U679 ( .A(SRAM_RDAT[2]), .B(n99), .C(n788), .Y(n1145) );
  OAI21BBX1 U680 ( .A(SRAM_RDAT[0]), .B(n97), .C(n790), .Y(sram_rdat[0]) );
  OAI21BBX1 U681 ( .A(SRAM_RDAT[1]), .B(n99), .C(n789), .Y(sram_rdat[1]) );
  MUX2IX1 U682 ( .D0(n156), .D1(n155), .S(r_i2crout[4]), .Y(n46) );
  NOR21XL U683 ( .B(r_do_ts[2]), .A(n86), .Y(DO_TS[2]) );
  OAI21BBX1 U684 ( .A(hit_ps), .B(mempsrd), .C(n14), .Y(n829) );
  MUX2IX1 U685 ( .D0(n155), .D1(n156), .S(r_i2crout[4]), .Y(n47) );
  NOR21XL U686 ( .B(bist_r_ctl[5]), .A(n72), .Y(SRAM_OEB) );
  NOR2X1 U687 ( .A(r_bck0[2]), .B(frc_hg_off), .Y(n889) );
  OAI22X1 U688 ( .A(mcuo_sda), .B(n303), .C(slvo_sda), .D(n297), .Y(n156) );
  OR2X1 U689 ( .A(r_gpio_ie[1]), .B(n91), .Y(GPIO_IE[1]) );
  AOI211X1 U690 ( .C(n1056), .D(n320), .A(r_dndo_sel[3]), .B(r_dndo_sel[2]), 
        .Y(n1055) );
  OAI21BBX1 U691 ( .A(n1057), .B(r_pwrctl[6]), .C(n1058), .Y(n1056) );
  OAI22X1 U692 ( .A(n295), .B(do_opt[6]), .C(do_opt[7]), .D(r_i2crout[5]), .Y(
        n1057) );
  OAI21BBX1 U693 ( .A(n1015), .B(r_dpdmctl[0]), .C(n323), .Y(n1058) );
  NAND21X1 U694 ( .B(r_otpi_gate), .A(n131), .Y(n884) );
  OA21X1 U695 ( .B(sdischg_duty), .C(n130), .A(r_srcctl[4]), .Y(n131) );
  INVX1 U696 ( .A(r_sdischg[6]), .Y(n130) );
  OAI21BBX1 U697 ( .A(r_xtm[7]), .B(n335), .C(r_aopt[5]), .Y(n979) );
  INVX1 U698 ( .A(r_ocdrv_enz), .Y(n335) );
  NOR2X1 U699 ( .A(n311), .B(r_dndo_sel[0]), .Y(n1063) );
  NOR2X1 U700 ( .A(r_dndo_sel[0]), .B(r_dndo_sel[1]), .Y(n1054) );
  NOR2X1 U701 ( .A(r_dpdo_sel[0]), .B(r_dpdmctl[2]), .Y(n1026) );
  NOR2X1 U702 ( .A(n325), .B(r_dpdo_sel[0]), .Y(n1027) );
  OAI221X1 U703 ( .A(r_pwrctl[7]), .B(n1011), .C(r_i2crout[5]), .D(n299), .E(
        n1012), .Y(n994) );
  OAI21X1 U704 ( .B(s0_rxdoe), .C(n295), .A(r_pwrctl[7]), .Y(n1012) );
  INVX1 U705 ( .A(n1013), .Y(n299) );
  AOI22X1 U706 ( .A(r_i2crout[5]), .B(n1014), .C(r_dpdmctl[3]), .D(n1015), .Y(
        n1011) );
  NAND2X1 U707 ( .A(r_dndo_sel[0]), .B(r_dndo_sel[1]), .Y(n1069) );
  NAND2X1 U708 ( .A(r_dpdo_sel[0]), .B(r_dpdmctl[2]), .Y(n1030) );
  NAND2X1 U709 ( .A(r_dpdo_sel[0]), .B(n325), .Y(n1029) );
  NAND2X1 U710 ( .A(r_dndo_sel[0]), .B(n311), .Y(n1065) );
  NAND2X1 U711 ( .A(r_i2cmcu_route[1]), .B(n306), .Y(n1049) );
  NAND2X1 U712 ( .A(r_i2cslv_route[1]), .B(n302), .Y(n1048) );
  OAI211X1 U713 ( .C(r_pwrctl[6]), .D(n1045), .A(n320), .B(n1046), .Y(n978) );
  AOI22X1 U714 ( .A(r_pwrctl[6]), .B(n1047), .C(r_i2crout[5]), .D(n1013), .Y(
        n1046) );
  AOI22X1 U715 ( .A(n1014), .B(n295), .C(r_dpdmctl[1]), .D(n1015), .Y(n1045)
         );
  NAND2X1 U716 ( .A(n338), .B(n295), .Y(n1047) );
  INVX1 U717 ( .A(r_dpdmctl[2]), .Y(n325) );
  NOR2X1 U718 ( .A(r_bck0[5]), .B(frc_lg_on), .Y(n895) );
  INVX1 U719 ( .A(r_dndo_sel[1]), .Y(n311) );
  AOI211X1 U720 ( .C(r_pwrctl[7]), .D(n1020), .A(r_dpdo_sel[0]), .B(n1021), 
        .Y(n1019) );
  OAI22X1 U721 ( .A(do_opt[7]), .B(n295), .C(r_i2crout[5]), .D(do_opt[6]), .Y(
        n1020) );
  AOI21X1 U722 ( .B(r_dpdmctl[2]), .C(n1015), .A(r_pwrctl[7]), .Y(n1021) );
  INVX1 U723 ( .A(r_bck0[4]), .Y(n319) );
  INVX1 U724 ( .A(r_sleep), .Y(n326) );
  INVX1 U725 ( .A(r_pwrdn), .Y(n336) );
  OAI22X1 U726 ( .A(slvo_sda), .B(n1048), .C(mcuo_sda), .D(n1049), .Y(n1013)
         );
  INVX1 U727 ( .A(r_i2crout[5]), .Y(n295) );
  INVX1 U728 ( .A(r_vpp0v_en), .Y(n318) );
  INVX1 U729 ( .A(r_pwrctl[6]), .Y(n323) );
  INVX1 U730 ( .A(PWREN_HOLD), .Y(n286) );
  NOR21XL U731 ( .B(esfrm_rrdy), .A(n26), .Y(sse_rdrdy) );
  INVX1 U732 ( .A(r_dpdo_sel[1]), .Y(n273) );
  INVX1 U733 ( .A(r_dndo_sel[2]), .Y(n308) );
  INVX1 U734 ( .A(r_dndo_sel[3]), .Y(n307) );
  OAI21BBX1 U735 ( .A(DI_GPIO[0]), .B(n100), .C(n790), .Y(di_gpio[0]) );
  NOR21XL U736 ( .B(r_vpp_en), .A(n72), .Y(VPP_SEL) );
  NOR21XL U737 ( .B(r_dpdmctl[6]), .A(n86), .Y(DO_DPDN[3]) );
  NOR21XL U738 ( .B(r_srcctl[5]), .A(n86), .Y(DO_SRCCTL[5]) );
  NOR21XL U739 ( .B(r_ccctl[0]), .A(n84), .Y(DO_CCCTL[0]) );
  NOR21XL U740 ( .B(r_regtrm[0]), .A(atpg_en), .Y(REGTRM[0]) );
  NOR21XL U741 ( .B(r_regtrm[1]), .A(n78), .Y(REGTRM[1]) );
  NOR21XL U742 ( .B(r_regtrm[3]), .A(n75), .Y(REGTRM[3]) );
  NOR21XL U743 ( .B(r_regtrm[4]), .A(n74), .Y(REGTRM[4]) );
  NOR21XL U744 ( .B(r_regtrm[5]), .A(n74), .Y(REGTRM[5]) );
  NOR21XL U745 ( .B(r_regtrm[6]), .A(n74), .Y(REGTRM[6]) );
  NOR21XL U746 ( .B(r_regtrm[7]), .A(n74), .Y(REGTRM[7]) );
  NOR21XL U747 ( .B(r_regtrm[8]), .A(n73), .Y(REGTRM[8]) );
  NOR21XL U748 ( .B(r_regtrm[9]), .A(n73), .Y(REGTRM[9]) );
  NOR21XL U749 ( .B(r_regtrm[11]), .A(atpg_en), .Y(REGTRM[11]) );
  NOR21XL U750 ( .B(r_regtrm[14]), .A(n78), .Y(REGTRM[14]) );
  NOR21XL U751 ( .B(r_regtrm[15]), .A(n78), .Y(REGTRM[15]) );
  NOR21XL U752 ( .B(r_regtrm[16]), .A(n78), .Y(REGTRM[16]) );
  NOR21XL U753 ( .B(r_regtrm[17]), .A(n78), .Y(REGTRM[17]) );
  NOR21XL U754 ( .B(r_regtrm[19]), .A(n78), .Y(REGTRM[19]) );
  NOR21XL U755 ( .B(r_regtrm[20]), .A(n78), .Y(REGTRM[20]) );
  NOR21XL U756 ( .B(r_regtrm[21]), .A(n77), .Y(REGTRM[21]) );
  NOR21XL U757 ( .B(r_regtrm[22]), .A(n77), .Y(REGTRM[22]) );
  NOR21XL U758 ( .B(r_regtrm[23]), .A(n77), .Y(REGTRM[23]) );
  NOR21XL U759 ( .B(r_regtrm[45]), .A(n75), .Y(REGTRM[45]) );
  NOR21XL U760 ( .B(r_regtrm[46]), .A(n75), .Y(REGTRM[46]) );
  NOR21XL U761 ( .B(r_regtrm[47]), .A(n75), .Y(REGTRM[47]) );
  NOR21XL U762 ( .B(r_regtrm[48]), .A(n75), .Y(REGTRM[48]) );
  NOR21XL U763 ( .B(r_regtrm[49]), .A(n75), .Y(REGTRM[49]) );
  NOR21XL U764 ( .B(r_sdischg[7]), .A(n79), .Y(LDO3P9V) );
  NOR21XL U765 ( .B(r_xtm[0]), .A(n71), .Y(XTM[0]) );
  NOR21XL U766 ( .B(r_xtm[1]), .A(n71), .Y(XTM[1]) );
  NOR21XL U767 ( .B(r_xana[0]), .A(n80), .Y(ANA_REGX[0]) );
  NOR21XL U768 ( .B(r_accctl[4]), .A(n85), .Y(DO_DPDN[0]) );
  NOR21XL U769 ( .B(x_daclsb[2]), .A(n83), .Y(DAC1_EN) );
  NOR21XL U770 ( .B(r_bck0[3]), .A(n83), .Y(BCK_REGX[3]) );
  NOR21XL U771 ( .B(r_xana[15]), .A(n81), .Y(ANA_REGX[15]) );
  NOR21XL U772 ( .B(r_xana[13]), .A(n81), .Y(ANA_REGX[13]) );
  NOR21XL U773 ( .B(r_xana[14]), .A(n81), .Y(ANA_REGX[14]) );
  NOR21XL U774 ( .B(r_xana[1]), .A(n81), .Y(ANA_REGX[1]) );
  NOR21XL U775 ( .B(r_xana[3]), .A(n81), .Y(ANA_REGX[3]) );
  NOR21XL U776 ( .B(r_regtrm[2]), .A(n77), .Y(REGTRM[2]) );
  NOR21XL U777 ( .B(r_regtrm[10]), .A(n91), .Y(REGTRM[10]) );
  NOR21XL U778 ( .B(r_regtrm[12]), .A(n78), .Y(REGTRM[12]) );
  NOR21XL U779 ( .B(r_regtrm[13]), .A(n78), .Y(REGTRM[13]) );
  NOR21XL U780 ( .B(r_regtrm[54]), .A(n74), .Y(REGTRM[54]) );
  NOR21XL U781 ( .B(r_dpdmctl[4]), .A(n85), .Y(DO_DPDN[1]) );
  NOR21XL U782 ( .B(r_regtrm[18]), .A(n78), .Y(REGTRM[18]) );
  NOR21XL U783 ( .B(r_regtrm[24]), .A(n77), .Y(REGTRM[24]) );
  NOR21XL U784 ( .B(r_regtrm[25]), .A(n77), .Y(REGTRM[25]) );
  NOR21XL U785 ( .B(r_regtrm[26]), .A(n77), .Y(REGTRM[26]) );
  NOR21XL U786 ( .B(r_regtrm[27]), .A(n77), .Y(REGTRM[27]) );
  NOR21XL U787 ( .B(r_regtrm[28]), .A(n77), .Y(REGTRM[28]) );
  NOR21XL U788 ( .B(r_regtrm[29]), .A(n77), .Y(REGTRM[29]) );
  NOR21XL U789 ( .B(r_regtrm[30]), .A(n76), .Y(REGTRM[30]) );
  NOR21XL U790 ( .B(r_regtrm[31]), .A(n76), .Y(REGTRM[31]) );
  NOR21XL U791 ( .B(r_regtrm[32]), .A(n76), .Y(REGTRM[32]) );
  NOR21XL U792 ( .B(r_regtrm[33]), .A(n76), .Y(REGTRM[33]) );
  NOR21XL U793 ( .B(r_regtrm[34]), .A(n76), .Y(REGTRM[34]) );
  NOR21XL U794 ( .B(r_regtrm[35]), .A(n76), .Y(REGTRM[35]) );
  NOR21XL U795 ( .B(r_regtrm[36]), .A(n76), .Y(REGTRM[36]) );
  NOR21XL U796 ( .B(r_regtrm[37]), .A(n76), .Y(REGTRM[37]) );
  NOR21XL U797 ( .B(r_regtrm[38]), .A(n76), .Y(REGTRM[38]) );
  NOR21XL U798 ( .B(r_regtrm[39]), .A(n76), .Y(REGTRM[39]) );
  NOR21XL U799 ( .B(r_regtrm[40]), .A(n75), .Y(REGTRM[40]) );
  NOR21XL U800 ( .B(r_regtrm[41]), .A(n75), .Y(REGTRM[41]) );
  NOR21XL U801 ( .B(r_regtrm[42]), .A(n84), .Y(REGTRM[42]) );
  NOR21XL U802 ( .B(r_regtrm[43]), .A(n75), .Y(REGTRM[43]) );
  NOR21XL U803 ( .B(r_regtrm[44]), .A(n75), .Y(REGTRM[44]) );
  NOR21XL U804 ( .B(r_regtrm[50]), .A(n74), .Y(REGTRM[50]) );
  NOR21XL U805 ( .B(r_regtrm[51]), .A(n74), .Y(REGTRM[51]) );
  NOR21XL U806 ( .B(r_regtrm[52]), .A(n74), .Y(REGTRM[52]) );
  NOR21XL U807 ( .B(r_regtrm[53]), .A(n74), .Y(REGTRM[53]) );
  NOR21XL U808 ( .B(r_regtrm[55]), .A(n74), .Y(REGTRM[55]) );
  NOR21XL U809 ( .B(r_aopt[0]), .A(n80), .Y(ANAOPT[0]) );
  NOR21XL U810 ( .B(r_aopt[2]), .A(n80), .Y(ANAOPT[2]) );
  NOR21XL U811 ( .B(r_aopt[6]), .A(n80), .Y(ANAOPT[6]) );
  NOR21XL U812 ( .B(r_aopt[7]), .A(n80), .Y(ANAOPT[7]) );
  NOR21XL U813 ( .B(r_accctl[3]), .A(n86), .Y(DO_DPDN[5]) );
  NOR21XL U814 ( .B(r_xana[5]), .A(n81), .Y(ANA_REGX[5]) );
  NOR21XL U815 ( .B(r_ana_tm[0]), .A(n82), .Y(ANA_TM[0]) );
  NOR21XL U816 ( .B(r_ana_tm[1]), .A(n82), .Y(ANA_TM[1]) );
  NOR21XL U817 ( .B(r_ana_tm[2]), .A(n82), .Y(ANA_TM[2]) );
  NOR21XL U818 ( .B(r_ana_tm[3]), .A(n82), .Y(ANA_TM[3]) );
  NOR21XL U819 ( .B(r_xana[7]), .A(n81), .Y(ANA_REGX[7]) );
  NOR21XL U820 ( .B(r_cctrx[3]), .A(n85), .Y(DO_CCTRX[3]) );
  NOR21XL U821 ( .B(r_xana_23), .A(n79), .Y(LFOSC_ENB) );
  NOR21XL U822 ( .B(r_dpdmctl[5]), .A(n85), .Y(DO_DPDN[2]) );
  NOR21XL U823 ( .B(r_xana[10]), .A(n80), .Y(ANA_REGX[10]) );
  NOR21XL U824 ( .B(r_xana[11]), .A(n80), .Y(ANA_REGX[11]) );
  NOR21XL U825 ( .B(r_dpdmctl[7]), .A(n85), .Y(DO_DPDN[4]) );
  NOR21XL U826 ( .B(r_cctrx[7]), .A(n85), .Y(DO_CCTRX[7]) );
  NOR21XL U827 ( .B(r_cctrx[6]), .A(n85), .Y(DO_CCTRX[6]) );
  NOR21XL U828 ( .B(r_cctrx[5]), .A(n85), .Y(DO_CCTRX[5]) );
  NOR21XL U829 ( .B(r_cctrx[4]), .A(n85), .Y(DO_CCTRX[4]) );
  NOR21XL U830 ( .B(r_xtm[2]), .A(n71), .Y(XTM[2]) );
  NOR21XL U831 ( .B(r_xtm[3]), .A(n71), .Y(XTM[3]) );
  NOR21XL U832 ( .B(r_cctrx[0]), .A(n84), .Y(DO_CCTRX[0]) );
  NOR21XL U833 ( .B(r_ccctl[7]), .A(n84), .Y(DO_CCCTL[7]) );
  NOR21XL U834 ( .B(r_ccctl[6]), .A(n84), .Y(DO_CCCTL[6]) );
  NOR21XL U835 ( .B(r_ccctl[4]), .A(n84), .Y(DO_CCCTL[4]) );
  NOR21XL U836 ( .B(r_ccctl[5]), .A(n84), .Y(DO_CCCTL[5]) );
  NOR21XL U837 ( .B(r_bck0[7]), .A(n83), .Y(BCK_REGX[7]) );
  NOR21XL U838 ( .B(r_bck1[7]), .A(n83), .Y(BCK_REGX[15]) );
  NOR21XL U839 ( .B(r_bck1[6]), .A(n83), .Y(BCK_REGX[14]) );
  NOR21XL U840 ( .B(r_bck1[5]), .A(n83), .Y(BCK_REGX[13]) );
  NOR21XL U841 ( .B(r_bck1[4]), .A(n82), .Y(BCK_REGX[12]) );
  NOR21XL U842 ( .B(r_bck1[3]), .A(n82), .Y(BCK_REGX[11]) );
  NOR21XL U843 ( .B(r_bck1[2]), .A(n82), .Y(BCK_REGX[10]) );
  NOR21XL U844 ( .B(r_bck1[0]), .A(n83), .Y(BCK_REGX[8]) );
  NOR21XL U845 ( .B(r_bck1[1]), .A(n83), .Y(BCK_REGX[9]) );
  NOR21XL U846 ( .B(r_bck0[6]), .A(n83), .Y(BCK_REGX[6]) );
  NOR21XL U847 ( .B(r_bck0[1]), .A(n83), .Y(BCK_REGX[1]) );
  NOR21XL U848 ( .B(r_bck0[0]), .A(n82), .Y(BCK_REGX[0]) );
  OAI21BBX1 U849 ( .A(DI_GPIO[1]), .B(n100), .C(n789), .Y(di_gpio[1]) );
  OR2X1 U850 ( .A(r_cctrx[1]), .B(n91), .Y(DO_CCTRX[1]) );
  OR2X1 U851 ( .A(r_cctrx[2]), .B(n90), .Y(DO_CCTRX[2]) );
  AND2X1 U852 ( .A(esfrm_rrdy), .B(n26), .Y(upd_rdrdy) );
  OR2X1 U853 ( .A(mcu_ram_r), .B(mcu_ram_w), .Y(ramacc) );
  OR2X1 U854 ( .A(r_gpio_ie[0]), .B(n90), .Y(GPIO_IE[0]) );
  INVX1 U857 ( .A(sfr_intr[2]), .Y(n687) );
  NOR21XL U858 ( .B(N262), .A(N261), .Y(n846) );
  NOR21XL U859 ( .B(i2c_ev_3), .A(sse_adr[7]), .Y(i2c_ev_2) );
  NOR21XL U860 ( .B(N268), .A(N267), .Y(n847) );
  INVX1 U861 ( .A(r_i2c_ninc), .Y(n686) );
  INVX1 U862 ( .A(N264), .Y(n332) );
  OAI21BBX1 U863 ( .A(PMEM_Q1[7]), .B(n96), .C(n783), .Y(pmem_q1[7]) );
  OAI21BBX1 U864 ( .A(PMEM_Q0[7]), .B(n97), .C(n791), .Y(pmem_q0[7]) );
  OAI21BBX1 U865 ( .A(PMEM_Q0[1]), .B(n97), .C(n797), .Y(pmem_q0[1]) );
  OAI21BBX1 U866 ( .A(PMEM_Q1[1]), .B(n96), .C(n789), .Y(pmem_q1[1]) );
  OAI21BBX1 U867 ( .A(PMEM_Q1[5]), .B(n96), .C(n785), .Y(pmem_q1[5]) );
  OAI21BBX1 U868 ( .A(PMEM_Q0[5]), .B(n96), .C(n793), .Y(pmem_q0[5]) );
  OAI21BBX1 U869 ( .A(PMEM_Q0[3]), .B(n97), .C(n795), .Y(pmem_q0[3]) );
  OAI21BBX1 U870 ( .A(PMEM_Q1[3]), .B(n96), .C(n787), .Y(pmem_q1[3]) );
  OAI21BBX1 U871 ( .A(PMEM_Q0[2]), .B(n98), .C(n796), .Y(pmem_q0[2]) );
  OAI21BBX1 U872 ( .A(PMEM_Q1[2]), .B(n96), .C(n788), .Y(pmem_q1[2]) );
  OAI21BBX1 U873 ( .A(PMEM_Q0[6]), .B(n97), .C(n792), .Y(pmem_q0[6]) );
  OAI21BBX1 U874 ( .A(PMEM_Q1[6]), .B(n96), .C(n784), .Y(pmem_q1[6]) );
  OAI21BBX1 U875 ( .A(PMEM_Q0[0]), .B(n98), .C(n798), .Y(pmem_q0[0]) );
  OAI21BBX1 U876 ( .A(PMEM_Q1[0]), .B(n97), .C(n790), .Y(pmem_q1[0]) );
  OAI21BBX1 U877 ( .A(PMEM_Q0[4]), .B(n97), .C(n794), .Y(pmem_q0[4]) );
  OAI21BBX1 U878 ( .A(PMEM_Q1[4]), .B(n96), .C(n786), .Y(pmem_q1[4]) );
  INVX1 U879 ( .A(sfr_intr[3]), .Y(n688) );
  INVX1 U880 ( .A(r_i2crout[4]), .Y(n296) );
  OAI21BBX1 U881 ( .A(t_di_gpio4), .B(n100), .C(n786), .Y(di_gpio[4]) );
  OAI21BBX1 U882 ( .A(XANAV[4]), .B(n99), .C(n786), .Y(di_xanav[4]) );
  NOR21X2 U883 ( .B(pmem_re), .A(n102), .Y(PMEM_RE) );
  NOR21X1 U884 ( .B(pmem_clk[0]), .A(n79), .Y(PMEM_CLK[0]) );
  NOR21X1 U885 ( .B(pmem_clk[1]), .A(n102), .Y(PMEM_CLK[1]) );
  NAND43X1 U886 ( .B(r_lt_gpi[1]), .C(n1120), .D(n270), .A(n110), .Y(n775) );
  NAND32X1 U887 ( .B(n1120), .C(r_lt_gpi[0]), .A(n158), .Y(n774) );
  NOR21XL U888 ( .B(r_do_ts[1]), .A(n87), .Y(DO_TS[1]) );
  NOR21XL U889 ( .B(r_do_ts[0]), .A(n86), .Y(DO_TS[0]) );
  NOR21XL U890 ( .B(r_pu_gpio[6]), .A(n79), .Y(GPIO_PU[6]) );
  NOR21XL U891 ( .B(r_pu_gpio[5]), .A(n79), .Y(GPIO_PU[5]) );
  NOR21XL U892 ( .B(r_pu_gpio[4]), .A(n79), .Y(GPIO_PU[4]) );
  NOR21XL U893 ( .B(r_pd_gpio[3]), .A(n86), .Y(GPIO_PD[3]) );
  NOR21XL U894 ( .B(r_pd_gpio[2]), .A(n87), .Y(GPIO_PD[2]) );
  NOR21XL U895 ( .B(r_pd_gpio[1]), .A(n87), .Y(GPIO_PD[1]) );
  NOR21XL U896 ( .B(r_pd_gpio[0]), .A(n87), .Y(GPIO_PD[0]) );
  NOR21XL U897 ( .B(r_pd_gpio[6]), .A(n87), .Y(GPIO_PD[6]) );
  NOR21XL U898 ( .B(r_pd_gpio[5]), .A(n87), .Y(GPIO_PD[5]) );
  NOR21XL U899 ( .B(r_pd_gpio[4]), .A(n86), .Y(GPIO_PD[4]) );
  NOR21XL U900 ( .B(r_pu_gpio[3]), .A(n79), .Y(GPIO_PU[3]) );
  NOR21XL U901 ( .B(r_pu_gpio[2]), .A(n79), .Y(GPIO_PU[2]) );
  NOR21XL U902 ( .B(r_pu_gpio[1]), .A(n79), .Y(GPIO_PU[1]) );
  NOR21XL U903 ( .B(r_pu_gpio[0]), .A(n79), .Y(GPIO_PU[0]) );
  NOR21XL U904 ( .B(di_tst), .A(n774), .Y(tm_atpg) );
  NAND21X1 U905 ( .B(i_rstz), .A(di_tst), .Y(n967) );
  NOR21XL U906 ( .B(r_lt_gpi[1]), .A(n71), .Y(lt_gpi[1]) );
  NAND21X1 U907 ( .B(n775), .A(x_clk), .Y(n200) );
  INVX1 U908 ( .A(r_lt_gpi[3]), .Y(n343) );
  INVX1 U909 ( .A(r_lt_gpi[1]), .Y(n158) );
  INVX1 U910 ( .A(n104), .Y(n110) );
  NAND21X1 U911 ( .B(n90), .A(di_tst), .Y(n104) );
  INVX1 U912 ( .A(r_lt_gpi[2]), .Y(n271) );
  INVX1 U913 ( .A(n106), .Y(n162) );
  NAND21X1 U914 ( .B(r_lt_gpi[2]), .A(r_lt_gpi[3]), .Y(n106) );
  INVX1 U915 ( .A(n108), .Y(n160) );
  NAND21X1 U916 ( .B(n271), .A(r_lt_gpi[3]), .Y(n108) );
  INVX1 U917 ( .A(r_lt_gpi[0]), .Y(n270) );
  AND2X1 U918 ( .A(r_lt_gpi[2]), .B(n343), .Y(n48) );
  INVX1 U919 ( .A(t_pmem_clk), .Y(n178) );
  INVX1 U920 ( .A(i_rstz), .Y(n246) );
  XOR3XL U921 ( .A(n47), .B(SRAM_A[4]), .C(DO_GPIO[4]), .Y(n224) );
  BUFXL U922 ( .A(n260), .Y(n50) );
  AO222X1 U923 ( .A(comp_smpl[1]), .B(n232), .C(n213), .D(n272), .E(t_pmem_csb), .F(n233), .Y(n220) );
  INVX2 U924 ( .A(wr_dacv[14]), .Y(n251) );
  NAND21X1 U925 ( .B(wr_dacv[15]), .A(n251), .Y(n259) );
endmodule


module SNPS_CLOCK_GATE_HIGH_core_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_1 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o, test_si, 
        test_se );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we, test_si, test_se;
  output pwm_o;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, net8870, n1, n2, n3, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [6:0] pwmcnt;

  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  glreg_a0_1 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm), .test_si(pwmcnt[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8870), .TE(test_se) );
  SDFFSQX1 pwmcnt_reg_6_ ( .D(N20), .SIN(pwmcnt[5]), .SMC(test_se), .C(net8870), .XS(n2), .Q(pwmcnt[6]) );
  SDFFSQX1 pwmcnt_reg_4_ ( .D(N18), .SIN(pwmcnt[3]), .SMC(test_se), .C(net8870), .XS(n2), .Q(pwmcnt[4]) );
  SDFFSQX1 pwmcnt_reg_5_ ( .D(N19), .SIN(pwmcnt[4]), .SMC(test_se), .C(net8870), .XS(n2), .Q(pwmcnt[5]) );
  SDFFSQX1 pwmcnt_reg_2_ ( .D(N16), .SIN(pwmcnt[1]), .SMC(test_se), .C(net8870), .XS(n2), .Q(pwmcnt[2]) );
  SDFFSQX1 pwmcnt_reg_1_ ( .D(N15), .SIN(pwmcnt[0]), .SMC(test_se), .C(net8870), .XS(n1), .Q(pwmcnt[1]) );
  SDFFSQX1 pwmcnt_reg_3_ ( .D(N17), .SIN(pwmcnt[2]), .SMC(test_se), .C(net8870), .XS(n2), .Q(pwmcnt[3]) );
  SDFFSQX1 pwmcnt_reg_0_ ( .D(N14), .SIN(test_si), .SMC(test_se), .C(net8870), 
        .XS(n1), .Q(pwmcnt[0]) );
  INVX1 U6 ( .A(n33), .Y(n4) );
  INVX1 U7 ( .A(n36), .Y(n13) );
  INVX1 U8 ( .A(n27), .Y(n8) );
  NOR21XL U9 ( .B(we), .A(wdat[7]), .Y(n33) );
  NAND2X1 U10 ( .A(n5), .B(n4), .Y(N13) );
  INVX1 U11 ( .A(n35), .Y(n12) );
  INVX1 U12 ( .A(n34), .Y(n11) );
  NOR2X1 U13 ( .A(n16), .B(r_pwm[3]), .Y(n27) );
  NOR2X1 U14 ( .A(pwmcnt[1]), .B(pwmcnt[0]), .Y(n36) );
  AOI21X1 U15 ( .B(n24), .C(n25), .A(n19), .Y(n23) );
  AOI32X1 U16 ( .A(n8), .B(n15), .C(r_pwm[2]), .D(r_pwm[3]), .E(n16), .Y(n24)
         );
  OAI221X1 U17 ( .A(n9), .B(n18), .C(r_pwm[2]), .D(n15), .E(n26), .Y(n25) );
  INVX1 U18 ( .A(pwmcnt[2]), .Y(n15) );
  AOI211X1 U19 ( .C(n13), .D(n7), .A(n27), .B(n28), .Y(n26) );
  INVX1 U20 ( .A(r_pwm[1]), .Y(n7) );
  AOI21X1 U21 ( .B(r_pwm[1]), .C(n18), .A(r_pwm[0]), .Y(n28) );
  OAI221X1 U22 ( .A(n19), .B(n20), .C(pwmcnt[6]), .D(n6), .E(n21), .Y(pwm_o)
         );
  AOI32X1 U23 ( .A(n22), .B(n14), .C(r_pwm[4]), .D(r_pwm[5]), .E(n17), .Y(n20)
         );
  OAI211X1 U24 ( .C(r_pwm[4]), .D(n14), .A(n22), .B(n23), .Y(n21) );
  INVX1 U25 ( .A(pwmcnt[4]), .Y(n14) );
  INVX1 U26 ( .A(pwmcnt[3]), .Y(n16) );
  INVX1 U27 ( .A(pwmcnt[1]), .Y(n18) );
  AND2X1 U28 ( .A(pwmcnt[6]), .B(n6), .Y(n19) );
  INVX1 U29 ( .A(r_pwm[6]), .Y(n6) );
  INVX1 U30 ( .A(pwmcnt[0]), .Y(n9) );
  GEN2XL U31 ( .D(pwmcnt[1]), .E(pwmcnt[0]), .C(n36), .B(r_pwm[7]), .A(n33), 
        .Y(N15) );
  GEN2XL U32 ( .D(pwmcnt[2]), .E(n13), .C(n35), .B(r_pwm[7]), .A(n33), .Y(N16)
         );
  GEN2XL U33 ( .D(pwmcnt[4]), .E(n11), .C(n31), .B(r_pwm[7]), .A(n33), .Y(N18)
         );
  GEN2XL U34 ( .D(pwmcnt[3]), .E(n12), .C(n34), .B(r_pwm[7]), .A(n33), .Y(N17)
         );
  NAND21X1 U35 ( .B(r_pwm[5]), .A(pwmcnt[5]), .Y(n22) );
  OAI21X1 U36 ( .B(n32), .C(n5), .A(n4), .Y(N19) );
  XNOR2XL U37 ( .A(n31), .B(pwmcnt[5]), .Y(n32) );
  OAI21X1 U38 ( .B(n29), .C(n5), .A(n4), .Y(N20) );
  XNOR2XL U39 ( .A(pwmcnt[6]), .B(n30), .Y(n29) );
  NOR2X1 U40 ( .A(pwmcnt[5]), .B(n10), .Y(n30) );
  INVX1 U41 ( .A(n31), .Y(n10) );
  OAI21X1 U42 ( .B(pwmcnt[0]), .C(n5), .A(n4), .Y(N14) );
  INVX1 U43 ( .A(pwmcnt[5]), .Y(n17) );
  NOR2X1 U44 ( .A(n11), .B(pwmcnt[4]), .Y(n31) );
  NOR2X1 U45 ( .A(n13), .B(pwmcnt[2]), .Y(n35) );
  NOR2X1 U46 ( .A(n12), .B(pwmcnt[3]), .Y(n34) );
  INVX1 U47 ( .A(r_pwm[7]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8888;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8888), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8888), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8888), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8888), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8888), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8888), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8888), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8888), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8888), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_0 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o, test_si, 
        test_se );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we, test_si, test_se;
  output pwm_o;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, net8906, n1, n2, n3, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [6:0] pwmcnt;

  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  glreg_a0_0 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm), .test_si(pwmcnt[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8906), .TE(test_se) );
  SDFFSQX1 pwmcnt_reg_6_ ( .D(N20), .SIN(pwmcnt[5]), .SMC(test_se), .C(net8906), .XS(n2), .Q(pwmcnt[6]) );
  SDFFSQX1 pwmcnt_reg_4_ ( .D(N18), .SIN(pwmcnt[3]), .SMC(test_se), .C(net8906), .XS(n2), .Q(pwmcnt[4]) );
  SDFFSQX1 pwmcnt_reg_5_ ( .D(N19), .SIN(pwmcnt[4]), .SMC(test_se), .C(net8906), .XS(n2), .Q(pwmcnt[5]) );
  SDFFSQX1 pwmcnt_reg_2_ ( .D(N16), .SIN(pwmcnt[1]), .SMC(test_se), .C(net8906), .XS(n2), .Q(pwmcnt[2]) );
  SDFFSQX1 pwmcnt_reg_3_ ( .D(N17), .SIN(pwmcnt[2]), .SMC(test_se), .C(net8906), .XS(n2), .Q(pwmcnt[3]) );
  SDFFSQX1 pwmcnt_reg_1_ ( .D(N15), .SIN(pwmcnt[0]), .SMC(test_se), .C(net8906), .XS(n1), .Q(pwmcnt[1]) );
  SDFFSQX1 pwmcnt_reg_0_ ( .D(N14), .SIN(test_si), .SMC(test_se), .C(net8906), 
        .XS(n1), .Q(pwmcnt[0]) );
  INVX1 U6 ( .A(n33), .Y(n4) );
  INVX1 U7 ( .A(n36), .Y(n15) );
  INVX1 U8 ( .A(n27), .Y(n8) );
  NOR21XL U9 ( .B(we), .A(wdat[7]), .Y(n33) );
  NAND2X1 U10 ( .A(n5), .B(n4), .Y(N13) );
  INVX1 U11 ( .A(n35), .Y(n13) );
  INVX1 U12 ( .A(n34), .Y(n12) );
  OAI221X1 U13 ( .A(n19), .B(n20), .C(pwmcnt[6]), .D(n6), .E(n21), .Y(pwm_o)
         );
  AOI32X1 U14 ( .A(n22), .B(n9), .C(r_pwm[4]), .D(r_pwm[5]), .E(n16), .Y(n20)
         );
  OAI211X1 U15 ( .C(r_pwm[4]), .D(n9), .A(n22), .B(n23), .Y(n21) );
  INVX1 U16 ( .A(pwmcnt[4]), .Y(n9) );
  NOR2X1 U17 ( .A(pwmcnt[1]), .B(pwmcnt[0]), .Y(n36) );
  AOI21X1 U18 ( .B(n24), .C(n25), .A(n19), .Y(n23) );
  AOI32X1 U19 ( .A(n8), .B(n11), .C(r_pwm[2]), .D(r_pwm[3]), .E(n18), .Y(n24)
         );
  OAI221X1 U20 ( .A(n14), .B(n17), .C(r_pwm[2]), .D(n11), .E(n26), .Y(n25) );
  INVX1 U21 ( .A(pwmcnt[2]), .Y(n11) );
  AOI211X1 U22 ( .C(n15), .D(n7), .A(n27), .B(n28), .Y(n26) );
  INVX1 U23 ( .A(r_pwm[1]), .Y(n7) );
  AOI21X1 U24 ( .B(r_pwm[1]), .C(n17), .A(r_pwm[0]), .Y(n28) );
  INVX1 U25 ( .A(pwmcnt[1]), .Y(n17) );
  NOR2X1 U26 ( .A(n18), .B(r_pwm[3]), .Y(n27) );
  INVX1 U27 ( .A(pwmcnt[3]), .Y(n18) );
  INVX1 U28 ( .A(pwmcnt[0]), .Y(n14) );
  GEN2XL U29 ( .D(pwmcnt[1]), .E(pwmcnt[0]), .C(n36), .B(r_pwm[7]), .A(n33), 
        .Y(N15) );
  GEN2XL U30 ( .D(pwmcnt[2]), .E(n15), .C(n35), .B(r_pwm[7]), .A(n33), .Y(N16)
         );
  GEN2XL U31 ( .D(pwmcnt[4]), .E(n12), .C(n31), .B(r_pwm[7]), .A(n33), .Y(N18)
         );
  GEN2XL U32 ( .D(pwmcnt[3]), .E(n13), .C(n34), .B(r_pwm[7]), .A(n33), .Y(N17)
         );
  NAND21X1 U33 ( .B(r_pwm[5]), .A(pwmcnt[5]), .Y(n22) );
  AND2X1 U34 ( .A(pwmcnt[6]), .B(n6), .Y(n19) );
  OAI21X1 U35 ( .B(n32), .C(n5), .A(n4), .Y(N19) );
  XNOR2XL U36 ( .A(n31), .B(pwmcnt[5]), .Y(n32) );
  OAI21X1 U37 ( .B(pwmcnt[0]), .C(n5), .A(n4), .Y(N14) );
  OAI21X1 U38 ( .B(n29), .C(n5), .A(n4), .Y(N20) );
  XNOR2XL U39 ( .A(pwmcnt[6]), .B(n30), .Y(n29) );
  NOR2X1 U40 ( .A(pwmcnt[5]), .B(n10), .Y(n30) );
  INVX1 U41 ( .A(n31), .Y(n10) );
  INVX1 U42 ( .A(r_pwm[6]), .Y(n6) );
  INVX1 U43 ( .A(pwmcnt[5]), .Y(n16) );
  NOR2X1 U44 ( .A(n12), .B(pwmcnt[4]), .Y(n31) );
  NOR2X1 U45 ( .A(n15), .B(pwmcnt[2]), .Y(n35) );
  NOR2X1 U46 ( .A(n13), .B(pwmcnt[3]), .Y(n34) );
  INVX1 U47 ( .A(r_pwm[7]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8924;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8924), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8924), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8924), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8924), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8924), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8924), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8924), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8924), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8924), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module divclk_a0 ( mclk, srstz, atpg_en, clk_1p0m, clk_500k, clk_100k, clk_50k, 
        clk_500, divff_o1, divff_o2, test_si, test_so, test_se );
  input mclk, srstz, atpg_en, test_si, test_se;
  output clk_1p0m, clk_500k, clk_100k, clk_50k, clk_500, divff_o1, divff_o2,
         test_so;
  wire   div500k_5_0, div1p0m_2, div100k_2, N23, N24, N25, N26, N37, N38, N39,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         n22, n23, n24, n1, n2, n3, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n25, n26, n27, n4, n5, n6, n7, n8, n9, n10;
  wire   [2:0] div12;
  wire   [6:0] div50k_100;

  CLKDLX1 U0_D1P0M_ICG ( .CK(mclk), .E(n22), .SE(atpg_en), .ECK(clk_1p0m) );
  CLKDLX1 U0_D500K_ICG ( .CK(clk_1p0m), .E(div1p0m_2), .SE(atpg_en), .ECK(
        clk_500k) );
  CLKDLX1 U0_D100K_ICG ( .CK(clk_500k), .E(n23), .SE(atpg_en), .ECK(clk_100k)
         );
  CLKDLX1 U0_D50K_ICG ( .CK(clk_100k), .E(div100k_2), .SE(atpg_en), .ECK(
        clk_50k) );
  CLKDLX1 U0_D0P5K_ICG ( .CK(clk_50k), .E(n24), .SE(atpg_en), .ECK(clk_500) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(srstz), .Y(n3) );
  divclk_a0_DW01_inc_0 add_60 ( .A(div50k_100), .SUM({N52, N51, N50, N49, N48, 
        N47, N46}) );
  SDFFRQX1 div1p0m_2_reg ( .D(n4), .SIN(test_si), .SMC(test_se), .C(clk_1p0m), 
        .XR(n1), .Q(div1p0m_2) );
  SDFFRQX1 div100k_2_reg ( .D(n5), .SIN(div50k_100[6]), .SMC(test_se), .C(
        clk_100k), .XR(n1), .Q(div100k_2) );
  SDFFRQX1 div50k_100_reg_6_ ( .D(N59), .SIN(div50k_100[5]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[6]) );
  SDFFRQX1 div50k_100_reg_5_ ( .D(N58), .SIN(div50k_100[4]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[5]) );
  SDFFRQX1 div50k_100_reg_4_ ( .D(N57), .SIN(div50k_100[3]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[4]) );
  SDFFRQX1 div50k_100_reg_3_ ( .D(N56), .SIN(div50k_100[2]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[3]) );
  SDFFRQX1 div500k_5_reg_1_ ( .D(N38), .SIN(div500k_5_0), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(divff_o2) );
  SDFFRQX1 div500k_5_reg_0_ ( .D(N37), .SIN(div100k_2), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(div500k_5_0) );
  SDFFRQX1 div12_reg_0_ ( .D(N23), .SIN(div1p0m_2), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(div12[0]) );
  SDFFRQX1 div50k_100_reg_1_ ( .D(N54), .SIN(div50k_100[0]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[1]) );
  SDFFRQX1 div50k_100_reg_2_ ( .D(N55), .SIN(div50k_100[1]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[2]) );
  SDFFRQX1 div500k_5_reg_2_ ( .D(N39), .SIN(divff_o2), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(test_so) );
  SDFFRQX1 div50k_100_reg_0_ ( .D(N53), .SIN(divff_o1), .SMC(test_se), .C(
        clk_50k), .XR(n1), .Q(div50k_100[0]) );
  SDFFRQX1 div12_reg_1_ ( .D(N24), .SIN(div12[0]), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(div12[1]) );
  SDFFRQX1 div12_reg_2_ ( .D(N25), .SIN(div12[1]), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(div12[2]) );
  SDFFRQX1 div12_reg_3_ ( .D(N26), .SIN(div12[2]), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(divff_o1) );
  XNOR2XL U6 ( .A(n19), .B(n18), .Y(n16) );
  XNOR2XL U7 ( .A(n14), .B(n16), .Y(N25) );
  INVX1 U8 ( .A(n26), .Y(n9) );
  NOR2X1 U9 ( .A(n25), .B(n26), .Y(n18) );
  NOR2X1 U10 ( .A(n15), .B(n20), .Y(N24) );
  XOR2X1 U11 ( .A(n16), .B(n21), .Y(n20) );
  XNOR2XL U12 ( .A(n9), .B(n25), .Y(n21) );
  NOR21XL U13 ( .B(n14), .A(n15), .Y(N26) );
  NOR21XL U14 ( .B(N48), .A(n24), .Y(N55) );
  NOR21XL U15 ( .B(N49), .A(n24), .Y(N56) );
  NOR21XL U16 ( .B(N47), .A(n24), .Y(N54) );
  NOR21XL U17 ( .B(N50), .A(n24), .Y(N57) );
  NOR21XL U18 ( .B(N51), .A(n24), .Y(N58) );
  NOR2X1 U19 ( .A(n11), .B(n10), .Y(n15) );
  NOR2X1 U20 ( .A(N23), .B(n11), .Y(n22) );
  XNOR2XL U21 ( .A(n19), .B(div12[1]), .Y(n26) );
  XNOR2XL U22 ( .A(n10), .B(div12[2]), .Y(n19) );
  XNOR2XL U23 ( .A(n9), .B(div12[0]), .Y(n25) );
  XNOR2XL U24 ( .A(n17), .B(divff_o1), .Y(n14) );
  NAND2X1 U25 ( .A(n18), .B(n19), .Y(n17) );
  INVX1 U26 ( .A(divff_o1), .Y(n10) );
  AND4X1 U27 ( .A(div50k_100[5]), .B(div50k_100[1]), .C(div50k_100[6]), .D(n12), .Y(n24) );
  NOR41XL U28 ( .D(div50k_100[0]), .A(div50k_100[4]), .B(div50k_100[3]), .C(
        div50k_100[2]), .Y(n12) );
  NOR21XL U29 ( .B(N46), .A(n24), .Y(N53) );
  NOR21XL U30 ( .B(N52), .A(n24), .Y(N59) );
  OAI32X1 U31 ( .A(n7), .B(test_so), .C(n8), .D(n13), .E(n6), .Y(N39) );
  INVX1 U32 ( .A(div500k_5_0), .Y(n8) );
  AOI21BBXL U33 ( .B(n23), .C(divff_o2), .A(N37), .Y(n13) );
  NOR3XL U34 ( .A(div500k_5_0), .B(divff_o2), .C(n6), .Y(n23) );
  NOR2X1 U35 ( .A(n23), .B(div500k_5_0), .Y(N37) );
  INVX1 U36 ( .A(test_so), .Y(n6) );
  NAND31X1 U37 ( .C(div12[0]), .A(div12[1]), .B(div12[2]), .Y(n11) );
  XOR2X1 U38 ( .A(n27), .B(div12[1]), .Y(N23) );
  XNOR2XL U39 ( .A(divff_o1), .B(div12[2]), .Y(n27) );
  XNOR2XL U40 ( .A(n7), .B(div500k_5_0), .Y(N38) );
  INVX1 U41 ( .A(divff_o2), .Y(n7) );
  INVX1 U42 ( .A(div100k_2), .Y(n5) );
  INVX1 U43 ( .A(div1p0m_2), .Y(n4) );
endmodule


module divclk_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module srambist_a0 ( clk, srstz, reg_hit, reg_w, reg_r, reg_wdat, iram_rdat, 
        xram_rdat, bist_en, bist_xram, bist_wr, bist_adr, bist_wdat, o_bistctl, 
        o_bistdat, test_si, test_se );
  input [1:0] reg_hit;
  input [7:0] reg_wdat;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  output [10:0] bist_adr;
  output [7:0] bist_wdat;
  output [6:0] o_bistctl;
  output [7:0] o_bistdat;
  input clk, srstz, reg_w, reg_r, test_si, test_se;
  output bist_en, bist_xram, bist_wr;
  wire   we_1_, bistctl_re, N21, busy_dly, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, r_bistfault, upd_fault, wd_fault, net8942, n110, n111, n10,
         n11, n12, n13, n25, n26, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n4, n6, n7, n8, n9, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n27, n28, n29, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140;
  wire   [1:0] rw_sta;

  INVX1 U11 ( .A(n13), .Y(n11) );
  INVX1 U12 ( .A(n13), .Y(n12) );
  INVX1 U13 ( .A(n13), .Y(n10) );
  INVX1 U14 ( .A(srstz), .Y(n13) );
  INVX8 U148 ( .A(n11), .Y(n25) );
  glreg_WIDTH1_0 u0_bistfault ( .clk(clk), .arstz(n11), .we(upd_fault), .wdat(
        wd_fault), .rdat(o_bistctl[3]), .test_si(o_bistdat[7]), .test_se(
        test_se) );
  glreg_WIDTH5_1 u0_bistctl ( .clk(clk), .arstz(n11), .we(n26), .wdat({
        reg_wdat[6:4], reg_wdat[2], n7}), .rdat({o_bistctl[6:4], 
        o_bistctl[2:1]}), .test_si(rw_sta[1]), .test_se(test_se) );
  glreg_a0_6 u0_bistdat ( .clk(clk), .arstz(n10), .we(we_1_), .wdat({
        reg_wdat[7:2], n7, reg_wdat[0]}), .rdat(o_bistdat), .test_si(
        o_bistctl[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_srambist_a0 clk_gate_adr_reg ( .CLK(clk), .EN(N86), 
        .ENCLK(net8942), .TE(test_se) );
  srambist_a0_DW01_inc_0 add_65 ( .A(bist_adr), .SUM({N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64}) );
  SDFFQX1 busy_dly_reg ( .D(o_bistctl[0]), .SIN(bistctl_re), .SMC(test_se), 
        .C(clk), .Q(busy_dly) );
  SDFFQX1 r_bistfault_reg ( .D(n110), .SIN(busy_dly), .SMC(test_se), .C(clk), 
        .Q(r_bistfault) );
  SDFFRQX1 bistctl_re_reg ( .D(N21), .SIN(bist_adr[10]), .SMC(test_se), .C(clk), .XR(n11), .Q(bistctl_re) );
  SDFFQX1 rw_sta_reg_1_ ( .D(n137), .SIN(rw_sta[0]), .SMC(test_se), .C(clk), 
        .Q(rw_sta[1]) );
  SDFFQX1 rw_sta_reg_0_ ( .D(n111), .SIN(r_bistfault), .SMC(test_se), .C(clk), 
        .Q(rw_sta[0]) );
  SDFFQX1 adr_reg_9_ ( .D(N96), .SIN(bist_adr[8]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[9]) );
  SDFFQX1 adr_reg_10_ ( .D(N97), .SIN(bist_adr[9]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[10]) );
  SDFFQX1 adr_reg_6_ ( .D(N93), .SIN(bist_adr[5]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[6]) );
  SDFFQX1 adr_reg_7_ ( .D(N94), .SIN(bist_adr[6]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[7]) );
  SDFFQX1 adr_reg_8_ ( .D(N95), .SIN(bist_adr[7]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[8]) );
  SDFFQX1 adr_reg_2_ ( .D(N89), .SIN(bist_adr[1]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[2]) );
  SDFFQX1 adr_reg_5_ ( .D(N92), .SIN(bist_adr[4]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[5]) );
  SDFFQX1 adr_reg_4_ ( .D(N91), .SIN(bist_adr[3]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[4]) );
  SDFFQX1 adr_reg_3_ ( .D(N90), .SIN(bist_adr[2]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[3]) );
  SDFFQX1 adr_reg_1_ ( .D(N88), .SIN(bist_adr[0]), .SMC(test_se), .C(net8942), 
        .Q(bist_adr[1]) );
  SDFFQX1 adr_reg_0_ ( .D(N87), .SIN(test_si), .SMC(test_se), .C(net8942), .Q(
        bist_adr[0]) );
  INVX1 U3 ( .A(1'b1), .Y(bist_xram) );
  INVX1 U5 ( .A(n138), .Y(bist_en) );
  INVX1 U6 ( .A(n19), .Y(n26) );
  INVX1 U7 ( .A(n82), .Y(n121) );
  INVX1 U8 ( .A(n83), .Y(n117) );
  NAND2X1 U9 ( .A(reg_hit[0]), .B(reg_w), .Y(n19) );
  INVX1 U10 ( .A(n105), .Y(n84) );
  AND2X1 U15 ( .A(reg_w), .B(reg_hit[1]), .Y(we_1_) );
  INVX1 U16 ( .A(n8), .Y(n7) );
  INVX1 U17 ( .A(n50), .Y(n130) );
  NAND21X1 U18 ( .B(n24), .A(n23), .Y(n83) );
  NAND2X1 U19 ( .A(n24), .B(n23), .Y(n82) );
  INVX1 U20 ( .A(n21), .Y(n23) );
  NAND21X1 U21 ( .B(n24), .A(n20), .Y(n105) );
  AND2X1 U22 ( .A(reg_r), .B(reg_hit[0]), .Y(N21) );
  INVX1 U23 ( .A(n119), .Y(n123) );
  INVX1 U24 ( .A(n104), .Y(n113) );
  INVX1 U25 ( .A(n100), .Y(n103) );
  INVX1 U26 ( .A(n97), .Y(n99) );
  INVX1 U27 ( .A(n94), .Y(n96) );
  INVX1 U28 ( .A(n91), .Y(n93) );
  INVX1 U29 ( .A(n88), .Y(n90) );
  INVX1 U30 ( .A(n85), .Y(n87) );
  INVX1 U31 ( .A(reg_wdat[1]), .Y(n8) );
  OAI21X1 U32 ( .B(n134), .C(n129), .A(n73), .Y(bist_wdat[0]) );
  NAND2X1 U33 ( .A(n134), .B(n129), .Y(n73) );
  INVX1 U34 ( .A(n78), .Y(n129) );
  XNOR2XL U35 ( .A(n134), .B(n80), .Y(bist_wdat[1]) );
  AOI21X1 U36 ( .B(n76), .C(n75), .A(n78), .Y(n80) );
  NAND2X1 U37 ( .A(n75), .B(n127), .Y(n76) );
  INVX1 U38 ( .A(n74), .Y(n127) );
  XNOR2XL U39 ( .A(n134), .B(n79), .Y(bist_wdat[2]) );
  AOI21X1 U40 ( .B(n76), .C(n127), .A(n78), .Y(n79) );
  XNOR2XL U41 ( .A(iram_rdat[2]), .B(n52), .Y(n45) );
  AOI21X1 U42 ( .B(n50), .C(n131), .A(n51), .Y(n52) );
  AOI31X1 U43 ( .A(iram_rdat[7]), .B(n43), .C(n44), .D(n135), .Y(n39) );
  AOI21X1 U44 ( .B(n130), .C(n140), .A(n45), .Y(n44) );
  INVX1 U45 ( .A(o_bistctl[0]), .Y(n138) );
  XOR2X1 U46 ( .A(iram_rdat[1]), .B(n49), .Y(n43) );
  AOI21X1 U47 ( .B(n50), .C(n42), .A(n51), .Y(n49) );
  XOR2X1 U48 ( .A(bist_wdat[3]), .B(iram_rdat[3]), .Y(n68) );
  XNOR2XL U49 ( .A(n134), .B(iram_rdat[7]), .Y(n70) );
  OAI22AX1 U50 ( .D(n76), .C(n73), .A(n134), .B(n76), .Y(bist_wdat[4]) );
  XNOR2XL U51 ( .A(iram_rdat[6]), .B(n61), .Y(n53) );
  OAI22X1 U52 ( .A(n133), .B(n131), .C(n62), .D(n135), .Y(n61) );
  XNOR2XL U53 ( .A(iram_rdat[0]), .B(n60), .Y(n54) );
  NAND2X1 U54 ( .A(n133), .B(n58), .Y(n60) );
  OAI22X1 U55 ( .A(n73), .B(n76), .C(n77), .D(n134), .Y(bist_wdat[3]) );
  NOR2X1 U56 ( .A(n78), .B(n76), .Y(n77) );
  INVX1 U57 ( .A(iram_rdat[4]), .Y(n140) );
  INVX1 U58 ( .A(iram_rdat[5]), .Y(n139) );
  NOR4XL U59 ( .A(n65), .B(n66), .C(n67), .D(n68), .Y(n64) );
  XOR2X1 U60 ( .A(bist_wdat[0]), .B(iram_rdat[0]), .Y(n66) );
  XNOR2XL U61 ( .A(bist_wdat[5]), .B(n139), .Y(n65) );
  XOR2X1 U62 ( .A(bist_wdat[6]), .B(iram_rdat[6]), .Y(n67) );
  NOR4XL U63 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(n63) );
  XNOR2XL U64 ( .A(n140), .B(bist_wdat[4]), .Y(n69) );
  XOR2X1 U65 ( .A(bist_wdat[1]), .B(iram_rdat[1]), .Y(n71) );
  XOR2X1 U66 ( .A(bist_wdat[2]), .B(iram_rdat[2]), .Y(n72) );
  OAI22X1 U67 ( .A(n73), .B(n127), .C(n74), .D(n134), .Y(bist_wdat[6]) );
  NAND2X1 U68 ( .A(n42), .B(n131), .Y(n50) );
  INVX1 U69 ( .A(n62), .Y(n131) );
  INVX1 U70 ( .A(n59), .Y(n133) );
  INVX1 U71 ( .A(n30), .Y(n17) );
  NAND32X1 U72 ( .B(n20), .C(n17), .A(n16), .Y(n21) );
  MUX2IX1 U73 ( .D0(rw_sta[1]), .D1(rw_sta[0]), .S(o_bistctl[2]), .Y(n16) );
  AO21X1 U74 ( .B(n117), .C(n109), .A(n108), .Y(N87) );
  AO21X1 U75 ( .B(N64), .C(n121), .A(n112), .Y(n108) );
  AO21X1 U76 ( .B(N69), .C(n121), .A(n95), .Y(N92) );
  GEN2XL U77 ( .D(bist_adr[5]), .E(n94), .C(n93), .B(n117), .A(n112), .Y(n95)
         );
  AO21X1 U78 ( .B(N65), .C(n121), .A(n114), .Y(N88) );
  GEN2XL U79 ( .D(bist_adr[0]), .E(bist_adr[1]), .C(n113), .B(n117), .A(n112), 
        .Y(n114) );
  AO21X1 U80 ( .B(N67), .C(n121), .A(n101), .Y(N90) );
  GEN2XL U81 ( .D(bist_adr[3]), .E(n100), .C(n99), .B(n117), .A(n112), .Y(n101) );
  AO21X1 U82 ( .B(N71), .C(n121), .A(n89), .Y(N94) );
  GEN2XL U83 ( .D(bist_adr[7]), .E(n88), .C(n87), .B(n117), .A(n112), .Y(n89)
         );
  AO21X1 U84 ( .B(N70), .C(n121), .A(n92), .Y(N93) );
  GEN2XL U85 ( .D(bist_adr[6]), .E(n91), .C(n90), .B(n117), .A(n112), .Y(n92)
         );
  AO21X1 U86 ( .B(N72), .C(n121), .A(n86), .Y(N95) );
  GEN2XL U87 ( .D(bist_adr[8]), .E(n85), .C(n123), .B(n117), .A(n112), .Y(n86)
         );
  AO21X1 U88 ( .B(N68), .C(n121), .A(n98), .Y(N91) );
  GEN2XL U89 ( .D(bist_adr[4]), .E(n97), .C(n96), .B(n117), .A(n112), .Y(n98)
         );
  AO21X1 U90 ( .B(N73), .C(n121), .A(n120), .Y(N96) );
  GEN2XL U91 ( .D(bist_adr[9]), .E(n119), .C(n118), .B(n117), .A(n116), .Y(
        n120) );
  INVX1 U92 ( .A(n115), .Y(n118) );
  INVX1 U93 ( .A(n15), .Y(n20) );
  NAND43X1 U94 ( .B(o_bistdat[6]), .C(n19), .D(n6), .A(o_bistdat[7]), .Y(n15)
         );
  INVX1 U95 ( .A(reg_wdat[0]), .Y(n6) );
  MUX2AXL U96 ( .D0(o_bistctl[1]), .D1(n8), .S(n26), .Y(n24) );
  NAND21X1 U97 ( .B(n84), .A(n12), .Y(n112) );
  NAND21X1 U98 ( .B(n82), .A(N74), .Y(n22) );
  NAND32X1 U99 ( .B(n107), .C(n106), .A(n105), .Y(N89) );
  AND2X1 U100 ( .A(N66), .B(n121), .Y(n107) );
  GEN2XL U101 ( .D(bist_adr[2]), .E(n104), .C(n103), .B(n117), .A(n102), .Y(
        n106) );
  NAND32X1 U102 ( .B(n81), .C(n29), .A(n28), .Y(N97) );
  NAND21X1 U103 ( .B(n83), .A(n27), .Y(n28) );
  NAND21X1 U104 ( .B(n84), .A(n22), .Y(n81) );
  XNOR2XL U105 ( .A(n115), .B(bist_adr[10]), .Y(n27) );
  NAND32X1 U106 ( .B(n20), .C(n18), .A(n21), .Y(N86) );
  NAND6XL U107 ( .A(bist_adr[4]), .B(bist_adr[8]), .C(bist_adr[6]), .D(
        bist_adr[3]), .E(bist_adr[7]), .F(n122), .Y(n124) );
  AND4X1 U108 ( .A(bist_adr[1]), .B(bist_adr[2]), .C(bist_adr[0]), .D(
        bist_adr[5]), .Y(n122) );
  NAND21X1 U109 ( .B(bist_adr[8]), .A(n87), .Y(n119) );
  NAND21X1 U110 ( .B(bist_adr[3]), .A(n103), .Y(n97) );
  NAND21X1 U111 ( .B(bist_adr[4]), .A(n99), .Y(n94) );
  NAND21X1 U112 ( .B(bist_adr[1]), .A(n109), .Y(n104) );
  NAND21X1 U113 ( .B(bist_adr[2]), .A(n113), .Y(n100) );
  NAND21X1 U114 ( .B(bist_adr[5]), .A(n96), .Y(n91) );
  NAND21X1 U115 ( .B(bist_adr[6]), .A(n93), .Y(n88) );
  NAND21X1 U116 ( .B(bist_adr[7]), .A(n90), .Y(n85) );
  INVX1 U117 ( .A(bist_adr[0]), .Y(n109) );
  NOR2X1 U118 ( .A(o_bistdat[2]), .B(o_bistdat[3]), .Y(n78) );
  INVX1 U119 ( .A(o_bistdat[5]), .Y(n134) );
  NOR2X1 U120 ( .A(n128), .B(o_bistdat[3]), .Y(n74) );
  INVX1 U121 ( .A(o_bistdat[2]), .Y(n128) );
  NAND2X1 U122 ( .A(o_bistdat[3]), .B(n128), .Y(n75) );
  OAI22X1 U123 ( .A(o_bistdat[4]), .B(n46), .C(n130), .D(n47), .Y(n38) );
  XNOR2XL U124 ( .A(n133), .B(n140), .Y(n47) );
  NOR32XL U125 ( .B(n48), .C(n45), .A(n43), .Y(n46) );
  AOI21X1 U126 ( .B(iram_rdat[4]), .C(n130), .A(iram_rdat[7]), .Y(n48) );
  NOR42XL U127 ( .C(n125), .D(n12), .A(n126), .B(n36), .Y(n35) );
  NOR4XL U128 ( .A(n37), .B(n38), .C(n39), .D(n40), .Y(n36) );
  NAND3X1 U129 ( .A(n53), .B(n54), .C(n55), .Y(n37) );
  XNOR2XL U130 ( .A(n41), .B(n139), .Y(n40) );
  ENOX1 U131 ( .A(bistctl_re), .B(n33), .C(wd_fault), .D(srstz), .Y(n110) );
  AOI31X1 U132 ( .A(busy_dly), .B(n17), .C(n34), .D(n35), .Y(n33) );
  AOI211X1 U133 ( .C(n63), .D(n64), .A(n136), .B(n25), .Y(n34) );
  NOR3XL U134 ( .A(n138), .B(rw_sta[1]), .C(n126), .Y(bist_wr) );
  XNOR2XL U135 ( .A(iram_rdat[3]), .B(n56), .Y(n55) );
  NAND2X1 U136 ( .A(n57), .B(n58), .Y(n56) );
  OAI22X1 U137 ( .A(o_bistdat[4]), .B(n130), .C(n59), .D(n50), .Y(n57) );
  ENOX1 U138 ( .A(n73), .B(n75), .C(n75), .D(o_bistdat[5]), .Y(bist_wdat[5])
         );
  NOR2X1 U139 ( .A(n132), .B(o_bistdat[1]), .Y(n62) );
  INVX1 U140 ( .A(o_bistdat[0]), .Y(n132) );
  NAND2X1 U141 ( .A(o_bistdat[1]), .B(n132), .Y(n42) );
  MUX2BXL U142 ( .D0(rw_sta[0]), .D1(n4), .S(n31), .Y(n111) );
  NAND2X1 U143 ( .A(n17), .B(n14), .Y(n4) );
  NOR2X1 U144 ( .A(n51), .B(o_bistdat[4]), .Y(n59) );
  OAI21X1 U145 ( .B(n138), .C(n32), .A(n12), .Y(n31) );
  NOR2X1 U146 ( .A(n126), .B(n125), .Y(n32) );
  NOR2X1 U147 ( .A(o_bistdat[0]), .B(o_bistdat[1]), .Y(n51) );
  OAI32X1 U149 ( .A(n136), .B(n18), .C(n9), .D(n31), .E(n125), .Y(n137) );
  INVX1 U150 ( .A(bist_wr), .Y(n9) );
  ENOX1 U151 ( .A(n133), .B(n42), .C(n42), .D(o_bistdat[4]), .Y(n41) );
  NAND2X1 U153 ( .A(n51), .B(o_bistdat[4]), .Y(n58) );
  INVX1 U154 ( .A(rw_sta[0]), .Y(n126) );
  NAND21X1 U155 ( .B(bist_adr[9]), .A(n123), .Y(n115) );
  INVX1 U156 ( .A(o_bistdat[4]), .Y(n135) );
  NAND21X1 U157 ( .B(rw_sta[0]), .A(n125), .Y(n30) );
  INVX1 U158 ( .A(rw_sta[1]), .Y(n125) );
  OR2X1 U159 ( .A(bistctl_re), .B(r_bistfault), .Y(upd_fault) );
  INVX1 U160 ( .A(o_bistctl[2]), .Y(n136) );
  NOR21XL U161 ( .B(r_bistfault), .A(bistctl_re), .Y(wd_fault) );
  OAI2B11X1 U162 ( .D(n124), .C(n123), .A(bist_adr[10]), .B(bist_adr[9]), .Y(
        o_bistctl[0]) );
  BUFX3 U163 ( .A(o_bistdat[5]), .Y(bist_wdat[7]) );
  INVX8 U164 ( .A(n11), .Y(n18) );
  INVX8 U165 ( .A(n25), .Y(n14) );
  INVX8 U166 ( .A(n10), .Y(n29) );
  INVX8 U167 ( .A(srstz), .Y(n102) );
  INVX8 U168 ( .A(n10), .Y(n116) );
endmodule


module srambist_a0_DW01_inc_0 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_srambist_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_6 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8960;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8960), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8960), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8960), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8960), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8960), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8960), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8960), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8960), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8960), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8978;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8978), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8978), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8978), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8978), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8978), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8978), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module regx_a0 ( regx_r, regx_w, di_drposc, di_imposc, di_rd_det, clk_500k, 
        r_imp_osc, regx_addr, regx_wdat, regx_rdat, regx_hitbst, regx_wrpwm, 
        regx_wrcvc, r_sdischg, r_bistctl, r_bistdat, r_vcomp, r_idacsh, 
        r_cvofsx, r_pwm, regx_wrdac, dac_r_vs, dac_comp, r_dac_en, r_sar_en, 
        r_aopt, r_xtm, r_adummyi, r_bck0, r_bck1, r_bck2, r_i2crout, r_xana, 
        di_xana, lt_gpi, di_tst, bkpt_pc, bkpt_ena, we_twlb, r_vpp_en, 
        r_vpp0v_en, r_otp_pwdn_en, r_otp_wpls, wd_twlb, r_sap, r_twlb, 
        upd_pwrv, ramacc, sse_idle, bus_idle, r_do_ts, r_dpdo_sel, r_dndo_sel, 
        di_ts, detclk, aswclk, atpg_en, di_aswk, clk, rrstz, test_si2, 
        test_si1, test_so1, test_se );
  input [6:0] regx_addr;
  input [7:0] regx_wdat;
  output [7:0] regx_rdat;
  output [1:0] regx_hitbst;
  output [1:0] regx_wrpwm;
  output [3:0] regx_wrcvc;
  input [7:0] r_sdischg;
  input [6:0] r_bistctl;
  input [7:0] r_bistdat;
  input [7:0] r_vcomp;
  input [7:0] r_idacsh;
  input [7:0] r_cvofsx;
  input [15:0] r_pwm;
  output [13:0] regx_wrdac;
  input [79:0] dac_r_vs;
  input [9:0] dac_comp;
  input [9:0] r_dac_en;
  input [9:0] r_sar_en;
  output [7:0] r_aopt;
  output [7:0] r_xtm;
  output [7:0] r_adummyi;
  output [7:0] r_bck0;
  output [7:0] r_bck1;
  output [7:0] r_bck2;
  output [5:0] r_i2crout;
  output [23:0] r_xana;
  input [4:0] di_xana;
  input [3:0] lt_gpi;
  output [14:0] bkpt_pc;
  output [1:0] wd_twlb;
  output [1:0] r_sap;
  input [1:0] r_twlb;
  output [6:0] r_do_ts;
  output [3:0] r_dpdo_sel;
  output [3:0] r_dndo_sel;
  input [4:0] di_aswk;
  input regx_r, regx_w, di_drposc, di_imposc, di_rd_det, clk_500k, di_tst,
         upd_pwrv, ramacc, sse_idle, bus_idle, di_ts, detclk, aswclk, atpg_en,
         clk, rrstz, test_si2, test_si1, test_se;
  output r_imp_osc, bkpt_ena, we_twlb, r_vpp_en, r_vpp0v_en, r_otp_pwdn_en,
         r_otp_wpls, test_so1;
  wire   we_19, we_7, we_6, we_5, we_4, reg1B_3_, reg10_7_, lt_drp,
         i2c_mode_upd, N8, d_we16, lt_reg1C_0, net8996, n132, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n60, n71, n72, n73, n74, n75, n1, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n23, n24, n25, n28, n29, n31, n32, n33, n59, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462,
         SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464,
         SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466,
         SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468,
         SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470,
         SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472,
         SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474,
         SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476,
         SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478,
         SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480,
         SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482,
         SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484,
         SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486,
         SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488,
         SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490,
         SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492,
         SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494,
         SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496,
         SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498,
         SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500,
         SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502,
         SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504,
         SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506,
         SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508,
         SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510,
         SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512,
         SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514,
         SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516,
         SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518,
         SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520,
         SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522,
         SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524,
         SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526,
         SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528,
         SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530,
         SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532,
         SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534,
         SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536,
         SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538,
         SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540,
         SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542,
         SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544,
         SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546,
         SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548,
         SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550,
         SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552,
         SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554,
         SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556,
         SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558,
         SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560,
         SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562,
         SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564,
         SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566,
         SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568,
         SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570,
         SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572,
         SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574,
         SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576,
         SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578,
         SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580,
         SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582,
         SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584,
         SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586,
         SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588,
         SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590,
         SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592,
         SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594,
         SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596,
         SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598,
         SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600,
         SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602,
         SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604,
         SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606,
         SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608,
         SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610,
         SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612,
         SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614,
         SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616,
         SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618,
         SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620,
         SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622,
         SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624,
         SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626,
         SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628,
         SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630,
         SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632,
         SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634,
         SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636,
         SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638,
         SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640,
         SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642,
         SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644,
         SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646,
         SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648,
         SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650,
         SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652,
         SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654,
         SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656,
         SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658,
         SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660,
         SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662,
         SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664,
         SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666,
         SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668,
         SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670,
         SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672,
         SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674,
         SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676,
         SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678,
         SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680,
         SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682,
         SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684,
         SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686,
         SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688,
         SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690,
         SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692,
         SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694,
         SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696,
         SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698,
         SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700,
         SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702,
         SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704,
         SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706,
         SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708,
         SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710,
         SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712,
         SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714,
         SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716,
         SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718,
         SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720,
         SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722,
         SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724,
         SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726,
         SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728,
         SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730,
         SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732,
         SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734,
         SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736,
         SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738,
         SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740,
         SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742,
         SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744,
         SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746,
         SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748,
         SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750,
         SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752,
         SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754,
         SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756,
         SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758,
         SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760,
         SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762,
         SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764,
         SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766,
         SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768,
         SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770,
         SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772,
         SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774,
         SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776,
         SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778,
         SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780,
         SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782,
         SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784,
         SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786,
         SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788,
         SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790,
         SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792,
         SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794,
         SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796,
         SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798,
         SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800,
         SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802,
         SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804,
         SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806,
         SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808,
         SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810,
         SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812,
         SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814,
         SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816,
         SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818,
         SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820,
         SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822,
         SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824,
         SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826,
         SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828,
         SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830,
         SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832,
         SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834,
         SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836,
         SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838,
         SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840,
         SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842,
         SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844,
         SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846,
         SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848,
         SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850,
         SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852,
         SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854,
         SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856,
         SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858,
         SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860,
         SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862,
         SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864,
         SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866,
         SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868,
         SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870,
         SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872,
         SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874,
         SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876,
         SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878,
         SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880,
         SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882,
         SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884,
         SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886,
         SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888,
         SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890,
         SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892,
         SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894,
         SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896,
         SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898,
         SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900,
         SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902,
         SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904,
         SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906,
         SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908,
         SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910,
         SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912,
         SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914,
         SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916,
         SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918,
         SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920,
         SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922,
         SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924,
         SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926,
         SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928,
         SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930,
         SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932,
         SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934,
         SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936,
         SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938,
         SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940,
         SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942,
         SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944,
         SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946,
         SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948,
         SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950,
         SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952,
         SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954,
         SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956,
         SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958,
         SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960,
         SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962,
         SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964,
         SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966,
         SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968,
         SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970,
         SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972,
         SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974,
         SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976,
         SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978,
         SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980,
         SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982,
         SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984,
         SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986,
         SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988,
         SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990,
         SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992,
         SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994,
         SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996,
         SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998,
         SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000,
         SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002,
         SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004,
         SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006,
         SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008,
         SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010,
         SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012,
         SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014,
         SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016;
  wire   [30:23] we;
  wire   [6:0] d_regx_addr;
  wire   [7:0] reg1F;
  wire   [3:2] reg1E;
  wire   [3:0] reg14;
  wire   [3:0] d_lt_gpi;
  wire   [5:0] lt_reg15_5_0;
  wire   [5:0] i2c_mode_wdat;
  wire   [5:0] d_lt_aswk;
  wire   [5:0] lt_aswk;
  wire   [7:0] wd18;

  INVX1 U68 ( .A(n56), .Y(n53) );
  INVX1 U69 ( .A(n56), .Y(n55) );
  INVX1 U70 ( .A(n57), .Y(n54) );
  INVX1 U71 ( .A(n57), .Y(n44) );
  INVX1 U72 ( .A(n57), .Y(n45) );
  INVX1 U73 ( .A(n57), .Y(n46) );
  INVX1 U74 ( .A(n57), .Y(n43) );
  INVX1 U75 ( .A(n58), .Y(n42) );
  INVX1 U76 ( .A(n58), .Y(n41) );
  INVX1 U77 ( .A(n58), .Y(n40) );
  INVX1 U78 ( .A(n57), .Y(n39) );
  INVX1 U79 ( .A(n57), .Y(n38) );
  INVX1 U80 ( .A(n57), .Y(n37) );
  INVX1 U81 ( .A(n56), .Y(n36) );
  INVX1 U82 ( .A(n56), .Y(n35) );
  INVX1 U83 ( .A(n56), .Y(n34) );
  INVX1 U84 ( .A(n56), .Y(n47) );
  INVX1 U85 ( .A(n56), .Y(n48) );
  INVX1 U86 ( .A(n56), .Y(n52) );
  INVX1 U87 ( .A(n56), .Y(n51) );
  INVX1 U88 ( .A(n57), .Y(n49) );
  INVX1 U89 ( .A(n57), .Y(n50) );
  INVX1 U90 ( .A(rrstz), .Y(n58) );
  INVX1 U91 ( .A(rrstz), .Y(n56) );
  INVX1 U92 ( .A(rrstz), .Y(n57) );
  glreg_a0_19 u0_reg04 ( .clk(clk), .arstz(n34), .we(we_4), .wdat({n62, n16, 
        n13, n9, n7, n59, wd_twlb}), .rdat(r_bck0), .test_si(r_xana[23]), 
        .test_se(test_se) );
  glreg_a0_18 u0_reg05 ( .clk(clk), .arstz(n35), .we(we_5), .wdat({n62, n15, 
        n13, n10, n6, n59, wd_twlb}), .rdat(r_bck1), .test_si(r_bck0[7]), 
        .test_se(test_se) );
  glreg_a0_17 u0_reg06 ( .clk(clk), .arstz(n36), .we(we_6), .wdat({n62, n16, 
        n12, n9, n6, n59, wd_twlb}), .rdat(r_bck2), .test_si(r_bck1[7]), 
        .test_se(test_se) );
  glreg_a0_16 u0_reg07 ( .clk(clk), .arstz(n37), .we(we_7), .wdat({n62, n15, 
        n12, n9, n7, n59, wd_twlb}), .rdat(r_adummyi), .test_si2(test_si2), 
        .test_si1(r_bck2[7]), .test_se(test_se) );
  glreg_WIDTH1_2 u0_reg10 ( .clk(clk), .arstz(n42), .we(1'b1), .wdat(ramacc), 
        .rdat(reg10_7_), .test_si(r_adummyi[6]), .test_se(test_se) );
  glreg_6_00000002 u0_reg12 ( .clk(clk), .arstz(n48), .we(we_twlb), .wdat({n62, 
        n16, n12, n10, n6, n59}), .rdat({r_vpp_en, r_vpp0v_en, r_otp_pwdn_en, 
        r_otp_wpls, r_sap}), .test_si(reg10_7_), .test_se(test_se) );
  glreg_a0_15 u0_reg13 ( .clk(clk), .arstz(n38), .we(we_19), .wdat({n62, n16, 
        n13, n10, n7, n33, wd_twlb}), .rdat({r_dpdo_sel, r_dndo_sel}), 
        .test_si(r_vpp_en), .test_se(test_se) );
  glreg_WIDTH6_1 u0_reg15 ( .clk(clk), .arstz(n50), .we(n75), .wdat({n12, n9, 
        n6, n33, wd_twlb}), .rdat(lt_reg15_5_0), .test_si(r_dpdo_sel[3]), 
        .test_se(test_se) );
  glreg_WIDTH6_0 u1_reg15 ( .clk(clk), .arstz(n49), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat({n132, r_i2crout[4:0]}), .test_si(r_xana[0]), 
        .test_se(test_se) );
  glreg_a0_14 u0_reg17 ( .clk(clk), .arstz(n39), .we(we[23]), .wdat({n62, n16, 
        n13, n10, n7, n33, wd_twlb[1], n28}), .rdat(r_aopt), .test_si(
        lt_reg15_5_0[5]), .test_se(test_se) );
  glreg_a0_13 u0_tmp18 ( .clk(clk), .arstz(n40), .we(we[24]), .wdat({n62, n15, 
        n13, n9, n7, n33, wd_twlb[1], n28}), .rdat(wd18), .test_si(bkpt_ena), 
        .test_se(test_se) );
  glreg_a0_12 u0_reg18 ( .clk(clk), .arstz(n41), .we(n74), .wdat(wd18), .rdat(
        bkpt_pc[7:0]), .test_si(r_aopt[7]), .test_se(test_se) );
  glreg_a0_11 u0_reg19 ( .clk(clk), .arstz(n42), .we(n74), .wdat({n62, n16, 
        n13, n10, n7, n33, n31, n28}), .rdat({bkpt_ena, bkpt_pc[14:8]}), 
        .test_si(bkpt_pc[7]), .test_se(test_se) );
  glreg_a0_10 u0_reg1A ( .clk(clk), .arstz(n43), .we(we[26]), .wdat({n63, n16, 
        n12, n9, n6, n33, n31, n28}), .rdat(r_xtm), .test_si(n115), .test_se(
        test_se) );
  dbnc_WIDTH2_TIMEOUT2_7 u0_ts_db ( .o_dbc(reg1B_3_), .o_chg(), .i_org(di_ts), 
        .clk(clk), .rstz(n55), .test_si(wd18[7]), .test_so(n114), .test_se(
        test_se) );
  glreg_WIDTH7_0 u0_reg1B ( .clk(clk), .arstz(n47), .we(we[27]), .wdat({n63, 
        n16, n13, regx_wdat[4], n33, n31, n28}), .rdat(r_do_ts), .test_si(
        r_xtm[7]), .test_se(test_se) );
  glreg_WIDTH1_1 u1_reg1C ( .clk(clk), .arstz(n41), .we(upd_pwrv), .wdat(
        lt_reg1C_0), .rdat(r_xana[0]), .test_si(n113), .test_se(test_se) );
  glreg_a0_9 u0_reg1C ( .clk(clk), .arstz(n46), .we(we[28]), .wdat({n63, n15, 
        n12, n10, n6, n33, n31, n28}), .rdat({r_xana[7:1], lt_reg1C_0}), 
        .test_si(r_do_ts[6]), .test_se(test_se) );
  glreg_a0_8 u0_reg1D ( .clk(clk), .arstz(n45), .we(we[29]), .wdat({n63, n16, 
        n13, n10, n7, n33, n31, wd_twlb[0]}), .rdat(r_xana[15:8]), .test_si(
        r_xana[7]), .test_se(test_se) );
  glreg_a0_7 u0_reg1E ( .clk(clk), .arstz(n44), .we(we[30]), .wdat({n63, n16, 
        n12, n9, n7, n33, wd_twlb}), .rdat({r_xana[23], r_imp_osc, 
        r_xana[21:20], reg1E, r_xana[17:16]}), .test_si(r_xana[15]), .test_se(
        test_se) );
  dbnc_WIDTH2_TIMEOUT2_6 u0_dosc_db ( .o_dbc(reg14[1]), .o_chg(), .i_org(
        di_imposc), .clk(clk), .rstz(n54), .test_si(lt_drp), .test_so(n117), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_5 u0_iosc_db ( .o_dbc(reg14[2]), .o_chg(), .i_org(
        di_drposc), .clk(clk), .rstz(n51), .test_si(n117), .test_so(n116), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_4 u0_xana_db ( .o_dbc(reg1F[0]), .o_chg(), .i_org(
        di_xana[0]), .clk(clk), .rstz(n48), .test_si(n114), .test_so(n113), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_3 u1_xana_db ( .o_dbc(reg1F[1]), .o_chg(), .i_org(
        di_xana[1]), .clk(clk), .rstz(n55), .test_si(n132), .test_so(n112), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_2 u2_xana_db ( .o_dbc(reg1F[2]), .o_chg(), .i_org(
        di_xana[2]), .clk(clk), .rstz(n53), .test_si(n112), .test_so(n111), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_1 u3_xana_db ( .o_dbc(reg1F[3]), .o_chg(), .i_org(
        di_xana[3]), .clk(clk), .rstz(n54), .test_si(n111), .test_so(n110), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_0 u4_xana_db ( .o_dbc(reg1F[4]), .o_chg(), .i_org(
        di_xana[4]), .clk(clk), .rstz(n49), .test_si(n110), .test_so(n109), 
        .test_se(test_se) );
  dbnc_a0_2 u5_xana_db ( .o_dbc(reg1F[5]), .o_chg(), .i_org(di_xana[0]), .clk(
        clk_500k), .rstz(n51), .test_si(n109), .test_so(n108), .test_se(
        test_se) );
  dbnc_a0_1 u6_xana_db ( .o_dbc(reg1F[6]), .o_chg(), .i_org(di_xana[1]), .clk(
        clk_500k), .rstz(n52), .test_si(n108), .test_so(test_so1), .test_se(
        test_se) );
  dbnc_a0_0 u0_rdet_db ( .o_dbc(reg1F[7]), .o_chg(), .i_org(di_rd_det), .clk(
        clk_500k), .rstz(n53), .test_si(n116), .test_so(n115), .test_se(
        test_se) );
  SNPS_CLOCK_GATE_HIGH_regx_a0 clk_gate_d_lt_gpi_reg ( .CLK(clk), .EN(n58), 
        .ENCLK(net8996), .TE(test_se) );
  regx_a0_DW_rightsh_0 srl_66 ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        dac_comp[9:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_sar_en[9:8], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_dac_en[9:8], 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_comp[7:0], r_sar_en[7:0], r_dac_en[7:0], dac_r_vs[63:0], 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_r_vs[79:64], reg1F, r_xana[23], r_imp_osc, r_xana[21:20], reg1E, 
        r_xana[17:0], r_do_ts[6:3], reg1B_3_, r_do_ts[2:0], r_xtm, bkpt_ena, 
        bkpt_pc, r_aopt, 1'b0, 1'b0, d_lt_aswk, sse_idle, 1'b0, r_i2crout, 
        d_lt_gpi, reg14, r_dpdo_sel, r_dndo_sel, r_vpp_en, r_vpp0v_en, 
        r_otp_pwdn_en, r_otp_wpls, r_sap, r_twlb, r_bistdat, reg10_7_, 
        r_bistctl, r_sdischg, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_pwm, r_adummyi, 
        r_bck2, r_bck1, r_bck0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_cvofsx, r_idacsh, r_vcomp}), .DATA_TC(1'b0), .SH({d_regx_addr[6:4], 
        n20, n18, d_regx_addr[1:0], 1'b0, 1'b0, 1'b0}), .B({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, 
        SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, 
        SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, 
        SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, 
        SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, 
        SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, 
        SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, 
        SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, 
        SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, 
        SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, 
        SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, 
        SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, 
        SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, 
        SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, 
        SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, 
        SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, 
        SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, 
        SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, 
        SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, 
        SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, 
        SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, 
        SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, 
        SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, 
        SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, 
        SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, 
        SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, 
        SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, 
        SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, 
        SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, 
        SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, 
        SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, 
        SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, 
        SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, 
        SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, 
        SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, 
        SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, 
        SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, 
        SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, 
        SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, 
        SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, 
        SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, 
        SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, 
        SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, 
        SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, 
        SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, 
        SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, 
        SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, 
        SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, 
        SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, 
        SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, 
        SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, 
        SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, 
        SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, 
        SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, 
        SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, 
        SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, 
        SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, 
        SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, 
        SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, 
        SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, 
        SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, 
        SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, 
        SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, 
        SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, 
        SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, 
        SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, 
        SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, 
        SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, 
        SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, 
        SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, 
        SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, 
        SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, 
        SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, 
        SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, 
        SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, 
        SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, 
        SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, 
        SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, 
        SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, 
        SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, 
        SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, 
        SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, 
        SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, 
        SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, 
        SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, 
        SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, 
        SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, 
        SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, 
        SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, 
        SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, 
        SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, 
        SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, 
        SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, 
        SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, 
        SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, 
        SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, 
        SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, 
        SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, 
        SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, 
        SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, 
        SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, 
        SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, 
        SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, 
        SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, 
        SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, 
        SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, 
        SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, 
        SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, 
        SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, 
        SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, 
        SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, 
        SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, 
        SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, 
        SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, 
        SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, 
        SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, 
        SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, 
        SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, 
        SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, 
        SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, 
        SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, 
        SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, 
        SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, 
        SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, 
        SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, 
        SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, 
        SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, 
        SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, 
        SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, 
        SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, 
        SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, 
        SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, 
        SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, 
        SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, 
        SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, 
        SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, 
        SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, 
        SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, 
        SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, 
        SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, 
        SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, 
        SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, 
        SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, 
        SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, 
        SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, 
        SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, 
        SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, 
        SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, 
        SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, 
        SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, 
        SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, 
        SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, 
        SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, 
        SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, 
        SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, 
        SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, 
        SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, 
        SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, 
        SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, 
        SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, 
        SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, 
        SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, 
        SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, 
        SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, 
        SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, 
        SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, 
        SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, 
        SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, 
        SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, 
        SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, 
        SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, 
        SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, 
        SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, 
        SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, 
        SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, 
        SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, 
        SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, 
        SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, 
        SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, 
        SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, 
        SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, 
        SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, 
        SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, 
        SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, 
        SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, 
        SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, 
        SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, 
        SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, 
        SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, 
        SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, 
        SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, 
        SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, 
        SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, 
        SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, 
        SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, 
        SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, 
        SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, 
        SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, 
        SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, 
        SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, 
        SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, 
        SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, 
        SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, 
        SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, 
        SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, 
        SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, 
        SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, 
        SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, 
        SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, 
        SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, 
        SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, 
        SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, 
        SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, 
        SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, 
        SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, 
        SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, 
        SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, 
        SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, 
        SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, 
        SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, 
        SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, 
        SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, 
        SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, 
        SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, 
        SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, 
        SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, 
        SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, 
        SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, 
        SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, 
        SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, 
        SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, 
        SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, 
        SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, 
        SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, 
        SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, 
        SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, 
        SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, 
        SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, 
        SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, 
        SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, 
        SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, 
        SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, 
        SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, 
        SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, 
        SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, 
        SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, 
        SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, 
        SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, 
        SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, 
        SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, 
        SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, 
        SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, 
        SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, 
        SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, 
        SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, 
        SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, 
        SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, 
        SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, 
        SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, 
        SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, 
        SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, 
        SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, 
        SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, 
        SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, 
        SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, 
        SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, 
        SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, 
        SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, 
        SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, 
        SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, 
        SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, 
        SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, 
        SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, 
        SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, 
        SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, 
        SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, 
        SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, 
        SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, 
        SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, 
        SYNOPSYS_UNCONNECTED_1016, regx_rdat}) );
  SDFFQX1 d_we16_reg ( .D(N8), .SIN(d_regx_addr[6]), .SMC(test_se), .C(clk), 
        .Q(d_we16) );
  SDFFQX1 d_lt_gpi_reg_2_ ( .D(lt_gpi[2]), .SIN(d_lt_gpi[1]), .SMC(test_se), 
        .C(net8996), .Q(d_lt_gpi[2]) );
  SDFFQX1 d_lt_drp_reg ( .D(lt_drp), .SIN(d_lt_aswk[5]), .SMC(test_se), .C(clk), .Q(reg14[0]) );
  SDFFQX1 d_di_tst_reg ( .D(di_tst), .SIN(test_si1), .SMC(test_se), .C(clk), 
        .Q(reg14[3]) );
  SDFFQX1 d_lt_gpi_reg_1_ ( .D(lt_gpi[1]), .SIN(d_lt_gpi[0]), .SMC(test_se), 
        .C(net8996), .Q(d_lt_gpi[1]) );
  SDFFQX1 d_lt_gpi_reg_0_ ( .D(lt_gpi[0]), .SIN(reg14[0]), .SMC(test_se), .C(
        net8996), .Q(d_lt_gpi[0]) );
  SDFFQX1 d_lt_aswk_reg_5_ ( .D(lt_aswk[5]), .SIN(d_lt_aswk[4]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[5]) );
  SDFFQX1 d_lt_aswk_reg_4_ ( .D(lt_aswk[4]), .SIN(d_lt_aswk[3]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[4]) );
  SDFFQX1 d_lt_aswk_reg_3_ ( .D(lt_aswk[3]), .SIN(d_lt_aswk[2]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[3]) );
  SDFFQX1 d_lt_aswk_reg_2_ ( .D(lt_aswk[2]), .SIN(d_lt_aswk[1]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[2]) );
  SDFFQX1 d_lt_aswk_reg_1_ ( .D(lt_aswk[1]), .SIN(d_lt_aswk[0]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[1]) );
  SDFFQX1 d_lt_aswk_reg_0_ ( .D(lt_aswk[0]), .SIN(reg14[3]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[0]) );
  SDFFQX1 d_regx_addr_reg_4_ ( .D(regx_addr[4]), .SIN(d_regx_addr[3]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[4]) );
  SDFFQX1 d_regx_addr_reg_3_ ( .D(regx_addr[3]), .SIN(d_regx_addr[2]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[3]) );
  SDFFQX1 d_regx_addr_reg_2_ ( .D(regx_addr[2]), .SIN(d_regx_addr[1]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[2]) );
  SDFFQX1 d_lt_gpi_reg_3_ ( .D(lt_gpi[3]), .SIN(d_lt_gpi[2]), .SMC(test_se), 
        .C(net8996), .Q(d_lt_gpi[3]) );
  SDFFQX1 d_regx_addr_reg_0_ ( .D(regx_addr[0]), .SIN(d_lt_gpi[3]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[0]) );
  SDFFQX1 d_regx_addr_reg_1_ ( .D(regx_addr[1]), .SIN(d_regx_addr[0]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[1]) );
  SDFFQX1 d_regx_addr_reg_6_ ( .D(regx_addr[6]), .SIN(d_regx_addr[5]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[6]) );
  SDFFQX1 d_regx_addr_reg_5_ ( .D(regx_addr[5]), .SIN(d_regx_addr[4]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[5]) );
  SDFFRQX1 lt_drp_reg ( .D(di_drposc), .SIN(lt_aswk[5]), .SMC(test_se), .C(
        detclk), .XR(n52), .Q(lt_drp) );
  SDFFRQX1 lt_aswk_reg_5_ ( .D(1'b1), .SIN(lt_aswk[4]), .SMC(test_se), .C(
        aswclk), .XR(n73), .Q(lt_aswk[5]) );
  SDFFRQX1 lt_aswk_reg_4_ ( .D(di_aswk[4]), .SIN(lt_aswk[3]), .SMC(test_se), 
        .C(aswclk), .XR(n73), .Q(lt_aswk[4]) );
  SDFFRQX1 lt_aswk_reg_3_ ( .D(di_aswk[3]), .SIN(lt_aswk[2]), .SMC(test_se), 
        .C(aswclk), .XR(n73), .Q(lt_aswk[3]) );
  SDFFRQX1 lt_aswk_reg_2_ ( .D(di_aswk[2]), .SIN(lt_aswk[1]), .SMC(test_se), 
        .C(aswclk), .XR(n73), .Q(lt_aswk[2]) );
  SDFFRQX1 lt_aswk_reg_1_ ( .D(di_aswk[1]), .SIN(lt_aswk[0]), .SMC(test_se), 
        .C(aswclk), .XR(n73), .Q(lt_aswk[1]) );
  SDFFRQX1 lt_aswk_reg_0_ ( .D(di_aswk[0]), .SIN(d_we16), .SMC(test_se), .C(
        aswclk), .XR(n73), .Q(lt_aswk[0]) );
  NAND32XL U4 ( .B(regx_addr[0]), .C(n68), .A(n76), .Y(n69) );
  INVX3 U7 ( .A(n101), .Y(n105) );
  INVX3 U8 ( .A(regx_addr[2]), .Y(n76) );
  AND3X1 U9 ( .A(n107), .B(n126), .C(n121), .Y(regx_wrdac[12]) );
  NAND32X1 U10 ( .B(regx_addr[1]), .C(n25), .A(n76), .Y(n97) );
  INVX1 U11 ( .A(regx_addr[3]), .Y(n121) );
  INVX2 U12 ( .A(n77), .Y(n126) );
  NAND32XL U13 ( .B(regx_addr[0]), .C(regx_addr[1]), .A(n76), .Y(n77) );
  INVX1 U14 ( .A(n100), .Y(n107) );
  INVX1 U15 ( .A(n67), .Y(n102) );
  NOR2XL U16 ( .A(regx_addr[0]), .B(n78), .Y(n1) );
  INVX2 U17 ( .A(regx_addr[0]), .Y(n25) );
  INVXL U18 ( .A(regx_wdat[3]), .Y(n5) );
  INVXL U19 ( .A(n5), .Y(n6) );
  INVXL U20 ( .A(n5), .Y(n7) );
  INVXL U21 ( .A(regx_wdat[4]), .Y(n8) );
  INVXL U22 ( .A(n8), .Y(n9) );
  INVXL U23 ( .A(n8), .Y(n10) );
  INVXL U24 ( .A(regx_wdat[5]), .Y(n11) );
  INVXL U25 ( .A(n11), .Y(n12) );
  INVXL U26 ( .A(n11), .Y(n13) );
  INVXL U27 ( .A(regx_wdat[6]), .Y(n14) );
  INVXL U28 ( .A(n14), .Y(n15) );
  INVXL U29 ( .A(n14), .Y(n16) );
  INVXL U30 ( .A(d_regx_addr[2]), .Y(n17) );
  INVXL U31 ( .A(n17), .Y(n18) );
  INVXL U32 ( .A(d_regx_addr[3]), .Y(n19) );
  INVXL U33 ( .A(n19), .Y(n20) );
  INVX1 U34 ( .A(n132), .Y(n21) );
  INVX1 U35 ( .A(n21), .Y(r_i2crout[5]) );
  BUFX3 U36 ( .A(r_imp_osc), .Y(r_xana[22]) );
  NAND43XL U37 ( .B(regx_addr[5]), .C(regx_addr[6]), .D(regx_addr[3]), .A(
        regx_addr[4]), .Y(n125) );
  INVX1 U38 ( .A(regx_addr[4]), .Y(n120) );
  AND2X2 U39 ( .A(n105), .B(n119), .Y(regx_wrdac[4]) );
  NOR2XL U40 ( .A(n78), .B(n25), .Y(n24) );
  INVX1 U41 ( .A(regx_addr[1]), .Y(n68) );
  AND2X1 U42 ( .A(n102), .B(n105), .Y(regx_wrdac[5]) );
  AND2X2 U43 ( .A(n105), .B(n128), .Y(regx_wrdac[3]) );
  INVXL U44 ( .A(n96), .Y(n106) );
  NAND21XL U45 ( .B(n92), .A(n104), .Y(n89) );
  AND2XL U46 ( .A(n124), .B(n128), .Y(regx_wrpwm[1]) );
  AND2XL U47 ( .A(n23), .B(n104), .Y(we[29]) );
  NAND32XL U48 ( .B(n120), .C(n98), .A(n95), .Y(n96) );
  AND3XL U49 ( .A(n107), .B(n128), .C(n121), .Y(regx_wrdac[13]) );
  AND2XL U50 ( .A(n105), .B(n24), .Y(regx_wrdac[9]) );
  AND2XL U51 ( .A(n103), .B(n105), .Y(regx_wrdac[6]) );
  AND3XL U52 ( .A(n106), .B(n128), .C(n121), .Y(regx_wrdac[1]) );
  AND2XL U53 ( .A(n105), .B(n126), .Y(regx_wrdac[2]) );
  INVXL U54 ( .A(n99), .Y(n95) );
  AND2XL U55 ( .A(n119), .B(n118), .Y(regx_wrcvc[2]) );
  NAND21XL U56 ( .B(n92), .A(n119), .Y(n93) );
  NAND32XL U57 ( .B(n122), .C(n121), .A(n120), .Y(n123) );
  AND2XL U58 ( .A(n23), .B(n119), .Y(we[26]) );
  AND2XL U59 ( .A(n104), .B(n118), .Y(we_5) );
  AND3XL U60 ( .A(regx_addr[3]), .B(n128), .C(n106), .Y(regx_wrdac[11]) );
  AND3XL U61 ( .A(regx_addr[3]), .B(n126), .C(n106), .Y(regx_wrdac[10]) );
  INVXL U62 ( .A(n66), .Y(n103) );
  NAND21XL U63 ( .B(regx_addr[5]), .A(n95), .Y(n122) );
  INVX1 U64 ( .A(n89), .Y(n75) );
  AND2X1 U65 ( .A(n104), .B(n105), .Y(regx_wrdac[7]) );
  INVX1 U66 ( .A(n92), .Y(n129) );
  AND2X1 U67 ( .A(n102), .B(n129), .Y(we_19) );
  AND2X1 U93 ( .A(n23), .B(n102), .Y(we[27]) );
  NAND32X1 U94 ( .B(n99), .C(n98), .A(n120), .Y(n100) );
  AND3XL U95 ( .A(n106), .B(n126), .C(n121), .Y(regx_wrdac[0]) );
  NAND21X2 U96 ( .B(n121), .A(n107), .Y(n101) );
  INVX1 U97 ( .A(n97), .Y(n128) );
  INVX1 U98 ( .A(n65), .Y(n104) );
  NAND32X1 U99 ( .B(n76), .C(n25), .A(n68), .Y(n65) );
  NAND32X1 U100 ( .B(n68), .C(n25), .A(n76), .Y(n67) );
  AND2XL U101 ( .A(n126), .B(n127), .Y(regx_hitbst[0]) );
  INVX1 U102 ( .A(n125), .Y(n127) );
  NAND21X1 U103 ( .B(n125), .A(regx_w), .Y(n92) );
  INVX1 U104 ( .A(n93), .Y(we_twlb) );
  AND2XL U105 ( .A(n118), .B(n126), .Y(regx_wrcvc[0]) );
  AND2X1 U106 ( .A(n24), .B(n124), .Y(regx_wrcvc[3]) );
  AND2XL U107 ( .A(n118), .B(n128), .Y(regx_wrcvc[1]) );
  AND2XL U108 ( .A(n124), .B(n126), .Y(regx_wrpwm[0]) );
  INVX1 U109 ( .A(n123), .Y(n124) );
  NOR3XL U110 ( .A(n120), .B(n121), .C(n122), .Y(n23) );
  AND2XL U111 ( .A(n128), .B(n127), .Y(regx_hitbst[1]) );
  AND2X1 U112 ( .A(n103), .B(n118), .Y(we_4) );
  AND2X1 U113 ( .A(n118), .B(n24), .Y(we_7) );
  AND2XL U114 ( .A(n118), .B(n1), .Y(we_6) );
  AND2X1 U115 ( .A(n24), .B(n129), .Y(we[23]) );
  AND2XL U116 ( .A(n23), .B(n1), .Y(we[30]) );
  AND2X1 U117 ( .A(n23), .B(n103), .Y(we[28]) );
  AND2XL U118 ( .A(n23), .B(n126), .Y(we[24]) );
  INVX1 U119 ( .A(n70), .Y(n74) );
  NAND21X1 U120 ( .B(n97), .A(n23), .Y(n70) );
  INVX1 U121 ( .A(n29), .Y(wd_twlb[0]) );
  INVX1 U122 ( .A(n32), .Y(wd_twlb[1]) );
  INVX1 U123 ( .A(n61), .Y(n33) );
  INVX1 U124 ( .A(n29), .Y(n28) );
  INVX1 U125 ( .A(n32), .Y(n31) );
  INVX1 U126 ( .A(n61), .Y(n59) );
  INVX1 U127 ( .A(n64), .Y(n62) );
  INVX1 U128 ( .A(n64), .Y(n63) );
  NAND21X1 U129 ( .B(regx_addr[6]), .A(regx_w), .Y(n99) );
  INVX1 U130 ( .A(n69), .Y(n119) );
  NAND32XL U131 ( .B(regx_addr[0]), .C(n76), .A(n68), .Y(n66) );
  INVX1 U132 ( .A(regx_addr[5]), .Y(n98) );
  AO21X1 U133 ( .B(bus_idle), .C(n91), .A(n90), .Y(i2c_mode_upd) );
  AND3X1 U134 ( .A(n75), .B(n62), .C(n14), .Y(n90) );
  NAND43X1 U135 ( .B(n88), .C(n87), .D(n86), .A(n85), .Y(n91) );
  NOR43XL U136 ( .B(n61), .C(n32), .D(n130), .A(n71), .Y(N8) );
  NAND3X1 U137 ( .A(n8), .B(n11), .C(n5), .Y(n71) );
  AND4XL U138 ( .A(n72), .B(wd_twlb[0]), .C(n1), .D(n129), .Y(n130) );
  NOR21XL U139 ( .B(n15), .A(n64), .Y(n72) );
  INVX1 U140 ( .A(n94), .Y(n118) );
  NAND32XL U141 ( .B(regx_addr[3]), .C(n122), .A(n120), .Y(n94) );
  INVX1 U142 ( .A(regx_wdat[2]), .Y(n61) );
  INVX1 U143 ( .A(regx_wdat[1]), .Y(n32) );
  INVX1 U144 ( .A(regx_wdat[0]), .Y(n29) );
  INVX1 U145 ( .A(regx_wdat[7]), .Y(n64) );
  XNOR2XL U146 ( .A(reg1E[3]), .B(n60), .Y(r_xana[19]) );
  XNOR2XL U147 ( .A(reg1E[2]), .B(n60), .Y(r_xana[18]) );
  NAND2X1 U148 ( .A(r_xana[20]), .B(di_drposc), .Y(n60) );
  AND4X1 U149 ( .A(n84), .B(n89), .C(n83), .D(n82), .Y(n85) );
  XOR2X1 U150 ( .A(n79), .B(r_i2crout[2]), .Y(n84) );
  XOR2X1 U151 ( .A(n80), .B(r_i2crout[1]), .Y(n83) );
  XOR2X1 U152 ( .A(n81), .B(r_i2crout[0]), .Y(n82) );
  MUX2X1 U153 ( .D0(lt_reg15_5_0[2]), .D1(n59), .S(n75), .Y(i2c_mode_wdat[2])
         );
  MUX2X1 U154 ( .D0(lt_reg15_5_0[0]), .D1(n28), .S(n75), .Y(i2c_mode_wdat[0])
         );
  MUX2X1 U155 ( .D0(lt_reg15_5_0[1]), .D1(n31), .S(n75), .Y(i2c_mode_wdat[1])
         );
  MUX2BXL U156 ( .D0(lt_reg15_5_0[3]), .D1(n5), .S(n75), .Y(i2c_mode_wdat[3])
         );
  MUX2BXL U157 ( .D0(lt_reg15_5_0[4]), .D1(n8), .S(n75), .Y(i2c_mode_wdat[4])
         );
  MUX2BXL U158 ( .D0(lt_reg15_5_0[5]), .D1(n11), .S(n75), .Y(i2c_mode_wdat[5])
         );
  XOR2X1 U159 ( .A(r_i2crout[4]), .B(lt_reg15_5_0[4]), .Y(n88) );
  XOR2X1 U160 ( .A(n132), .B(lt_reg15_5_0[5]), .Y(n87) );
  XOR2X1 U161 ( .A(r_i2crout[3]), .B(lt_reg15_5_0[3]), .Y(n86) );
  INVX1 U162 ( .A(lt_reg15_5_0[0]), .Y(n81) );
  INVX1 U163 ( .A(lt_reg15_5_0[1]), .Y(n80) );
  INVX1 U164 ( .A(lt_reg15_5_0[2]), .Y(n79) );
  OA21X1 U165 ( .B(n131), .C(atpg_en), .A(n50), .Y(n73) );
  INVX1 U166 ( .A(d_we16), .Y(n131) );
  AND2X2 U167 ( .A(n105), .B(n1), .Y(regx_wrdac[8]) );
  NAND21X1 U168 ( .B(n76), .A(regx_addr[1]), .Y(n78) );
endmodule


module regx_a0_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745;

  BUFXL U2149 ( .A(SH[5]), .Y(n3667) );
  BUFXL U2150 ( .A(SH[6]), .Y(n3668) );
  INVX1 U2151 ( .A(n3702), .Y(n3689) );
  INVX1 U2152 ( .A(n3702), .Y(n3690) );
  INVX1 U2153 ( .A(n3699), .Y(n3697) );
  INVX1 U2154 ( .A(n3738), .Y(n3728) );
  INVX1 U2155 ( .A(n3740), .Y(n3729) );
  INVX1 U2156 ( .A(n3740), .Y(n3727) );
  INVX1 U2157 ( .A(n3699), .Y(n3698) );
  INVX1 U2158 ( .A(n3702), .Y(n3688) );
  INVX1 U2159 ( .A(n3738), .Y(n3720) );
  INVX1 U2160 ( .A(n3738), .Y(n3719) );
  INVX1 U2161 ( .A(n3738), .Y(n3718) );
  INVX1 U2162 ( .A(n3739), .Y(n3722) );
  INVX1 U2163 ( .A(n3701), .Y(n3691) );
  INVX1 U2164 ( .A(n3700), .Y(n3694) );
  INVX1 U2165 ( .A(n3740), .Y(n3732) );
  INVX1 U2166 ( .A(n3740), .Y(n3725) );
  INVX1 U2167 ( .A(n3739), .Y(n3735) );
  INVX1 U2168 ( .A(n3737), .Y(n3736) );
  NOR3XL U2169 ( .A(A[175]), .B(n3728), .C(n3697), .Y(n3279) );
  INVX1 U2170 ( .A(n3703), .Y(n3686) );
  INVX1 U2171 ( .A(n3703), .Y(n3687) );
  INVX1 U2172 ( .A(n3704), .Y(n3684) );
  INVX1 U2173 ( .A(n3703), .Y(n3685) );
  INVX1 U2174 ( .A(n3738), .Y(n3721) );
  INVX1 U2175 ( .A(n3739), .Y(n3723) );
  INVX1 U2176 ( .A(n3699), .Y(n3696) );
  INVX1 U2177 ( .A(n3701), .Y(n3692) );
  INVX1 U2178 ( .A(n3705), .Y(n3695) );
  INVX1 U2179 ( .A(n3700), .Y(n3693) );
  INVX1 U2180 ( .A(n3740), .Y(n3731) );
  INVX1 U2181 ( .A(n3740), .Y(n3733) );
  INVX1 U2182 ( .A(n3738), .Y(n3730) );
  INVX1 U2183 ( .A(n3738), .Y(n3726) );
  INVX1 U2184 ( .A(n3739), .Y(n3724) );
  INVX1 U2185 ( .A(n3740), .Y(n3734) );
  INVX1 U2186 ( .A(n3713), .Y(n3702) );
  INVX1 U2187 ( .A(n3714), .Y(n3699) );
  INVX1 U2188 ( .A(n3743), .Y(n3737) );
  INVX1 U2189 ( .A(n3742), .Y(n3738) );
  INVX1 U2190 ( .A(n3741), .Y(n3740) );
  INVX1 U2191 ( .A(n3742), .Y(n3739) );
  INVX1 U2192 ( .A(n3711), .Y(n3706) );
  INVX1 U2193 ( .A(n3713), .Y(n3701) );
  INVX1 U2194 ( .A(n3714), .Y(n3700) );
  INVX1 U2195 ( .A(n3713), .Y(n3703) );
  INVX1 U2196 ( .A(n3712), .Y(n3704) );
  INVX1 U2197 ( .A(n3712), .Y(n3705) );
  MUX4X1 U2198 ( .D0(n3301), .D1(n3302), .D2(n3303), .D3(n3304), .S0(n3669), 
        .S1(n3682), .Y(n3289) );
  NOR3XL U2199 ( .A(n3707), .B(n3729), .C(A[343]), .Y(n3303) );
  NOR3XL U2200 ( .A(n3706), .B(n3729), .C(A[351]), .Y(n3304) );
  NOR21XL U2201 ( .B(n3306), .A(n3720), .Y(n3301) );
  MUX4X1 U2202 ( .D0(n3292), .D1(n3293), .D2(n3294), .D3(n3295), .S0(n3677), 
        .S1(n3673), .Y(n3291) );
  NOR3XL U2203 ( .A(n3708), .B(n3728), .C(A[367]), .Y(n3294) );
  NOR3XL U2204 ( .A(n3708), .B(n3728), .C(A[359]), .Y(n3292) );
  NOR3XL U2205 ( .A(n3706), .B(n3728), .C(A[375]), .Y(n3293) );
  MUX4X1 U2206 ( .D0(n3549), .D1(n3550), .D2(n3551), .D3(n3552), .S0(n3669), 
        .S1(n3681), .Y(n3537) );
  NOR3XL U2207 ( .A(n3716), .B(n3736), .C(A[338]), .Y(n3551) );
  NOR3XL U2208 ( .A(n3707), .B(n3743), .C(A[346]), .Y(n3552) );
  NOR21XL U2209 ( .B(n3554), .A(n3722), .Y(n3549) );
  MUX4X1 U2210 ( .D0(n3399), .D1(n3400), .D2(n3401), .D3(n3402), .S0(n3670), 
        .S1(n3681), .Y(n3387) );
  NOR3XL U2211 ( .A(n3716), .B(n3732), .C(A[341]), .Y(n3401) );
  NOR3XL U2212 ( .A(n3705), .B(n3732), .C(A[349]), .Y(n3402) );
  NOR21XL U2213 ( .B(n3404), .A(n3744), .Y(n3399) );
  MUX4X1 U2214 ( .D0(n3602), .D1(n3603), .D2(n3604), .D3(n3605), .S0(n3670), 
        .S1(n3682), .Y(n3590) );
  NOR3XL U2215 ( .A(n3703), .B(n3742), .C(A[337]), .Y(n3604) );
  NOR3XL U2216 ( .A(n3705), .B(n3741), .C(A[345]), .Y(n3605) );
  NOR21XL U2217 ( .B(n3607), .A(n3720), .Y(n3602) );
  MUX4X1 U2218 ( .D0(n3449), .D1(n3450), .D2(n3451), .D3(n3452), .S0(n3670), 
        .S1(n3681), .Y(n3437) );
  NOR3XL U2219 ( .A(n3704), .B(n3734), .C(A[340]), .Y(n3451) );
  NOR3XL U2220 ( .A(n3716), .B(SH[9]), .C(A[348]), .Y(n3452) );
  NOR21XL U2221 ( .B(n3454), .A(n3720), .Y(n3449) );
  MUX4X1 U2222 ( .D0(n3349), .D1(n3350), .D2(n3351), .D3(n3352), .S0(n3670), 
        .S1(n3681), .Y(n3337) );
  NOR3XL U2223 ( .A(n3704), .B(n3730), .C(A[342]), .Y(n3351) );
  NOR3XL U2224 ( .A(n3706), .B(n3730), .C(A[350]), .Y(n3352) );
  NOR21XL U2225 ( .B(n3354), .A(n3721), .Y(n3349) );
  MUX4X1 U2226 ( .D0(n3655), .D1(n3656), .D2(n3657), .D3(n3658), .S0(n3670), 
        .S1(n3682), .Y(n3643) );
  NOR3XL U2227 ( .A(n3707), .B(n3723), .C(A[336]), .Y(n3657) );
  NOR3XL U2228 ( .A(n3704), .B(n3727), .C(A[344]), .Y(n3658) );
  NOR21XL U2229 ( .B(n3660), .A(n3718), .Y(n3655) );
  MUX4X1 U2230 ( .D0(n3499), .D1(n3500), .D2(n3501), .D3(n3502), .S0(n3670), 
        .S1(n3681), .Y(n3487) );
  NOR3XL U2231 ( .A(n3703), .B(n3723), .C(A[339]), .Y(n3501) );
  NOR3XL U2232 ( .A(n3704), .B(n3725), .C(A[347]), .Y(n3502) );
  NOR21XL U2233 ( .B(n3504), .A(n3719), .Y(n3499) );
  MUX4X1 U2234 ( .D0(n3390), .D1(n3391), .D2(n3392), .D3(n3393), .S0(SH[4]), 
        .S1(n3671), .Y(n3389) );
  NOR3XL U2235 ( .A(n3704), .B(n3731), .C(A[365]), .Y(n3392) );
  NOR3XL U2236 ( .A(n3705), .B(n3732), .C(A[357]), .Y(n3390) );
  NOR3XL U2237 ( .A(n3704), .B(n3732), .C(A[373]), .Y(n3391) );
  MUX4X1 U2238 ( .D0(n3593), .D1(n3594), .D2(n3595), .D3(n3596), .S0(n3682), 
        .S1(n3674), .Y(n3592) );
  NOR3XL U2239 ( .A(n3708), .B(SH[9]), .C(A[361]), .Y(n3595) );
  NOR3XL U2240 ( .A(n3705), .B(n3741), .C(A[353]), .Y(n3593) );
  NOR3XL U2241 ( .A(n3705), .B(n3741), .C(A[369]), .Y(n3594) );
  MUX4X1 U2242 ( .D0(n3440), .D1(n3441), .D2(n3442), .D3(n3443), .S0(SH[4]), 
        .S1(n3673), .Y(n3439) );
  NOR3XL U2243 ( .A(n3708), .B(n3741), .C(A[364]), .Y(n3442) );
  NOR3XL U2244 ( .A(n3707), .B(n3741), .C(A[356]), .Y(n3440) );
  NOR3XL U2245 ( .A(n3708), .B(SH[9]), .C(A[372]), .Y(n3441) );
  MUX4X1 U2246 ( .D0(n3340), .D1(n3341), .D2(n3342), .D3(n3343), .S0(n3678), 
        .S1(n3673), .Y(n3339) );
  NOR3XL U2247 ( .A(n3707), .B(n3730), .C(A[366]), .Y(n3342) );
  NOR3XL U2248 ( .A(n3707), .B(n3730), .C(A[358]), .Y(n3340) );
  NOR3XL U2249 ( .A(n3703), .B(n3730), .C(A[374]), .Y(n3341) );
  MUX4X1 U2250 ( .D0(n3646), .D1(n3647), .D2(n3648), .D3(n3649), .S0(n3677), 
        .S1(n3674), .Y(n3645) );
  NOR3XL U2251 ( .A(n3703), .B(n3727), .C(A[360]), .Y(n3648) );
  NOR3XL U2252 ( .A(n3704), .B(n3727), .C(A[352]), .Y(n3646) );
  NOR3XL U2253 ( .A(n3705), .B(n3727), .C(A[368]), .Y(n3647) );
  MUX4X1 U2254 ( .D0(n3490), .D1(n3491), .D2(n3492), .D3(n3493), .S0(n3679), 
        .S1(n3673), .Y(n3489) );
  NOR3XL U2255 ( .A(n3703), .B(n3724), .C(A[363]), .Y(n3492) );
  NOR3XL U2256 ( .A(n3704), .B(n3723), .C(A[355]), .Y(n3490) );
  NOR3XL U2257 ( .A(n3703), .B(n3724), .C(A[371]), .Y(n3491) );
  MUX4X1 U2258 ( .D0(n3540), .D1(n3541), .D2(n3542), .D3(n3543), .S0(n3680), 
        .S1(SH[3]), .Y(n3539) );
  NOR3XL U2259 ( .A(n3716), .B(n3725), .C(A[362]), .Y(n3542) );
  NOR3XL U2260 ( .A(n3706), .B(n3725), .C(A[354]), .Y(n3540) );
  NOR3XL U2261 ( .A(n3706), .B(n3725), .C(A[370]), .Y(n3541) );
  INVX1 U2262 ( .A(n3715), .Y(n3713) );
  INVX1 U2263 ( .A(n3715), .Y(n3714) );
  INVX1 U2264 ( .A(n3737), .Y(n3741) );
  INVX1 U2265 ( .A(n3676), .Y(n3669) );
  INVX1 U2266 ( .A(n3710), .Y(n3707) );
  INVX1 U2267 ( .A(n3710), .Y(n3708) );
  INVX1 U2268 ( .A(n3745), .Y(n3743) );
  INVX1 U2269 ( .A(n3716), .Y(n3711) );
  INVX1 U2270 ( .A(n3737), .Y(n3742) );
  INVX1 U2271 ( .A(n3710), .Y(n3709) );
  INVX1 U2272 ( .A(n3676), .Y(n3670) );
  INVX1 U2273 ( .A(n3683), .Y(n3681) );
  INVX1 U2274 ( .A(n3676), .Y(n3672) );
  INVX1 U2275 ( .A(n3676), .Y(n3674) );
  INVX1 U2276 ( .A(n3676), .Y(n3673) );
  INVX1 U2277 ( .A(n3683), .Y(n3682) );
  INVX1 U2278 ( .A(n3715), .Y(n3712) );
  INVX1 U2279 ( .A(n3676), .Y(n3675) );
  INVX1 U2280 ( .A(n3745), .Y(n3744) );
  INVX1 U2281 ( .A(n3683), .Y(n3678) );
  INVX1 U2282 ( .A(n3683), .Y(n3679) );
  INVX1 U2283 ( .A(n3683), .Y(n3680) );
  INVX1 U2284 ( .A(n3676), .Y(n3671) );
  MUX2IX1 U2285 ( .D0(A[15]), .D1(A[271]), .S(n3690), .Y(n3311) );
  MUX2IX1 U2286 ( .D0(n3264), .D1(n3265), .S(SH[7]), .Y(B[7]) );
  MUX4X1 U2287 ( .D0(n3266), .D1(n3267), .D2(n3268), .D3(n3269), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3265) );
  MUX4X1 U2288 ( .D0(n3288), .D1(n3289), .D2(n3290), .D3(n3291), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3264) );
  MUX3X1 U2289 ( .D0(n3278), .D1(n3279), .D2(n3280), .S0(n3675), .S1(n3682), 
        .Y(n3267) );
  MUX2IX1 U2290 ( .D0(A[71]), .D1(A[327]), .S(n3690), .Y(n3306) );
  NOR21XL U2291 ( .B(n3296), .A(n3718), .Y(n3295) );
  MUX2IX1 U2292 ( .D0(A[127]), .D1(A[383]), .S(n3689), .Y(n3296) );
  NOR21XL U2293 ( .B(n3305), .A(n3719), .Y(n3302) );
  MUX2IX1 U2294 ( .D0(A[79]), .D1(A[335]), .S(n3689), .Y(n3305) );
  MUX2X1 U2295 ( .D0(n3307), .D1(n3308), .S(n3681), .Y(n3288) );
  NOR4XL U2296 ( .A(n3722), .B(n3691), .C(n3670), .D(A[23]), .Y(n3308) );
  MUX2IX1 U2297 ( .D0(n3309), .D1(n3310), .S(n3669), .Y(n3307) );
  NAND2X1 U2298 ( .A(n3311), .B(n3737), .Y(n3310) );
  NAND2X1 U2299 ( .A(n3312), .B(n3737), .Y(n3309) );
  MUX2IX1 U2300 ( .D0(A[7]), .D1(A[263]), .S(n3688), .Y(n3312) );
  MUX2IX1 U2301 ( .D0(n3313), .D1(n3314), .S(SH[7]), .Y(B[6]) );
  MUX4X1 U2302 ( .D0(n3315), .D1(n3316), .D2(n3317), .D3(n3318), .S0(SH[5]), 
        .S1(n3668), .Y(n3314) );
  MUX4X1 U2303 ( .D0(n3336), .D1(n3337), .D2(n3338), .D3(n3339), .S0(SH[6]), 
        .S1(n3667), .Y(n3313) );
  MUX2X1 U2304 ( .D0(n3327), .D1(n3328), .S(n3681), .Y(n3316) );
  MUX2IX1 U2305 ( .D0(A[13]), .D1(A[269]), .S(n3686), .Y(n3409) );
  MUX2IX1 U2306 ( .D0(A[9]), .D1(A[265]), .S(n3688), .Y(n3612) );
  MUX2IX1 U2307 ( .D0(A[12]), .D1(A[268]), .S(n3688), .Y(n3459) );
  MUX2IX1 U2308 ( .D0(A[11]), .D1(A[267]), .S(n3684), .Y(n3509) );
  MUX2IX1 U2309 ( .D0(A[10]), .D1(A[266]), .S(n3685), .Y(n3559) );
  MUX2IX1 U2310 ( .D0(n3361), .D1(n3362), .S(SH[7]), .Y(B[5]) );
  MUX4X1 U2311 ( .D0(n3363), .D1(n3364), .D2(n3365), .D3(n3366), .S0(n3667), 
        .S1(n3668), .Y(n3362) );
  MUX4X1 U2312 ( .D0(n3386), .D1(n3387), .D2(n3388), .D3(n3389), .S0(n3668), 
        .S1(n3667), .Y(n3361) );
  MUX4X1 U2313 ( .D0(n3371), .D1(n3372), .D2(n3373), .D3(n3374), .S0(n3678), 
        .S1(n3672), .Y(n3365) );
  MUX2IX1 U2314 ( .D0(n3561), .D1(n3562), .S(SH[7]), .Y(B[1]) );
  MUX4X1 U2315 ( .D0(n3563), .D1(n3564), .D2(n3565), .D3(n3566), .S0(SH[5]), 
        .S1(n3668), .Y(n3562) );
  MUX4X1 U2316 ( .D0(n3589), .D1(n3590), .D2(n3591), .D3(n3592), .S0(SH[6]), 
        .S1(n3667), .Y(n3561) );
  MUX4X1 U2317 ( .D0(n3567), .D1(n3568), .D2(n3569), .D3(n3570), .S0(n3680), 
        .S1(n3675), .Y(n3566) );
  MUX2IX1 U2318 ( .D0(n3411), .D1(n3412), .S(SH[7]), .Y(B[4]) );
  MUX4X1 U2319 ( .D0(n3413), .D1(n3414), .D2(n3415), .D3(n3416), .S0(n3667), 
        .S1(n3668), .Y(n3412) );
  MUX4X1 U2320 ( .D0(n3436), .D1(n3437), .D2(n3438), .D3(n3439), .S0(n3668), 
        .S1(n3667), .Y(n3411) );
  MUX4X1 U2321 ( .D0(n3421), .D1(n3422), .D2(n3423), .D3(n3424), .S0(n3682), 
        .S1(n3672), .Y(n3415) );
  MUX2IX1 U2322 ( .D0(n3614), .D1(n3615), .S(SH[7]), .Y(B[0]) );
  MUX4X1 U2323 ( .D0(n3616), .D1(n3617), .D2(n3618), .D3(n3619), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3615) );
  MUX4X1 U2324 ( .D0(n3642), .D1(n3643), .D2(n3644), .D3(n3645), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3614) );
  MUX4X1 U2325 ( .D0(n3620), .D1(n3621), .D2(n3622), .D3(n3623), .S0(n3678), 
        .S1(n3674), .Y(n3619) );
  MUX2IX1 U2326 ( .D0(n3461), .D1(n3462), .S(SH[7]), .Y(B[3]) );
  MUX4X1 U2327 ( .D0(n3463), .D1(n3464), .D2(n3465), .D3(n3466), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3462) );
  MUX4X1 U2328 ( .D0(n3486), .D1(n3487), .D2(n3488), .D3(n3489), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3461) );
  MUX4X1 U2329 ( .D0(n3471), .D1(n3472), .D2(n3473), .D3(n3474), .S0(n3679), 
        .S1(n3673), .Y(n3465) );
  MUX2IX1 U2330 ( .D0(n3511), .D1(n3512), .S(SH[7]), .Y(B[2]) );
  MUX4X1 U2331 ( .D0(n3513), .D1(n3514), .D2(n3515), .D3(n3516), .S0(SH[5]), 
        .S1(n3668), .Y(n3512) );
  MUX4X1 U2332 ( .D0(n3536), .D1(n3537), .D2(n3538), .D3(n3539), .S0(SH[6]), 
        .S1(n3667), .Y(n3511) );
  MUX4X1 U2333 ( .D0(n3521), .D1(n3522), .D2(n3523), .D3(n3524), .S0(n3680), 
        .S1(n3675), .Y(n3515) );
  MUX2IX1 U2334 ( .D0(A[69]), .D1(A[325]), .S(n3687), .Y(n3404) );
  MUX2IX1 U2335 ( .D0(A[65]), .D1(A[321]), .S(n3688), .Y(n3607) );
  MUX2IX1 U2336 ( .D0(A[68]), .D1(A[324]), .S(n3685), .Y(n3454) );
  MUX2IX1 U2337 ( .D0(A[70]), .D1(A[326]), .S(n3688), .Y(n3354) );
  MUX2IX1 U2338 ( .D0(A[64]), .D1(A[320]), .S(n3690), .Y(n3660) );
  MUX2IX1 U2339 ( .D0(A[67]), .D1(A[323]), .S(n3684), .Y(n3504) );
  MUX2IX1 U2340 ( .D0(A[66]), .D1(A[322]), .S(n3685), .Y(n3554) );
  NOR21XL U2341 ( .B(n3403), .A(n3722), .Y(n3400) );
  MUX2IX1 U2342 ( .D0(A[77]), .D1(A[333]), .S(n3687), .Y(n3403) );
  NOR21XL U2343 ( .B(n3606), .A(n3720), .Y(n3603) );
  MUX2IX1 U2344 ( .D0(A[73]), .D1(A[329]), .S(n3687), .Y(n3606) );
  NOR21XL U2345 ( .B(n3453), .A(n3720), .Y(n3450) );
  MUX2IX1 U2346 ( .D0(A[76]), .D1(A[332]), .S(n3685), .Y(n3453) );
  NOR21XL U2347 ( .B(n3353), .A(n3721), .Y(n3350) );
  MUX2IX1 U2348 ( .D0(A[78]), .D1(A[334]), .S(n3689), .Y(n3353) );
  NOR21XL U2349 ( .B(n3659), .A(n3718), .Y(n3656) );
  MUX2IX1 U2350 ( .D0(A[72]), .D1(A[328]), .S(n3689), .Y(n3659) );
  NOR21XL U2351 ( .B(n3503), .A(n3719), .Y(n3500) );
  MUX2IX1 U2352 ( .D0(A[75]), .D1(A[331]), .S(n3684), .Y(n3503) );
  NOR21XL U2353 ( .B(n3553), .A(n3720), .Y(n3550) );
  MUX2IX1 U2354 ( .D0(A[74]), .D1(A[330]), .S(n3685), .Y(n3553) );
  NOR21XL U2355 ( .B(n3394), .A(n3720), .Y(n3393) );
  MUX2IX1 U2356 ( .D0(A[125]), .D1(A[381]), .S(n3687), .Y(n3394) );
  NOR21XL U2357 ( .B(n3597), .A(n3721), .Y(n3596) );
  MUX2IX1 U2358 ( .D0(A[121]), .D1(A[377]), .S(n3687), .Y(n3597) );
  NOR21XL U2359 ( .B(n3444), .A(n3721), .Y(n3443) );
  MUX2IX1 U2360 ( .D0(A[124]), .D1(A[380]), .S(n3686), .Y(n3444) );
  NOR21XL U2361 ( .B(n3344), .A(n3721), .Y(n3343) );
  MUX2IX1 U2362 ( .D0(A[126]), .D1(A[382]), .S(n3689), .Y(n3344) );
  NOR21XL U2363 ( .B(n3650), .A(n3718), .Y(n3649) );
  MUX2IX1 U2364 ( .D0(A[120]), .D1(A[376]), .S(n3689), .Y(n3650) );
  NOR21XL U2365 ( .B(n3494), .A(n3718), .Y(n3493) );
  MUX2IX1 U2366 ( .D0(A[123]), .D1(A[379]), .S(n3684), .Y(n3494) );
  NOR21XL U2367 ( .B(n3544), .A(n3722), .Y(n3543) );
  MUX2IX1 U2368 ( .D0(A[122]), .D1(A[378]), .S(n3685), .Y(n3544) );
  MUX2X1 U2369 ( .D0(n3405), .D1(n3406), .S(n3681), .Y(n3386) );
  NOR4XL U2370 ( .A(n3723), .B(n3691), .C(n3670), .D(A[21]), .Y(n3406) );
  MUX2IX1 U2371 ( .D0(n3407), .D1(n3408), .S(n3669), .Y(n3405) );
  NAND2X1 U2372 ( .A(n3409), .B(n3745), .Y(n3408) );
  MUX2X1 U2373 ( .D0(n3608), .D1(n3609), .S(n3680), .Y(n3589) );
  NOR4XL U2374 ( .A(n3722), .B(n3691), .C(n3670), .D(A[17]), .Y(n3609) );
  MUX2IX1 U2375 ( .D0(n3610), .D1(n3611), .S(n3669), .Y(n3608) );
  NAND2X1 U2376 ( .A(n3612), .B(n3745), .Y(n3611) );
  MUX2X1 U2377 ( .D0(n3455), .D1(n3456), .S(n3681), .Y(n3436) );
  NOR4XL U2378 ( .A(n3722), .B(n3691), .C(n3671), .D(A[20]), .Y(n3456) );
  MUX2IX1 U2379 ( .D0(n3457), .D1(n3458), .S(n3669), .Y(n3455) );
  NAND2X1 U2380 ( .A(n3459), .B(n3745), .Y(n3458) );
  MUX2X1 U2381 ( .D0(n3661), .D1(n3662), .S(n3680), .Y(n3642) );
  NOR4XL U2382 ( .A(n3723), .B(n3691), .C(n3671), .D(A[16]), .Y(n3662) );
  MUX2IX1 U2383 ( .D0(n3663), .D1(n3664), .S(n3669), .Y(n3661) );
  NAND2X1 U2384 ( .A(n3665), .B(n3739), .Y(n3664) );
  MUX2X1 U2385 ( .D0(n3505), .D1(n3506), .S(n3680), .Y(n3486) );
  NOR4XL U2386 ( .A(n3722), .B(n3691), .C(n3671), .D(A[19]), .Y(n3506) );
  MUX2IX1 U2387 ( .D0(n3507), .D1(n3508), .S(n3669), .Y(n3505) );
  NAND2X1 U2388 ( .A(n3509), .B(n3739), .Y(n3508) );
  MUX2X1 U2389 ( .D0(n3555), .D1(n3556), .S(n3680), .Y(n3536) );
  NOR4XL U2390 ( .A(n3722), .B(n3691), .C(n3671), .D(A[18]), .Y(n3556) );
  MUX2IX1 U2391 ( .D0(n3557), .D1(n3558), .S(n3669), .Y(n3555) );
  NAND2X1 U2392 ( .A(n3559), .B(n3745), .Y(n3558) );
  MUX2IX1 U2393 ( .D0(A[8]), .D1(A[264]), .S(n3690), .Y(n3665) );
  NAND2X1 U2394 ( .A(n3666), .B(n3745), .Y(n3663) );
  MUX2IX1 U2395 ( .D0(A[0]), .D1(A[256]), .S(n3684), .Y(n3666) );
  NAND2X1 U2396 ( .A(n3410), .B(n3739), .Y(n3407) );
  MUX2IX1 U2397 ( .D0(A[5]), .D1(A[261]), .S(n3686), .Y(n3410) );
  NAND2X1 U2398 ( .A(n3613), .B(n3739), .Y(n3610) );
  MUX2IX1 U2399 ( .D0(A[1]), .D1(A[257]), .S(n3688), .Y(n3613) );
  NAND2X1 U2400 ( .A(n3460), .B(n3739), .Y(n3457) );
  MUX2IX1 U2401 ( .D0(A[4]), .D1(A[260]), .S(n3685), .Y(n3460) );
  NAND2X1 U2402 ( .A(n3510), .B(n3745), .Y(n3507) );
  MUX2IX1 U2403 ( .D0(A[3]), .D1(A[259]), .S(n3684), .Y(n3510) );
  NAND2X1 U2404 ( .A(n3560), .B(n3745), .Y(n3557) );
  MUX2IX1 U2405 ( .D0(A[2]), .D1(A[258]), .S(n3685), .Y(n3560) );
  MUX2IX1 U2406 ( .D0(A[6]), .D1(A[262]), .S(n3688), .Y(n3360) );
  NAND2X1 U2407 ( .A(n3359), .B(n3739), .Y(n3358) );
  MUX2IX1 U2408 ( .D0(A[14]), .D1(A[270]), .S(n3688), .Y(n3359) );
  MUX2X1 U2409 ( .D0(n3355), .D1(n3356), .S(n3681), .Y(n3336) );
  NOR4XL U2410 ( .A(n3722), .B(n3691), .C(n3670), .D(A[22]), .Y(n3356) );
  MUX2IX1 U2411 ( .D0(n3357), .D1(n3358), .S(n3669), .Y(n3355) );
  NAND2X1 U2412 ( .A(n3360), .B(n3745), .Y(n3357) );
  MUX2IX1 U2413 ( .D0(A[135]), .D1(A[391]), .S(n3690), .Y(n3287) );
  MUX2IX1 U2414 ( .D0(A[143]), .D1(A[399]), .S(n3690), .Y(n3285) );
  MUX4X1 U2415 ( .D0(n3297), .D1(n3298), .D2(n3299), .D3(n3300), .S0(n3677), 
        .S1(n3672), .Y(n3290) );
  NOR3XL U2416 ( .A(A[47]), .B(n3728), .C(n3697), .Y(n3299) );
  NOR3XL U2417 ( .A(A[63]), .B(n3728), .C(n3697), .Y(n3300) );
  NOR3XL U2418 ( .A(A[39]), .B(n3729), .C(n3697), .Y(n3297) );
  MUX4X1 U2419 ( .D0(n3281), .D1(n3282), .D2(n3283), .D3(n3284), .S0(n3677), 
        .S1(n3673), .Y(n3266) );
  NOR3XL U2420 ( .A(A[159]), .B(n3728), .C(n3697), .Y(n3284) );
  NOR21XL U2421 ( .B(n3285), .A(n3718), .Y(n3283) );
  NOR21XL U2422 ( .B(n3287), .A(n3719), .Y(n3281) );
  MUX4X1 U2423 ( .D0(n3635), .D1(n3636), .D2(n3637), .D3(n3638), .S0(n3677), 
        .S1(n3674), .Y(n3616) );
  NOR3XL U2424 ( .A(A[152]), .B(n3726), .C(n3714), .Y(n3638) );
  NOR21XL U2425 ( .B(n3639), .A(n3719), .Y(n3637) );
  NOR21XL U2426 ( .B(n3640), .A(n3719), .Y(n3636) );
  MUX4X1 U2427 ( .D0(n3270), .D1(n3271), .D2(n3272), .D3(n3273), .S0(n3677), 
        .S1(n3674), .Y(n3269) );
  NOR3XL U2428 ( .A(A[239]), .B(n3732), .C(n3694), .Y(n3272) );
  NOR3XL U2429 ( .A(A[255]), .B(n3725), .C(n3694), .Y(n3273) );
  NOR3XL U2430 ( .A(A[231]), .B(n3728), .C(n3698), .Y(n3270) );
  NOR21XL U2431 ( .B(n3641), .A(n3719), .Y(n3635) );
  MUX2IX1 U2432 ( .D0(A[128]), .D1(A[384]), .S(n3690), .Y(n3641) );
  NOR21XL U2433 ( .B(n3286), .A(n3718), .Y(n3282) );
  MUX2IX1 U2434 ( .D0(A[151]), .D1(A[407]), .S(n3689), .Y(n3286) );
  NOR3XL U2435 ( .A(A[247]), .B(n3727), .C(n3698), .Y(n3271) );
  NOR3XL U2436 ( .A(A[55]), .B(n3729), .C(n3697), .Y(n3298) );
  INVX1 U2437 ( .A(SH[8]), .Y(n3715) );
  MUX4X1 U2438 ( .D0(n3274), .D1(n3275), .D2(n3276), .D3(n3277), .S0(n3677), 
        .S1(n3674), .Y(n3268) );
  AOI21X1 U2439 ( .B(A[207]), .C(n3709), .A(n3736), .Y(n3276) );
  AOI21X1 U2440 ( .B(A[199]), .C(n3709), .A(n3736), .Y(n3274) );
  AOI21X1 U2441 ( .B(A[215]), .C(n3709), .A(n3736), .Y(n3275) );
  INVX1 U2442 ( .A(n3683), .Y(n3677) );
  INVX1 U2443 ( .A(SH[4]), .Y(n3683) );
  AOI211X1 U2444 ( .C(n3675), .D(A[191]), .A(n3735), .B(n3698), .Y(n3280) );
  NOR3XL U2445 ( .A(A[167]), .B(n3728), .C(n3698), .Y(n3278) );
  NOR3XL U2446 ( .A(A[223]), .B(n3728), .C(n3698), .Y(n3277) );
  INVX1 U2447 ( .A(n3717), .Y(n3710) );
  INVX1 U2448 ( .A(SH[8]), .Y(n3717) );
  INVX1 U2449 ( .A(SH[9]), .Y(n3745) );
  INVX1 U2450 ( .A(SH[8]), .Y(n3716) );
  MUX2IX1 U2451 ( .D0(A[129]), .D1(A[385]), .S(n3687), .Y(n3588) );
  MUX2IX1 U2452 ( .D0(A[137]), .D1(A[393]), .S(n3686), .Y(n3586) );
  MUX2IX1 U2453 ( .D0(A[193]), .D1(A[449]), .S(n3686), .Y(n3577) );
  MUX2IX1 U2454 ( .D0(A[201]), .D1(A[457]), .S(n3686), .Y(n3575) );
  MUX2IX1 U2455 ( .D0(A[144]), .D1(A[400]), .S(n3690), .Y(n3640) );
  MUX2IX1 U2456 ( .D0(A[130]), .D1(A[386]), .S(n3684), .Y(n3535) );
  MUX2IX1 U2457 ( .D0(A[138]), .D1(A[394]), .S(n3684), .Y(n3533) );
  MUX4X1 U2458 ( .D0(n3571), .D1(n3572), .D2(n3573), .D3(n3574), .S0(n3679), 
        .S1(SH[3]), .Y(n3565) );
  NOR3XL U2459 ( .A(A[217]), .B(n3742), .C(SH[8]), .Y(n3574) );
  NOR21XL U2460 ( .B(n3575), .A(n3744), .Y(n3573) );
  NOR21XL U2461 ( .B(n3577), .A(n3720), .Y(n3571) );
  MUX4X1 U2462 ( .D0(n3582), .D1(n3583), .D2(n3584), .D3(n3585), .S0(n3679), 
        .S1(n3675), .Y(n3563) );
  NOR3XL U2463 ( .A(A[153]), .B(n3741), .C(n3693), .Y(n3585) );
  NOR21XL U2464 ( .B(n3586), .A(n3721), .Y(n3584) );
  NOR21XL U2465 ( .B(n3588), .A(n3744), .Y(n3582) );
  MUX4X1 U2466 ( .D0(n3479), .D1(n3480), .D2(n3481), .D3(n3482), .S0(n3679), 
        .S1(n3673), .Y(n3463) );
  NOR3XL U2467 ( .A(A[155]), .B(n3744), .C(n3698), .Y(n3482) );
  NOR21XL U2468 ( .B(n3483), .A(n3718), .Y(n3481) );
  NOR21XL U2469 ( .B(n3485), .A(n3718), .Y(n3479) );
  MUX4X1 U2470 ( .D0(n3529), .D1(n3530), .D2(n3531), .D3(n3532), .S0(n3680), 
        .S1(n3675), .Y(n3513) );
  NOR3XL U2471 ( .A(A[154]), .B(n3724), .C(n3693), .Y(n3532) );
  NOR21XL U2472 ( .B(n3533), .A(n3721), .Y(n3531) );
  NOR21XL U2473 ( .B(n3535), .A(n3744), .Y(n3529) );
  NOR21XL U2474 ( .B(n3587), .A(n3719), .Y(n3583) );
  MUX2IX1 U2475 ( .D0(A[145]), .D1(A[401]), .S(n3687), .Y(n3587) );
  NOR21XL U2476 ( .B(n3576), .A(n3744), .Y(n3572) );
  MUX2IX1 U2477 ( .D0(A[209]), .D1(A[465]), .S(n3686), .Y(n3576) );
  NOR21XL U2478 ( .B(n3484), .A(n3718), .Y(n3480) );
  MUX2IX1 U2479 ( .D0(A[147]), .D1(A[403]), .S(n3685), .Y(n3484) );
  NOR21XL U2480 ( .B(n3534), .A(n3722), .Y(n3530) );
  MUX2IX1 U2481 ( .D0(A[146]), .D1(A[402]), .S(n3684), .Y(n3534) );
  INVX1 U2482 ( .A(SH[3]), .Y(n3676) );
  MUX2IX1 U2483 ( .D0(A[133]), .D1(A[389]), .S(n3687), .Y(n3385) );
  MUX2IX1 U2484 ( .D0(A[141]), .D1(A[397]), .S(n3687), .Y(n3383) );
  MUX2IX1 U2485 ( .D0(A[132]), .D1(A[388]), .S(n3686), .Y(n3435) );
  MUX2IX1 U2486 ( .D0(A[140]), .D1(A[396]), .S(n3686), .Y(n3433) );
  MUX2IX1 U2487 ( .D0(A[134]), .D1(A[390]), .S(n3688), .Y(n3335) );
  MUX2IX1 U2488 ( .D0(A[142]), .D1(A[398]), .S(n3689), .Y(n3333) );
  MUX2IX1 U2489 ( .D0(A[136]), .D1(A[392]), .S(n3690), .Y(n3639) );
  MUX2IX1 U2490 ( .D0(A[192]), .D1(A[448]), .S(n3690), .Y(n3630) );
  MUX2IX1 U2491 ( .D0(A[200]), .D1(A[456]), .S(n3688), .Y(n3628) );
  MUX2IX1 U2492 ( .D0(A[131]), .D1(A[387]), .S(n3684), .Y(n3485) );
  MUX2IX1 U2493 ( .D0(A[139]), .D1(A[395]), .S(n3685), .Y(n3483) );
  NOR21XL U2494 ( .B(n3334), .A(n3720), .Y(n3330) );
  MUX2IX1 U2495 ( .D0(A[150]), .D1(A[406]), .S(n3689), .Y(n3334) );
  MUX4X1 U2496 ( .D0(n3395), .D1(n3396), .D2(n3397), .D3(n3398), .S0(SH[4]), 
        .S1(n3672), .Y(n3388) );
  NOR3XL U2497 ( .A(A[45]), .B(n3732), .C(n3710), .Y(n3397) );
  NOR3XL U2498 ( .A(A[61]), .B(n3732), .C(n3710), .Y(n3398) );
  NOR3XL U2499 ( .A(A[37]), .B(n3732), .C(n3710), .Y(n3395) );
  MUX4X1 U2500 ( .D0(n3598), .D1(n3599), .D2(n3600), .D3(n3601), .S0(n3682), 
        .S1(n3674), .Y(n3591) );
  NOR3XL U2501 ( .A(A[41]), .B(SH[9]), .C(n3692), .Y(n3600) );
  NOR3XL U2502 ( .A(A[57]), .B(SH[9]), .C(n3713), .Y(n3601) );
  NOR3XL U2503 ( .A(A[49]), .B(SH[9]), .C(n3692), .Y(n3599) );
  MUX4X1 U2504 ( .D0(n3445), .D1(n3446), .D2(n3447), .D3(n3448), .S0(SH[4]), 
        .S1(n3672), .Y(n3438) );
  NOR3XL U2505 ( .A(A[44]), .B(n3734), .C(n3695), .Y(n3447) );
  NOR3XL U2506 ( .A(A[60]), .B(n3733), .C(n3695), .Y(n3448) );
  NOR3XL U2507 ( .A(A[36]), .B(n3734), .C(n3695), .Y(n3445) );
  MUX4X1 U2508 ( .D0(n3345), .D1(n3346), .D2(n3347), .D3(n3348), .S0(n3678), 
        .S1(n3671), .Y(n3338) );
  NOR3XL U2509 ( .A(A[46]), .B(n3730), .C(n3696), .Y(n3347) );
  NOR3XL U2510 ( .A(A[62]), .B(n3730), .C(n3696), .Y(n3348) );
  NOR3XL U2511 ( .A(A[38]), .B(n3730), .C(n3696), .Y(n3345) );
  MUX4X1 U2512 ( .D0(n3323), .D1(n3324), .D2(n3325), .D3(n3326), .S0(n3677), 
        .S1(n3671), .Y(n3317) );
  AOI21X1 U2513 ( .B(A[206]), .C(n3708), .A(n3736), .Y(n3325) );
  AOI21X1 U2514 ( .B(A[198]), .C(n3708), .A(n3735), .Y(n3323) );
  AOI21X1 U2515 ( .B(A[214]), .C(n3707), .A(n3735), .Y(n3324) );
  MUX4X1 U2516 ( .D0(n3651), .D1(n3652), .D2(n3653), .D3(n3654), .S0(n3677), 
        .S1(n3674), .Y(n3644) );
  NOR3XL U2517 ( .A(A[40]), .B(n3727), .C(n3694), .Y(n3653) );
  NOR3XL U2518 ( .A(A[56]), .B(n3727), .C(n3693), .Y(n3654) );
  NOR3XL U2519 ( .A(A[32]), .B(n3727), .C(n3694), .Y(n3651) );
  MUX4X1 U2520 ( .D0(n3624), .D1(n3625), .D2(n3626), .D3(n3627), .S0(n3678), 
        .S1(n3674), .Y(n3618) );
  NOR3XL U2521 ( .A(A[216]), .B(n3726), .C(n3692), .Y(n3627) );
  NOR21XL U2522 ( .B(n3628), .A(n3720), .Y(n3626) );
  NOR21XL U2523 ( .B(n3630), .A(n3719), .Y(n3624) );
  MUX4X1 U2524 ( .D0(n3495), .D1(n3496), .D2(n3497), .D3(n3498), .S0(n3679), 
        .S1(n3673), .Y(n3488) );
  NOR3XL U2525 ( .A(A[59]), .B(n3724), .C(n3714), .Y(n3498) );
  NOR3XL U2526 ( .A(A[43]), .B(n3723), .C(n3714), .Y(n3497) );
  NOR3XL U2527 ( .A(A[35]), .B(n3723), .C(n3714), .Y(n3495) );
  MUX4X1 U2528 ( .D0(n3545), .D1(n3546), .D2(n3547), .D3(n3548), .S0(n3680), 
        .S1(SH[3]), .Y(n3538) );
  NOR3XL U2529 ( .A(A[42]), .B(n3725), .C(n3693), .Y(n3547) );
  NOR3XL U2530 ( .A(A[58]), .B(n3725), .C(n3693), .Y(n3548) );
  NOR3XL U2531 ( .A(A[34]), .B(n3725), .C(SH[8]), .Y(n3545) );
  MUX4X1 U2532 ( .D0(n3375), .D1(n3376), .D2(n3377), .D3(n3378), .S0(n3678), 
        .S1(n3671), .Y(n3364) );
  NOR3XL U2533 ( .A(A[173]), .B(n3731), .C(n3710), .Y(n3377) );
  NOR3XL U2534 ( .A(A[189]), .B(n3731), .C(n3710), .Y(n3378) );
  NOR3XL U2535 ( .A(A[165]), .B(n3731), .C(n3711), .Y(n3375) );
  MUX4X1 U2536 ( .D0(n3578), .D1(n3579), .D2(n3580), .D3(n3581), .S0(n3679), 
        .S1(n3675), .Y(n3564) );
  NOR3XL U2537 ( .A(A[169]), .B(n3742), .C(n3692), .Y(n3580) );
  NOR3XL U2538 ( .A(A[185]), .B(n3743), .C(SH[8]), .Y(n3581) );
  NOR3XL U2539 ( .A(A[161]), .B(n3743), .C(n3692), .Y(n3578) );
  MUX4X1 U2540 ( .D0(n3425), .D1(n3426), .D2(n3427), .D3(n3428), .S0(n3682), 
        .S1(n3672), .Y(n3414) );
  NOR3XL U2541 ( .A(A[172]), .B(n3733), .C(n3712), .Y(n3427) );
  NOR3XL U2542 ( .A(A[188]), .B(n3733), .C(n3712), .Y(n3428) );
  NOR3XL U2543 ( .A(A[164]), .B(n3733), .C(n3712), .Y(n3425) );
  MUX4X1 U2544 ( .D0(n3631), .D1(n3632), .D2(n3633), .D3(n3634), .S0(n3678), 
        .S1(n3674), .Y(n3617) );
  NOR3XL U2545 ( .A(A[168]), .B(n3726), .C(n3693), .Y(n3633) );
  NOR3XL U2546 ( .A(A[184]), .B(n3726), .C(n3692), .Y(n3634) );
  NOR3XL U2547 ( .A(A[160]), .B(n3726), .C(n3692), .Y(n3631) );
  MUX4X1 U2548 ( .D0(n3475), .D1(n3476), .D2(n3477), .D3(n3478), .S0(n3679), 
        .S1(n3673), .Y(n3464) );
  NOR3XL U2549 ( .A(A[171]), .B(n3734), .C(n3698), .Y(n3477) );
  NOR3XL U2550 ( .A(A[187]), .B(n3734), .C(n3695), .Y(n3478) );
  NOR3XL U2551 ( .A(A[163]), .B(n3734), .C(n3698), .Y(n3475) );
  MUX4X1 U2552 ( .D0(n3525), .D1(n3526), .D2(n3527), .D3(n3528), .S0(n3679), 
        .S1(n3675), .Y(n3514) );
  NOR3XL U2553 ( .A(A[170]), .B(n3724), .C(n3694), .Y(n3527) );
  NOR3XL U2554 ( .A(A[186]), .B(n3724), .C(n3693), .Y(n3528) );
  NOR3XL U2555 ( .A(A[162]), .B(n3724), .C(n3694), .Y(n3525) );
  MUX4X1 U2556 ( .D0(n3379), .D1(n3380), .D2(n3381), .D3(n3382), .S0(n3678), 
        .S1(n3672), .Y(n3363) );
  NOR3XL U2557 ( .A(A[157]), .B(n3731), .C(n3711), .Y(n3382) );
  NOR21XL U2558 ( .B(n3383), .A(n3743), .Y(n3381) );
  NOR21XL U2559 ( .B(n3385), .A(n3743), .Y(n3379) );
  MUX4X1 U2560 ( .D0(n3429), .D1(n3430), .D2(n3431), .D3(n3432), .S0(n3682), 
        .S1(n3672), .Y(n3413) );
  NOR3XL U2561 ( .A(A[156]), .B(n3733), .C(n3711), .Y(n3432) );
  NOR21XL U2562 ( .B(n3433), .A(n3721), .Y(n3431) );
  NOR21XL U2563 ( .B(n3435), .A(n3743), .Y(n3429) );
  MUX4X1 U2564 ( .D0(n3329), .D1(n3330), .D2(n3331), .D3(n3332), .S0(n3678), 
        .S1(n3671), .Y(n3315) );
  NOR3XL U2565 ( .A(A[158]), .B(n3729), .C(n3696), .Y(n3332) );
  NOR21XL U2566 ( .B(n3333), .A(n3721), .Y(n3331) );
  NOR21XL U2567 ( .B(n3335), .A(n3721), .Y(n3329) );
  MUX4X1 U2568 ( .D0(n3367), .D1(n3368), .D2(n3369), .D3(n3370), .S0(n3678), 
        .S1(n3671), .Y(n3366) );
  NOR3XL U2569 ( .A(A[237]), .B(n3731), .C(n3696), .Y(n3369) );
  NOR3XL U2570 ( .A(A[253]), .B(n3730), .C(n3696), .Y(n3370) );
  NOR3XL U2571 ( .A(A[229]), .B(n3731), .C(n3696), .Y(n3367) );
  MUX4X1 U2572 ( .D0(n3417), .D1(n3418), .D2(n3419), .D3(n3420), .S0(n3682), 
        .S1(n3672), .Y(n3416) );
  NOR3XL U2573 ( .A(A[236]), .B(n3733), .C(n3711), .Y(n3419) );
  NOR3XL U2574 ( .A(A[252]), .B(n3732), .C(n3711), .Y(n3420) );
  NOR3XL U2575 ( .A(A[228]), .B(n3733), .C(n3711), .Y(n3417) );
  MUX4X1 U2576 ( .D0(n3319), .D1(n3320), .D2(n3321), .D3(n3322), .S0(n3677), 
        .S1(n3672), .Y(n3318) );
  NOR3XL U2577 ( .A(A[238]), .B(n3729), .C(n3697), .Y(n3321) );
  NOR3XL U2578 ( .A(A[254]), .B(n3729), .C(n3697), .Y(n3322) );
  NOR3XL U2579 ( .A(A[230]), .B(n3729), .C(n3696), .Y(n3319) );
  MUX4X1 U2580 ( .D0(n3467), .D1(n3468), .D2(n3469), .D3(n3470), .S0(n3679), 
        .S1(n3673), .Y(n3466) );
  NOR3XL U2581 ( .A(A[235]), .B(n3742), .C(n3695), .Y(n3469) );
  NOR3XL U2582 ( .A(A[251]), .B(n3742), .C(n3695), .Y(n3470) );
  NOR3XL U2583 ( .A(A[227]), .B(n3734), .C(n3695), .Y(n3467) );
  MUX4X1 U2584 ( .D0(n3517), .D1(n3518), .D2(n3519), .D3(n3520), .S0(n3680), 
        .S1(n3675), .Y(n3516) );
  NOR3XL U2585 ( .A(A[250]), .B(n3724), .C(n3714), .Y(n3520) );
  NOR3XL U2586 ( .A(A[234]), .B(n3723), .C(n3714), .Y(n3519) );
  NOR3XL U2587 ( .A(A[226]), .B(n3724), .C(n3694), .Y(n3517) );
  NOR21XL U2588 ( .B(n3384), .A(n3744), .Y(n3380) );
  MUX2IX1 U2589 ( .D0(A[149]), .D1(A[405]), .S(n3687), .Y(n3384) );
  NOR21XL U2590 ( .B(n3434), .A(n3744), .Y(n3430) );
  MUX2IX1 U2591 ( .D0(A[148]), .D1(A[404]), .S(n3686), .Y(n3434) );
  NOR21XL U2592 ( .B(n3629), .A(n3719), .Y(n3625) );
  MUX2IX1 U2593 ( .D0(A[208]), .D1(A[464]), .S(n3689), .Y(n3629) );
  AOI21X1 U2594 ( .B(A[205]), .C(n3707), .A(n3736), .Y(n3373) );
  AOI21X1 U2595 ( .B(A[204]), .C(n3706), .A(n3735), .Y(n3423) );
  AOI21X1 U2596 ( .B(A[203]), .C(n3705), .A(n3736), .Y(n3473) );
  AOI21X1 U2597 ( .B(A[202]), .C(n3704), .A(n3736), .Y(n3523) );
  AOI21X1 U2598 ( .B(A[213]), .C(n3707), .A(n3735), .Y(n3372) );
  AOI21X1 U2599 ( .B(A[212]), .C(n3708), .A(n3735), .Y(n3422) );
  AOI21X1 U2600 ( .B(A[211]), .C(n3709), .A(n3736), .Y(n3472) );
  AOI21X1 U2601 ( .B(A[210]), .C(n3708), .A(n3735), .Y(n3522) );
  AOI21X1 U2602 ( .B(A[197]), .C(n3705), .A(n3735), .Y(n3371) );
  AOI21X1 U2603 ( .B(A[196]), .C(n3703), .A(n3735), .Y(n3421) );
  AOI21X1 U2604 ( .B(A[195]), .C(n3708), .A(n3736), .Y(n3471) );
  AOI21X1 U2605 ( .B(A[194]), .C(n3705), .A(n3735), .Y(n3521) );
  NOR3XL U2606 ( .A(A[48]), .B(n3727), .C(n3693), .Y(n3652) );
  NOR3XL U2607 ( .A(A[240]), .B(n3726), .C(n3714), .Y(n3621) );
  NOR3XL U2608 ( .A(A[246]), .B(n3729), .C(n3697), .Y(n3320) );
  NOR3XL U2609 ( .A(A[221]), .B(n3731), .C(n3710), .Y(n3374) );
  NOR3XL U2610 ( .A(A[220]), .B(n3733), .C(n3711), .Y(n3424) );
  NOR3XL U2611 ( .A(A[244]), .B(n3733), .C(n3712), .Y(n3418) );
  NOR3XL U2612 ( .A(A[222]), .B(n3729), .C(n3697), .Y(n3326) );
  NOR3XL U2613 ( .A(A[243]), .B(n3744), .C(n3695), .Y(n3468) );
  NOR3XL U2614 ( .A(A[242]), .B(n3723), .C(n3694), .Y(n3518) );
  NOR3XL U2615 ( .A(A[233]), .B(n3727), .C(n3713), .Y(n3569) );
  NOR3XL U2616 ( .A(A[232]), .B(n3726), .C(n3693), .Y(n3622) );
  NOR3XL U2617 ( .A(A[53]), .B(n3732), .C(n3711), .Y(n3396) );
  NOR3XL U2618 ( .A(A[245]), .B(n3731), .C(n3696), .Y(n3368) );
  NOR3XL U2619 ( .A(A[241]), .B(n3743), .C(SH[8]), .Y(n3568) );
  NOR3XL U2620 ( .A(A[52]), .B(n3741), .C(n3695), .Y(n3446) );
  NOR3XL U2621 ( .A(A[54]), .B(n3730), .C(n3696), .Y(n3346) );
  NOR3XL U2622 ( .A(A[51]), .B(n3723), .C(n3714), .Y(n3496) );
  NOR3XL U2623 ( .A(A[50]), .B(n3725), .C(n3693), .Y(n3546) );
  NOR3XL U2624 ( .A(A[181]), .B(n3731), .C(n3710), .Y(n3376) );
  NOR3XL U2625 ( .A(A[177]), .B(n3743), .C(SH[8]), .Y(n3579) );
  NOR3XL U2626 ( .A(A[180]), .B(n3733), .C(n3712), .Y(n3426) );
  NOR3XL U2627 ( .A(A[176]), .B(n3726), .C(n3692), .Y(n3632) );
  NOR3XL U2628 ( .A(A[179]), .B(n3734), .C(n3711), .Y(n3476) );
  NOR3XL U2629 ( .A(A[178]), .B(n3725), .C(n3694), .Y(n3526) );
  NOR3XL U2630 ( .A(A[224]), .B(n3726), .C(n3692), .Y(n3620) );
  NOR3XL U2631 ( .A(A[33]), .B(SH[9]), .C(n3691), .Y(n3598) );
  NOR3XL U2632 ( .A(A[225]), .B(n3743), .C(n3692), .Y(n3567) );
  NOR3XL U2633 ( .A(A[249]), .B(n3742), .C(SH[8]), .Y(n3570) );
  NOR3XL U2634 ( .A(A[248]), .B(n3726), .C(n3691), .Y(n3623) );
  NOR3XL U2635 ( .A(A[219]), .B(n3742), .C(n3695), .Y(n3474) );
  NOR3XL U2636 ( .A(A[218]), .B(n3724), .C(n3694), .Y(n3524) );
  AOI211X1 U2637 ( .C(A[166]), .D(n3676), .A(n3734), .B(n3698), .Y(n3327) );
  AOI211X1 U2638 ( .C(n3675), .D(A[190]), .A(n3734), .B(n3698), .Y(n3328) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regx_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N16, N17, N18, N19, N20,
         net9014, n12, n3, n4, n5, n6, n7, n8, n9, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9014), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N20), .SIN(db_cnt_2_), .SMC(test_se), .C(net9014), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N18), .SIN(db_cnt_0_), .SMC(test_se), .C(net9014), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N17), .SIN(o_dbc), .SMC(test_se), .C(net9014), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N19), .SIN(db_cnt_1_), .SMC(test_se), .C(net9014), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n12), .SIN(d_org_0_), .SMC(test_se), .C(net9014), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n6), .Y(n1) );
  NOR21XL U4 ( .B(n3), .A(n4), .Y(n6) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  OAI22X1 U6 ( .A(db_cnt_2_), .B(n5), .C(n7), .D(n2), .Y(N19) );
  AOI21BBXL U7 ( .B(n1), .C(db_cnt_1_), .A(N17), .Y(n7) );
  AO22AXL U8 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR2X1 U9 ( .A(n3), .B(n4), .Y(o_chg) );
  NOR2X1 U10 ( .A(n1), .B(db_cnt_0_), .Y(N17) );
  NAND4X1 U11 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(db_cnt_0_), .Y(
        n3) );
  NAND3X1 U12 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(n6), .Y(n5) );
  ENOX1 U13 ( .A(n2), .B(n5), .C(test_so), .D(n6), .Y(N20) );
  NOR2X1 U14 ( .A(n8), .B(n1), .Y(N18) );
  XNOR2XL U15 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n8) );
  NAND31X1 U16 ( .C(db_cnt_0_), .A(n4), .B(n9), .Y(N16) );
  NOR3XL U17 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n9) );
  INVX1 U18 ( .A(db_cnt_2_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N16, N17, N18, N19, N20,
         net9032, n12, n3, n4, n5, n6, n7, n8, n9, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9032), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N20), .SIN(db_cnt_2_), .SMC(test_se), .C(net9032), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N18), .SIN(db_cnt_0_), .SMC(test_se), .C(net9032), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N17), .SIN(o_dbc), .SMC(test_se), .C(net9032), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N19), .SIN(db_cnt_1_), .SMC(test_se), .C(net9032), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n12), .SIN(d_org_0_), .SMC(test_se), .C(net9032), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n6), .Y(n1) );
  NOR21XL U4 ( .B(n3), .A(n4), .Y(n6) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  OAI22X1 U6 ( .A(db_cnt_2_), .B(n5), .C(n7), .D(n2), .Y(N19) );
  AOI21BBXL U7 ( .B(n1), .C(db_cnt_1_), .A(N17), .Y(n7) );
  AO22AXL U8 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR2X1 U9 ( .A(n3), .B(n4), .Y(o_chg) );
  NOR2X1 U10 ( .A(n1), .B(db_cnt_0_), .Y(N17) );
  NAND4X1 U11 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(db_cnt_0_), .Y(
        n3) );
  NAND3X1 U12 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(n6), .Y(n5) );
  ENOX1 U13 ( .A(n2), .B(n5), .C(test_so), .D(n6), .Y(N20) );
  NOR2X1 U14 ( .A(n8), .B(n1), .Y(N18) );
  XNOR2XL U15 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n8) );
  NAND31X1 U16 ( .C(db_cnt_0_), .A(n4), .B(n9), .Y(N16) );
  NOR3XL U17 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n9) );
  INVX1 U18 ( .A(db_cnt_2_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N16, N17, N18, N19, N20,
         net9050, n12, n3, n4, n5, n6, n7, n8, n9, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_2 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9050), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N20), .SIN(db_cnt_2_), .SMC(test_se), .C(net9050), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N18), .SIN(db_cnt_0_), .SMC(test_se), .C(net9050), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N17), .SIN(o_dbc), .SMC(test_se), .C(net9050), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N19), .SIN(db_cnt_1_), .SMC(test_se), .C(net9050), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n12), .SIN(d_org_0_), .SMC(test_se), .C(net9050), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n6), .Y(n1) );
  NOR21XL U4 ( .B(n3), .A(n4), .Y(n6) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  OAI22X1 U6 ( .A(db_cnt_2_), .B(n5), .C(n7), .D(n2), .Y(N19) );
  AOI21BBXL U7 ( .B(n1), .C(db_cnt_1_), .A(N17), .Y(n7) );
  AO22AXL U8 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR2X1 U9 ( .A(n3), .B(n4), .Y(o_chg) );
  NOR2X1 U10 ( .A(n1), .B(db_cnt_0_), .Y(N17) );
  NAND4X1 U11 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(db_cnt_0_), .Y(
        n3) );
  NAND3X1 U12 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(n6), .Y(n5) );
  ENOX1 U13 ( .A(n2), .B(n5), .C(test_so), .D(n6), .Y(N20) );
  NOR2X1 U14 ( .A(n8), .B(n1), .Y(N18) );
  XNOR2XL U15 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n8) );
  NAND31X1 U16 ( .C(db_cnt_0_), .A(n4), .B(n9), .Y(N16) );
  NOR3XL U17 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n9) );
  INVX1 U18 ( .A(db_cnt_2_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_4 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_5 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_6 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module glreg_a0_7 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9068;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_7 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9068), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9068), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9068), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9068), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9068), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9068), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9068), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9068), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9068), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_8 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9086;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_8 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9086), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9086), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9086), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9086), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9086), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9086), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9086), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9086), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9086), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_9 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9104;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_9 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9104), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9104), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9104), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9104), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9104), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9104), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9104), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9104), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9104), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH7_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9122;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9122), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9122), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9122), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9122), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9122), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9122), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9122), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9122), 
        .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_7 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module glreg_a0_10 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9140;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_10 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9140), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9140), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9140), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9140), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9140), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9140), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9140), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9140), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9140), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_11 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9158;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_11 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9158), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9158), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9158), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9158), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9158), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9158), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9158), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9158), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9158), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_12 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9176;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_12 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9176), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9176), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9176), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9176), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9176), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9176), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9176), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9176), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9176), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_13 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9194;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_13 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9194), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9194), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9194), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9194), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9194), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9194), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9194), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9194), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9194), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_14 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9212;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_14 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9212), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9212), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9212), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9212), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9212), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9212), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9212), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9212), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9212), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9230;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9230), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9230), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9230), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9230), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9230), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9230), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9230), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9248;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9248), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9248), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9248), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9248), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9248), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9248), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9248), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_15 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9266;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_15 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9266), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9266), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9266), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9266), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9266), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9266), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9266), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9266), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9266), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_6_00000002 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9284;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9284), .TE(test_se) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9284), 
        .XS(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9284), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9284), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9284), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9284), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9284), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_a0_16 ( clk, arstz, we, wdat, rdat, test_si2, test_si1, test_se
 );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si2, test_si1, test_se;
  wire   net9302;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_16 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9302), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9302), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9302), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9302), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9302), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9302), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9302), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si1), .SMC(test_se), .C(net9302), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(test_si2), .SMC(test_se), .C(net9302), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_17 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9320;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_17 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9320), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9320), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9320), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9320), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9320), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9320), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9320), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9320), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9320), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_18 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9338;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_18 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9338), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9338), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9338), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9338), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9338), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9338), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9338), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9338), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9338), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_19 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9356;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_19 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9356), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9356), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9356), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9356), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9356), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9356), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9356), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9356), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9356), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module cvctl_a0 ( r_cvcwr, wdat, r_sdischg, r_vcomp, r_idacsh, r_cvofsx, 
        r_cvofs, sdischg_duty, r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, 
        r_fw_pwrv, r_dac0, r_dac3, clk_100k, clk, srstz, test_si, test_se );
  input [5:0] r_cvcwr;
  input [7:0] wdat;
  output [7:0] r_sdischg;
  output [7:0] r_vcomp;
  output [7:0] r_idacsh;
  output [7:0] r_cvofsx;
  output [15:0] r_cvofs;
  input [11:0] r_fw_pwrv;
  output [10:0] r_dac0;
  output [5:0] r_dac3;
  input r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, clk_100k, clk, srstz,
         test_si, test_se;
  output sdischg_duty;
  wire   clk_5k, N29, N34, N35, N36, N38, N39, N40, N41, N42, N47, N84, N94,
         N95, N96, N97, N98, N99, N106, N107, N108, N109, N115, N121, N122,
         N123, N126, N127, N128, N129, N130, net9374, n81, N68, N67, N66, N65,
         N64, N63, N62, N61, N60, n2, n4, n5, n6, n7, n8, n9, N83, N82, N81,
         N80, N79, N78, N77, N76, N75, N74, N73, N72, N59, N58, N57, N56, N55,
         N54, N53, N52, N51, N50, N49, N48, n34, n35, n36, n37, n38, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, add_62_carry_1_, add_62_carry_2_, add_62_carry_3_,
         add_62_carry_4_, add_62_carry_5_, n3, n12, n17, n18, n19, n20, n21,
         n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33;
  wire   [4:0] div20_cnt;
  wire   [10:1] cv_code;
  wire   [4:0] sdischg_cnt;
  wire   [4:2] add_81_carry;
  wire   [4:2] add_41_carry;
  wire   [2:1] add_3_root_sub_0_root_add_46_3_carry;

  HAD1X1 add_81_U1_1_1 ( .A(sdischg_cnt[1]), .B(sdischg_cnt[0]), .CO(
        add_81_carry[2]), .SO(N121) );
  HAD1X1 add_81_U1_1_2 ( .A(sdischg_cnt[2]), .B(add_81_carry[2]), .CO(
        add_81_carry[3]), .SO(N122) );
  HAD1X1 add_81_U1_1_3 ( .A(sdischg_cnt[3]), .B(add_81_carry[3]), .CO(
        add_81_carry[4]), .SO(N123) );
  HAD1X1 add_41_U1_1_1 ( .A(div20_cnt[1]), .B(div20_cnt[0]), .CO(
        add_41_carry[2]), .SO(N34) );
  HAD1X1 add_41_U1_1_2 ( .A(div20_cnt[2]), .B(add_41_carry[2]), .CO(
        add_41_carry[3]), .SO(N35) );
  HAD1X1 add_41_U1_1_3 ( .A(div20_cnt[3]), .B(add_41_carry[3]), .CO(
        add_41_carry[4]), .SO(N36) );
  FAD1X1 add_3_root_sub_0_root_add_46_3_U1_1 ( .A(N47), .B(r_vcomp[1]), .CI(
        add_3_root_sub_0_root_add_46_3_carry[1]), .CO(
        add_3_root_sub_0_root_add_46_3_carry[2]), .SO(N61) );
  INVX1 U4 ( .A(n9), .Y(n8) );
  INVX1 U5 ( .A(n9), .Y(n4) );
  INVX1 U6 ( .A(n9), .Y(n5) );
  INVX1 U7 ( .A(n9), .Y(n6) );
  INVX1 U8 ( .A(n9), .Y(n7) );
  INVX1 U9 ( .A(n9), .Y(n2) );
  INVX1 U10 ( .A(srstz), .Y(n9) );
  glreg_a0_25 u0_v_comp ( .clk(clk), .arstz(n8), .we(r_cvcwr[3]), .wdat(wdat), 
        .rdat(r_vcomp), .test_si(r_sdischg[7]), .test_se(test_se) );
  glreg_a0_24 u0_idac_shift ( .clk(clk), .arstz(n7), .we(r_cvcwr[4]), .wdat(
        wdat), .rdat(r_idacsh), .test_si(r_cvofs[15]), .test_se(test_se) );
  glreg_a0_23 u0_cv_ofsx ( .clk(clk), .arstz(n6), .we(r_cvcwr[5]), .wdat(wdat), 
        .rdat(r_cvofsx), .test_si(sdischg_duty), .test_se(test_se) );
  glreg_a0_22 u0_cvofs01 ( .clk(clk), .arstz(n5), .we(r_cvcwr[0]), .wdat(wdat), 
        .rdat(r_cvofs[7:0]), .test_si(r_cvofsx[7]), .test_se(test_se) );
  glreg_a0_21 u0_cvofs23 ( .clk(clk), .arstz(n4), .we(r_cvcwr[1]), .wdat(wdat), 
        .rdat(r_cvofs[15:8]), .test_si(r_cvofs[7]), .test_se(test_se) );
  glreg_a0_20 u0_sdischg ( .clk(clk), .arstz(n2), .we(r_cvcwr[2]), .wdat(wdat), 
        .rdat(r_sdischg), .test_si(r_idacsh[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_cvctl_a0 clk_gate_sdischg_cnt_reg ( .CLK(clk_100k), 
        .EN(N115), .ENCLK(net9374), .TE(test_se) );
  cvctl_a0_DW01_sub_1 sub_2_root_sub_0_root_add_46_3 ( .A(r_fw_pwrv), .B({1'b0, 
        1'b0, 1'b0, 1'b0, r_idacsh}), .CI(1'b0), .DIFF({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .CO() );
  cvctl_a0_DW01_add_2 add_1_root_sub_0_root_add_46_3 ( .A({r_cvofsx[7], 
        r_cvofsx[7], r_cvofsx[7], r_cvofsx[7], r_cvofsx}), .B({1'b0, 1'b0, 
        1'b0, N68, N67, N66, N65, N64, N63, N62, N61, N60}), .CI(1'b0), .SUM({
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}), .CO() );
  cvctl_a0_DW01_add_1 add_0_root_sub_0_root_add_46_3 ( .A({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .B({N83, N82, N81, N80, N79, 
        N78, N77, N76, N75, N74, N73, N72}), .CI(1'b0), .SUM({N84, cv_code, 
        r_dac0[0]}), .CO() );
  FAD1X1 add_62_U1_1 ( .A(N95), .B(N107), .CI(add_62_carry_1_), .CO(
        add_62_carry_2_), .SO(r_dac3[1]) );
  FAD1X1 add_62_U1_2 ( .A(N96), .B(N108), .CI(add_62_carry_2_), .CO(
        add_62_carry_3_), .SO(r_dac3[2]) );
  FAD1X1 add_62_U1_3 ( .A(N97), .B(N109), .CI(add_62_carry_3_), .CO(
        add_62_carry_4_), .SO(r_dac3[3]) );
  SDFFRQX1 sdischg_cnt_reg_0_ ( .D(N126), .SIN(div20_cnt[4]), .SMC(test_se), 
        .C(net9374), .XR(srstz), .Q(sdischg_cnt[0]) );
  SDFFRQX1 sdischg_cnt_reg_4_ ( .D(N130), .SIN(sdischg_cnt[3]), .SMC(test_se), 
        .C(net9374), .XR(n6), .Q(sdischg_cnt[4]) );
  SDFFRQX1 sdischg_cnt_reg_1_ ( .D(N127), .SIN(sdischg_cnt[0]), .SMC(test_se), 
        .C(net9374), .XR(srstz), .Q(sdischg_cnt[1]) );
  SDFFRQX1 sdischg_cnt_reg_2_ ( .D(N128), .SIN(sdischg_cnt[1]), .SMC(test_se), 
        .C(net9374), .XR(n4), .Q(sdischg_cnt[2]) );
  SDFFRQX1 div20_cnt_reg_2_ ( .D(N40), .SIN(div20_cnt[1]), .SMC(test_se), .C(
        clk_100k), .XR(n2), .Q(div20_cnt[2]) );
  SDFFRQX1 div20_cnt_reg_1_ ( .D(N39), .SIN(div20_cnt[0]), .SMC(test_se), .C(
        clk_100k), .XR(n5), .Q(div20_cnt[1]) );
  SDFFRQX1 div20_cnt_reg_3_ ( .D(N41), .SIN(div20_cnt[2]), .SMC(test_se), .C(
        clk_100k), .XR(n4), .Q(div20_cnt[3]) );
  SDFFRQX1 div20_cnt_reg_0_ ( .D(N38), .SIN(clk_5k), .SMC(test_se), .C(
        clk_100k), .XR(n8), .Q(div20_cnt[0]) );
  SDFFRQX1 div20_cnt_reg_4_ ( .D(N42), .SIN(div20_cnt[3]), .SMC(test_se), .C(
        clk_100k), .XR(n8), .Q(div20_cnt[4]) );
  SDFFRQX1 sdischg_cnt_reg_3_ ( .D(N129), .SIN(sdischg_cnt[2]), .SMC(test_se), 
        .C(net9374), .XR(n6), .Q(sdischg_cnt[3]) );
  SDFFRQX1 sdischg_reg ( .D(n81), .SIN(sdischg_cnt[4]), .SMC(test_se), .C(
        net9374), .XR(n7), .Q(sdischg_duty) );
  SDFFRQX1 clk_5k_reg ( .D(N29), .SIN(test_si), .SMC(test_se), .C(clk_100k), 
        .XR(n5), .Q(clk_5k) );
  INVX1 U11 ( .A(N84), .Y(n3) );
  INVX1 U14 ( .A(N98), .Y(n12) );
  NOR2X1 U19 ( .A(n26), .B(n52), .Y(n50) );
  NOR2X1 U20 ( .A(n72), .B(r_dac0[10]), .Y(n75) );
  NOR2X1 U21 ( .A(n76), .B(r_dac0[9]), .Y(n73) );
  INVX1 U22 ( .A(n76), .Y(r_dac0[10]) );
  NOR2X1 U23 ( .A(n23), .B(cv_code[1]), .Y(N94) );
  NOR2X1 U24 ( .A(n51), .B(n23), .Y(N98) );
  XNOR2XL U25 ( .A(cv_code[5]), .B(n50), .Y(n51) );
  NAND2X1 U26 ( .A(n25), .B(n3), .Y(r_dac0[6]) );
  NAND2X1 U27 ( .A(n28), .B(n23), .Y(r_dac0[1]) );
  NAND2X1 U28 ( .A(n27), .B(n23), .Y(r_dac0[2]) );
  NAND2X1 U29 ( .A(n26), .B(n3), .Y(r_dac0[4]) );
  INVX1 U30 ( .A(cv_code[6]), .Y(n25) );
  INVX1 U31 ( .A(cv_code[2]), .Y(n27) );
  INVX1 U32 ( .A(cv_code[4]), .Y(n26) );
  XNOR2XL U33 ( .A(cv_code[2]), .B(cv_code[1]), .Y(n55) );
  NAND3X1 U34 ( .A(cv_code[2]), .B(cv_code[1]), .C(cv_code[3]), .Y(n52) );
  NAND2X1 U35 ( .A(cv_code[5]), .B(n50), .Y(n49) );
  INVX1 U36 ( .A(cv_code[1]), .Y(n28) );
  INVX1 U37 ( .A(N84), .Y(n23) );
  XOR2X1 U38 ( .A(N99), .B(add_62_carry_5_), .Y(r_dac3[5]) );
  NOR2X1 U39 ( .A(n48), .B(n23), .Y(N99) );
  NOR21XL U40 ( .B(add_62_carry_4_), .A(n12), .Y(add_62_carry_5_) );
  XNOR2XL U41 ( .A(n49), .B(n25), .Y(n48) );
  NOR2X1 U42 ( .A(N84), .B(cv_code[10]), .Y(n76) );
  NAND21X1 U43 ( .B(cv_code[9]), .A(n23), .Y(r_dac0[9]) );
  XOR2X1 U44 ( .A(add_62_carry_4_), .B(N98), .Y(r_dac3[4]) );
  OAI21BBX1 U45 ( .A(cv_code[10]), .B(cv_code[9]), .C(n23), .Y(n74) );
  INVX1 U46 ( .A(N106), .Y(n17) );
  NOR2X1 U47 ( .A(r_dac0[10]), .B(cv_code[9]), .Y(n72) );
  NOR3XL U48 ( .A(n30), .B(n58), .C(n29), .Y(n56) );
  XOR2X1 U49 ( .A(N94), .B(N106), .Y(r_dac3[0]) );
  OR2X1 U50 ( .A(cv_code[8]), .B(N84), .Y(r_dac0[8]) );
  OR2X1 U51 ( .A(cv_code[7]), .B(N84), .Y(r_dac0[7]) );
  OR2X1 U52 ( .A(cv_code[5]), .B(N84), .Y(r_dac0[5]) );
  OR2X1 U53 ( .A(cv_code[3]), .B(N84), .Y(r_dac0[3]) );
  NOR21XL U54 ( .B(N35), .A(n62), .Y(N40) );
  NOR21XL U55 ( .B(N36), .A(n62), .Y(N41) );
  NOR21XL U56 ( .B(N34), .A(n62), .Y(N39) );
  INVX1 U57 ( .A(n37), .Y(n19) );
  NOR21XL U58 ( .B(N123), .A(n37), .Y(N129) );
  NOR21XL U59 ( .B(N122), .A(n37), .Y(N128) );
  NOR21XL U60 ( .B(N121), .A(n37), .Y(N127) );
  NOR2X1 U61 ( .A(n53), .B(n23), .Y(N97) );
  AO2222XL U62 ( .A(r_cvofs[7]), .B(n72), .C(r_cvofs[15]), .D(n73), .E(
        r_cvofs[14]), .F(n74), .G(r_cvofs[6]), .H(n75), .Y(N109) );
  XNOR2XL U63 ( .A(n52), .B(n26), .Y(n53) );
  XNOR2XL U64 ( .A(r_vcomp[3]), .B(n60), .Y(N63) );
  NAND2X1 U65 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .Y(n60) );
  XNOR2XL U66 ( .A(r_vcomp[4]), .B(n58), .Y(N64) );
  XNOR2XL U67 ( .A(n59), .B(n29), .Y(N65) );
  NOR2X1 U68 ( .A(n58), .B(n30), .Y(n59) );
  XNOR2XL U69 ( .A(r_vcomp[7]), .B(n57), .Y(N67) );
  NAND2X1 U70 ( .A(r_vcomp[6]), .B(n56), .Y(n57) );
  GEN2XL U71 ( .D(N84), .E(n27), .C(N94), .B(cv_code[3]), .A(n54), .Y(N96) );
  AO2222XL U72 ( .A(r_cvofs[2]), .B(n72), .C(r_cvofs[10]), .D(n73), .E(
        r_cvofs[13]), .F(n74), .G(r_cvofs[5]), .H(n75), .Y(N108) );
  NOR4XL U73 ( .A(cv_code[3]), .B(n28), .C(n27), .D(n23), .Y(n54) );
  XOR2X1 U74 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .Y(N62) );
  XOR2X1 U75 ( .A(n56), .B(r_vcomp[6]), .Y(N66) );
  AND3X1 U76 ( .A(r_vcomp[7]), .B(n56), .C(r_vcomp[6]), .Y(N68) );
  AO2222XL U77 ( .A(r_cvofs[0]), .B(n72), .C(r_cvofs[8]), .D(n73), .E(
        r_cvofs[11]), .F(n74), .G(r_cvofs[3]), .H(n75), .Y(N106) );
  NOR32XL U78 ( .B(r_hlsb_en), .C(clk_5k), .A(r_hlsb_sel), .Y(N47) );
  NOR21XL U79 ( .B(r_vcomp[0]), .A(n47), .Y(
        add_3_root_sub_0_root_add_46_3_carry[1]) );
  NOR2X1 U80 ( .A(n55), .B(n23), .Y(N95) );
  AO2222XL U81 ( .A(r_cvofs[1]), .B(n72), .C(r_cvofs[9]), .D(n73), .E(
        r_cvofs[12]), .F(n74), .G(r_cvofs[4]), .H(n75), .Y(N107) );
  NOR21XL U82 ( .B(N94), .A(n17), .Y(add_62_carry_1_) );
  XNOR2XL U83 ( .A(r_vcomp[0]), .B(n47), .Y(N60) );
  NAND3X1 U84 ( .A(r_hlsb_en), .B(clk_5k), .C(r_hlsb_sel), .Y(n47) );
  NAND3X1 U85 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .C(r_vcomp[3]), .Y(n58) );
  INVX1 U86 ( .A(r_vcomp[4]), .Y(n30) );
  INVX1 U87 ( .A(r_vcomp[5]), .Y(n29) );
  NOR21XL U88 ( .B(sdischg_cnt[3]), .A(r_sdischg[3]), .Y(n46) );
  OAI32X1 U89 ( .A(n22), .B(sdischg_cnt[2]), .C(n46), .D(sdischg_cnt[3]), .E(
        n21), .Y(n44) );
  INVX1 U90 ( .A(r_sdischg[3]), .Y(n21) );
  AO222X1 U91 ( .A(n34), .B(n19), .C(n35), .D(n36), .E(sdischg_duty), .F(n37), 
        .Y(n81) );
  AOI22BXL U92 ( .B(N126), .A(n38), .D(r_sdischg[1]), .C(sdischg_cnt[1]), .Y(
        n35) );
  OAI22AX1 U93 ( .D(n36), .C(n43), .A(sdischg_cnt[4]), .B(n20), .Y(n34) );
  EORX1 U94 ( .A(n20), .B(sdischg_cnt[4]), .C(n45), .D(n44), .Y(n36) );
  AOI21X1 U95 ( .B(sdischg_cnt[2]), .C(n22), .A(n46), .Y(n45) );
  AOI21BX1 U96 ( .C(sdischg_cnt[1]), .B(r_sdischg[1]), .A(n44), .Y(n43) );
  OAI221X1 U97 ( .A(n63), .B(n18), .C(n64), .D(n33), .E(r_hlsb_en), .Y(n62) );
  INVX1 U98 ( .A(r_hlsb_freq), .Y(n18) );
  AOI211X1 U99 ( .C(div20_cnt[1]), .D(div20_cnt[0]), .A(div20_cnt[3]), .B(
        div20_cnt[2]), .Y(n64) );
  AOI21X1 U100 ( .B(div20_cnt[0]), .C(div20_cnt[3]), .A(n65), .Y(n63) );
  NOR2X1 U101 ( .A(r_sdischg[6]), .B(r_sdischg[5]), .Y(n37) );
  NAND2X1 U102 ( .A(n33), .B(n68), .Y(n65) );
  OAI21X1 U103 ( .B(div20_cnt[1]), .C(div20_cnt[2]), .A(div20_cnt[3]), .Y(n68)
         );
  INVX1 U104 ( .A(div20_cnt[4]), .Y(n33) );
  INVX1 U105 ( .A(r_sdischg[4]), .Y(n20) );
  NOR2X1 U106 ( .A(n37), .B(sdischg_cnt[0]), .Y(N126) );
  INVX1 U107 ( .A(r_sdischg[2]), .Y(n22) );
  NAND2X1 U108 ( .A(r_sdischg[0]), .B(n19), .Y(n38) );
  NOR2X1 U109 ( .A(n61), .B(n62), .Y(N42) );
  XNOR2XL U110 ( .A(div20_cnt[4]), .B(add_41_carry[4]), .Y(n61) );
  NOR2X1 U111 ( .A(div20_cnt[0]), .B(n62), .Y(N38) );
  NOR2X1 U112 ( .A(n37), .B(n70), .Y(N130) );
  XNOR2XL U113 ( .A(sdischg_cnt[4]), .B(add_81_carry[4]), .Y(n70) );
  OAI21BX1 U114 ( .C(n69), .B(div20_cnt[3]), .A(r_hlsb_freq), .Y(n66) );
  OAI31XL U115 ( .A(div20_cnt[1]), .B(r_hlsb_duty), .C(div20_cnt[0]), .D(
        div20_cnt[2]), .Y(n69) );
  AOI31X1 U116 ( .A(n66), .B(n67), .C(n32), .D(n31), .Y(N29) );
  INVX1 U117 ( .A(r_hlsb_en), .Y(n31) );
  NAND3X1 U118 ( .A(div20_cnt[0]), .B(div20_cnt[3]), .C(r_hlsb_duty), .Y(n67)
         );
  INVX1 U119 ( .A(n65), .Y(n32) );
  NAND42X1 U120 ( .C(sdischg_cnt[0]), .D(sdischg_cnt[1]), .A(n37), .B(n71), 
        .Y(N115) );
  NOR3XL U121 ( .A(sdischg_cnt[2]), .B(sdischg_cnt[4]), .C(sdischg_cnt[3]), 
        .Y(n71) );
endmodule


module cvctl_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module cvctl_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  XOR2X1 U2 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U4 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  XOR2X1 U5 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U6 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  AND2X1 U7 ( .A(carry[10]), .B(A[10]), .Y(carry[11]) );
endmodule


module cvctl_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n11, n12, n13, n14, n15, n16, n17, n18, n19;
  wire   [10:1] carry;

  FAD1X1 U2_7 ( .A(A[7]), .B(n11), .CI(carry[7]), .CO(carry[8]), .SO(DIFF[7])
         );
  FAD1X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n13), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n14), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n16), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n17), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR2X1 U1 ( .A(n1), .B(A[11]), .Y(DIFF[11]) );
  NOR2X1 U2 ( .A(A[10]), .B(carry[10]), .Y(n1) );
  XNOR2XL U3 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2XL U4 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2XL U5 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  INVX1 U6 ( .A(B[3]), .Y(n15) );
  INVX1 U7 ( .A(B[4]), .Y(n14) );
  INVX1 U8 ( .A(B[5]), .Y(n13) );
  INVX1 U9 ( .A(B[6]), .Y(n12) );
  INVX1 U10 ( .A(B[1]), .Y(n17) );
  NAND21X1 U11 ( .B(n18), .A(n19), .Y(carry[1]) );
  INVX1 U12 ( .A(A[0]), .Y(n19) );
  INVX1 U13 ( .A(B[2]), .Y(n16) );
  INVX1 U14 ( .A(B[7]), .Y(n11) );
  XNOR2XL U15 ( .A(n18), .B(A[0]), .Y(DIFF[0]) );
  OR2X1 U16 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  INVX1 U17 ( .A(B[0]), .Y(n18) );
  OR2X1 U18 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_cvctl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_20 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9392;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_20 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9392), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9392), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9392), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9392), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9392), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9392), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9392), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9392), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9392), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_21 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9410;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_21 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9410), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9410), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9410), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9410), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9410), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9410), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9410), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9410), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9410), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_22 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9428;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_22 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9428), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9428), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9428), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9428), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9428), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9428), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9428), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9428), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9428), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_23 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9446;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_23 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9446), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9446), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9446), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9446), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9446), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9446), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9446), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9446), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9446), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_24 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9464;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_24 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9464), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9464), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9464), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9464), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9464), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9464), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9464), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9464), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9464), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_25 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9482;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_25 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9482), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9482), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9482), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9482), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9482), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9482), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9482), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9482), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9482), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcp_a0 ( dp_comp, dm_comp, id_comp, intr, tx_en, tx_dat, r_dat, r_sta, 
        r_ctl, r_msk, r_crc, r_acc, r_dpdmsta, r_wdat, r_wr, r_re, clk, srstz, 
        r_tui, test_si, test_so, test_se );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  output [7:0] r_crc;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input [7:0] r_wdat;
  input [6:0] r_wr;
  output [7:0] r_tui;
  input dp_comp, dm_comp, id_comp, r_re, clk, srstz, test_si, test_se;
  output intr, tx_en, tx_dat, test_so;
  wire   r_dm, r_dmchg, r_acc_int, r_wr_last, r_wr_other, n3, n4, n1;

  INVX1 U3 ( .A(n4), .Y(n3) );
  INVX1 U4 ( .A(srstz), .Y(n4) );
  dpdmacc_a0 u0_dpdmacc ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(
        id_comp), .r_re_0(r_re), .r_wr_1(r_wr[6]), .r_wdat(r_wdat), .r_acc(
        r_acc), .r_dpdmsta(r_dpdmsta), .r_dm(r_dm), .r_dmchg(r_dmchg), .r_int(
        r_acc_int), .clk(clk), .rstz(srstz), .test_si(test_si), .test_se(
        test_se) );
  fcpegn_a0 u0_fcpegn ( .intr(intr), .tx_en(tx_en), .tx_dat(tx_dat), .r_dat(
        r_dat), .r_sta(r_sta), .r_ctl(r_ctl), .r_msk(r_msk), .r_wr(r_wr[4:0]), 
        .r_wdat(r_wdat), .ff_idn(r_dm), .ff_chg(n1), .r_acc_int(r_acc_int), 
        .clk(clk), .srstz(n3), .r_tui(r_tui), .test_si(r_crc[7]), .test_so(
        test_so), .test_se(test_se) );
  fcpcrc_a0 u0_fcpcrc ( .tx_crc(r_crc), .crc_din(r_wdat), .crc_en(r_ctl[2]), 
        .crc_shfi(r_wr_other), .crc_shfl(r_wr_last), .clk(clk), .srstz(n3), 
        .test_si(r_dpdmsta[5]), .test_se(test_se) );
  BUFX3 U1 ( .A(r_dmchg), .Y(n1) );
  AND2X1 U2 ( .A(r_wr[5]), .B(r_ctl[3]), .Y(r_wr_last) );
  NOR21XL U5 ( .B(r_wr[5]), .A(r_ctl[3]), .Y(r_wr_other) );
endmodule


module fcpcrc_a0 ( tx_crc, crc_din, crc_en, crc_shfi, crc_shfl, clk, srstz, 
        test_si, test_se );
  output [7:0] tx_crc;
  input [7:0] crc_din;
  input crc_en, crc_shfi, crc_shfl, clk, srstz, test_si, test_se;
  wire   N81, N82, N83, N84, N85, N86, N87, N88, N89, net9500, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n1;

  SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 clk_gate_crc8_r_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net9500), .TE(test_se) );
  SDFFRQX1 crc8_r_reg_1_ ( .D(N83), .SIN(tx_crc[0]), .SMC(test_se), .C(net9500), .XR(srstz), .Q(tx_crc[1]) );
  SDFFRQX1 crc8_r_reg_0_ ( .D(N82), .SIN(test_si), .SMC(test_se), .C(net9500), 
        .XR(srstz), .Q(tx_crc[0]) );
  SDFFRQX1 crc8_r_reg_4_ ( .D(N86), .SIN(tx_crc[3]), .SMC(test_se), .C(net9500), .XR(srstz), .Q(tx_crc[4]) );
  SDFFRQX1 crc8_r_reg_3_ ( .D(N85), .SIN(tx_crc[2]), .SMC(test_se), .C(net9500), .XR(srstz), .Q(tx_crc[3]) );
  SDFFRQX1 crc8_r_reg_2_ ( .D(N84), .SIN(tx_crc[1]), .SMC(test_se), .C(net9500), .XR(srstz), .Q(tx_crc[2]) );
  SDFFRQX1 crc8_r_reg_6_ ( .D(N88), .SIN(tx_crc[5]), .SMC(test_se), .C(net9500), .XR(srstz), .Q(tx_crc[6]) );
  SDFFRQX1 crc8_r_reg_7_ ( .D(N89), .SIN(tx_crc[6]), .SMC(test_se), .C(net9500), .XR(srstz), .Q(tx_crc[7]) );
  SDFFRQX1 crc8_r_reg_5_ ( .D(N87), .SIN(tx_crc[4]), .SMC(test_se), .C(net9500), .XR(srstz), .Q(tx_crc[5]) );
  XNOR2XL U3 ( .A(n36), .B(n37), .Y(n15) );
  XNOR2XL U4 ( .A(n35), .B(n34), .Y(n19) );
  XNOR2XL U5 ( .A(n8), .B(n1), .Y(n35) );
  XNOR2XL U6 ( .A(n28), .B(n24), .Y(n13) );
  XNOR2XL U7 ( .A(n13), .B(n23), .Y(n8) );
  XNOR2XL U8 ( .A(n2), .B(n9), .Y(n28) );
  OAI22X1 U9 ( .A(n15), .B(n3), .C(n16), .D(n5), .Y(N87) );
  XNOR2XL U10 ( .A(n17), .B(n18), .Y(n16) );
  XNOR2XL U11 ( .A(n6), .B(n15), .Y(n18) );
  XNOR2XL U12 ( .A(n19), .B(n14), .Y(n17) );
  OAI22X1 U13 ( .A(n24), .B(n3), .C(n25), .D(n5), .Y(N85) );
  XNOR2XL U14 ( .A(n19), .B(n13), .Y(n25) );
  OAI22X1 U15 ( .A(n20), .B(n3), .C(n21), .D(n5), .Y(N86) );
  XOR2X1 U16 ( .A(n19), .B(n22), .Y(n21) );
  XNOR2XL U17 ( .A(n14), .B(n23), .Y(n22) );
  XNOR2XL U18 ( .A(n31), .B(n32), .Y(n14) );
  XNOR2XL U19 ( .A(n1), .B(n30), .Y(n32) );
  XNOR2XL U20 ( .A(n23), .B(n9), .Y(n31) );
  XOR2X1 U21 ( .A(n20), .B(n2), .Y(n23) );
  XNOR2XL U22 ( .A(n27), .B(n26), .Y(n6) );
  XNOR2XL U23 ( .A(n15), .B(n28), .Y(n27) );
  XNOR2XL U24 ( .A(n41), .B(n42), .Y(n24) );
  XNOR2XL U25 ( .A(crc_din[3]), .B(n43), .Y(n42) );
  XNOR2XL U26 ( .A(n38), .B(n39), .Y(n20) );
  XNOR2XL U27 ( .A(crc_din[4]), .B(n40), .Y(n39) );
  OAI22X1 U28 ( .A(n2), .B(n3), .C(n4), .D(n5), .Y(N89) );
  XOR2X1 U29 ( .A(n6), .B(n7), .Y(n4) );
  XNOR2XL U30 ( .A(n8), .B(n2), .Y(n7) );
  OAI22X1 U31 ( .A(n34), .B(n3), .C(n19), .D(n5), .Y(N82) );
  OAI22X1 U32 ( .A(n9), .B(n3), .C(n10), .D(n5), .Y(N88) );
  XNOR2XL U33 ( .A(n11), .B(n12), .Y(n10) );
  XNOR2XL U34 ( .A(n13), .B(n9), .Y(n12) );
  XNOR2XL U35 ( .A(n14), .B(n6), .Y(n11) );
  INVX1 U36 ( .A(n15), .Y(n1) );
  OAI22X1 U37 ( .A(n26), .B(n3), .C(n6), .D(n5), .Y(N84) );
  XNOR2XL U38 ( .A(crc_din[1]), .B(n33), .Y(n30) );
  XNOR2XL U39 ( .A(crc_din[2]), .B(n29), .Y(n26) );
  XNOR2XL U40 ( .A(crc_din[0]), .B(n41), .Y(n34) );
  OAI22X1 U41 ( .A(n30), .B(n3), .C(n14), .D(n5), .Y(N83) );
  XOR2X1 U42 ( .A(n41), .B(n33), .Y(n38) );
  XNOR2XL U43 ( .A(n43), .B(n40), .Y(n51) );
  XNOR2XL U44 ( .A(n44), .B(n45), .Y(n9) );
  XNOR2XL U45 ( .A(n33), .B(n43), .Y(n45) );
  XNOR2XL U46 ( .A(n29), .B(n48), .Y(n44) );
  XNOR2XL U47 ( .A(tx_crc[6]), .B(crc_din[6]), .Y(n48) );
  XNOR2XL U48 ( .A(n49), .B(n50), .Y(n2) );
  XOR2X1 U49 ( .A(n51), .B(n29), .Y(n49) );
  XNOR2XL U50 ( .A(tx_crc[7]), .B(crc_din[7]), .Y(n50) );
  XNOR2XL U51 ( .A(n38), .B(n29), .Y(n36) );
  XNOR2XL U52 ( .A(tx_crc[5]), .B(crc_din[5]), .Y(n37) );
  NAND21X1 U53 ( .B(crc_shfl), .A(crc_en), .Y(n3) );
  NAND2X1 U54 ( .A(crc_shfl), .B(crc_en), .Y(n5) );
  OR2X1 U55 ( .A(crc_shfi), .B(n3), .Y(N81) );
  XOR2X1 U56 ( .A(n46), .B(n47), .Y(n33) );
  XOR2X1 U57 ( .A(tx_crc[5]), .B(tx_crc[6]), .Y(n46) );
  XNOR2XL U58 ( .A(tx_crc[1]), .B(n40), .Y(n47) );
  XNOR2XL U59 ( .A(tx_crc[3]), .B(n53), .Y(n43) );
  XNOR2XL U60 ( .A(tx_crc[7]), .B(tx_crc[4]), .Y(n40) );
  XNOR2XL U61 ( .A(n51), .B(n54), .Y(n41) );
  XOR2X1 U62 ( .A(tx_crc[0]), .B(tx_crc[5]), .Y(n54) );
  XOR2X1 U63 ( .A(tx_crc[7]), .B(tx_crc[6]), .Y(n53) );
  XNOR2XL U64 ( .A(n52), .B(n53), .Y(n29) );
  XNOR2XL U65 ( .A(tx_crc[5]), .B(tx_crc[2]), .Y(n52) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcpegn_a0 ( intr, tx_en, tx_dat, r_dat, r_sta, r_ctl, r_msk, r_wr, 
        r_wdat, ff_idn, ff_chg, r_acc_int, clk, srstz, r_tui, test_si, test_so, 
        test_se );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  input [4:0] r_wr;
  input [7:0] r_wdat;
  output [7:0] r_tui;
  input ff_idn, ff_chg, r_acc_int, clk, srstz, test_si, test_se;
  output intr, tx_en, tx_dat, test_so;
  wire   N22, upd_dbuf_en, us_cnt_2_, us_cnt_1_, us_cnt_0_, N85, N87, N88,
         N141, N142, N144, N145, N172, N173, adp_tx_ui_7_, adp_tx_ui_6_, N205,
         N221, N222, N223, N224, N225, N226, N227, N228, N260, N261, N348,
         N349, N356, N362, N363, N444, rx_trans_8_chg, N1005, N1006, N1007,
         N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1043,
         net9522, net9526, net9529, net9530, net9531, net9532, net9533,
         net9534, net9537, net9540, net9545, net9550, net9555, n26, n27, n28,
         n29, n30, n31, n32, n516, n525, n526, N1259, N1258, N1257, N1256,
         N1255, N1254, N1253, N1252, N161, N160, N159, N108, N107, n41, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n461, n464, n4, n83, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n463, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n517, n518, n519, n520, n521, n522,
         n523, n524, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n20, n21, n22, n23, n24, n25, n33, n34, n35, n36, n37, n38, n39,
         n40, n42, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3;
  wire   [6:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;
  wire   [7:0] upd_dbuf;
  wire   [10:0] rxtx_buf;
  wire   [4:1] rx_ui_3_8;
  wire   [4:1] rx_ui_5_8;
  wire   [5:0] catch_sync;
  wire   [7:0] ui_intv_cnt;
  wire   [6:2] symb_cnt;
  wire   [6:0] adp_tx_1_4;
  wire   [7:0] tui_wdat;
  wire   [11:0] trans_buf;
  wire   [1:0] new_rx_sync_cnt;
  wire   [3:0] fcp_state;
  wire   [5:1] add_264_carry;
  wire   [5:1] add_263_carry;
  wire   [8:6] add_274_2_carry;
  wire   [8:6] add_274_carry;

  FAD1X1 add_264_U1_1 ( .A(n69), .B(n72), .CI(add_264_carry[1]), .CO(
        add_264_carry[2]), .SO(rx_ui_5_8[1]) );
  FAD1X1 add_264_U1_2 ( .A(n71), .B(n73), .CI(add_264_carry[2]), .CO(
        add_264_carry[3]), .SO(rx_ui_5_8[2]) );
  FAD1X1 add_264_U1_3 ( .A(n72), .B(n67), .CI(add_264_carry[3]), .CO(
        add_264_carry[4]), .SO(rx_ui_5_8[3]) );
  FAD1X1 add_264_U1_4 ( .A(n73), .B(n68), .CI(add_264_carry[4]), .CO(
        add_264_carry[5]), .SO(rx_ui_5_8[4]) );
  FAD1X1 add_263_U1_1 ( .A(n71), .B(n72), .CI(add_263_carry[1]), .CO(
        add_263_carry[2]), .SO(rx_ui_3_8[1]) );
  FAD1X1 add_263_U1_2 ( .A(n72), .B(n73), .CI(add_263_carry[2]), .CO(
        add_263_carry[3]), .SO(rx_ui_3_8[2]) );
  FAD1X1 add_263_U1_3 ( .A(n73), .B(n67), .CI(add_263_carry[3]), .CO(
        add_263_carry[4]), .SO(rx_ui_3_8[3]) );
  FAD1X1 add_263_U1_4 ( .A(n67), .B(n6), .CI(add_263_carry[4]), .CO(
        add_263_carry[5]), .SO(rx_ui_3_8[4]) );
  FAD1X1 add_274_2_U1_6 ( .A(N160), .B(ui_intv_cnt[6]), .CI(add_274_2_carry[6]), .CO(add_274_2_carry[7]), .SO(N172) );
  FAD1X1 add_274_2_U1_7 ( .A(N161), .B(ui_intv_cnt[7]), .CI(add_274_2_carry[7]), .CO(add_274_2_carry[8]), .SO(N173) );
  FAD1X1 add_274_U1_6 ( .A(N107), .B(ui_intv_cnt[6]), .CI(add_274_carry[6]), 
        .CO(add_274_carry[7]), .SO(N144) );
  FAD1X1 add_274_U1_7 ( .A(N108), .B(ui_intv_cnt[7]), .CI(add_274_carry[7]), 
        .CO(add_274_carry[8]), .SO(N145) );
  INVX1 U23 ( .A(n51), .Y(n46) );
  INVX1 U24 ( .A(n51), .Y(n47) );
  INVX1 U25 ( .A(n51), .Y(n48) );
  INVX1 U26 ( .A(n51), .Y(n49) );
  INVX1 U27 ( .A(n51), .Y(n50) );
  INVX1 U28 ( .A(n51), .Y(n45) );
  INVX1 U29 ( .A(n51), .Y(n43) );
  INVX1 U30 ( .A(n51), .Y(n44) );
  INVX1 U31 ( .A(n51), .Y(n41) );
  INVX1 U32 ( .A(srstz), .Y(n51) );
  MAJ3X1 U619 ( .A(rx_ui_3_8[1]), .B(n447), .C(n117), .Y(n446) );
  glreg_8_00000000 u0_fcpctl ( .clk(clk), .arstz(n46), .we(r_wr[0]), .wdat({
        r_wdat[7:3], n23, r_wdat[1:0]}), .rdat({n464, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, r_ctl[4:0]}), .test_si(r_ctl[7]), .test_se(
        test_se) );
  glsta_a0_0 u0_fcpsta ( .clk(clk), .arstz(n45), .rst0(1'b0), .set2({r_acc_int, 
        setsta[6:5], n536, setsta[3], n525, n4, setsta[0]}), .clr1(clrsta), 
        .rdat(r_sta), .irq(r_irq), .test_si(r_msk[7]), .test_se(test_se) );
  glreg_a0_4 u0_fcpmsk ( .clk(clk), .arstz(n44), .we(r_wr[2]), .wdat({
        r_wdat[7:3], n23, r_wdat[1:0]}), .rdat(r_msk), .test_si(r_dat[7]), 
        .test_se(test_se) );
  glreg_a0_3 u0_fcpdat ( .clk(clk), .arstz(n43), .we(upd_dbuf_en), .wdat(
        upd_dbuf), .rdat(r_dat), .test_si(n464), .test_se(test_se) );
  glreg_a0_2 u0_fcptui ( .clk(clk), .arstz(n41), .we(n83), .wdat(tui_wdat), 
        .rdat(r_tui), .test_si(r_sta[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 clk_gate_catch_sync_reg ( .CLK(clk), .EN(
        n526), .ENCLK(net9522), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 clk_gate_ui_intv_cnt_reg ( .CLK(clk), .EN(
        N205), .ENCLK(net9540), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 clk_gate_rxtx_buf_reg ( .CLK(clk), .EN(N22), 
        .ENCLK(net9545), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 clk_gate_fcp_state_reg ( .CLK(clk), .EN(
        N1005), .ENCLK(net9550), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 clk_gate_symb_cnt_reg ( .CLK(clk), .EN(
        N1043), .ENCLK(net9555), .TE(test_se) );
  fcpegn_a0_DW01_inc_0 r611 ( .A({symb_cnt[6:4], n14, n12, n8, n16}), .SUM({
        n26, n27, n28, n29, n30, n31, n32}) );
  fcpegn_a0_DW01_inc_1 add_283_round ( .A({1'b0, adp_tx_ui_7_, adp_tx_ui_6_, 
        n75, r_tui[4:1]}), .SUM({adp_tx_1_4, SYNOPSYS_UNCONNECTED_3}) );
  fcpegn_a0_DW01_inc_2 add_316_aco ( .A({N1259, N1258, N1257, N1256, N1255, 
        N1254, N1253, N1252}), .SUM({N228, N227, N226, N225, N224, N223, N222, 
        N221}) );
  SDFFRQX1 rxtx_buf_reg_8_ ( .D(trans_buf[8]), .SIN(rxtx_buf[7]), .SMC(test_se), .C(net9545), .XR(n47), .Q(rxtx_buf[8]) );
  SDFFRQX1 rxtx_buf_reg_10_ ( .D(trans_buf[10]), .SIN(rxtx_buf[9]), .SMC(
        test_se), .C(net9545), .XR(n47), .Q(rxtx_buf[10]) );
  SDFFRQX1 rxtx_buf_reg_9_ ( .D(trans_buf[9]), .SIN(rxtx_buf[8]), .SMC(test_se), .C(net9545), .XR(n47), .Q(rxtx_buf[9]) );
  SDFFRQX1 rxtx_buf_reg_0_ ( .D(trans_buf[0]), .SIN(rx_trans_8_chg), .SMC(
        test_se), .C(net9545), .XR(n48), .Q(rxtx_buf[0]) );
  SDFFRQX1 rxtx_buf_reg_4_ ( .D(trans_buf[4]), .SIN(rxtx_buf[3]), .SMC(test_se), .C(net9545), .XR(n47), .Q(rxtx_buf[4]) );
  SDFFRQX1 rxtx_buf_reg_6_ ( .D(trans_buf[6]), .SIN(rxtx_buf[5]), .SMC(test_se), .C(net9545), .XR(n47), .Q(rxtx_buf[6]) );
  SDFFRQX1 rxtx_buf_reg_7_ ( .D(trans_buf[7]), .SIN(rxtx_buf[6]), .SMC(test_se), .C(net9545), .XR(n47), .Q(rxtx_buf[7]) );
  SDFFRQX1 rxtx_buf_reg_3_ ( .D(trans_buf[3]), .SIN(rxtx_buf[2]), .SMC(test_se), .C(net9545), .XR(n48), .Q(rxtx_buf[3]) );
  SDFFRQX1 rxtx_buf_reg_5_ ( .D(trans_buf[5]), .SIN(rxtx_buf[4]), .SMC(test_se), .C(net9545), .XR(n47), .Q(rxtx_buf[5]) );
  SDFFRQX1 rxtx_buf_reg_1_ ( .D(trans_buf[1]), .SIN(rxtx_buf[0]), .SMC(test_se), .C(net9545), .XR(n49), .Q(rxtx_buf[1]) );
  SDFFRQX1 rx_byte_pchk_reg ( .D(N356), .SIN(new_rx_sync_cnt[1]), .SMC(test_se), .C(clk), .XR(n50), .Q(setsta[5]) );
  SDFFRQX1 rxtx_buf_reg_2_ ( .D(trans_buf[2]), .SIN(rxtx_buf[1]), .SMC(test_se), .C(net9545), .XR(n47), .Q(rxtx_buf[2]) );
  SDFFRQX1 new_rx_sync_cnt_reg_1_ ( .D(N349), .SIN(new_rx_sync_cnt[0]), .SMC(
        test_se), .C(clk), .XR(n44), .Q(new_rx_sync_cnt[1]) );
  SDFFRQX1 new_rx_sync_cnt_reg_0_ ( .D(N348), .SIN(fcp_state[3]), .SMC(test_se), .C(clk), .XR(n41), .Q(new_rx_sync_cnt[0]) );
  SDFFQX1 rx_trans_8_chg_reg ( .D(n516), .SIN(setsta[5]), .SMC(test_se), .C(
        clk), .Q(rx_trans_8_chg) );
  SDFFRQX1 us_cnt_reg_3_ ( .D(N88), .SIN(us_cnt_2_), .SMC(test_se), .C(clk), 
        .XR(n43), .Q(test_so) );
  SDFFRQX1 us_cnt_reg_2_ ( .D(N87), .SIN(us_cnt_1_), .SMC(test_se), .C(clk), 
        .XR(n45), .Q(us_cnt_2_) );
  SDFFRQX1 us_cnt_reg_1_ ( .D(n461), .SIN(us_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(srstz), .Q(us_cnt_1_) );
  SDFFRQX1 us_cnt_reg_0_ ( .D(N85), .SIN(ui_intv_cnt[7]), .SMC(test_se), .C(
        clk), .XR(n47), .Q(us_cnt_0_) );
  SDFFRQX1 ui_intv_cnt_reg_6_ ( .D(net9529), .SIN(n11), .SMC(test_se), .C(
        net9540), .XR(n49), .Q(ui_intv_cnt[6]) );
  SDFFRQX1 ui_intv_cnt_reg_7_ ( .D(net9526), .SIN(ui_intv_cnt[6]), .SMC(
        test_se), .C(net9540), .XR(n49), .Q(ui_intv_cnt[7]) );
  SDFFRQX1 ui_intv_cnt_reg_4_ ( .D(net9531), .SIN(N141), .SMC(test_se), .C(
        net9540), .XR(n49), .Q(N142) );
  SDFFRQX1 ui_intv_cnt_reg_1_ ( .D(net9534), .SIN(ui_intv_cnt[0]), .SMC(
        test_se), .C(net9540), .XR(n48), .Q(ui_intv_cnt[1]) );
  SDFFRQX1 ui_intv_cnt_reg_3_ ( .D(net9532), .SIN(ui_intv_cnt[2]), .SMC(
        test_se), .C(net9540), .XR(n48), .Q(N141) );
  SDFFRQX1 ui_intv_cnt_reg_0_ ( .D(net9537), .SIN(r_tui[7]), .SMC(test_se), 
        .C(net9540), .XR(n48), .Q(ui_intv_cnt[0]) );
  SDFFRQX1 ui_intv_cnt_reg_2_ ( .D(net9533), .SIN(ui_intv_cnt[1]), .SMC(
        test_se), .C(net9540), .XR(n48), .Q(ui_intv_cnt[2]) );
  SDFFRQX1 ui_intv_cnt_reg_5_ ( .D(net9530), .SIN(n3), .SMC(test_se), .C(
        net9540), .XR(n49), .Q(ui_intv_cnt[5]) );
  SDFFSQX1 catch_sync_reg_5_ ( .D(n11), .SIN(catch_sync[4]), .SMC(test_se), 
        .C(net9522), .XS(n46), .Q(catch_sync[5]) );
  SDFFRQX1 catch_sync_reg_4_ ( .D(n3), .SIN(catch_sync[3]), .SMC(test_se), .C(
        net9522), .XR(n48), .Q(catch_sync[4]) );
  SDFFRQX1 sync_length_reg_1_ ( .D(N261), .SIN(N362), .SMC(test_se), .C(
        net9540), .XR(n49), .Q(N363) );
  SDFFRQX1 symb_cnt_reg_4_ ( .D(N1014), .SIN(n14), .SMC(test_se), .C(net9555), 
        .XR(n50), .Q(symb_cnt[4]) );
  SDFFRQX1 symb_cnt_reg_5_ ( .D(N1015), .SIN(symb_cnt[4]), .SMC(test_se), .C(
        net9555), .XR(n50), .Q(symb_cnt[5]) );
  SDFFRQX1 symb_cnt_reg_6_ ( .D(N1016), .SIN(symb_cnt[5]), .SMC(test_se), .C(
        net9555), .XR(n49), .Q(symb_cnt[6]) );
  SDFFRQX1 sync_length_reg_0_ ( .D(N260), .SIN(symb_cnt[6]), .SMC(test_se), 
        .C(net9540), .XR(n49), .Q(N362) );
  SDFFRQX1 symb_cnt_reg_3_ ( .D(N1013), .SIN(n12), .SMC(test_se), .C(net9555), 
        .XR(n50), .Q(symb_cnt[3]) );
  SDFFSQX1 catch_sync_reg_3_ ( .D(N141), .SIN(catch_sync[2]), .SMC(test_se), 
        .C(net9522), .XS(n46), .Q(catch_sync[3]) );
  SDFFRQX1 symb_cnt_reg_1_ ( .D(N1011), .SIN(n16), .SMC(test_se), .C(net9555), 
        .XR(n50), .Q(N160) );
  SDFFRQX1 symb_cnt_reg_2_ ( .D(N1012), .SIN(n8), .SMC(test_se), .C(net9555), 
        .XR(n50), .Q(symb_cnt[2]) );
  SDFFRQX1 symb_cnt_reg_0_ ( .D(N1010), .SIN(tx_dat), .SMC(test_se), .C(
        net9555), .XR(n50), .Q(N159) );
  SDFFRQX1 catch_sync_reg_1_ ( .D(ui_intv_cnt[1]), .SIN(catch_sync[0]), .SMC(
        test_se), .C(net9522), .XR(n48), .Q(catch_sync[1]) );
  SDFFRQX1 catch_sync_reg_2_ ( .D(ui_intv_cnt[2]), .SIN(catch_sync[1]), .SMC(
        test_se), .C(net9522), .XR(n48), .Q(catch_sync[2]) );
  SDFFRQX1 catch_sync_reg_0_ ( .D(ui_intv_cnt[0]), .SIN(test_si), .SMC(test_se), .C(net9522), .XR(n48), .Q(catch_sync[0]) );
  SDFFSQX1 tx_dbuf_keep_empty_reg ( .D(N444), .SIN(N363), .SMC(test_se), .C(
        clk), .XS(n47), .Q(r_ctl[7]) );
  SDFFRQX1 rxtx_buf_reg_11_ ( .D(trans_buf[11]), .SIN(rxtx_buf[10]), .SMC(
        test_se), .C(net9545), .XR(n49), .Q(tx_dat) );
  SDFFRQX1 fcp_state_reg_3_ ( .D(N1009), .SIN(fcp_state[2]), .SMC(test_se), 
        .C(net9550), .XR(n49), .Q(fcp_state[3]) );
  SDFFRQX1 fcp_state_reg_1_ ( .D(N1007), .SIN(fcp_state[0]), .SMC(test_se), 
        .C(net9550), .XR(n50), .Q(fcp_state[1]) );
  SDFFRQX1 fcp_state_reg_2_ ( .D(N1008), .SIN(fcp_state[1]), .SMC(test_se), 
        .C(net9550), .XR(n50), .Q(fcp_state[2]) );
  SDFFRQX1 fcp_state_reg_0_ ( .D(N1006), .SIN(catch_sync[5]), .SMC(test_se), 
        .C(net9550), .XR(n50), .Q(fcp_state[0]) );
  BUFX3 U4 ( .A(n270), .Y(n2) );
  BUFX3 U5 ( .A(N142), .Y(n3) );
  INVX1 U6 ( .A(ff_idn), .Y(n5) );
  INVX1 U7 ( .A(n333), .Y(n6) );
  INVX1 U8 ( .A(n122), .Y(n7) );
  INVX1 U9 ( .A(n131), .Y(n8) );
  INVX1 U10 ( .A(n100), .Y(n9) );
  INVX1 U11 ( .A(n58), .Y(n10) );
  INVX1 U12 ( .A(n123), .Y(n11) );
  INVX1 U13 ( .A(n128), .Y(n12) );
  INVX1 U14 ( .A(r_ctl[0]), .Y(n13) );
  INVX1 U15 ( .A(n126), .Y(n14) );
  INVX1 U16 ( .A(r_wr[3]), .Y(n15) );
  BUFX3 U17 ( .A(N159), .Y(n16) );
  INVX1 U18 ( .A(N141), .Y(n17) );
  XNOR2XL U19 ( .A(n186), .B(n187), .Y(n157) );
  XNOR2XL U20 ( .A(n184), .B(n185), .Y(n159) );
  INVX1 U21 ( .A(r_wr[3]), .Y(n80) );
  INVX1 U22 ( .A(r_wr[4]), .Y(n81) );
  NOR2X1 U33 ( .A(n22), .B(n78), .Y(clrsta[1]) );
  NOR2X1 U34 ( .A(n33), .B(n78), .Y(clrsta[4]) );
  NOR2X1 U35 ( .A(n21), .B(n78), .Y(clrsta[0]) );
  NOR2X1 U36 ( .A(n35), .B(n78), .Y(clrsta[6]) );
  NOR2X1 U37 ( .A(n24), .B(n78), .Y(clrsta[2]) );
  NOR2X1 U38 ( .A(n36), .B(n78), .Y(clrsta[7]) );
  NOR2X1 U39 ( .A(n25), .B(n78), .Y(clrsta[3]) );
  INVX1 U40 ( .A(n24), .Y(n23) );
  INVX1 U41 ( .A(n295), .Y(n542) );
  INVX1 U42 ( .A(r_wr[1]), .Y(n78) );
  INVX1 U43 ( .A(r_wdat[6]), .Y(n35) );
  INVX1 U44 ( .A(r_wdat[3]), .Y(n25) );
  INVX1 U45 ( .A(r_wdat[4]), .Y(n33) );
  INVX1 U46 ( .A(r_wdat[2]), .Y(n24) );
  INVX1 U47 ( .A(r_wdat[7]), .Y(n36) );
  INVX1 U48 ( .A(r_wdat[0]), .Y(n21) );
  INVX1 U49 ( .A(r_wdat[1]), .Y(n22) );
  NOR2X1 U50 ( .A(n542), .B(n541), .Y(n264) );
  NOR2X1 U51 ( .A(n549), .B(n543), .Y(n295) );
  INVX1 U52 ( .A(n269), .Y(n79) );
  INVX1 U53 ( .A(n257), .Y(n42) );
  NOR2X1 U54 ( .A(n34), .B(n78), .Y(clrsta[5]) );
  OAI221X1 U55 ( .A(n103), .B(n155), .C(n34), .D(n81), .E(n158), .Y(
        tui_wdat[5]) );
  OAI221X1 U56 ( .A(n155), .B(n104), .C(n33), .D(n81), .E(n158), .Y(
        tui_wdat[4]) );
  OAI221X1 U57 ( .A(n105), .B(n155), .C(n25), .D(n81), .E(n158), .Y(
        tui_wdat[3]) );
  INVX1 U58 ( .A(n159), .Y(n105) );
  INVX1 U59 ( .A(n167), .Y(n101) );
  INVX1 U60 ( .A(n157), .Y(n103) );
  INVX1 U61 ( .A(n173), .Y(n104) );
  INVX1 U62 ( .A(n316), .Y(n66) );
  NAND2X1 U63 ( .A(n159), .B(n160), .Y(n179) );
  INVX1 U64 ( .A(n505), .Y(n113) );
  INVX1 U65 ( .A(n377), .Y(n543) );
  INVX1 U66 ( .A(n420), .Y(n541) );
  INVX1 U67 ( .A(n348), .Y(n549) );
  NOR2X1 U68 ( .A(n293), .B(n80), .Y(n269) );
  INVX1 U69 ( .A(n256), .Y(n52) );
  NAND2X1 U70 ( .A(n253), .B(n58), .Y(n257) );
  INVX1 U71 ( .A(n249), .Y(n58) );
  OAI222XL U72 ( .A(r_wr[4]), .B(n154), .C(n155), .D(n156), .E(n35), .F(n81), 
        .Y(tui_wdat[6]) );
  XNOR2XL U73 ( .A(n101), .B(n157), .Y(n156) );
  AND2X1 U74 ( .A(N224), .B(n279), .Y(net9532) );
  AND2X1 U75 ( .A(N226), .B(n279), .Y(net9530) );
  AND2X1 U76 ( .A(N223), .B(n279), .Y(net9533) );
  AND2X1 U77 ( .A(N222), .B(n279), .Y(net9534) );
  OAI2B11X1 U78 ( .D(N221), .C(n90), .A(n278), .B(n38), .Y(net9537) );
  OAI2B11X1 U79 ( .D(n160), .C(n155), .A(n158), .B(n161), .Y(tui_wdat[2]) );
  EORX1 U80 ( .A(r_wr[4]), .B(n23), .C(n154), .D(r_wr[4]), .Y(n161) );
  ENOX1 U81 ( .A(n280), .B(n278), .C(N225), .D(n279), .Y(net9531) );
  ENOX1 U82 ( .A(n280), .B(n278), .C(N227), .D(n279), .Y(net9529) );
  INVX1 U83 ( .A(n280), .Y(n38) );
  NAND3X1 U84 ( .A(n278), .B(n90), .C(n38), .Y(N205) );
  NAND31X1 U85 ( .C(n162), .A(n81), .B(n154), .Y(n155) );
  XNOR2XL U86 ( .A(n36), .B(n54), .Y(n342) );
  NAND2X1 U87 ( .A(n162), .B(n81), .Y(n158) );
  INVX1 U88 ( .A(r_wdat[5]), .Y(n34) );
  XNOR2XL U89 ( .A(n68), .B(add_263_carry[5]), .Y(n449) );
  XNOR2XL U90 ( .A(n177), .B(n176), .Y(n167) );
  AOI21X1 U91 ( .B(n176), .C(n177), .A(n175), .Y(n169) );
  OAI21BBX1 U92 ( .A(n216), .B(n233), .C(n239), .Y(n231) );
  OAI21X1 U93 ( .B(n216), .C(n233), .A(n235), .Y(n239) );
  NOR32XL U94 ( .B(n186), .C(n181), .A(n180), .Y(n177) );
  NOR21XL U95 ( .B(n181), .A(n180), .Y(n187) );
  XNOR2XL U96 ( .A(n180), .B(n181), .Y(n173) );
  XNOR2XL U97 ( .A(n233), .B(n234), .Y(n196) );
  XOR2X1 U98 ( .A(n235), .B(n216), .Y(n234) );
  NOR2X1 U99 ( .A(n132), .B(n114), .Y(n505) );
  AOI211X1 U100 ( .C(n111), .D(n309), .A(n245), .B(n307), .Y(n308) );
  NAND2X1 U101 ( .A(n132), .B(n130), .Y(N107) );
  INVX1 U102 ( .A(n418), .Y(n130) );
  INVX1 U103 ( .A(n339), .Y(n70) );
  NOR21XL U104 ( .B(n183), .A(n182), .Y(n185) );
  NAND32X1 U105 ( .B(n184), .C(n182), .A(n183), .Y(n180) );
  XNOR2XL U106 ( .A(n341), .B(n68), .Y(n316) );
  NAND2X1 U107 ( .A(n73), .B(n67), .Y(n341) );
  XNOR2XL U108 ( .A(n73), .B(n67), .Y(n318) );
  NOR2X1 U109 ( .A(n545), .B(n245), .Y(n393) );
  INVX1 U110 ( .A(n307), .Y(n37) );
  XNOR2XL U111 ( .A(n182), .B(n183), .Y(n160) );
  OAI21X1 U112 ( .B(n73), .C(n67), .A(n68), .Y(n321) );
  NOR2X1 U113 ( .A(n491), .B(n54), .Y(n427) );
  AOI32X1 U114 ( .A(n545), .B(n112), .C(n492), .D(n283), .E(n548), .Y(n491) );
  NAND2X1 U115 ( .A(n67), .B(add_264_carry[5]), .Y(n142) );
  INVX1 U116 ( .A(n309), .Y(n109) );
  INVX1 U117 ( .A(n509), .Y(n55) );
  INVX1 U118 ( .A(n492), .Y(n111) );
  INVX1 U119 ( .A(n486), .Y(n57) );
  NOR4XL U120 ( .A(n283), .B(n284), .C(n40), .D(n54), .Y(n525) );
  NAND2X1 U121 ( .A(n285), .B(n548), .Y(n284) );
  OAI211X1 U122 ( .C(n549), .D(n113), .A(n110), .B(n542), .Y(N1043) );
  INVX1 U123 ( .A(n293), .Y(n546) );
  NAND2X1 U124 ( .A(n493), .B(n544), .Y(n377) );
  NOR2X1 U125 ( .A(n550), .B(n352), .Y(n420) );
  NOR2X1 U126 ( .A(n533), .B(n551), .Y(n493) );
  NAND2X1 U127 ( .A(n535), .B(n551), .Y(n348) );
  INVX1 U128 ( .A(n376), .Y(n550) );
  BUFX3 U129 ( .A(ff_idn), .Y(r_ctl[5]) );
  XNOR2XL U130 ( .A(n265), .B(n266), .Y(n261) );
  XNOR2XL U131 ( .A(n271), .B(n272), .Y(n265) );
  XNOR2XL U132 ( .A(n267), .B(n268), .Y(n266) );
  XNOR2XL U133 ( .A(n252), .B(n251), .Y(n271) );
  AO33X1 U134 ( .A(n249), .B(n264), .C(ff_idn), .D(n261), .E(n260), .F(n52), 
        .Y(trans_buf[0]) );
  XNOR2XL U135 ( .A(n263), .B(n255), .Y(n267) );
  XNOR2XL U136 ( .A(n250), .B(n248), .Y(n272) );
  XNOR2XL U137 ( .A(n258), .B(n254), .Y(n268) );
  OAI21X1 U138 ( .B(n85), .C(n58), .A(n259), .Y(trans_buf[1]) );
  AOI32X1 U139 ( .A(n42), .B(n260), .C(n261), .D(n52), .E(n61), .Y(n259) );
  OAI211X1 U140 ( .C(n2), .D(n342), .A(n58), .B(n343), .Y(n256) );
  AOI21X1 U141 ( .B(n344), .C(n79), .A(n77), .Y(n343) );
  NOR2X1 U142 ( .A(n269), .B(n270), .Y(n249) );
  AOI22X1 U143 ( .A(n52), .B(n263), .C(n59), .D(n253), .Y(n247) );
  NOR2X1 U144 ( .A(n77), .B(n52), .Y(n253) );
  OAI222XL U145 ( .A(n255), .B(n256), .C(n254), .D(n257), .E(n86), .F(n58), 
        .Y(trans_buf[3]) );
  OAI222XL U146 ( .A(n254), .B(n256), .C(n258), .D(n257), .E(n82), .F(n58), 
        .Y(trans_buf[2]) );
  INVX1 U147 ( .A(n495), .Y(n39) );
  INVX1 U148 ( .A(n258), .Y(n61) );
  NOR32XL U149 ( .B(n281), .C(n278), .A(n280), .Y(n279) );
  OAI2B11X1 U150 ( .D(n264), .C(n40), .A(n79), .B(n346), .Y(n280) );
  AND2X1 U151 ( .A(N228), .B(n279), .Y(net9526) );
  NOR2X1 U152 ( .A(n383), .B(n121), .Y(N1259) );
  OAI22X1 U153 ( .A(n100), .B(n58), .C(n345), .D(n13), .Y(N260) );
  EORX1 U154 ( .A(n2), .B(n344), .C(n342), .D(n79), .Y(n345) );
  INVX1 U155 ( .A(n263), .Y(n59) );
  INVX1 U156 ( .A(n255), .Y(n60) );
  INVX1 U157 ( .A(n243), .Y(n83) );
  AOI31X1 U158 ( .A(ff_chg), .B(n244), .C(n245), .D(r_wr[4]), .Y(n243) );
  OAI22X1 U159 ( .A(r_wr[3]), .B(n85), .C(n80), .D(n21), .Y(upd_dbuf[0]) );
  OAI22X1 U160 ( .A(r_wr[3]), .B(n82), .C(n80), .D(n22), .Y(upd_dbuf[1]) );
  OAI22X1 U161 ( .A(r_wr[3]), .B(n86), .C(n80), .D(n24), .Y(upd_dbuf[2]) );
  OAI22X1 U162 ( .A(n36), .B(n81), .C(r_wr[4]), .D(n74), .Y(tui_wdat[7]) );
  OAI22X1 U163 ( .A(n21), .B(n81), .C(n166), .D(n155), .Y(tui_wdat[0]) );
  XNOR2XL U164 ( .A(n125), .B(n17), .Y(n166) );
  OAI211X1 U165 ( .C(n110), .D(n305), .A(n10), .B(n346), .Y(N22) );
  OAI21X1 U166 ( .B(n133), .C(n134), .A(n15), .Y(upd_dbuf_en) );
  NAND4X1 U167 ( .A(n146), .B(n147), .C(n148), .D(n149), .Y(n133) );
  NAND4X1 U168 ( .A(n135), .B(n136), .C(n137), .D(n138), .Y(n134) );
  NOR3XL U169 ( .A(n150), .B(n151), .C(n90), .Y(n149) );
  AOI21X1 U170 ( .B(n538), .C(n277), .A(r_wr[3]), .Y(N444) );
  INVX1 U171 ( .A(n334), .Y(n73) );
  INVX1 U172 ( .A(n153), .Y(n67) );
  AOI31X1 U173 ( .A(n543), .B(n126), .C(n276), .D(n408), .Y(n406) );
  INVX1 U174 ( .A(n330), .Y(n72) );
  INVX1 U175 ( .A(n291), .Y(n71) );
  OAI221X1 U176 ( .A(n56), .B(n423), .C(n424), .D(n54), .E(n425), .Y(n408) );
  AOI221XL U177 ( .A(n415), .B(n541), .C(n543), .D(n405), .E(n549), .Y(n423)
         );
  AOI221XL U178 ( .A(n473), .B(n474), .C(n421), .D(n419), .E(n475), .Y(n424)
         );
  AOI31X1 U179 ( .A(n296), .B(n541), .C(n98), .D(n426), .Y(n425) );
  OAI31XL U180 ( .A(n151), .B(n422), .C(n409), .D(n53), .Y(n426) );
  INVX1 U181 ( .A(n427), .Y(n53) );
  NOR2X1 U182 ( .A(n340), .B(n291), .Y(add_263_carry[1]) );
  AOI22X1 U183 ( .A(rx_ui_3_8[3]), .B(n124), .C(rx_ui_3_8[2]), .D(n122), .Y(
        n443) );
  ENOX1 U184 ( .A(n406), .B(n119), .C(n27), .D(n407), .Y(N1015) );
  ENOX1 U185 ( .A(n406), .B(n116), .C(n28), .D(n407), .Y(N1014) );
  ENOX1 U186 ( .A(n406), .B(n128), .C(n30), .D(n407), .Y(N1012) );
  ENOX1 U187 ( .A(n406), .B(n131), .C(n31), .D(n407), .Y(N1011) );
  INVX1 U188 ( .A(n445), .Y(n63) );
  NOR32XL U189 ( .B(n204), .C(n205), .A(n208), .Y(n213) );
  NAND31X1 U190 ( .C(n172), .A(n171), .B(n174), .Y(n162) );
  AOI33X1 U191 ( .A(n175), .B(n176), .C(n177), .D(n101), .E(n102), .F(n178), 
        .Y(n174) );
  AOI22X1 U192 ( .A(n157), .B(n179), .C(n104), .D(n157), .Y(n178) );
  INVX1 U193 ( .A(n169), .Y(n102) );
  XNOR2XL U194 ( .A(n218), .B(n238), .Y(n204) );
  XNOR2XL U195 ( .A(n231), .B(n232), .Y(n238) );
  OAI22X1 U196 ( .A(n206), .B(n20), .C(n106), .D(n207), .Y(n175) );
  AOI21X1 U197 ( .B(n203), .C(n202), .A(n210), .Y(n206) );
  XNOR2XL U198 ( .A(n208), .B(n209), .Y(n207) );
  NAND2X1 U199 ( .A(n205), .B(n204), .Y(n209) );
  OAI211X1 U200 ( .C(n409), .D(n305), .A(n410), .B(n411), .Y(n407) );
  AOI31X1 U201 ( .A(ff_idn), .B(n419), .C(n89), .D(n363), .Y(n410) );
  AOI22AXL U202 ( .A(n412), .B(n413), .D(n414), .C(n56), .Y(n411) );
  INVX1 U203 ( .A(n421), .Y(n89) );
  OAI211X1 U204 ( .C(n167), .D(n168), .A(n169), .B(n170), .Y(n154) );
  OAI31XL U205 ( .A(n173), .B(n159), .C(n160), .D(n103), .Y(n168) );
  NOR21XL U206 ( .B(n171), .A(n172), .Y(n170) );
  OAI21X1 U207 ( .B(n232), .C(n237), .A(n240), .Y(n233) );
  OAI21BBX1 U208 ( .A(n237), .B(n232), .C(N107), .Y(n240) );
  OAI22X1 U209 ( .A(n106), .B(n200), .C(n20), .D(n201), .Y(n176) );
  XNOR2XL U210 ( .A(n202), .B(n203), .Y(n201) );
  XNOR2XL U211 ( .A(n204), .B(n205), .Y(n200) );
  NAND2X1 U212 ( .A(n129), .B(n404), .Y(n235) );
  INVX1 U213 ( .A(n375), .Y(n132) );
  NAND2X1 U214 ( .A(n235), .B(n537), .Y(n237) );
  INVX1 U215 ( .A(n405), .Y(n129) );
  NOR32XL U216 ( .B(add_274_carry[8]), .C(n193), .A(n196), .Y(n205) );
  NOR21XL U217 ( .B(n231), .A(n232), .Y(n215) );
  XNOR2XL U218 ( .A(N107), .B(n236), .Y(n193) );
  XNOR2XL U219 ( .A(n232), .B(n237), .Y(n236) );
  OAI21X1 U220 ( .B(n241), .C(n116), .A(n230), .Y(n216) );
  INVX1 U221 ( .A(n333), .Y(n68) );
  NOR2X1 U222 ( .A(n504), .B(n505), .Y(n492) );
  NOR2X1 U223 ( .A(n131), .B(n537), .Y(n418) );
  OAI22X1 U224 ( .A(n106), .B(n190), .C(n20), .D(n191), .Y(n181) );
  XNOR2XL U225 ( .A(add_274_2_carry[8]), .B(n192), .Y(n191) );
  XNOR2XL U226 ( .A(add_274_carry[8]), .B(n193), .Y(n190) );
  NOR2X1 U227 ( .A(n107), .B(n71), .Y(n339) );
  OAI22X1 U228 ( .A(n20), .B(n194), .C(n106), .D(n195), .Y(n186) );
  XNOR2XL U229 ( .A(n198), .B(n199), .Y(n194) );
  XNOR2XL U230 ( .A(n196), .B(n197), .Y(n195) );
  NAND2X1 U231 ( .A(add_274_2_carry[8]), .B(n192), .Y(n199) );
  NAND2X1 U232 ( .A(n382), .B(n100), .Y(n372) );
  OAI21X1 U233 ( .B(n126), .C(n372), .A(n380), .Y(n369) );
  AOI21X1 U234 ( .B(n117), .C(n69), .A(add_263_carry[1]), .Y(n327) );
  INVX1 U235 ( .A(n340), .Y(n69) );
  INVX1 U236 ( .A(n380), .Y(n115) );
  NAND2X1 U237 ( .A(n241), .B(n116), .Y(n230) );
  NAND2X1 U238 ( .A(n119), .B(n116), .Y(n274) );
  OAI221X1 U239 ( .A(n275), .B(n112), .C(n40), .D(n293), .E(n310), .Y(n307) );
  NAND4X1 U240 ( .A(n311), .B(n121), .C(n312), .D(n313), .Y(n310) );
  AOI32X1 U241 ( .A(n319), .B(n120), .C(n320), .D(n151), .E(n282), .Y(n312) );
  NOR3XL U242 ( .A(n309), .B(n314), .C(n40), .Y(n313) );
  INVX1 U243 ( .A(n518), .Y(n114) );
  NAND2X1 U244 ( .A(add_274_carry[8]), .B(n193), .Y(n197) );
  NAND2X1 U245 ( .A(n382), .B(n130), .Y(n373) );
  NOR2X1 U246 ( .A(n115), .B(n360), .Y(n351) );
  INVX1 U247 ( .A(n347), .Y(n95) );
  OAI31XL U248 ( .A(n348), .B(n96), .C(n349), .D(n350), .Y(n347) );
  AOI33X1 U249 ( .A(n351), .B(n352), .C(n353), .D(n354), .E(n355), .F(n99), 
        .Y(n350) );
  INVX1 U250 ( .A(n356), .Y(n99) );
  NOR32XL U251 ( .B(n494), .C(n552), .A(n551), .Y(n245) );
  NOR32XL U252 ( .B(add_274_2_carry[8]), .C(n192), .A(n198), .Y(n203) );
  XNOR2XL U253 ( .A(n225), .B(n126), .Y(n202) );
  XNOR2XL U254 ( .A(n20), .B(n189), .Y(n164) );
  AOI21X1 U255 ( .B(n537), .C(n123), .A(add_274_2_carry[6]), .Y(n189) );
  XNOR2XL U256 ( .A(adp_tx_1_4[5]), .B(n123), .Y(n469) );
  NOR2X1 U257 ( .A(n383), .B(n122), .Y(N1254) );
  NOR2X1 U258 ( .A(n383), .B(n17), .Y(N1255) );
  NOR2X1 U259 ( .A(n383), .B(n125), .Y(N1256) );
  NOR2X1 U260 ( .A(n383), .B(n123), .Y(N1257) );
  NOR2X1 U261 ( .A(n383), .B(n117), .Y(N1253) );
  XNOR2XL U262 ( .A(adp_tx_1_4[6]), .B(n120), .Y(n470) );
  XNOR2XL U263 ( .A(adp_tx_1_4[4]), .B(n125), .Y(n468) );
  XNOR2XL U264 ( .A(adp_tx_1_4[3]), .B(n124), .Y(n467) );
  AOI22X1 U265 ( .A(N172), .B(n106), .C(N144), .D(n20), .Y(n182) );
  NOR2X1 U266 ( .A(n383), .B(n120), .Y(N1258) );
  XNOR2XL U267 ( .A(n120), .B(adp_tx_ui_6_), .Y(n528) );
  NOR3XL U268 ( .A(n538), .B(n95), .C(n276), .Y(setsta[0]) );
  NAND3X1 U269 ( .A(n552), .B(n551), .C(n494), .Y(n293) );
  INVX1 U270 ( .A(n151), .Y(n545) );
  NOR2X1 U271 ( .A(n383), .B(n107), .Y(N1252) );
  NOR3XL U272 ( .A(n124), .B(n125), .C(n164), .Y(n183) );
  AND2X1 U273 ( .A(n230), .B(n119), .Y(n218) );
  AOI22X1 U274 ( .A(N173), .B(n106), .C(N145), .D(n20), .Y(n184) );
  INVX1 U275 ( .A(n277), .Y(n4) );
  AOI221XL U276 ( .A(n73), .B(n545), .C(n393), .D(n75), .E(n245), .Y(n396) );
  NOR31X1 U277 ( .C(n357), .A(n358), .B(n359), .Y(n353) );
  INVX1 U278 ( .A(n504), .Y(n110) );
  NOR2X1 U279 ( .A(n537), .B(n123), .Y(add_274_2_carry[6]) );
  NOR2X1 U280 ( .A(n100), .B(n537), .Y(n358) );
  NAND2X1 U281 ( .A(n376), .B(n377), .Y(n354) );
  NOR2X1 U282 ( .A(n291), .B(n144), .Y(add_264_carry[1]) );
  XNOR2XL U283 ( .A(n220), .B(n127), .Y(n198) );
  XNOR2XL U284 ( .A(n116), .B(n128), .Y(n220) );
  NOR21XL U285 ( .B(n459), .A(n460), .Y(n454) );
  XNOR2XL U286 ( .A(n124), .B(n72), .Y(n460) );
  XNOR2XL U287 ( .A(n120), .B(n68), .Y(n141) );
  XNOR2XL U288 ( .A(n145), .B(n121), .Y(n135) );
  NAND21X1 U289 ( .B(n142), .A(n68), .Y(n145) );
  XNOR2XL U290 ( .A(n125), .B(n73), .Y(n458) );
  XNOR2XL U291 ( .A(adp_tx_1_4[1]), .B(n117), .Y(n471) );
  XNOR2XL U292 ( .A(adp_tx_ui_7_), .B(n121), .Y(n530) );
  XNOR2XL U293 ( .A(n123), .B(n75), .Y(n529) );
  NOR2X1 U294 ( .A(n305), .B(n150), .Y(n536) );
  NAND2X1 U295 ( .A(n366), .B(n131), .Y(n309) );
  NAND4X1 U296 ( .A(n122), .B(n123), .C(n17), .D(n480), .Y(n421) );
  NOR2X1 U297 ( .A(n120), .B(n478), .Y(n480) );
  NAND2X1 U298 ( .A(n56), .B(n349), .Y(n509) );
  NOR3XL U299 ( .A(n333), .B(n153), .C(n334), .Y(n315) );
  ENOX1 U300 ( .A(n153), .B(n151), .C(adp_tx_ui_6_), .D(n393), .Y(n401) );
  NOR3XL U301 ( .A(n415), .B(n420), .C(n296), .Y(n363) );
  INVX1 U302 ( .A(n20), .Y(n106) );
  INVX1 U303 ( .A(n276), .Y(n56) );
  NOR3XL U304 ( .A(n282), .B(n476), .C(n413), .Y(n475) );
  NAND2X1 U305 ( .A(n422), .B(n545), .Y(n305) );
  NOR2X1 U306 ( .A(n355), .B(n276), .Y(n487) );
  NAND2X1 U307 ( .A(n334), .B(n17), .Y(n328) );
  NOR2X1 U308 ( .A(n139), .B(n140), .Y(n137) );
  XNOR2XL U309 ( .A(rx_ui_5_8[3]), .B(n17), .Y(n139) );
  XNOR2XL U310 ( .A(n141), .B(n142), .Y(n140) );
  INVX1 U311 ( .A(n281), .Y(n90) );
  NAND2X1 U312 ( .A(n116), .B(n217), .Y(n210) );
  INVX1 U313 ( .A(n227), .Y(n127) );
  INVX1 U314 ( .A(n428), .Y(n112) );
  INVX1 U315 ( .A(n415), .Y(n98) );
  INVX1 U316 ( .A(ff_chg), .Y(n40) );
  XNOR2XL U317 ( .A(adp_tx_1_4[0]), .B(n107), .Y(n472) );
  XNOR2XL U318 ( .A(n117), .B(n69), .Y(n456) );
  NOR4XL U319 ( .A(n130), .B(n110), .C(n276), .D(n128), .Y(n486) );
  AND2X1 U320 ( .A(n534), .B(n115), .Y(n283) );
  NAND4X1 U321 ( .A(n404), .B(n126), .C(n119), .D(n118), .Y(n534) );
  OAI22X1 U322 ( .A(n479), .B(n283), .C(n473), .D(n539), .Y(n419) );
  INVX1 U323 ( .A(n479), .Y(n548) );
  INVX1 U324 ( .A(n217), .Y(n108) );
  NOR21XL U325 ( .B(n496), .A(n497), .Y(n488) );
  INVX1 U326 ( .A(ff_idn), .Y(n54) );
  OAI21X1 U327 ( .B(n126), .C(n128), .A(n380), .Y(n285) );
  NOR2X1 U328 ( .A(n377), .B(n150), .Y(n497) );
  OAI211X1 U329 ( .C(n55), .D(n376), .A(n502), .B(n503), .Y(n484) );
  NAND4X1 U330 ( .A(ff_idn), .B(n492), .C(n545), .D(n112), .Y(n503) );
  OAI31XL U331 ( .A(n276), .B(n504), .C(n113), .D(n543), .Y(n502) );
  NOR3XL U332 ( .A(n54), .B(n476), .C(n282), .Y(n412) );
  NAND2X1 U333 ( .A(ff_chg), .B(n545), .Y(n275) );
  OAI21BBX1 U334 ( .A(n56), .B(n497), .C(n496), .Y(n513) );
  INVX1 U335 ( .A(n474), .Y(n539) );
  NAND21X1 U336 ( .B(n285), .A(n222), .Y(n244) );
  NAND3X1 U337 ( .A(n545), .B(n244), .C(ff_idn), .Y(n278) );
  INVX1 U338 ( .A(n282), .Y(n547) );
  OAI21X1 U339 ( .B(n94), .C(n93), .A(n293), .Y(n286) );
  INVX1 U340 ( .A(n352), .Y(n540) );
  AOI21X1 U341 ( .B(n93), .C(n94), .A(n286), .Y(n461) );
  NOR2X1 U342 ( .A(n40), .B(n282), .Y(n526) );
  NOR3XL U343 ( .A(n533), .B(fcp_state[1]), .C(n544), .Y(n352) );
  INVX1 U344 ( .A(fcp_state[0]), .Y(n552) );
  NAND2X1 U345 ( .A(fcp_state[3]), .B(n552), .Y(n533) );
  NOR32XL U346 ( .B(fcp_state[0]), .C(fcp_state[3]), .A(fcp_state[2]), .Y(n535) );
  NAND2X1 U347 ( .A(n535), .B(fcp_state[1]), .Y(n376) );
  INVX1 U348 ( .A(fcp_state[1]), .Y(n551) );
  INVX1 U349 ( .A(fcp_state[2]), .Y(n544) );
  AOI22X1 U350 ( .A(r_wdat[1]), .B(n269), .C(r_dat[1]), .D(n270), .Y(n254) );
  AOI22X1 U351 ( .A(r_wdat[7]), .B(n269), .C(n270), .D(r_dat[7]), .Y(n263) );
  AOI22X1 U352 ( .A(r_wdat[0]), .B(n269), .C(r_dat[0]), .D(n270), .Y(n258) );
  AOI22X1 U353 ( .A(n23), .B(n269), .C(r_dat[2]), .D(n270), .Y(n255) );
  ENOX1 U354 ( .A(n35), .B(n79), .C(r_dat[6]), .D(n270), .Y(n251) );
  ENOX1 U355 ( .A(n33), .B(n79), .C(r_dat[4]), .D(n270), .Y(n250) );
  ENOX1 U356 ( .A(n25), .B(n79), .C(r_dat[3]), .D(n270), .Y(n252) );
  ENOX1 U357 ( .A(n34), .B(n79), .C(r_dat[5]), .D(n270), .Y(n248) );
  OAI32X1 U358 ( .A(n76), .B(n512), .C(n79), .D(r_ctl[7]), .E(n514), .Y(n495)
         );
  INVX1 U359 ( .A(r_ctl[4]), .Y(n76) );
  AOI22X1 U360 ( .A(n487), .B(n352), .C(n55), .D(n550), .Y(n514) );
  AO2222XL U361 ( .A(n249), .B(rxtx_buf[5]), .C(n52), .D(n248), .E(n60), .F(
        n77), .G(n253), .H(n250), .Y(trans_buf[6]) );
  AO2222XL U362 ( .A(n249), .B(rxtx_buf[4]), .C(n52), .D(n250), .E(n62), .F(
        n77), .G(n253), .H(n252), .Y(trans_buf[5]) );
  INVX1 U363 ( .A(n254), .Y(n62) );
  AO2222XL U364 ( .A(n249), .B(rxtx_buf[7]), .C(n250), .D(n77), .E(n52), .F(
        n59), .G(n42), .H(n251), .Y(trans_buf[8]) );
  AO2222XL U365 ( .A(n249), .B(rxtx_buf[6]), .C(n252), .D(n77), .E(n52), .F(
        n251), .G(n253), .H(n248), .Y(trans_buf[7]) );
  AO2222XL U366 ( .A(rxtx_buf[9]), .B(n249), .C(n251), .D(n77), .E(n52), .F(
        n59), .G(n42), .H(n263), .Y(trans_buf[10]) );
  AO2222XL U367 ( .A(n249), .B(rxtx_buf[3]), .C(n52), .D(n252), .E(n61), .F(
        n77), .G(n253), .H(n60), .Y(trans_buf[4]) );
  NAND32X1 U368 ( .B(n498), .C(n484), .A(n499), .Y(N1007) );
  AOI32X1 U369 ( .A(n547), .B(ff_idn), .C(n476), .D(n500), .E(n501), .Y(n499)
         );
  OAI21BBX1 U370 ( .A(n77), .B(r_ctl[1]), .C(n260), .Y(n501) );
  GEN2XL U371 ( .D(n486), .E(n549), .C(n497), .B(n538), .A(n495), .Y(n500) );
  NAND4X1 U372 ( .A(n287), .B(n288), .C(n289), .D(n290), .Y(intr) );
  AOI22X1 U373 ( .A(r_msk[2]), .B(r_irq[2]), .C(r_msk[3]), .D(r_irq[3]), .Y(
        n289) );
  AOI22X1 U374 ( .A(r_msk[4]), .B(r_irq[4]), .C(r_msk[5]), .D(r_irq[5]), .Y(
        n288) );
  AOI22X1 U375 ( .A(r_msk[6]), .B(r_irq[6]), .C(r_msk[7]), .D(r_irq[7]), .Y(
        n287) );
  OAI221X1 U376 ( .A(n487), .B(n540), .C(n54), .D(n539), .E(n489), .Y(N1008)
         );
  AOI31X1 U377 ( .A(r_ctl[0]), .B(n490), .C(r_ctl[1]), .D(n427), .Y(n489) );
  OAI31XL U378 ( .A(n276), .B(r_ctl[7]), .C(n488), .D(n39), .Y(n490) );
  OAI211X1 U379 ( .C(r_ctl[1]), .D(n506), .A(n507), .B(n508), .Y(N1006) );
  AOI31X1 U380 ( .A(r_ctl[4]), .B(n546), .C(n512), .D(n412), .Y(n507) );
  AOI221XL U381 ( .A(n549), .B(n57), .C(n550), .D(n509), .E(n498), .Y(n508) );
  AOI21X1 U382 ( .B(n513), .C(n538), .A(n495), .Y(n506) );
  NAND2X1 U383 ( .A(n262), .B(n247), .Y(trans_buf[11]) );
  AOI22X1 U384 ( .A(n59), .B(n13), .C(rxtx_buf[10]), .D(n249), .Y(n262) );
  NAND2X1 U385 ( .A(n246), .B(n247), .Y(trans_buf[9]) );
  AOI22X1 U386 ( .A(n248), .B(n13), .C(rxtx_buf[8]), .D(n249), .Y(n246) );
  NAND31X1 U387 ( .C(n484), .A(n39), .B(n485), .Y(N1009) );
  OA222X1 U388 ( .A(n348), .B(n486), .C(n540), .D(n487), .E(n488), .F(r_ctl[7]), .Y(n485) );
  OAI21BBX1 U389 ( .A(N363), .B(n10), .C(n256), .Y(N261) );
  OAI22X1 U390 ( .A(n22), .B(n81), .C(n155), .D(n163), .Y(tui_wdat[1]) );
  XNOR2XL U391 ( .A(n164), .B(n165), .Y(n163) );
  NAND2X1 U392 ( .A(N141), .B(N142), .Y(n165) );
  ENOX1 U393 ( .A(n15), .B(n34), .C(n80), .D(rxtx_buf[5]), .Y(upd_dbuf[5]) );
  ENOX1 U394 ( .A(n15), .B(n25), .C(n80), .D(rxtx_buf[3]), .Y(upd_dbuf[3]) );
  ENOX1 U395 ( .A(n15), .B(n33), .C(n80), .D(rxtx_buf[4]), .Y(upd_dbuf[4]) );
  ENOX1 U396 ( .A(n15), .B(n35), .C(n80), .D(rxtx_buf[6]), .Y(upd_dbuf[6]) );
  ENOX1 U397 ( .A(n36), .B(n80), .C(n80), .D(rxtx_buf[7]), .Y(upd_dbuf[7]) );
  OAI22X1 U398 ( .A(r_tui[7]), .B(n75), .C(catch_sync[3]), .D(n74), .Y(n334)
         );
  OAI22X1 U399 ( .A(r_tui[7]), .B(r_tui[3]), .C(catch_sync[1]), .D(n74), .Y(
        n291) );
  OAI22X1 U400 ( .A(catch_sync[4]), .B(n74), .C(r_tui[7]), .D(adp_tx_ui_6_), 
        .Y(n153) );
  OAI22X1 U401 ( .A(r_tui[7]), .B(r_tui[4]), .C(catch_sync[2]), .D(n74), .Y(
        n330) );
  OAI22X1 U402 ( .A(r_tui[7]), .B(r_tui[2]), .C(catch_sync[0]), .D(n74), .Y(
        n340) );
  OAI21X1 U403 ( .B(r_tui[6]), .C(n75), .A(adp_tx_ui_7_), .Y(adp_tx_ui_6_) );
  AO22X1 U404 ( .A(n408), .B(n14), .C(n29), .D(n407), .Y(N1013) );
  INVX1 U405 ( .A(r_tui[7]), .Y(n74) );
  INVX1 U406 ( .A(r_tui[5]), .Y(n75) );
  NAND2X1 U407 ( .A(n449), .B(ui_intv_cnt[5]), .Y(n445) );
  NAND2X1 U408 ( .A(r_tui[6]), .B(n75), .Y(adp_tx_ui_7_) );
  OAI221X1 U409 ( .A(rx_ui_3_8[3]), .B(n124), .C(rx_ui_3_8[2]), .D(n122), .E(
        n446), .Y(n444) );
  NOR2X1 U410 ( .A(ui_intv_cnt[0]), .B(n448), .Y(n447) );
  XNOR2XL U411 ( .A(n69), .B(n71), .Y(n448) );
  AOI32X1 U412 ( .A(n428), .B(n88), .C(n87), .D(n111), .E(n429), .Y(n409) );
  OR4X1 U413 ( .A(n430), .B(n431), .C(n40), .D(n84), .Y(n429) );
  OAI31XL U414 ( .A(n432), .B(ui_intv_cnt[6]), .C(ui_intv_cnt[5]), .D(n110), 
        .Y(n431) );
  AOI21BX1 U415 ( .C(n439), .B(n440), .A(n441), .Y(n430) );
  OAI21X1 U416 ( .B(ui_intv_cnt[5]), .C(n449), .A(n450), .Y(n440) );
  AOI33X1 U417 ( .A(n445), .B(n125), .C(rx_ui_3_8[4]), .D(n68), .E(n120), .F(
        add_263_carry[5]), .Y(n450) );
  AOI211X1 U418 ( .C(N142), .D(n64), .A(n442), .B(n439), .Y(n441) );
  INVX1 U419 ( .A(rx_ui_3_8[4]), .Y(n64) );
  GEN2XL U420 ( .D(N141), .E(n65), .C(n443), .B(n444), .A(n63), .Y(n442) );
  INVX1 U421 ( .A(rx_ui_3_8[3]), .Y(n65) );
  ENOX1 U422 ( .A(n406), .B(n118), .C(n26), .D(n407), .Y(N1016) );
  ENOX1 U423 ( .A(n406), .B(n537), .C(n32), .D(n407), .Y(N1010) );
  NOR21XL U424 ( .B(n211), .A(n212), .Y(n171) );
  OAI31XL U425 ( .A(n213), .B(n106), .C(n214), .D(n118), .Y(n212) );
  AOI33X1 U426 ( .A(n106), .B(n108), .C(symb_cnt[4]), .D(n214), .E(n20), .F(
        n213), .Y(n211) );
  NAND2X1 U427 ( .A(n215), .B(n216), .Y(n214) );
  AOI21X1 U428 ( .B(n129), .C(symb_cnt[3]), .A(n241), .Y(n232) );
  NOR2X1 U429 ( .A(n132), .B(symb_cnt[2]), .Y(n405) );
  NOR2X1 U430 ( .A(N159), .B(N160), .Y(n375) );
  NAND2X1 U431 ( .A(n121), .B(n451), .Y(n439) );
  OAI21BBX1 U432 ( .A(n68), .B(add_263_carry[5]), .C(ui_intv_cnt[6]), .Y(n451)
         );
  NOR2X1 U433 ( .A(n129), .B(symb_cnt[3]), .Y(n241) );
  NAND2X1 U434 ( .A(symb_cnt[2]), .B(n132), .Y(n404) );
  XNOR2XL U435 ( .A(N159), .B(n235), .Y(N108) );
  GEN2XL U436 ( .D(n515), .E(n373), .C(symb_cnt[2]), .B(symb_cnt[3]), .A(n369), 
        .Y(n349) );
  NAND21X1 U437 ( .B(n358), .A(n131), .Y(n515) );
  XNOR2XL U438 ( .A(N363), .B(n9), .Y(n382) );
  OAI22X1 U439 ( .A(catch_sync[5]), .B(n74), .C(r_tui[7]), .D(adp_tx_ui_7_), 
        .Y(n333) );
  XOR2X1 U440 ( .A(n215), .B(n229), .Y(n208) );
  OAI21X1 U441 ( .B(n230), .C(symb_cnt[5]), .A(n216), .Y(n229) );
  INVX1 U442 ( .A(N159), .Y(n537) );
  AOI21BBXL U443 ( .B(n337), .C(n72), .A(n338), .Y(n336) );
  AOI21X1 U444 ( .B(n72), .C(n337), .A(n122), .Y(n338) );
  OAI221X1 U445 ( .A(ui_intv_cnt[1]), .B(n339), .C(ui_intv_cnt[0]), .D(n291), 
        .E(n327), .Y(n337) );
  INVX1 U446 ( .A(N160), .Y(n131) );
  OAI32X1 U447 ( .A(n218), .B(n106), .C(n213), .D(n219), .E(n20), .Y(n172) );
  AOI31X1 U448 ( .A(n202), .B(n210), .C(n203), .D(symb_cnt[5]), .Y(n219) );
  NOR3XL U449 ( .A(n95), .B(r_ctl[7]), .C(n276), .Y(n270) );
  INVX1 U450 ( .A(n367), .Y(n96) );
  GEN2XL U451 ( .D(n97), .E(symb_cnt[2]), .C(symb_cnt[3]), .B(n368), .A(n369), 
        .Y(n367) );
  INVX1 U452 ( .A(n372), .Y(n97) );
  NAND2X1 U453 ( .A(n370), .B(n371), .Y(n368) );
  NOR2X1 U454 ( .A(n274), .B(symb_cnt[6]), .Y(n380) );
  NOR2X1 U455 ( .A(n115), .B(symb_cnt[2]), .Y(n518) );
  INVX1 U456 ( .A(symb_cnt[4]), .Y(n116) );
  OAI211X1 U457 ( .C(n517), .D(n114), .A(n378), .B(n492), .Y(n355) );
  AOI22X1 U458 ( .A(N363), .B(n130), .C(N362), .D(n131), .Y(n517) );
  OAI21X1 U459 ( .B(N160), .C(symb_cnt[2]), .A(n372), .Y(n371) );
  OAI21X1 U460 ( .B(N362), .C(N159), .A(n373), .Y(n370) );
  INVX1 U461 ( .A(symb_cnt[5]), .Y(n119) );
  OAI32X1 U462 ( .A(n87), .B(new_rx_sync_cnt[1]), .C(n37), .D(n306), .E(n88), 
        .Y(N349) );
  AOI21X1 U463 ( .B(n307), .C(n87), .A(n308), .Y(n306) );
  OAI22X1 U464 ( .A(N141), .B(n153), .C(ui_intv_cnt[2]), .D(n334), .Y(n437) );
  OAI21BBX1 U465 ( .A(n331), .B(n315), .C(n332), .Y(n311) );
  OAI21X1 U466 ( .B(n315), .C(n331), .A(n120), .Y(n332) );
  OAI221X1 U467 ( .A(N142), .B(n318), .C(ui_intv_cnt[5]), .D(n66), .E(n335), 
        .Y(n331) );
  OAI22AX1 U468 ( .D(n328), .C(n336), .A(n17), .B(n334), .Y(n335) );
  OAI21X1 U469 ( .B(n68), .C(n125), .A(n433), .Y(n432) );
  OAI22X1 U470 ( .A(N142), .B(n333), .C(n434), .D(n435), .Y(n433) );
  AOI21X1 U471 ( .B(n67), .C(n124), .A(n436), .Y(n435) );
  AOI211X1 U472 ( .C(n72), .D(n70), .A(n437), .B(n438), .Y(n434) );
  NAND3X1 U473 ( .A(n110), .B(n378), .C(n379), .Y(n360) );
  NAND41X1 U474 ( .D(n359), .A(n380), .B(n381), .C(n357), .Y(n379) );
  OAI22X1 U475 ( .A(N362), .B(N159), .C(N160), .D(n382), .Y(n381) );
  AOI22X1 U476 ( .A(N141), .B(n153), .C(ui_intv_cnt[2]), .D(n334), .Y(n436) );
  AOI21X1 U477 ( .B(n339), .C(n330), .A(ui_intv_cnt[1]), .Y(n438) );
  NAND3X1 U478 ( .A(N362), .B(n518), .C(N363), .Y(n378) );
  NAND2X1 U479 ( .A(n382), .B(N160), .Y(n357) );
  XNOR2XL U480 ( .A(n537), .B(symb_cnt[2]), .Y(N161) );
  NOR2X1 U481 ( .A(N159), .B(n123), .Y(add_274_carry[6]) );
  AND4X1 U482 ( .A(n384), .B(n385), .C(n386), .D(n387), .Y(n383) );
  XNOR2XL U483 ( .A(n402), .B(n107), .Y(n384) );
  XNOR2XL U484 ( .A(ui_intv_cnt[6]), .B(n401), .Y(n385) );
  NOR2X1 U485 ( .A(n397), .B(n398), .Y(n386) );
  OAI21X1 U486 ( .B(n228), .C(n221), .A(n222), .Y(n227) );
  NOR2X1 U487 ( .A(N160), .B(symb_cnt[3]), .Y(n228) );
  OAI31XL U488 ( .A(n114), .B(n365), .C(n374), .D(n110), .Y(n356) );
  AOI21X1 U489 ( .B(N362), .C(n537), .A(n131), .Y(n374) );
  OAI211X1 U490 ( .C(n56), .D(n541), .A(n109), .B(n294), .Y(n277) );
  AOI211X1 U491 ( .C(n295), .D(n296), .A(n16), .B(n264), .Y(n294) );
  INVX1 U492 ( .A(N141), .Y(n124) );
  NAND3X1 U493 ( .A(fcp_state[0]), .B(n494), .C(fcp_state[1]), .Y(n151) );
  INVX1 U494 ( .A(ui_intv_cnt[5]), .Y(n123) );
  XNOR2XL U495 ( .A(n392), .B(n122), .Y(n391) );
  ENOX1 U496 ( .A(n151), .B(n340), .C(r_tui[2]), .D(n393), .Y(n392) );
  NOR3XL U497 ( .A(n292), .B(us_cnt_2_), .C(n91), .Y(n281) );
  NAND4X1 U498 ( .A(n519), .B(n281), .C(n520), .D(n521), .Y(n276) );
  XNOR2XL U499 ( .A(n7), .B(r_tui[2]), .Y(n519) );
  NOR4XL U500 ( .A(n522), .B(n523), .C(n524), .D(n527), .Y(n521) );
  NOR3XL U501 ( .A(n528), .B(n529), .C(n530), .Y(n520) );
  OAI21X1 U502 ( .B(n221), .C(n222), .A(n223), .Y(n192) );
  AOI32X1 U503 ( .A(n221), .B(n131), .C(symb_cnt[3]), .D(n224), .E(n126), .Y(
        n223) );
  XNOR2XL U504 ( .A(N160), .B(n221), .Y(n224) );
  NOR2X1 U505 ( .A(n115), .B(symb_cnt[3]), .Y(n504) );
  INVX1 U506 ( .A(symb_cnt[2]), .Y(n128) );
  INVX1 U507 ( .A(ui_intv_cnt[1]), .Y(n117) );
  BUFX3 U508 ( .A(n188), .Y(n20) );
  GEN2XL U509 ( .D(N142), .E(n242), .C(ui_intv_cnt[5]), .B(ui_intv_cnt[6]), 
        .A(ui_intv_cnt[7]), .Y(n188) );
  NAND4X1 U510 ( .A(n124), .B(n107), .C(n117), .D(n122), .Y(n242) );
  INVX1 U511 ( .A(ui_intv_cnt[2]), .Y(n122) );
  OAI22X1 U512 ( .A(n127), .B(n128), .C(n226), .D(n116), .Y(n225) );
  NOR2X1 U513 ( .A(symb_cnt[2]), .B(n227), .Y(n226) );
  INVX1 U514 ( .A(ui_intv_cnt[0]), .Y(n107) );
  INVX1 U515 ( .A(N362), .Y(n100) );
  AOI22X1 U516 ( .A(r_msk[0]), .B(r_irq[0]), .C(r_msk[1]), .D(r_irq[1]), .Y(
        n290) );
  AOI21X1 U517 ( .B(N362), .C(N363), .A(n128), .Y(n359) );
  AOI21X1 U518 ( .B(n375), .C(N362), .A(N363), .Y(n365) );
  ENOX1 U519 ( .A(n144), .B(n151), .C(r_tui[1]), .D(n393), .Y(n395) );
  ENOX1 U520 ( .A(n291), .B(n151), .C(r_tui[3]), .D(n393), .Y(n394) );
  NOR2X1 U521 ( .A(fcp_state[2]), .B(fcp_state[3]), .Y(n494) );
  NOR4XL U522 ( .A(n388), .B(n389), .C(n390), .D(n391), .Y(n387) );
  XNOR2XL U523 ( .A(ui_intv_cnt[5]), .B(n396), .Y(n388) );
  XNOR2XL U524 ( .A(n395), .B(n117), .Y(n389) );
  XNOR2XL U525 ( .A(n394), .B(n124), .Y(n390) );
  NAND2X1 U526 ( .A(symb_cnt[2]), .B(N159), .Y(n221) );
  NAND4X1 U527 ( .A(n463), .B(n459), .C(n465), .D(n466), .Y(n296) );
  XNOR2XL U528 ( .A(ui_intv_cnt[2]), .B(adp_tx_1_4[2]), .Y(n463) );
  NOR2X1 U529 ( .A(n471), .B(n472), .Y(n465) );
  NOR4XL U530 ( .A(n467), .B(n468), .C(n469), .D(n470), .Y(n466) );
  AOI221XL U531 ( .A(n315), .B(n120), .C(n316), .D(n123), .E(n317), .Y(n314)
         );
  AOI22X1 U532 ( .A(n66), .B(ui_intv_cnt[5]), .C(n318), .D(N142), .Y(n317) );
  ENOX1 U533 ( .A(new_rx_sync_cnt[0]), .B(n37), .C(new_rx_sync_cnt[0]), .D(
        n308), .Y(N348) );
  NAND3X1 U534 ( .A(us_cnt_0_), .B(n293), .C(us_cnt_1_), .Y(n292) );
  NOR43XL U535 ( .B(n477), .C(n120), .D(ui_intv_cnt[2]), .A(n478), .Y(n413) );
  XNOR2XL U536 ( .A(n123), .B(n124), .Y(n477) );
  AOI22AXL U537 ( .A(n482), .B(n109), .D(n483), .C(N363), .Y(n415) );
  AOI21X1 U538 ( .B(n366), .C(n482), .A(n109), .Y(n483) );
  NAND2X1 U539 ( .A(N159), .B(n100), .Y(n482) );
  XNOR2XL U540 ( .A(n152), .B(n153), .Y(n148) );
  XNOR2XL U541 ( .A(n11), .B(add_264_carry[5]), .Y(n152) );
  AND4X1 U542 ( .A(n452), .B(n453), .C(n454), .D(n455), .Y(n422) );
  XNOR2XL U543 ( .A(n71), .B(ui_intv_cnt[2]), .Y(n453) );
  XNOR2XL U544 ( .A(n67), .B(ui_intv_cnt[5]), .Y(n452) );
  NOR4XL U545 ( .A(n456), .B(n457), .C(n458), .D(n141), .Y(n455) );
  XNOR2XL U546 ( .A(n117), .B(r_tui[1]), .Y(n524) );
  XNOR2XL U547 ( .A(ui_intv_cnt[7]), .B(n399), .Y(n398) );
  AOI221XL U548 ( .A(n545), .B(n68), .C(n393), .D(adp_tx_ui_7_), .E(n245), .Y(
        n399) );
  XNOR2XL U549 ( .A(n125), .B(r_tui[4]), .Y(n527) );
  XNOR2XL U550 ( .A(n400), .B(n125), .Y(n397) );
  ENOX1 U551 ( .A(n151), .B(n330), .C(r_tui[4]), .D(n393), .Y(n400) );
  XNOR2XL U552 ( .A(n107), .B(r_tui[0]), .Y(n523) );
  XNOR2XL U553 ( .A(n124), .B(r_tui[3]), .Y(n522) );
  INVX1 U554 ( .A(symb_cnt[3]), .Y(n126) );
  NOR4XL U555 ( .A(n537), .B(n126), .C(n114), .D(N160), .Y(n428) );
  INVX1 U556 ( .A(N142), .Y(n125) );
  NAND21X1 U557 ( .B(n403), .A(r_tui[0]), .Y(n402) );
  AOI21X1 U558 ( .B(n74), .C(n545), .A(n393), .Y(n403) );
  INVX1 U559 ( .A(ui_intv_cnt[6]), .Y(n120) );
  INVX1 U560 ( .A(ui_intv_cnt[7]), .Y(n121) );
  NAND2X1 U561 ( .A(symb_cnt[3]), .B(n225), .Y(n217) );
  NOR2X1 U562 ( .A(n110), .B(n12), .Y(n366) );
  NOR2X1 U563 ( .A(n90), .B(ui_intv_cnt[7]), .Y(n459) );
  NAND4X1 U564 ( .A(n459), .B(N142), .C(n107), .D(n117), .Y(n478) );
  OAI22X1 U565 ( .A(n322), .B(n323), .C(ui_intv_cnt[5]), .D(n321), .Y(n319) );
  NOR2X1 U566 ( .A(n324), .B(n318), .Y(n323) );
  AOI21X1 U567 ( .B(n324), .C(n318), .A(n125), .Y(n322) );
  AND2X1 U568 ( .A(n325), .B(n326), .Y(n324) );
  NAND2X1 U569 ( .A(r_tui[1]), .B(n74), .Y(n144) );
  AOI31X1 U570 ( .A(n56), .B(n361), .C(n362), .D(n363), .Y(n346) );
  AO21X1 U571 ( .B(n309), .C(n364), .A(n365), .Y(n362) );
  AO222X1 U572 ( .A(n352), .B(n360), .C(n354), .D(n356), .E(n96), .F(n549), 
        .Y(n361) );
  NAND3X1 U573 ( .A(N362), .B(n537), .C(n366), .Y(n364) );
  AOI32X1 U574 ( .A(n330), .B(n328), .C(ui_intv_cnt[2]), .D(n73), .E(N141), 
        .Y(n325) );
  NAND2X1 U575 ( .A(N160), .B(symb_cnt[3]), .Y(n222) );
  OAI211X1 U576 ( .C(ui_intv_cnt[0]), .D(n327), .A(n328), .B(n329), .Y(n326)
         );
  AOI22X1 U577 ( .A(n72), .B(n122), .C(n71), .D(n117), .Y(n329) );
  AOI221XL U578 ( .A(n543), .B(n126), .C(n415), .D(n416), .E(n417), .Y(n414)
         );
  AOI21X1 U579 ( .B(n418), .C(n12), .A(n348), .Y(n417) );
  ENOX1 U580 ( .A(n349), .B(n376), .C(n355), .D(n352), .Y(n416) );
  NAND2X1 U581 ( .A(n11), .B(n321), .Y(n320) );
  NOR32XL U582 ( .B(n8), .C(n366), .A(N159), .Y(n476) );
  AOI21X1 U583 ( .B(n493), .C(fcp_state[2]), .A(n245), .Y(n479) );
  XNOR2XL U584 ( .A(rx_ui_5_8[4]), .B(N142), .Y(n146) );
  XNOR2XL U585 ( .A(n144), .B(ui_intv_cnt[0]), .Y(n457) );
  NOR3XL U586 ( .A(n40), .B(n16), .C(n309), .Y(n512) );
  INVX1 U587 ( .A(test_so), .Y(n91) );
  NOR21XL U588 ( .B(n536), .A(n297), .Y(N356) );
  XNOR2XL U589 ( .A(rxtx_buf[0]), .B(n298), .Y(n297) );
  XNOR2XL U590 ( .A(n299), .B(n300), .Y(n298) );
  XNOR2XL U591 ( .A(n301), .B(n302), .Y(n300) );
  XNOR2XL U592 ( .A(ui_intv_cnt[2]), .B(rx_ui_5_8[2]), .Y(n147) );
  XNOR2XL U593 ( .A(r_dat[7]), .B(n5), .Y(n344) );
  NOR4XL U594 ( .A(n544), .B(fcp_state[0]), .C(fcp_state[1]), .D(fcp_state[3]), 
        .Y(n474) );
  NAND3X1 U595 ( .A(n494), .B(n551), .C(fcp_state[0]), .Y(n282) );
  NOR3XL U596 ( .A(n88), .B(new_rx_sync_cnt[0]), .C(n275), .Y(setsta[3]) );
  AND3X1 U597 ( .A(symb_cnt[5]), .B(n481), .C(symb_cnt[6]), .Y(n473) );
  NAND3X1 U598 ( .A(n126), .B(n116), .C(n128), .Y(n481) );
  NAND2X1 U599 ( .A(n14), .B(n505), .Y(n150) );
  INVX1 U600 ( .A(symb_cnt[6]), .Y(n118) );
  NAND4X1 U601 ( .A(n418), .B(n504), .C(n549), .D(n12), .Y(n496) );
  NAND2X1 U602 ( .A(n510), .B(n511), .Y(n498) );
  NAND4X1 U603 ( .A(n547), .B(n109), .C(n16), .D(n54), .Y(n511) );
  OAI21X1 U604 ( .B(n428), .C(n111), .A(n545), .Y(n510) );
  INVX1 U605 ( .A(rx_trans_8_chg), .Y(n84) );
  NOR3XL U606 ( .A(n273), .B(n54), .C(n539), .Y(setsta[6]) );
  NAND3X1 U607 ( .A(symb_cnt[6]), .B(n274), .C(ff_chg), .Y(n273) );
  XNOR2XL U608 ( .A(ui_intv_cnt[1]), .B(rx_ui_5_8[1]), .Y(n138) );
  XNOR2XL U609 ( .A(n143), .B(n144), .Y(n136) );
  XNOR2XL U610 ( .A(n71), .B(ui_intv_cnt[0]), .Y(n143) );
  XNOR2XL U611 ( .A(n303), .B(n304), .Y(n299) );
  XNOR2XL U612 ( .A(rxtx_buf[3]), .B(rxtx_buf[2]), .Y(n304) );
  XNOR2XL U613 ( .A(n82), .B(n54), .Y(n303) );
  INVX1 U614 ( .A(r_ctl[0]), .Y(n77) );
  OAI32X1 U615 ( .A(n292), .B(us_cnt_2_), .C(n281), .D(n286), .E(n92), .Y(N87)
         );
  INVX1 U616 ( .A(r_ctl[7]), .Y(n538) );
  INVX1 U617 ( .A(new_rx_sync_cnt[0]), .Y(n87) );
  INVX1 U618 ( .A(new_rx_sync_cnt[1]), .Y(n88) );
  XNOR2XL U620 ( .A(rxtx_buf[5]), .B(rxtx_buf[4]), .Y(n301) );
  XNOR2XL U621 ( .A(rxtx_buf[7]), .B(rxtx_buf[6]), .Y(n302) );
  OAI32X1 U622 ( .A(n275), .B(rx_trans_8_chg), .C(n150), .D(ff_chg), .E(n84), 
        .Y(n516) );
  OAI32X1 U623 ( .A(n92), .B(test_so), .C(n292), .D(n91), .E(n286), .Y(N88) );
  OR2X1 U624 ( .A(r_ctl[1]), .B(n77), .Y(n260) );
  INVX1 U625 ( .A(rxtx_buf[1]), .Y(n82) );
  NAND4X1 U626 ( .A(n151), .B(n264), .C(n531), .D(n532), .Y(N1005) );
  AOI211X1 U627 ( .C(ff_chg), .D(n285), .A(n54), .B(n551), .Y(n532) );
  AOI21X1 U628 ( .B(fcp_state[2]), .C(n533), .A(n283), .Y(n531) );
  INVX1 U629 ( .A(us_cnt_0_), .Y(n94) );
  INVX1 U630 ( .A(rxtx_buf[2]), .Y(n86) );
  INVX1 U631 ( .A(us_cnt_1_), .Y(n93) );
  NOR2X1 U632 ( .A(us_cnt_0_), .B(n546), .Y(N85) );
  INVX1 U633 ( .A(us_cnt_2_), .Y(n92) );
  INVX1 U634 ( .A(rxtx_buf[0]), .Y(n85) );
  BUFX3 U635 ( .A(tx_en), .Y(r_ctl[6]) );
  INVX1 U636 ( .A(n264), .Y(tx_en) );
endmodule


module fcpegn_a0_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module fcpegn_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(SUM[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
endmodule


module fcpegn_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9572;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9572), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9572), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9572), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9572), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9572), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9572), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9572), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9572), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9572), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9590;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9590), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9590), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9590), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9590), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9590), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9590), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9590), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9590), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9590), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9608;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9608), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9608), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9608), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9608), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9608), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9608), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9608), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9608), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9608), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_0 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_0 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[2]), .Y(n2) );
  INVX1 U4 ( .A(set2[0]), .Y(n14) );
  INVX1 U5 ( .A(set2[1]), .Y(n13) );
  INVX1 U6 ( .A(set2[4]), .Y(n15) );
  NAND3X1 U7 ( .A(n4), .B(n1), .C(n16), .Y(n21) );
  INVX1 U8 ( .A(set2[3]), .Y(n3) );
  INVX1 U9 ( .A(set2[7]), .Y(n1) );
  NOR2X1 U10 ( .A(rdat[6]), .B(n4), .Y(irq[6]) );
  NOR2X1 U11 ( .A(rdat[7]), .B(n1), .Y(irq[7]) );
  NAND4X1 U12 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U13 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U14 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U15 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U16 ( .C(n13), .D(n12), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U17 ( .A(rdat[1]), .Y(n12) );
  AOI211X1 U18 ( .C(n3), .D(n11), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U19 ( .A(rdat[3]), .Y(n11) );
  AOI211X1 U20 ( .C(n15), .D(n10), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U21 ( .A(rdat[4]), .Y(n10) );
  AOI211X1 U22 ( .C(n16), .D(n9), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U23 ( .A(rdat[5]), .Y(n9) );
  AOI211X1 U24 ( .C(n14), .D(n8), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U25 ( .A(rdat[0]), .Y(n8) );
  AOI211X1 U26 ( .C(n2), .D(n7), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U27 ( .A(rdat[2]), .Y(n7) );
  AOI211X1 U28 ( .C(n4), .D(n6), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U29 ( .A(rdat[6]), .Y(n6) );
  AOI211X1 U30 ( .C(n1), .D(n5), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U31 ( .A(rdat[7]), .Y(n5) );
  NOR2X1 U32 ( .A(rdat[0]), .B(n14), .Y(irq[0]) );
  NOR2X1 U33 ( .A(rdat[1]), .B(n13), .Y(irq[1]) );
  NOR2X1 U34 ( .A(rdat[4]), .B(n15), .Y(irq[4]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n2), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[3]), .B(n3), .Y(irq[3]) );
  INVX1 U37 ( .A(set2[6]), .Y(n4) );
  INVX1 U38 ( .A(set2[5]), .Y(n16) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9626;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9626), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9626), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9626), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9626), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9626), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9626), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9626), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9626), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9626), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000000 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9644;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9644), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9644), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9644), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9644), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9644), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9644), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9644), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9644), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9644), 
        .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dpdmacc_a0 ( dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, r_wdat, r_acc, 
        r_dpdmsta, r_dm, r_dmchg, r_int, clk, rstz, test_si, test_se );
  input [7:0] r_wdat;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, clk, rstz, test_si, test_se;
  output r_dm, r_dmchg, r_int;
  wire   dp_chg, dp_rise, dm_fall, dp_active_acc, dp_inacti_acc, dm_active_acc,
         dm_inacti_acc, upd00, n3, n4, n5, n6, n28, n29, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n30, n31,
         n32, n33, n34, n35, n36, n37, n2, n7, n8, n9, n10, n11, n38;
  wire   [7:0] wd00;

  INVX1 U4 ( .A(n6), .Y(n4) );
  INVX1 U5 ( .A(n6), .Y(n3) );
  INVX1 U6 ( .A(n6), .Y(n5) );
  INVX1 U7 ( .A(rstz), .Y(n6) );
  ff_sync_2 u0_dpsync ( .i_org(dp_comp), .o_dbc(r_dpdmsta[6]), .o_chg(dp_chg), 
        .clk(clk), .rstz(n4), .test_si(n28), .test_se(test_se) );
  ff_sync_1 u0_dmsync ( .i_org(dm_comp), .o_dbc(r_dpdmsta[7]), .o_chg(r_dmchg), 
        .clk(clk), .rstz(n4), .test_si(n29), .test_se(test_se) );
  ff_sync_0 u0_idsync ( .i_org(id_comp), .o_dbc(r_dpdmsta[5]), .o_chg(), .clk(
        clk), .rstz(n5), .test_si(r_dpdmsta[6]), .test_se(test_se) );
  filter150us_a0_1 u0_dpfltr ( .active_hit(dp_active_acc), .inacti_hit(
        dp_inacti_acc), .start_edge(dp_rise), .any_edge(dp_chg), .clk(clk), 
        .rstz(n5), .test_si(r_dpdmsta[4]), .test_so(n28), .test_se(test_se) );
  filter150us_a0_0 u0_dmfltr ( .active_hit(dm_active_acc), .inacti_hit(
        dm_inacti_acc), .start_edge(dm_fall), .any_edge(r_dmchg), .clk(clk), 
        .rstz(n5), .test_si(r_acc[7]), .test_so(n29), .test_se(test_se) );
  glreg_a0_5 u0_accmltr ( .clk(clk), .arstz(n3), .we(upd00), .wdat(wd00), 
        .rdat(r_acc), .test_si(test_si), .test_se(test_se) );
  glreg_WIDTH5_0 u0_dpdmsta ( .clk(clk), .arstz(n4), .we(r_wr_1), .wdat(
        r_wdat[4:0]), .rdat(r_dpdmsta[4:0]), .test_si(r_dpdmsta[7]), .test_se(
        test_se) );
  INVX1 U3 ( .A(r_re_0), .Y(n38) );
  NAND2X1 U8 ( .A(n32), .B(n38), .Y(upd00) );
  NOR2X1 U9 ( .A(n2), .B(n8), .Y(n32) );
  OAI22X1 U10 ( .A(n38), .B(n27), .C(r_re_0), .D(n30), .Y(wd00[0]) );
  XNOR2XL U11 ( .A(n26), .B(n11), .Y(n30) );
  OAI22X1 U12 ( .A(n18), .B(n38), .C(r_re_0), .D(n19), .Y(wd00[4]) );
  XNOR2XL U13 ( .A(n17), .B(n10), .Y(n19) );
  INVX1 U14 ( .A(n27), .Y(n8) );
  INVX1 U15 ( .A(n18), .Y(n2) );
  NOR2X1 U16 ( .A(n17), .B(n10), .Y(n15) );
  NOR2X1 U17 ( .A(n26), .B(n11), .Y(n24) );
  OAI21X1 U18 ( .B(n32), .C(n38), .A(n33), .Y(r_int) );
  AOI33X1 U19 ( .A(n8), .B(n11), .C(n34), .D(n2), .E(n10), .F(n35), .Y(n33) );
  NOR3XL U20 ( .A(r_acc[5]), .B(r_acc[7]), .C(r_acc[6]), .Y(n35) );
  AOI21BX1 U21 ( .C(r_acc[7]), .B(n12), .A(r_re_0), .Y(wd00[7]) );
  NAND21X1 U22 ( .B(n13), .A(r_acc[6]), .Y(n12) );
  AOI21BX1 U23 ( .C(r_acc[3]), .B(n21), .A(r_re_0), .Y(wd00[3]) );
  NAND21X1 U24 ( .B(n22), .A(r_acc[2]), .Y(n21) );
  NOR2X1 U25 ( .A(r_re_0), .B(n16), .Y(wd00[5]) );
  XNOR2XL U26 ( .A(r_acc[5]), .B(n15), .Y(n16) );
  NOR2X1 U27 ( .A(r_re_0), .B(n25), .Y(wd00[1]) );
  XNOR2XL U28 ( .A(r_acc[1]), .B(n24), .Y(n25) );
  NOR2X1 U29 ( .A(r_re_0), .B(n23), .Y(wd00[2]) );
  XOR2X1 U30 ( .A(n22), .B(r_acc[2]), .Y(n23) );
  NOR2X1 U31 ( .A(r_re_0), .B(n14), .Y(wd00[6]) );
  XOR2X1 U32 ( .A(n13), .B(r_acc[6]), .Y(n14) );
  OAI21X1 U33 ( .B(dm_inacti_acc), .C(n7), .A(n37), .Y(n18) );
  OAI21BX1 U34 ( .C(dm_active_acc), .B(r_dpdmsta[7]), .A(n7), .Y(n37) );
  INVX1 U35 ( .A(r_dpdmsta[1]), .Y(n7) );
  OAI21X1 U36 ( .B(dp_inacti_acc), .C(n9), .A(n36), .Y(n27) );
  OAI21BBX1 U37 ( .A(r_dpdmsta[6]), .B(dp_active_acc), .C(n9), .Y(n36) );
  INVX1 U38 ( .A(r_dpdmsta[0]), .Y(n9) );
  NOR21XL U39 ( .B(dp_chg), .A(r_dpdmsta[6]), .Y(dp_rise) );
  AND2X1 U40 ( .A(r_dmchg), .B(r_dpdmsta[7]), .Y(dm_fall) );
  NAND2X1 U41 ( .A(n2), .B(n20), .Y(n17) );
  NAND4X1 U42 ( .A(r_acc[6]), .B(r_acc[5]), .C(r_acc[4]), .D(r_acc[7]), .Y(n20) );
  NAND2X1 U43 ( .A(n15), .B(r_acc[5]), .Y(n13) );
  NOR3XL U44 ( .A(r_acc[1]), .B(r_acc[3]), .C(r_acc[2]), .Y(n34) );
  NAND2X1 U45 ( .A(n8), .B(n31), .Y(n26) );
  NAND4X1 U46 ( .A(r_acc[2]), .B(r_acc[1]), .C(r_acc[0]), .D(r_acc[3]), .Y(n31) );
  NAND2X1 U47 ( .A(n24), .B(r_acc[1]), .Y(n22) );
  INVX1 U48 ( .A(r_acc[4]), .Y(n10) );
  INVX1 U49 ( .A(r_acc[0]), .Y(n11) );
  BUFX3 U50 ( .A(r_dpdmsta[7]), .Y(r_dm) );
endmodule


module glreg_WIDTH5_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9662;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9662), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9662), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9662), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9662), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9662), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9662), 
        .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9680;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9680), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9680), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9680), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9680), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9680), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9680), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9680), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9680), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9680), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_0 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz, test_si, test_so, test_se );
  input start_edge, any_edge, clk, rstz, test_si, test_se;
  output active_hit, inacti_hit, test_so;
  wire   dbcnt_10_, dbcnt_9_, dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_,
         dbcnt_3_, dbcnt_2_, dbcnt_1_, dbcnt_0_, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, net9698, n2, n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n4, n14;

  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9698), .TE(test_se) );
  filter150us_a0_0_DW01_inc_0 add_76 ( .A({test_so, dbcnt_10_, dbcnt_9_, 
        dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_, dbcnt_3_, dbcnt_2_, 
        dbcnt_1_, dbcnt_0_}), .SUM({N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12}) );
  SDFFRQX1 dbcnt_reg_4_ ( .D(N29), .SIN(dbcnt_3_), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_4_) );
  SDFFRQX1 dbcnt_reg_3_ ( .D(N28), .SIN(dbcnt_2_), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_3_) );
  SDFFRQX1 dbcnt_reg_11_ ( .D(N36), .SIN(dbcnt_10_), .SMC(test_se), .C(net9698), .XR(n2), .Q(test_so) );
  SDFFRQX1 dbcnt_reg_2_ ( .D(N27), .SIN(dbcnt_1_), .SMC(test_se), .C(net9698), 
        .XR(rstz), .Q(dbcnt_2_) );
  SDFFRQX1 dbcnt_reg_1_ ( .D(N26), .SIN(dbcnt_0_), .SMC(test_se), .C(net9698), 
        .XR(rstz), .Q(dbcnt_1_) );
  SDFFRQX1 dbcnt_reg_0_ ( .D(N25), .SIN(test_si), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_0_) );
  SDFFRQX1 dbcnt_reg_7_ ( .D(N32), .SIN(dbcnt_6_), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_7_) );
  SDFFRQX1 dbcnt_reg_5_ ( .D(N30), .SIN(dbcnt_4_), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_5_) );
  SDFFRQX1 dbcnt_reg_6_ ( .D(N31), .SIN(dbcnt_5_), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_6_) );
  SDFFRQX1 dbcnt_reg_9_ ( .D(N34), .SIN(dbcnt_8_), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_9_) );
  SDFFRQX1 dbcnt_reg_8_ ( .D(N33), .SIN(dbcnt_7_), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_8_) );
  SDFFRQX1 dbcnt_reg_10_ ( .D(N35), .SIN(dbcnt_9_), .SMC(test_se), .C(net9698), 
        .XR(n2), .Q(dbcnt_10_) );
  BUFX3 U3 ( .A(n9), .Y(n1) );
  INVX1 U6 ( .A(any_edge), .Y(n4) );
  AND2X1 U7 ( .A(N22), .B(n9), .Y(N35) );
  AND2X1 U8 ( .A(N20), .B(n9), .Y(N33) );
  AND2X1 U9 ( .A(N21), .B(n9), .Y(N34) );
  NOR3XL U10 ( .A(n11), .B(any_edge), .C(n14), .Y(n9) );
  AND2X1 U11 ( .A(N16), .B(n9), .Y(N29) );
  AND2X1 U12 ( .A(N15), .B(n9), .Y(N28) );
  AND2X1 U13 ( .A(N19), .B(n9), .Y(N32) );
  AND2X1 U14 ( .A(N17), .B(n9), .Y(N30) );
  AND2X1 U15 ( .A(N18), .B(n9), .Y(N31) );
  AND2X1 U16 ( .A(N14), .B(n1), .Y(N27) );
  AND2X1 U17 ( .A(N13), .B(n1), .Y(N26) );
  INVX1 U18 ( .A(n5), .Y(n14) );
  OR2X1 U19 ( .A(n1), .B(any_edge), .Y(N24) );
  AOI211X1 U20 ( .C(n5), .D(n6), .A(n4), .B(start_edge), .Y(inacti_hit) );
  AOI21X1 U21 ( .B(n7), .C(n8), .A(test_so), .Y(n5) );
  NAND32X1 U22 ( .B(dbcnt_4_), .C(dbcnt_3_), .A(n13), .Y(n7) );
  NOR3XL U23 ( .A(dbcnt_5_), .B(dbcnt_7_), .C(dbcnt_6_), .Y(n13) );
  AND3X1 U24 ( .A(dbcnt_8_), .B(dbcnt_10_), .C(dbcnt_9_), .Y(n8) );
  NOR3XL U25 ( .A(n6), .B(test_so), .C(n7), .Y(active_hit) );
  NAND4X1 U26 ( .A(dbcnt_2_), .B(dbcnt_1_), .C(dbcnt_0_), .D(n8), .Y(n6) );
  AND2X1 U27 ( .A(N23), .B(n1), .Y(N36) );
  NOR4XL U28 ( .A(dbcnt_0_), .B(dbcnt_10_), .C(n7), .D(n12), .Y(n11) );
  OR4X1 U29 ( .A(dbcnt_9_), .B(dbcnt_8_), .C(dbcnt_2_), .D(dbcnt_1_), .Y(n12)
         );
  OAI21BBX1 U30 ( .A(N12), .B(n9), .C(n10), .Y(N25) );
  OAI21X1 U31 ( .B(n11), .C(n14), .A(any_edge), .Y(n10) );
endmodule


module filter150us_a0_0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_1 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz, test_si, test_so, test_se );
  input start_edge, any_edge, clk, rstz, test_si, test_se;
  output active_hit, inacti_hit, test_so;
  wire   dbcnt_10_, dbcnt_9_, dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_,
         dbcnt_3_, dbcnt_2_, dbcnt_1_, dbcnt_0_, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, net9716, n2, n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n4, n14;

  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9716), .TE(test_se) );
  filter150us_a0_1_DW01_inc_0 add_76 ( .A({test_so, dbcnt_10_, dbcnt_9_, 
        dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_, dbcnt_3_, dbcnt_2_, 
        dbcnt_1_, dbcnt_0_}), .SUM({N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12}) );
  SDFFRQX1 dbcnt_reg_4_ ( .D(N29), .SIN(dbcnt_3_), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_4_) );
  SDFFRQX1 dbcnt_reg_3_ ( .D(N28), .SIN(dbcnt_2_), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_3_) );
  SDFFRQX1 dbcnt_reg_11_ ( .D(N36), .SIN(dbcnt_10_), .SMC(test_se), .C(net9716), .XR(n2), .Q(test_so) );
  SDFFRQX1 dbcnt_reg_2_ ( .D(N27), .SIN(dbcnt_1_), .SMC(test_se), .C(net9716), 
        .XR(rstz), .Q(dbcnt_2_) );
  SDFFRQX1 dbcnt_reg_1_ ( .D(N26), .SIN(dbcnt_0_), .SMC(test_se), .C(net9716), 
        .XR(rstz), .Q(dbcnt_1_) );
  SDFFRQX1 dbcnt_reg_0_ ( .D(N25), .SIN(test_si), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_0_) );
  SDFFRQX1 dbcnt_reg_7_ ( .D(N32), .SIN(dbcnt_6_), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_7_) );
  SDFFRQX1 dbcnt_reg_5_ ( .D(N30), .SIN(dbcnt_4_), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_5_) );
  SDFFRQX1 dbcnt_reg_6_ ( .D(N31), .SIN(dbcnt_5_), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_6_) );
  SDFFRQX1 dbcnt_reg_9_ ( .D(N34), .SIN(dbcnt_8_), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_9_) );
  SDFFRQX1 dbcnt_reg_8_ ( .D(N33), .SIN(dbcnt_7_), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_8_) );
  SDFFRQX1 dbcnt_reg_10_ ( .D(N35), .SIN(dbcnt_9_), .SMC(test_se), .C(net9716), 
        .XR(n2), .Q(dbcnt_10_) );
  BUFX3 U3 ( .A(n9), .Y(n1) );
  INVX1 U6 ( .A(any_edge), .Y(n14) );
  AND2X1 U7 ( .A(N22), .B(n9), .Y(N35) );
  AND2X1 U8 ( .A(N20), .B(n9), .Y(N33) );
  AND2X1 U9 ( .A(N21), .B(n9), .Y(N34) );
  NOR3XL U10 ( .A(n11), .B(any_edge), .C(n4), .Y(n9) );
  AND2X1 U11 ( .A(N15), .B(n9), .Y(N28) );
  AND2X1 U12 ( .A(N19), .B(n9), .Y(N32) );
  AND2X1 U13 ( .A(N17), .B(n9), .Y(N30) );
  AND2X1 U14 ( .A(N18), .B(n9), .Y(N31) );
  AND2X1 U15 ( .A(N14), .B(n9), .Y(N27) );
  AND2X1 U16 ( .A(N13), .B(n1), .Y(N26) );
  AND2X1 U17 ( .A(N16), .B(n1), .Y(N29) );
  INVX1 U18 ( .A(n5), .Y(n4) );
  OR2X1 U19 ( .A(n1), .B(any_edge), .Y(N24) );
  AOI211X1 U20 ( .C(n5), .D(n6), .A(n14), .B(start_edge), .Y(inacti_hit) );
  AOI21X1 U21 ( .B(n7), .C(n8), .A(test_so), .Y(n5) );
  NAND32X1 U22 ( .B(dbcnt_4_), .C(dbcnt_3_), .A(n13), .Y(n7) );
  NOR3XL U23 ( .A(dbcnt_5_), .B(dbcnt_7_), .C(dbcnt_6_), .Y(n13) );
  AND3X1 U24 ( .A(dbcnt_8_), .B(dbcnt_10_), .C(dbcnt_9_), .Y(n8) );
  NOR3XL U25 ( .A(n6), .B(test_so), .C(n7), .Y(active_hit) );
  NAND4X1 U26 ( .A(dbcnt_2_), .B(dbcnt_1_), .C(dbcnt_0_), .D(n8), .Y(n6) );
  AND2X1 U27 ( .A(N23), .B(n1), .Y(N36) );
  NOR4XL U28 ( .A(dbcnt_0_), .B(dbcnt_10_), .C(n7), .D(n12), .Y(n11) );
  OR4X1 U29 ( .A(dbcnt_9_), .B(dbcnt_8_), .C(dbcnt_2_), .D(dbcnt_1_), .Y(n12)
         );
  OAI21BBX1 U30 ( .A(N12), .B(n9), .C(n10), .Y(N25) );
  OAI21X1 U31 ( .B(n11), .C(n4), .A(any_edge), .Y(n10) );
endmodule


module filter150us_a0_1_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ff_sync_0 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg;
  wire   d_org_0_;

  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_1 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg;
  wire   d_org_0_;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_2 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg;
  wire   d_org_0_;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module dacmux_a0 ( clk, srstz, i_comp, r_comp_opt, r_wdat, r_adofs, r_isofs, 
        r_wr, dacv_wr, o_dacv, o_shrst, o_hold, o_dac1, o_daci_sel, o_dat, 
        r_dac_en, r_sar_en, o_dactl, o_cmpsta, x_daclsb, o_intr, o_smpl, 
        test_si2, test_si1, test_so1, test_se );
  input [2:0] r_comp_opt;
  input [7:0] r_wdat;
  output [7:0] r_adofs;
  output [7:0] r_isofs;
  input [10:0] r_wr;
  input [17:0] dacv_wr;
  output [143:0] o_dacv;
  output [9:0] o_dac1;
  output [17:0] o_daci_sel;
  output [17:0] o_dat;
  output [17:0] r_dac_en;
  output [17:0] r_sar_en;
  output [7:0] o_dactl;
  output [7:0] o_cmpsta;
  output [5:0] x_daclsb;
  output [4:0] o_smpl;
  input clk, srstz, i_comp, test_si2, test_si1, test_se;
  output o_shrst, o_hold, o_intr, test_so1;
  wire   dacyc_done, updcmp, semi_start, sacyc_done, sar_ini, sar_nxt,
         sampl_begn, sampl_done, ps_md4ch, updlsb, wda_6_, N1239, N1240, N1241,
         N1242, N1243, N1244, N1245, N1246, N1247, N1250, N1251, N1252, N1253,
         N1254, N1255, N1256, N1257, N1258, N1261, N1262, N1263, N1264, N1265,
         N1266, N1267, N1268, N1269, N1272, N1273, N1274, N1275, N1276, N1277,
         N1278, N1279, N1280, N1283, N1284, N1285, N1286, N1287, N1288, N1289,
         N1290, N1291, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301,
         N1302, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313,
         N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1327,
         N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1338, N1339,
         N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1349, N1350, N1351,
         N1352, N1353, N1354, N1355, N1356, N1357, N1360, N1361, N1362, N1363,
         N1364, N1365, N1366, N1367, N1368, N1371, N1372, N1373, N1374, N1375,
         N1376, N1377, N1378, N1379, N1382, N1383, N1384, N1385, N1386, N1387,
         N1388, N1389, N1390, N1393, N1394, N1395, N1396, N1397, N1398, N1399,
         N1400, N1401, N1404, N1405, N1406, N1407, N1408, N1409, N1410, N1411,
         N1412, N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423,
         N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434, n571,
         n563, n568, n569, n564, n567, n570, n100, n562, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n565, n566, n64, n94, n95, n96, n137,
         n138, n139, n140, n141, n143, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n207, n208, n209, n210, n211, n212, n213, n214, n215, n217,
         n218, n219, n220, n221, n301, n302, n304, n305, n306, n308, n309,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n330, n333, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n414, n415, n416, n417, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n456, n457, n458, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n84, n86, n88, n90, n92, n97, n98, n99, n101,
         n102, n103, n104, n105, n106, n107, n109, n110, n111, n112, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n142, n144, n145, n205, n206, n216, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n303, n307, n310,
         n311, n312, n313, n314, n315, n329, n331, n332, n334, n413, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n455, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561;
  wire   [1:0] syn_comp;
  wire   [4:0] cs_ptr;
  wire   [17:0] datcmp;
  wire   [4:0] ps_ptr;
  wire   [9:0] r_dac1v;
  wire   [9:0] r_rpt_v;
  wire   [17:0] app_dacis;
  wire   [17:0] pos_dacis;
  wire   [5:0] wdlsb;
  wire   [17:0] upd;
  wire   [143:0] r_dacvs;
  wire   [7:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;

  INVX1 U172 ( .A(n190), .Y(n189) );
  INVX1 U175 ( .A(n190), .Y(n183) );
  INVX1 U176 ( .A(n190), .Y(n182) );
  INVX1 U177 ( .A(n191), .Y(n181) );
  INVX1 U178 ( .A(n192), .Y(n180) );
  INVX1 U179 ( .A(n192), .Y(n179) );
  INVX1 U180 ( .A(n191), .Y(n178) );
  INVX1 U181 ( .A(n190), .Y(n177) );
  INVX1 U182 ( .A(n191), .Y(n175) );
  INVX1 U183 ( .A(n191), .Y(n174) );
  INVX1 U184 ( .A(n192), .Y(n173) );
  INVX1 U185 ( .A(n190), .Y(n172) );
  INVX1 U186 ( .A(n191), .Y(n171) );
  INVX1 U187 ( .A(n192), .Y(n170) );
  INVX1 U188 ( .A(n191), .Y(n169) );
  INVX1 U189 ( .A(n191), .Y(n168) );
  INVX1 U190 ( .A(n192), .Y(n167) );
  INVX1 U191 ( .A(n192), .Y(n166) );
  INVX1 U192 ( .A(n192), .Y(n176) );
  INVX1 U193 ( .A(n192), .Y(n165) );
  INVX1 U194 ( .A(n191), .Y(n187) );
  INVX1 U195 ( .A(n191), .Y(n186) );
  INVX1 U196 ( .A(n191), .Y(n185) );
  INVX1 U197 ( .A(n190), .Y(n184) );
  INVX1 U198 ( .A(n192), .Y(n164) );
  INVX1 U199 ( .A(n190), .Y(n188) );
  INVX1 U201 ( .A(srstz), .Y(n190) );
  INVX1 U224 ( .A(n192), .Y(n163) );
  INVX1 U225 ( .A(srstz), .Y(n192) );
  INVX1 U226 ( .A(srstz), .Y(n191) );
  glreg_00000012 u0_compi ( .clk(clk), .arstz(n189), .we(updcmp), .wdat(datcmp), .rdat(o_dat), .test_si(o_cmpsta[7]), .test_se(test_se) );
  dac2sar_a0 u0_dac2sar ( .r_dac_t(o_dactl[3:2]), .r_dacyc(o_dactl[7]), 
        .r_sar10(n64), .sar_ini(sar_ini), .sar_nxt(sar_nxt), .semi_nxt(n94), 
        .auto_sar(n456), .busy(o_dactl[0]), .stop(n458), .sync_i(syn_comp[1]), 
        .sampl_begn(sampl_begn), .sampl_done(sampl_done), .sh_rst(o_shrst), 
        .dacyc_done(dacyc_done), .sacyc_done(sacyc_done), .ps_sample(), 
        .dac_v(r_dac1v), .rpt_v(r_rpt_v), .clk(clk), .srstz(n189), .test_si2(
        o_dat[17]), .test_si1(test_si1), .test_so1(n566), .test_se(test_se) );
  shmux_00000005_00000012_00000012 u0_shmux ( .ps_md4ch(ps_md4ch), 
        .r_comp_swtch(r_comp_opt[2]), .r_semi(n96), .r_loop(o_dactl[1]), 
        .r_dac_en(r_dac_en), .wr_dacv(dacv_wr), .busy(o_dactl[0]), .sh_hold(
        o_hold), .stop(n458), .semi_start(semi_start), .auto_start(n457), 
        .mxcyc_done(n100), .sampl_begn(sampl_begn), .sampl_done(sampl_done), 
        .app_dacis(app_dacis), .pos_dacis(pos_dacis), .cs_ptr(cs_ptr), 
        .ps_ptr(ps_ptr), .clk(clk), .srstz(n189), .test_si2(r_sar_en[7]), 
        .test_si1(o_shrst), .test_so1(test_so1), .test_se(test_se) );
  glreg_WIDTH7_1 u0_dactl ( .clk(clk), .arstz(n188), .we(n95), .wdat({
        r_wdat[7], n6, n9, r_wdat[4:3], n4, r_wdat[1]}), .rdat(o_dactl[7:1]), 
        .test_si(x_daclsb[5]), .test_se(test_se) );
  glreg_a0_49 u0_dacen ( .clk(clk), .arstz(n163), .we(r_wr[1]), .wdat({
        r_wdat[7], n6, n9, r_wdat[4:3], n4, n60, n50}), .rdat(r_dac_en[7:0]), 
        .test_si(n566), .test_se(test_se) );
  glreg_a0_48 u0_saren ( .clk(clk), .arstz(n164), .we(r_wr[2]), .wdat({
        r_wdat[7], n6, n9, r_wdat[4:3], n4, n60, n51}), .rdat(r_sar_en[7:0]), 
        .test_si(r_isofs[7]), .test_se(test_se) );
  glreg_WIDTH6_2 u0_daclsb ( .clk(clk), .arstz(srstz), .we(updlsb), .wdat(
        wdlsb), .rdat(x_daclsb), .test_si(r_dac_en[7]), .test_se(test_se) );
  glreg_a0_47 dacvs_0__u0 ( .clk(clk), .arstz(n165), .we(upd[0]), .wdat({n58, 
        n12, n17, n38, n41, n45, n49, n14}), .rdat(r_dacvs[7:0]), .test_si(
        test_si2), .test_se(test_se) );
  glreg_a0_46 dacvs_1__u0 ( .clk(clk), .arstz(n176), .we(upd[1]), .wdat({n57, 
        n13, n17, n38, n41, n45, n49, n15}), .rdat(r_dacvs[15:8]), .test_si(
        r_dacvs[7]), .test_se(test_se) );
  glreg_a0_45 dacvs_2__u0 ( .clk(clk), .arstz(n166), .we(upd[2]), .wdat({n58, 
        n13, n17, n38, n41, n45, n49, n15}), .rdat(r_dacvs[23:16]), .test_si(
        r_dacvs[15]), .test_se(test_se) );
  glreg_a0_44 dacvs_3__u0 ( .clk(clk), .arstz(n167), .we(upd[3]), .wdat({n58, 
        n12, n69, n68, n67, n66, n65, n14}), .rdat(r_dacvs[31:24]), .test_si(
        r_dacvs[23]), .test_se(test_se) );
  glreg_a0_43 dacvs_4__u0 ( .clk(clk), .arstz(n168), .we(upd[4]), .wdat({n57, 
        n13, n69, n68, n67, n66, n65, n15}), .rdat(r_dacvs[39:32]), .test_si(
        r_dacvs[31]), .test_se(test_se) );
  glreg_a0_42 dacvs_5__u0 ( .clk(clk), .arstz(n169), .we(upd[5]), .wdat({n57, 
        n12, n17, n38, n41, n45, n49, n14}), .rdat(r_dacvs[47:40]), .test_si(
        r_dacvs[39]), .test_se(test_se) );
  glreg_a0_41 dacvs_6__u0 ( .clk(clk), .arstz(n170), .we(upd[6]), .wdat({n58, 
        n13, n17, n38, n41, n45, n49, n15}), .rdat(r_dacvs[55:48]), .test_si(
        r_dacvs[47]), .test_se(test_se) );
  glreg_a0_40 dacvs_7__u0 ( .clk(clk), .arstz(n171), .we(upd[7]), .wdat({n57, 
        n13, n17, n38, n41, n45, n49, n15}), .rdat(r_dacvs[63:56]), .test_si(
        r_dacvs[55]), .test_se(test_se) );
  glreg_a0_39 dacvs_8__u0 ( .clk(clk), .arstz(n172), .we(upd[8]), .wdat({n57, 
        n13, n69, n68, n67, n66, n65, n15}), .rdat(r_dacvs[71:64]), .test_si(
        r_dacvs[63]), .test_se(test_se) );
  glreg_a0_38 dacvs_9__u0 ( .clk(clk), .arstz(n173), .we(upd[9]), .wdat({n58, 
        n13, n17, n38, n41, n45, n49, n15}), .rdat(r_dacvs[79:72]), .test_si(
        r_dacvs[71]), .test_se(test_se) );
  glreg_a0_37 dacvs_10__u0 ( .clk(clk), .arstz(n174), .we(upd[10]), .wdat({n58, 
        n13, n69, n68, n67, n66, n65, n15}), .rdat(r_dacvs[87:80]), .test_si(
        r_dacvs[79]), .test_se(test_se) );
  glreg_a0_36 dacvs_11__u0 ( .clk(clk), .arstz(n175), .we(upd[11]), .wdat({n57, 
        n12, n69, n68, n67, n66, n65, n14}), .rdat(r_dacvs[95:88]), .test_si(
        r_dacvs[87]), .test_se(test_se) );
  glreg_a0_35 dacvs_12__u0 ( .clk(clk), .arstz(n177), .we(upd[12]), .wdat({n58, 
        n12, n17, n38, n41, n45, n49, n14}), .rdat(r_dacvs[103:96]), .test_si(
        r_dacvs[95]), .test_se(test_se) );
  glreg_a0_34 dacvs_13__u0 ( .clk(clk), .arstz(n178), .we(upd[13]), .wdat({n58, 
        n13, n69, n68, n67, n66, n65, n15}), .rdat(r_dacvs[111:104]), 
        .test_si(r_dacvs[103]), .test_se(test_se) );
  glreg_a0_33 dacvs_14__u0 ( .clk(clk), .arstz(n179), .we(upd[14]), .wdat({n57, 
        n12, n69, n68, n67, n66, n65, n14}), .rdat(r_dacvs[119:112]), 
        .test_si(r_dacvs[111]), .test_se(test_se) );
  glreg_a0_32 dacvs_15__u0 ( .clk(clk), .arstz(n180), .we(upd[15]), .wdat({n58, 
        n12, n17, n38, n41, n45, n49, n14}), .rdat(r_dacvs[127:120]), 
        .test_si(r_dacvs[119]), .test_se(test_se) );
  glreg_a0_31 dacvs_16__u0 ( .clk(clk), .arstz(n181), .we(upd[16]), .wdat({n57, 
        n12, n69, n68, n67, n66, n65, n14}), .rdat(r_dacvs[135:128]), 
        .test_si(r_dacvs[127]), .test_se(test_se) );
  glreg_a0_30 dacvs_17__u0 ( .clk(clk), .arstz(n182), .we(upd[17]), .wdat({n57, 
        n12, n69, n68, n67, n66, n65, n14}), .rdat(r_dacvs[143:136]), 
        .test_si(r_dacvs[135]), .test_se(test_se) );
  glsta_a0_1 u0_cmpsta ( .clk(clk), .arstz(n183), .rst0(1'b0), .set2(setsta), 
        .clr1(clrsta), .rdat(o_cmpsta), .irq(r_irq), .test_si(r_adofs[7]), 
        .test_se(test_se) );
  glreg_a0_29 u0_adofs ( .clk(clk), .arstz(n184), .we(r_wr[5]), .wdat({
        r_wdat[7], n6, n8, r_wdat[4:3], n4, n60, n51}), .rdat({n562, n563, 
        n564, n567, n568, n569, n570, n571}), .test_si(syn_comp[1]), .test_se(
        test_se) );
  glreg_a0_28 u0_isofs ( .clk(clk), .arstz(n185), .we(r_wr[6]), .wdat({
        r_wdat[7], n6, n9, r_wdat[4:3], n4, r_wdat[1], n51}), .rdat(r_isofs), 
        .test_si(o_dactl[7]), .test_se(test_se) );
  glreg_a0_27 u1_dacen ( .clk(clk), .arstz(n186), .we(r_wr[7]), .wdat({
        r_wdat[7], n6, n9, r_wdat[4:3], n4, n60, n50}), .rdat(r_dac_en[15:8]), 
        .test_si(pos_dacis[17]), .test_se(test_se) );
  glreg_a0_26 u1_saren ( .clk(clk), .arstz(n187), .we(r_wr[8]), .wdat({
        r_wdat[7], n6, n9, r_wdat[4:3], n4, n60, n51}), .rdat(r_sar_en[15:8]), 
        .test_si(r_dac_en[15]), .test_se(test_se) );
  glreg_WIDTH2_1 u2_dacen ( .clk(clk), .arstz(n172), .we(r_wr[9]), .wdat({n60, 
        n51}), .rdat(r_dac_en[17:16]), .test_si(r_sar_en[15]), .test_so(n565), 
        .test_se(test_se) );
  glreg_WIDTH2_0 u2_saren ( .clk(clk), .arstz(n188), .we(r_wr[10]), .wdat({n60, 
        n51}), .rdat(r_sar_en[17:16]), .test_si(n565), .test_se(test_se) );
  dacmux_a0_DW01_add_0 add_235_I18 ( .A({1'b0, r_dacvs[143:136]}), .B({
        r_adofs[7], n110, n92, n90, n88, n86, n84, n82, r_adofs[0]}), .CI(1'b0), .SUM({N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426}), .CO()
         );
  dacmux_a0_DW01_add_1 add_235_I17 ( .A({1'b0, r_dacvs[135:128]}), .B({
        r_adofs[7], n110, r_adofs[6:0]}), .CI(1'b0), .SUM({N1423, N1422, N1421, 
        N1420, N1419, N1418, N1417, N1416, N1415}), .CO() );
  dacmux_a0_DW01_add_2 add_235_I16 ( .A({1'b0, r_dacvs[127:120]}), .B({n112, 
        n110, n92, n90, n88, n86, n84, n82, n107}), .CI(1'b0), .SUM({N1412, 
        N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404}), .CO() );
  dacmux_a0_DW01_add_3 add_235_I15 ( .A({1'b0, r_dacvs[119:112]}), .B({n112, 
        n110, r_adofs[6:1], n107}), .CI(1'b0), .SUM({N1401, N1400, N1399, 
        N1398, N1397, N1396, N1395, N1394, N1393}), .CO() );
  dacmux_a0_DW01_add_4 add_235_I14 ( .A({1'b0, r_dacvs[111:104]}), .B({n112, 
        n110, n92, n90, n88, n86, n84, n82, n107}), .CI(1'b0), .SUM({N1390, 
        N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382}), .CO() );
  dacmux_a0_DW01_add_5 add_235_I13 ( .A({1'b0, r_dacvs[103:96]}), .B({n112, 
        n110, r_adofs[6:1], n107}), .CI(1'b0), .SUM({N1379, N1378, N1377, 
        N1376, N1375, N1374, N1373, N1372, N1371}), .CO() );
  dacmux_a0_DW01_add_6 add_235_I12 ( .A({1'b0, r_dacvs[95:88]}), .B({n112, 
        n110, n92, n90, n88, n86, n84, n82, n107}), .CI(1'b0), .SUM({N1368, 
        N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360}), .CO() );
  dacmux_a0_DW01_add_7 add_235_I11 ( .A({1'b0, r_dacvs[87:80]}), .B({n112, 
        n110, r_adofs[6:1], n106}), .CI(1'b0), .SUM({N1357, N1356, N1355, 
        N1354, N1353, N1352, N1351, N1350, N1349}), .CO() );
  dacmux_a0_DW01_add_8 add_235_I10 ( .A({1'b0, r_dacvs[79:72]}), .B({n111, 
        n110, n92, n90, n88, n86, n84, n82, n106}), .CI(1'b0), .SUM({N1346, 
        N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338}), .CO() );
  dacmux_a0_DW01_add_9 add_235_I9 ( .A({1'b0, r_dacvs[71:64]}), .B({n111, n110, 
        r_adofs[6:1], n106}), .CI(1'b0), .SUM({N1335, N1334, N1333, N1332, 
        N1331, N1330, N1329, N1328, N1327}), .CO() );
  dacmux_a0_DW01_add_10 add_235_I8 ( .A({1'b0, r_dacvs[63:56]}), .B({n111, 
        n111, n92, n90, n88, n86, n84, n82, n106}), .CI(1'b0), .SUM({N1324, 
        N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316}), .CO() );
  dacmux_a0_DW01_add_11 add_235_I7 ( .A({1'b0, r_dacvs[55:48]}), .B({n112, 
        n111, r_adofs[6:1], n106}), .CI(1'b0), .SUM({N1313, N1312, N1311, 
        N1310, N1309, N1308, N1307, N1306, N1305}), .CO() );
  dacmux_a0_DW01_add_12 add_235_I6 ( .A({1'b0, r_dacvs[47:40]}), .B({n112, 
        n111, n92, n90, n88, n86, n84, n82, r_adofs[0]}), .CI(1'b0), .SUM({
        N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294}), .CO()
         );
  dacmux_a0_DW01_add_13 add_235_I5 ( .A({1'b0, r_dacvs[39:32]}), .B({n112, 
        n111, r_adofs[6:1], n571}), .CI(1'b0), .SUM({N1291, N1290, N1289, 
        N1288, N1287, N1286, N1285, N1284, N1283}), .CO() );
  dacmux_a0_DW01_add_14 add_235_I4 ( .A({1'b0, r_dacvs[31:24]}), .B({
        r_adofs[7], n111, n92, n90, n88, n86, n84, n82, r_adofs[0]}), .CI(1'b0), .SUM({N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272}), .CO()
         );
  dacmux_a0_DW01_add_15 add_235_I3 ( .A({1'b0, r_dacvs[23:16]}), .B({
        r_isofs[7], r_isofs}), .CI(1'b0), .SUM({N1269, N1268, N1267, N1266, 
        N1265, N1264, N1263, N1262, N1261}), .CO() );
  dacmux_a0_DW01_add_16 add_235_I2 ( .A({1'b0, r_dacvs[15:8]}), .B({n112, n111, 
        r_adofs[6:1], n571}), .CI(1'b0), .SUM({N1258, N1257, N1256, N1255, 
        N1254, N1253, N1252, N1251, N1250}), .CO() );
  dacmux_a0_DW01_add_17 add_235 ( .A({1'b0, r_dacvs[7:0]}), .B({r_adofs[7], 
        n111, n92, n90, n88, n86, n84, n82, n571}), .CI(1'b0), .SUM({N1247, 
        N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239}), .CO() );
  SDFFQX1 syn_comp_reg_1_ ( .D(syn_comp[0]), .SIN(syn_comp[0]), .SMC(test_se), 
        .C(clk), .Q(syn_comp[1]) );
  SDFFQX1 syn_comp_reg_0_ ( .D(i_comp), .SIN(r_dacvs[143]), .SMC(test_se), .C(
        clk), .Q(syn_comp[0]) );
  BUFX3 U21 ( .A(n431), .Y(n1) );
  INVX3 U22 ( .A(n234), .Y(n458) );
  NAND21XL U23 ( .B(ps_ptr[2]), .A(ps_ptr[1]), .Y(n244) );
  NAND21XL U24 ( .B(n241), .A(ps_ptr[2]), .Y(n240) );
  NAND21XL U25 ( .B(ps_ptr[1]), .A(ps_ptr[2]), .Y(n245) );
  NAND21X1 U26 ( .B(n253), .A(n252), .Y(n254) );
  INVX2 U27 ( .A(n242), .Y(n262) );
  NAND21X1 U28 ( .B(ps_ptr[2]), .A(n241), .Y(n242) );
  MUX2IX1 U29 ( .D0(n251), .D1(n250), .S(ps_ptr[3]), .Y(n252) );
  MUX2IX1 U30 ( .D0(n247), .D1(n246), .S(ps_ptr[3]), .Y(n248) );
  MUX2IX1 U31 ( .D0(n257), .D1(n256), .S(ps_ptr[3]), .Y(n258) );
  MUX2IX1 U32 ( .D0(n266), .D1(n265), .S(ps_ptr[3]), .Y(n267) );
  AO21X1 U33 ( .B(N1321), .C(n525), .A(n524), .Y(o_dacv[61]) );
  GEN2XL U34 ( .D(n470), .E(n469), .C(n468), .B(n478), .A(n467), .Y(n489) );
  AO21X1 U35 ( .B(N1306), .C(n522), .A(n521), .Y(o_dacv[49]) );
  AO21X1 U36 ( .B(N1289), .C(n516), .A(n515), .Y(o_dacv[38]) );
  AO21X1 U37 ( .B(N1274), .C(n513), .A(n512), .Y(o_dacv[26]) );
  INVX1 U38 ( .A(ps_ptr[1]), .Y(n241) );
  AO21X1 U39 ( .B(N1305), .C(n522), .A(n521), .Y(o_dacv[48]) );
  NAND21X1 U40 ( .B(n249), .A(n248), .Y(n255) );
  NAND21X1 U41 ( .B(n268), .A(n267), .Y(n269) );
  NAND21X1 U42 ( .B(n259), .A(n258), .Y(n270) );
  INVX2 U43 ( .A(n239), .Y(n457) );
  MUX2X1 U44 ( .D0(n481), .D1(n482), .S(pos_dacis[16]), .Y(n494) );
  MUX2BXL U45 ( .D0(n473), .D1(n472), .S(pos_dacis[14]), .Y(n480) );
  BUFX3 U46 ( .A(r_wdat[0]), .Y(n50) );
  BUFX3 U47 ( .A(r_wdat[1]), .Y(n60) );
  BUFXL U48 ( .A(r_wdat[0]), .Y(n51) );
  AND3X1 U49 ( .A(n537), .B(n538), .C(n543), .Y(n2) );
  INVXL U50 ( .A(r_wdat[2]), .Y(n3) );
  INVXL U51 ( .A(n3), .Y(n4) );
  INVXL U52 ( .A(r_wdat[6]), .Y(n5) );
  INVXL U53 ( .A(n5), .Y(n6) );
  INVXL U54 ( .A(r_wdat[5]), .Y(n7) );
  INVXL U55 ( .A(n7), .Y(n8) );
  INVXL U56 ( .A(n7), .Y(n9) );
  INVXL U57 ( .A(n412), .Y(n10) );
  INVXL U58 ( .A(n412), .Y(n11) );
  BUFX3 U59 ( .A(n126), .Y(wda_6_) );
  INVX1 U60 ( .A(wda_6_), .Y(n12) );
  INVX1 U61 ( .A(wda_6_), .Y(n13) );
  BUFX3 U62 ( .A(n125), .Y(n454) );
  INVX1 U63 ( .A(n454), .Y(n14) );
  INVX1 U64 ( .A(n454), .Y(n15) );
  INVX1 U65 ( .A(n69), .Y(n16) );
  INVX1 U66 ( .A(n16), .Y(n17) );
  INVX1 U67 ( .A(n530), .Y(n18) );
  INVX1 U68 ( .A(n68), .Y(n37) );
  INVX1 U69 ( .A(n37), .Y(n38) );
  NOR2X1 U70 ( .A(n156), .B(n102), .Y(n39) );
  INVX1 U71 ( .A(n67), .Y(n40) );
  INVX1 U72 ( .A(n40), .Y(n41) );
  INVX1 U73 ( .A(n203), .Y(n42) );
  NOR2X1 U74 ( .A(n104), .B(n143), .Y(n43) );
  INVX1 U75 ( .A(n66), .Y(n44) );
  INVX1 U76 ( .A(n44), .Y(n45) );
  BUFX3 U77 ( .A(n337), .Y(n46) );
  NOR2X1 U78 ( .A(n104), .B(n156), .Y(n47) );
  INVX1 U79 ( .A(n65), .Y(n48) );
  INVX1 U80 ( .A(n48), .Y(n49) );
  BUFX3 U81 ( .A(n335), .Y(n52) );
  BUFX3 U82 ( .A(n336), .Y(n53) );
  NOR2X1 U83 ( .A(o_dactl[0]), .B(semi_start), .Y(n290) );
  INVX1 U84 ( .A(n290), .Y(n54) );
  INVX1 U85 ( .A(n290), .Y(n55) );
  NOR2X1 U86 ( .A(n104), .B(n151), .Y(n56) );
  MUX2IX1 U87 ( .D0(r_rpt_v[9]), .D1(r_wdat[7]), .S(n137), .Y(n70) );
  INVX1 U88 ( .A(n70), .Y(n57) );
  INVX1 U89 ( .A(n70), .Y(n58) );
  INVX1 U90 ( .A(n529), .Y(n59) );
  NAND21X2 U91 ( .B(n276), .A(n275), .Y(sar_ini) );
  NOR2X1 U92 ( .A(n143), .B(n102), .Y(n61) );
  NOR2X1 U93 ( .A(n104), .B(n148), .Y(n62) );
  INVX1 U94 ( .A(n231), .Y(n63) );
  INVXL U95 ( .A(dacv_wr[13]), .Y(n284) );
  NAND21XL U96 ( .B(n276), .A(n237), .Y(semi_start) );
  AND2XL U97 ( .A(r_wr[4]), .B(n6), .Y(clrsta[6]) );
  AND2XL U98 ( .A(r_wdat[4]), .B(r_wr[4]), .Y(clrsta[4]) );
  MUX2XL U99 ( .D0(n9), .D1(o_dactl[5]), .S(n236), .Y(ps_md4ch) );
  MUX2IX1 U100 ( .D0(n480), .D1(n81), .S(pos_dacis[15]), .Y(n500) );
  OAI31XL U101 ( .A(n303), .B(pos_dacis[0]), .C(n300), .D(n464), .Y(n431) );
  MUX2X1 U102 ( .D0(n332), .D1(n80), .S(pos_dacis[7]), .Y(n462) );
  INVX1 U103 ( .A(pos_dacis[3]), .Y(n298) );
  INVX1 U104 ( .A(pos_dacis[0]), .Y(n295) );
  MUX2BXL U105 ( .D0(r_rpt_v[3]), .D1(n206), .S(n137), .Y(n65) );
  MUX2BXL U106 ( .D0(r_rpt_v[4]), .D1(n3), .S(n137), .Y(n66) );
  MUX2BXL U107 ( .D0(r_rpt_v[5]), .D1(n223), .S(n137), .Y(n67) );
  MUX2BXL U108 ( .D0(r_rpt_v[6]), .D1(n205), .S(n137), .Y(n68) );
  MUX2BXL U109 ( .D0(r_rpt_v[7]), .D1(n7), .S(n137), .Y(n69) );
  MUX2XL U110 ( .D0(x_daclsb[5]), .D1(n6), .S(r_wr[3]), .Y(wdlsb[5]) );
  MUX2XL U111 ( .D0(x_daclsb[4]), .D1(n8), .S(r_wr[3]), .Y(wdlsb[4]) );
  MUX2XL U112 ( .D0(r_rpt_v[1]), .D1(n60), .S(r_wr[3]), .Y(wdlsb[1]) );
  MUX2XL U113 ( .D0(x_daclsb[2]), .D1(n4), .S(r_wr[3]), .Y(wdlsb[2]) );
  MUX2XL U114 ( .D0(x_daclsb[3]), .D1(r_wdat[4]), .S(r_wr[3]), .Y(wdlsb[3]) );
  OAI222XL U115 ( .A(n209), .B(n535), .C(n210), .D(n536), .E(cs_ptr[4]), .F(
        n435), .Y(n140) );
  INVX1 U116 ( .A(dacv_wr[7]), .Y(n228) );
  INVX1 U117 ( .A(dacv_wr[4]), .Y(n232) );
  INVX1 U118 ( .A(dacv_wr[5]), .Y(n230) );
  INVX1 U119 ( .A(dacv_wr[6]), .Y(n229) );
  INVX1 U120 ( .A(n162), .Y(n530) );
  INVX1 U121 ( .A(dacv_wr[9]), .Y(n288) );
  NAND21X1 U122 ( .B(n102), .A(n99), .Y(n162) );
  NAND2X1 U123 ( .A(n102), .B(n99), .Y(n159) );
  INVX1 U124 ( .A(n193), .Y(n529) );
  NAND21X1 U125 ( .B(n99), .A(n73), .Y(n150) );
  NAND21X1 U126 ( .B(n99), .A(n71), .Y(n158) );
  NAND21X1 U127 ( .B(n99), .A(n72), .Y(n155) );
  INVXL U128 ( .A(dacv_wr[16]), .Y(n280) );
  INVX1 U129 ( .A(dacv_wr[17]), .Y(n278) );
  INVX1 U130 ( .A(dacv_wr[15]), .Y(n282) );
  INVX1 U131 ( .A(dacv_wr[8]), .Y(n291) );
  INVXL U132 ( .A(dacv_wr[14]), .Y(n283) );
  INVX1 U133 ( .A(dacv_wr[12]), .Y(n285) );
  NAND21X1 U134 ( .B(n99), .A(n103), .Y(n193) );
  INVX1 U135 ( .A(n101), .Y(n99) );
  NOR2X1 U136 ( .A(n101), .B(n11), .Y(n321) );
  INVX1 U137 ( .A(n103), .Y(n102) );
  NOR2X1 U138 ( .A(n10), .B(n99), .Y(n323) );
  NAND2X1 U139 ( .A(n102), .B(n101), .Y(n161) );
  NOR2X1 U140 ( .A(n104), .B(n143), .Y(n71) );
  NOR2X1 U141 ( .A(n104), .B(n156), .Y(n72) );
  NOR2X1 U142 ( .A(n156), .B(n102), .Y(n330) );
  NOR2X1 U143 ( .A(n104), .B(n151), .Y(n73) );
  NOR2X1 U144 ( .A(n151), .B(n102), .Y(n337) );
  NOR2X1 U145 ( .A(n143), .B(n102), .Y(n333) );
  NAND21X1 U146 ( .B(n101), .A(n56), .Y(n149) );
  NAND21X1 U147 ( .B(n101), .A(n74), .Y(n146) );
  NAND21X1 U148 ( .B(n99), .A(n62), .Y(n147) );
  NAND21X1 U149 ( .B(n101), .A(n47), .Y(n154) );
  NAND21X1 U150 ( .B(n101), .A(n43), .Y(n157) );
  NAND32X1 U151 ( .B(n96), .C(n458), .A(n95), .Y(n239) );
  AO21X1 U152 ( .B(r_wr[0]), .C(n235), .A(n458), .Y(n95) );
  NAND21X1 U153 ( .B(n50), .A(r_wr[0]), .Y(n234) );
  INVX3 U154 ( .A(n245), .Y(n264) );
  INVX2 U155 ( .A(n244), .Y(n261) );
  INVX1 U156 ( .A(n482), .Y(n488) );
  INVX1 U157 ( .A(n428), .Y(n455) );
  NAND21X1 U158 ( .B(n427), .A(n426), .Y(n428) );
  INVX1 U159 ( .A(n60), .Y(n206) );
  INVX1 U160 ( .A(r_wdat[4]), .Y(n205) );
  INVX1 U161 ( .A(n238), .Y(n100) );
  INVX1 U162 ( .A(r_wdat[3]), .Y(n223) );
  OAI22AX1 U163 ( .D(dacv_wr[1]), .C(n55), .A(n151), .B(n289), .Y(upd[1]) );
  OAI22AX1 U164 ( .D(dacv_wr[0]), .C(n55), .A(n151), .B(n292), .Y(upd[0]) );
  OAI22X1 U165 ( .A(n148), .B(n289), .C(n230), .D(n54), .Y(upd[5]) );
  OAI22X1 U166 ( .A(n143), .B(n292), .C(n291), .D(n54), .Y(upd[8]) );
  OAI22X1 U167 ( .A(n148), .B(n292), .C(n232), .D(n54), .Y(upd[4]) );
  OAI22X1 U168 ( .A(n156), .B(n289), .C(n284), .D(n54), .Y(upd[13]) );
  OAI22X1 U169 ( .A(n156), .B(n292), .C(n285), .D(n54), .Y(upd[12]) );
  OAI22X1 U170 ( .A(n143), .B(n289), .C(n288), .D(n54), .Y(upd[9]) );
  OAI22X1 U171 ( .A(n278), .B(n54), .C(n152), .D(n137), .Y(upd[17]) );
  OAI22X1 U173 ( .A(n280), .B(n54), .C(n153), .D(n137), .Y(upd[16]) );
  OAI22X1 U174 ( .A(n282), .B(n55), .C(n154), .D(n63), .Y(upd[15]) );
  OAI22X1 U200 ( .A(n283), .B(n55), .C(n155), .D(n63), .Y(upd[14]) );
  OAI22X1 U202 ( .A(n286), .B(n55), .C(n157), .D(n63), .Y(upd[11]) );
  OAI22X1 U203 ( .A(n287), .B(n55), .C(n158), .D(n63), .Y(upd[10]) );
  OAI22X1 U204 ( .A(n228), .B(n55), .C(n146), .D(n63), .Y(upd[7]) );
  OAI22X1 U205 ( .A(n229), .B(n55), .C(n147), .D(n63), .Y(upd[6]) );
  OAI22AX1 U206 ( .D(dacv_wr[3]), .C(n55), .A(n149), .B(n63), .Y(upd[3]) );
  OAI22AX1 U207 ( .D(dacv_wr[2]), .C(n55), .A(n150), .B(n63), .Y(upd[2]) );
  INVX1 U208 ( .A(n237), .Y(n94) );
  INVX1 U209 ( .A(N1423), .Y(n552) );
  INVX1 U210 ( .A(N1434), .Y(n553) );
  INVX1 U211 ( .A(N1346), .Y(n545) );
  INVX1 U212 ( .A(N1335), .Y(n544) );
  INVX1 U213 ( .A(N1412), .Y(n551) );
  INVX1 U214 ( .A(N1368), .Y(n547) );
  INVX1 U215 ( .A(N1357), .Y(n546) );
  INVX1 U216 ( .A(N1401), .Y(n550) );
  INVX1 U217 ( .A(N1379), .Y(n548) );
  INVX1 U218 ( .A(N1390), .Y(n549) );
  INVX1 U219 ( .A(n514), .Y(n515) );
  NAND21X1 U220 ( .B(n562), .A(N1291), .Y(n514) );
  AND2X1 U221 ( .A(n60), .B(r_wr[4]), .Y(clrsta[1]) );
  AND2X1 U222 ( .A(r_wr[4]), .B(n9), .Y(clrsta[5]) );
  AND2X1 U223 ( .A(r_wr[4]), .B(r_wdat[3]), .Y(clrsta[3]) );
  INVX1 U227 ( .A(N1280), .Y(n513) );
  INVX1 U228 ( .A(N1324), .Y(n525) );
  INVX1 U229 ( .A(N1291), .Y(n516) );
  INVX1 U230 ( .A(N1247), .Y(n504) );
  INVX1 U231 ( .A(N1302), .Y(n519) );
  INVX1 U232 ( .A(N1313), .Y(n522) );
  INVX1 U233 ( .A(N1258), .Y(n507) );
  INVX1 U234 ( .A(n511), .Y(n512) );
  NAND21X1 U235 ( .B(r_adofs[7]), .A(N1280), .Y(n511) );
  INVX1 U236 ( .A(n523), .Y(n524) );
  NAND21X1 U237 ( .B(r_adofs[7]), .A(N1324), .Y(n523) );
  INVX1 U238 ( .A(n502), .Y(n503) );
  NAND21X1 U239 ( .B(n562), .A(N1247), .Y(n502) );
  INVX1 U240 ( .A(n517), .Y(n518) );
  NAND21X1 U241 ( .B(r_adofs[7]), .A(N1302), .Y(n517) );
  INVX1 U242 ( .A(n505), .Y(n506) );
  NAND21X1 U243 ( .B(n562), .A(N1258), .Y(n505) );
  AND2X1 U244 ( .A(r_wr[4]), .B(n4), .Y(clrsta[2]) );
  AND2X1 U245 ( .A(r_wr[4]), .B(r_wdat[7]), .Y(clrsta[7]) );
  INVX1 U246 ( .A(cs_ptr[1]), .Y(n103) );
  INVX1 U247 ( .A(cs_ptr[0]), .Y(n101) );
  NAND21X1 U248 ( .B(cs_ptr[4]), .A(n528), .Y(n151) );
  NAND21X1 U249 ( .B(cs_ptr[4]), .A(n527), .Y(n156) );
  NAND21X1 U250 ( .B(cs_ptr[4]), .A(n526), .Y(n143) );
  NOR2X1 U251 ( .A(n104), .B(n148), .Y(n74) );
  NOR2X1 U252 ( .A(n148), .B(n102), .Y(n335) );
  INVX1 U253 ( .A(n227), .Y(n531) );
  NAND21X1 U254 ( .B(cs_ptr[4]), .A(n533), .Y(n227) );
  INVX1 U255 ( .A(cs_ptr[1]), .Y(n104) );
  NAND2X1 U256 ( .A(cs_ptr[4]), .B(n101), .Y(n210) );
  NAND2X1 U257 ( .A(cs_ptr[4]), .B(n99), .Y(n209) );
  INVX1 U258 ( .A(dacyc_done), .Y(n558) );
  NOR2X1 U259 ( .A(n162), .B(n160), .Y(setsta[5]) );
  NOR2X1 U260 ( .A(n162), .B(n195), .Y(setsta[1]) );
  NOR2X1 U261 ( .A(n161), .B(n160), .Y(setsta[6]) );
  NOR2X1 U262 ( .A(n193), .B(n195), .Y(setsta[0]) );
  NOR2X1 U263 ( .A(n161), .B(n195), .Y(setsta[2]) );
  NOR2X1 U264 ( .A(n159), .B(n160), .Y(setsta[7]) );
  NOR2X1 U265 ( .A(n159), .B(n195), .Y(setsta[3]) );
  NOR2X1 U266 ( .A(n193), .B(n160), .Y(setsta[4]) );
  INVX1 U267 ( .A(n231), .Y(n137) );
  NAND21X1 U268 ( .B(n162), .A(n231), .Y(n289) );
  NAND21X1 U269 ( .B(n193), .A(n231), .Y(n292) );
  NAND21X1 U270 ( .B(n162), .A(n279), .Y(n152) );
  NAND21X1 U271 ( .B(n193), .A(n279), .Y(n153) );
  INVX1 U272 ( .A(n329), .Y(n331) );
  AO21X1 U273 ( .B(N1243), .C(n504), .A(n503), .Y(o_dacv[4]) );
  AO21X1 U274 ( .B(N1242), .C(n504), .A(n503), .Y(o_dacv[3]) );
  AO21X1 U275 ( .B(N1246), .C(n504), .A(n503), .Y(o_dacv[7]) );
  AO21X1 U276 ( .B(N1266), .C(n510), .A(n509), .Y(o_dacv[21]) );
  AO21X1 U277 ( .B(N1253), .C(n507), .A(n506), .Y(o_dacv[11]) );
  NAND21X2 U278 ( .B(n274), .A(n273), .Y(n275) );
  AND2XL U279 ( .A(n239), .B(n238), .Y(n274) );
  GEN2XL U280 ( .D(n460), .E(n459), .C(n478), .B(n455), .A(n434), .Y(n479) );
  AND3X1 U281 ( .A(n433), .B(n478), .C(n432), .Y(n434) );
  AO21X1 U282 ( .B(N1241), .C(n504), .A(n503), .Y(o_dacv[2]) );
  NAND21X1 U283 ( .B(n500), .A(n483), .Y(n482) );
  AO21X1 U284 ( .B(N1255), .C(n507), .A(n506), .Y(o_dacv[13]) );
  AO21X1 U285 ( .B(N1263), .C(n510), .A(n509), .Y(o_dacv[18]) );
  OAI211X1 U286 ( .C(n313), .D(n311), .A(n310), .B(n307), .Y(n329) );
  AO21X1 U287 ( .B(n461), .C(n462), .A(n475), .Y(n460) );
  OR2X1 U288 ( .A(n418), .B(n75), .Y(n427) );
  AOI21X1 U289 ( .B(n462), .C(n420), .A(n470), .Y(n75) );
  NAND32X1 U290 ( .B(n1), .C(n329), .A(n463), .Y(n314) );
  AO21X1 U291 ( .B(N1244), .C(n504), .A(n503), .Y(o_dacv[5]) );
  INVX1 U292 ( .A(n413), .Y(n433) );
  OAI22X1 U293 ( .A(n459), .B(n495), .C(n478), .D(n429), .Y(n467) );
  AND2X1 U294 ( .A(n455), .B(n460), .Y(n429) );
  OAI211X1 U295 ( .C(n488), .D(n487), .A(n486), .B(n485), .Y(n499) );
  OAI211X1 U296 ( .C(n311), .D(n307), .A(n310), .B(n313), .Y(n465) );
  AO21X1 U297 ( .B(N1245), .C(n504), .A(n503), .Y(o_dacv[6]) );
  AO21X1 U298 ( .B(N1240), .C(n504), .A(n503), .Y(o_dacv[1]) );
  AO21X1 U299 ( .B(N1265), .C(n510), .A(n509), .Y(o_dacv[20]) );
  AO21X1 U300 ( .B(N1262), .C(n510), .A(n509), .Y(o_dacv[17]) );
  AO21X1 U301 ( .B(N1264), .C(n510), .A(n509), .Y(o_dacv[19]) );
  AO21X1 U302 ( .B(N1261), .C(n510), .A(n509), .Y(o_dacv[16]) );
  AO21X1 U303 ( .B(N1267), .C(n510), .A(n509), .Y(o_dacv[22]) );
  AO21X1 U304 ( .B(N1268), .C(n510), .A(n509), .Y(o_dacv[23]) );
  AND2X1 U305 ( .A(n494), .B(n488), .Y(n76) );
  INVX1 U306 ( .A(n474), .Y(n483) );
  OAI211X1 U307 ( .C(n480), .D(n484), .A(n479), .B(n486), .Y(n474) );
  INVX1 U308 ( .A(n1), .Y(n313) );
  INVX1 U309 ( .A(n224), .Y(n276) );
  INVX1 U310 ( .A(n334), .Y(n470) );
  NAND2X1 U311 ( .A(n77), .B(n461), .Y(n476) );
  NAND4X1 U312 ( .A(n463), .B(n1), .C(n430), .D(n466), .Y(n77) );
  NAND6XL U313 ( .A(n9), .B(r_wdat[3]), .C(n4), .D(n226), .E(n225), .F(n5), 
        .Y(n237) );
  INVX1 U314 ( .A(n423), .Y(n426) );
  INVX1 U315 ( .A(n294), .Y(n461) );
  NAND21X1 U316 ( .B(n334), .A(n426), .Y(n294) );
  AO21X1 U317 ( .B(N1285), .C(n516), .A(n515), .Y(o_dacv[34]) );
  INVX1 U318 ( .A(n109), .Y(n106) );
  INVX1 U319 ( .A(n109), .Y(n107) );
  NAND2X1 U320 ( .A(N1423), .B(n114), .Y(n317) );
  NAND2X1 U321 ( .A(N1434), .B(n114), .Y(n316) );
  NAND2X1 U322 ( .A(N1346), .B(n114), .Y(n308) );
  NAND2X1 U323 ( .A(N1335), .B(n114), .Y(n309) );
  NAND2X1 U324 ( .A(N1412), .B(n114), .Y(n318) );
  NAND2X1 U325 ( .A(N1368), .B(n114), .Y(n305) );
  NAND2X1 U326 ( .A(N1357), .B(n114), .Y(n306) );
  NAND2X1 U327 ( .A(N1401), .B(n114), .Y(n319) );
  NAND2X1 U328 ( .A(N1379), .B(n114), .Y(n304) );
  NAND2X1 U329 ( .A(N1390), .B(n114), .Y(n320) );
  INVX1 U330 ( .A(n109), .Y(r_adofs[0]) );
  OAI21BBX1 U331 ( .A(N1367), .B(n547), .C(n305), .Y(o_dacv[95]) );
  OAI21BBX1 U332 ( .A(N1356), .B(n546), .C(n306), .Y(o_dacv[87]) );
  OAI21BBX1 U333 ( .A(N1400), .B(n550), .C(n319), .Y(o_dacv[119]) );
  OAI21BBX1 U334 ( .A(N1378), .B(n548), .C(n304), .Y(o_dacv[103]) );
  OAI21BBX1 U335 ( .A(N1389), .B(n549), .C(n320), .Y(o_dacv[111]) );
  AO21X1 U336 ( .B(N1295), .C(n519), .A(n518), .Y(o_dacv[41]) );
  AO21X1 U337 ( .B(N1284), .C(n516), .A(n515), .Y(o_dacv[33]) );
  AO21X1 U338 ( .B(N1297), .C(n519), .A(n518), .Y(o_dacv[43]) );
  AO21X1 U339 ( .B(N1275), .C(n513), .A(n512), .Y(o_dacv[27]) );
  AO21X1 U340 ( .B(N1276), .C(n513), .A(n512), .Y(o_dacv[28]) );
  AO21X1 U341 ( .B(N1277), .C(n513), .A(n512), .Y(o_dacv[29]) );
  AO21X1 U342 ( .B(N1279), .C(n513), .A(n512), .Y(o_dacv[31]) );
  AO21X1 U343 ( .B(N1273), .C(n513), .A(n512), .Y(o_dacv[25]) );
  AO21X1 U344 ( .B(N1254), .C(n507), .A(n506), .Y(o_dacv[12]) );
  AO21X1 U345 ( .B(N1257), .C(n507), .A(n506), .Y(o_dacv[15]) );
  AO21X1 U346 ( .B(N1310), .C(n522), .A(n521), .Y(o_dacv[53]) );
  AO21X1 U347 ( .B(N1322), .C(n525), .A(n524), .Y(o_dacv[62]) );
  AO21X1 U348 ( .B(N1323), .C(n525), .A(n524), .Y(o_dacv[63]) );
  AO21X1 U349 ( .B(N1307), .C(n522), .A(n521), .Y(o_dacv[50]) );
  INVX1 U350 ( .A(n520), .Y(n521) );
  NAND21X1 U351 ( .B(r_adofs[7]), .A(N1313), .Y(n520) );
  AO21X1 U352 ( .B(N1300), .C(n519), .A(n518), .Y(o_dacv[46]) );
  AO21X1 U353 ( .B(N1256), .C(n507), .A(n506), .Y(o_dacv[14]) );
  INVX1 U354 ( .A(N1269), .Y(n510) );
  OAI21BBX1 U355 ( .A(N1365), .B(n547), .C(n305), .Y(o_dacv[93]) );
  OAI21BBX1 U356 ( .A(N1354), .B(n546), .C(n306), .Y(o_dacv[85]) );
  OAI21BBX1 U357 ( .A(N1398), .B(n550), .C(n319), .Y(o_dacv[117]) );
  OAI21BBX1 U358 ( .A(N1376), .B(n548), .C(n304), .Y(o_dacv[101]) );
  OAI21BBX1 U359 ( .A(N1387), .B(n549), .C(n320), .Y(o_dacv[109]) );
  OAI21BBX1 U360 ( .A(N1361), .B(n547), .C(n305), .Y(o_dacv[89]) );
  OAI21BBX1 U361 ( .A(N1350), .B(n546), .C(n306), .Y(o_dacv[81]) );
  OAI21BBX1 U362 ( .A(N1394), .B(n550), .C(n319), .Y(o_dacv[113]) );
  OAI21BBX1 U363 ( .A(N1372), .B(n548), .C(n304), .Y(o_dacv[97]) );
  OAI21BBX1 U364 ( .A(N1383), .B(n549), .C(n320), .Y(o_dacv[105]) );
  OAI21BBX1 U365 ( .A(N1364), .B(n547), .C(n305), .Y(o_dacv[92]) );
  OAI21BBX1 U366 ( .A(N1353), .B(n546), .C(n306), .Y(o_dacv[84]) );
  OAI21BBX1 U367 ( .A(N1397), .B(n550), .C(n319), .Y(o_dacv[116]) );
  OAI21BBX1 U368 ( .A(N1375), .B(n548), .C(n304), .Y(o_dacv[100]) );
  OAI21BBX1 U369 ( .A(N1386), .B(n549), .C(n320), .Y(o_dacv[108]) );
  OAI21BBX1 U370 ( .A(N1363), .B(n547), .C(n305), .Y(o_dacv[91]) );
  OAI21BBX1 U371 ( .A(N1352), .B(n546), .C(n306), .Y(o_dacv[83]) );
  OAI21BBX1 U372 ( .A(N1396), .B(n550), .C(n319), .Y(o_dacv[115]) );
  OAI21BBX1 U373 ( .A(N1374), .B(n548), .C(n304), .Y(o_dacv[99]) );
  OAI21BBX1 U374 ( .A(N1385), .B(n549), .C(n320), .Y(o_dacv[107]) );
  OAI21BBX1 U375 ( .A(N1362), .B(n547), .C(n305), .Y(o_dacv[90]) );
  OAI21BBX1 U376 ( .A(N1351), .B(n546), .C(n306), .Y(o_dacv[82]) );
  OAI21BBX1 U377 ( .A(N1395), .B(n550), .C(n319), .Y(o_dacv[114]) );
  OAI21BBX1 U378 ( .A(N1373), .B(n548), .C(n304), .Y(o_dacv[98]) );
  OAI21BBX1 U379 ( .A(N1384), .B(n549), .C(n320), .Y(o_dacv[106]) );
  OAI21BBX1 U380 ( .A(N1366), .B(n547), .C(n305), .Y(o_dacv[94]) );
  OAI21BBX1 U381 ( .A(N1355), .B(n546), .C(n306), .Y(o_dacv[86]) );
  OAI21BBX1 U382 ( .A(N1399), .B(n550), .C(n319), .Y(o_dacv[118]) );
  OAI21BBX1 U383 ( .A(N1377), .B(n548), .C(n304), .Y(o_dacv[102]) );
  OAI21BBX1 U384 ( .A(N1388), .B(n549), .C(n320), .Y(o_dacv[110]) );
  INVX1 U385 ( .A(n115), .Y(n110) );
  INVX1 U386 ( .A(n501), .Y(n490) );
  INVX1 U387 ( .A(n115), .Y(n111) );
  INVX1 U388 ( .A(n115), .Y(n112) );
  INVX1 U389 ( .A(n203), .Y(n528) );
  INVX1 U390 ( .A(n281), .Y(n527) );
  NAND21X1 U391 ( .B(n534), .A(cs_ptr[3]), .Y(n281) );
  NAND2X1 U392 ( .A(o_dactl[0]), .B(n140), .Y(n412) );
  INVX1 U393 ( .A(n218), .Y(n526) );
  INVX1 U394 ( .A(cs_ptr[3]), .Y(n533) );
  OAI22X1 U395 ( .A(n218), .B(n540), .C(n204), .D(n555), .Y(n443) );
  INVX1 U396 ( .A(n204), .Y(n559) );
  NAND21X1 U397 ( .B(n534), .A(n531), .Y(n148) );
  NOR32XL U398 ( .B(cs_ptr[4]), .C(n103), .A(n203), .Y(n336) );
  OAI21AX1 U399 ( .B(n63), .C(n138), .A(r_wr[3]), .Y(updlsb) );
  INVX1 U400 ( .A(n207), .Y(n96) );
  AND3X1 U401 ( .A(n541), .B(n542), .C(n557), .Y(n78) );
  MUX2BXL U402 ( .D0(n558), .D1(sacyc_done), .S(n456), .Y(n238) );
  INVX1 U403 ( .A(n233), .Y(n456) );
  NAND21X1 U404 ( .B(n96), .A(n140), .Y(n233) );
  INVX1 U405 ( .A(o_dactl[0]), .Y(n235) );
  INVX1 U406 ( .A(n138), .Y(n64) );
  NAND21X1 U407 ( .B(n148), .A(n194), .Y(n160) );
  NAND21X1 U408 ( .B(n151), .A(n194), .Y(n195) );
  NAND2X1 U409 ( .A(n301), .B(n302), .Y(o_intr) );
  NOR4XL U410 ( .A(r_irq[3]), .B(r_irq[2]), .C(r_irq[1]), .D(r_irq[0]), .Y(
        n301) );
  NOR4XL U411 ( .A(r_irq[7]), .B(r_irq[6]), .C(r_irq[5]), .D(r_irq[4]), .Y(
        n302) );
  AO21X1 U412 ( .B(n96), .C(dacyc_done), .A(sacyc_done), .Y(n231) );
  AOI21X1 U413 ( .B(n207), .C(n208), .A(n558), .Y(sar_nxt) );
  NAND2X1 U414 ( .A(n141), .B(n140), .Y(n208) );
  NOR2X1 U415 ( .A(n139), .B(n558), .Y(updcmp) );
  XNOR2XL U416 ( .A(n140), .B(n141), .Y(n139) );
  OAI22X1 U417 ( .A(n151), .B(n444), .C(n450), .D(n561), .Y(datcmp[1]) );
  NOR2X1 U418 ( .A(n162), .B(n151), .Y(n450) );
  OAI22X1 U419 ( .A(n148), .B(n444), .C(n448), .D(n560), .Y(datcmp[5]) );
  NOR2X1 U420 ( .A(n162), .B(n148), .Y(n448) );
  INVX1 U421 ( .A(n277), .Y(n279) );
  NAND21X1 U422 ( .B(n203), .A(cs_ptr[4]), .Y(n277) );
  NAND21X1 U423 ( .B(n501), .A(n500), .Y(o_smpl[4]) );
  AO21X1 U424 ( .B(N1312), .C(n522), .A(n521), .Y(o_dacv[55]) );
  AO21X1 U425 ( .B(N1311), .C(n522), .A(n521), .Y(o_dacv[54]) );
  AO21X1 U426 ( .B(N1251), .C(n507), .A(n506), .Y(o_dacv[9]) );
  AO21X1 U427 ( .B(N1288), .C(n516), .A(n515), .Y(o_dacv[37]) );
  AO21X1 U428 ( .B(N1287), .C(n516), .A(n515), .Y(o_dacv[36]) );
  AO21X1 U429 ( .B(N1286), .C(n516), .A(n515), .Y(o_dacv[35]) );
  AO21X1 U430 ( .B(N1299), .C(n519), .A(n518), .Y(o_dacv[45]) );
  AO21X1 U431 ( .B(N1320), .C(n525), .A(n524), .Y(o_dacv[60]) );
  AO21X1 U432 ( .B(N1278), .C(n513), .A(n512), .Y(o_dacv[30]) );
  AO21X1 U433 ( .B(N1298), .C(n519), .A(n518), .Y(o_dacv[44]) );
  AO21X1 U434 ( .B(N1294), .C(n519), .A(n518), .Y(o_dacv[40]) );
  NAND31X1 U435 ( .C(n423), .A(n422), .B(n421), .Y(n468) );
  NAND21X1 U436 ( .B(n420), .A(pos_dacis[9]), .Y(n421) );
  NAND21X1 U437 ( .B(n470), .A(n419), .Y(n422) );
  AO21X1 U438 ( .B(N1290), .C(n516), .A(n515), .Y(o_dacv[39]) );
  AO2222X1 U439 ( .A(n263), .B(r_sar_en[6]), .C(n260), .D(r_sar_en[0]), .E(
        n261), .F(r_sar_en[2]), .G(n264), .H(r_sar_en[4]), .Y(n247) );
  AO2222X1 U440 ( .A(r_dac_en[12]), .B(n264), .C(r_dac_en[14]), .D(n263), .E(
        r_dac_en[8]), .F(n262), .G(r_dac_en[10]), .H(n261), .Y(n250) );
  AO2222X1 U441 ( .A(r_dac_en[13]), .B(n264), .C(n263), .D(r_dac_en[15]), .E(
        r_dac_en[9]), .F(n262), .G(r_dac_en[11]), .H(n261), .Y(n256) );
  AO21X1 U442 ( .B(N1296), .C(n519), .A(n518), .Y(o_dacv[42]) );
  AO21X1 U443 ( .B(N1283), .C(n516), .A(n515), .Y(o_dacv[32]) );
  AO21X1 U444 ( .B(N1301), .C(n519), .A(n518), .Y(o_dacv[47]) );
  NAND31X1 U445 ( .C(pos_dacis[6]), .A(n79), .B(n466), .Y(n469) );
  MUX2IX1 U446 ( .D0(n465), .D1(n464), .S(n463), .Y(n79) );
  NAND2X1 U447 ( .A(n315), .B(n430), .Y(n80) );
  MUX3X1 U448 ( .D0(n465), .D1(n313), .D2(n314), .S0(n463), .S1(pos_dacis[6]), 
        .Y(n332) );
  AO21X1 U449 ( .B(N1239), .C(n504), .A(n503), .Y(o_dacv[0]) );
  AO21X1 U450 ( .B(N1319), .C(n525), .A(n524), .Y(o_dacv[59]) );
  NAND3X1 U451 ( .A(n480), .B(n479), .C(n486), .Y(n81) );
  XOR2X1 U452 ( .A(n298), .B(pos_dacis[2]), .Y(n300) );
  NAND21X1 U453 ( .B(n499), .A(n498), .Y(o_smpl[3]) );
  NAND21X1 U454 ( .B(n501), .A(n497), .Y(n498) );
  NAND21X1 U455 ( .B(n496), .A(n495), .Y(n497) );
  AO21X1 U456 ( .B(N1252), .C(n507), .A(n506), .Y(o_dacv[10]) );
  OAI22X1 U457 ( .A(n432), .B(n425), .C(n433), .D(n424), .Y(n475) );
  INVX1 U458 ( .A(pos_dacis[11]), .Y(n425) );
  INVX1 U459 ( .A(n468), .Y(n424) );
  AO21X1 U460 ( .B(n490), .C(n489), .A(n499), .Y(o_smpl[1]) );
  AO21X1 U461 ( .B(N1309), .C(n522), .A(n521), .Y(o_dacv[52]) );
  NAND5XL U462 ( .A(n478), .B(n477), .C(n476), .D(n486), .E(n484), .Y(n481) );
  INVX1 U463 ( .A(n475), .Y(n477) );
  INVX1 U464 ( .A(n476), .Y(n471) );
  INVX1 U465 ( .A(n297), .Y(n310) );
  OAI211XL U466 ( .C(n299), .D(n298), .A(n296), .B(n295), .Y(n297) );
  INVX1 U467 ( .A(pos_dacis[2]), .Y(n296) );
  AO21XL U468 ( .B(n494), .C(n493), .A(n492), .Y(o_smpl[2]) );
  INVX1 U469 ( .A(pos_dacis[17]), .Y(n493) );
  AO21X1 U470 ( .B(N1318), .C(n525), .A(n524), .Y(o_dacv[58]) );
  AO21X1 U471 ( .B(N1317), .C(n525), .A(n524), .Y(o_dacv[57]) );
  AO21X1 U472 ( .B(N1308), .C(n522), .A(n521), .Y(o_dacv[51]) );
  AO21X1 U473 ( .B(N1316), .C(n525), .A(n524), .Y(o_dacv[56]) );
  INVX1 U474 ( .A(n312), .Y(n463) );
  NAND21X1 U475 ( .B(pos_dacis[4]), .A(n311), .Y(n312) );
  AO21XL U476 ( .B(n483), .C(n490), .A(n76), .Y(o_smpl[0]) );
  INVX1 U477 ( .A(pos_dacis[5]), .Y(n311) );
  INVX1 U478 ( .A(pos_dacis[4]), .Y(n307) );
  NOR21XL U479 ( .B(app_dacis[10]), .A(n98), .Y(o_daci_sel[10]) );
  NOR21XL U480 ( .B(app_dacis[7]), .A(n98), .Y(o_daci_sel[7]) );
  NOR21XL U481 ( .B(app_dacis[8]), .A(n97), .Y(o_daci_sel[8]) );
  NOR21XL U482 ( .B(app_dacis[11]), .A(n97), .Y(o_daci_sel[11]) );
  NOR21XL U483 ( .B(app_dacis[16]), .A(n98), .Y(o_daci_sel[16]) );
  NOR21XL U484 ( .B(app_dacis[3]), .A(n98), .Y(o_daci_sel[3]) );
  NOR21XL U485 ( .B(app_dacis[4]), .A(n97), .Y(o_daci_sel[4]) );
  NOR21XL U486 ( .B(app_dacis[6]), .A(n97), .Y(o_daci_sel[6]) );
  NOR21XL U487 ( .B(app_dacis[5]), .A(n98), .Y(o_daci_sel[5]) );
  NOR21XL U488 ( .B(app_dacis[2]), .A(n97), .Y(o_daci_sel[2]) );
  NOR21XL U489 ( .B(app_dacis[0]), .A(n97), .Y(o_daci_sel[0]) );
  NOR21XL U490 ( .B(app_dacis[1]), .A(n98), .Y(o_daci_sel[1]) );
  NOR21XL U491 ( .B(app_dacis[17]), .A(n97), .Y(o_daci_sel[17]) );
  NOR21XL U492 ( .B(app_dacis[14]), .A(n98), .Y(o_daci_sel[14]) );
  INVX1 U493 ( .A(n222), .Y(n226) );
  NAND6XL U494 ( .A(r_wdat[7]), .B(n96), .C(n235), .D(n216), .E(n206), .F(n205), .Y(n222) );
  NAND43X1 U495 ( .B(n145), .C(n144), .D(n142), .A(n136), .Y(n216) );
  AO2222XL U496 ( .A(r_sar_en[2]), .B(dacv_wr[2]), .C(r_sar_en[3]), .D(
        dacv_wr[3]), .E(r_sar_en[0]), .F(dacv_wr[0]), .G(r_sar_en[1]), .H(
        dacv_wr[1]), .Y(n145) );
  NOR21XL U497 ( .B(app_dacis[15]), .A(n97), .Y(o_daci_sel[15]) );
  NOR21XL U498 ( .B(app_dacis[9]), .A(n98), .Y(o_daci_sel[9]) );
  INVX1 U499 ( .A(pos_dacis[6]), .Y(n430) );
  NOR21XL U500 ( .B(app_dacis[13]), .A(n97), .Y(o_daci_sel[13]) );
  NOR21XL U501 ( .B(app_dacis[12]), .A(n98), .Y(o_daci_sel[12]) );
  NAND21X1 U502 ( .B(pos_dacis[9]), .A(n420), .Y(n334) );
  NAND21X1 U503 ( .B(pos_dacis[11]), .A(n432), .Y(n423) );
  INVX1 U504 ( .A(pos_dacis[7]), .Y(n466) );
  OAI221X1 U505 ( .A(n230), .B(n129), .C(n556), .D(n232), .E(n128), .Y(n144)
         );
  INVX1 U506 ( .A(r_sar_en[5]), .Y(n129) );
  OA222X1 U507 ( .A(n555), .B(n229), .C(n291), .D(n127), .E(n554), .F(n228), 
        .Y(n128) );
  INVX1 U508 ( .A(r_sar_en[8]), .Y(n127) );
  OAI221X1 U509 ( .A(n283), .B(n133), .C(n284), .D(n132), .E(n131), .Y(n142)
         );
  INVX1 U510 ( .A(r_sar_en[14]), .Y(n133) );
  INVX1 U511 ( .A(r_sar_en[13]), .Y(n132) );
  OA222X1 U512 ( .A(n282), .B(n130), .C(n536), .D(n280), .E(n535), .F(n278), 
        .Y(n131) );
  INVX1 U513 ( .A(pos_dacis[8]), .Y(n420) );
  INVX1 U514 ( .A(pos_dacis[10]), .Y(n432) );
  OA2222XL U515 ( .A(n540), .B(n287), .C(n539), .D(n288), .E(n285), .F(n135), 
        .G(n286), .H(n134), .Y(n136) );
  INVX1 U516 ( .A(r_sar_en[12]), .Y(n135) );
  INVX1 U517 ( .A(r_sar_en[11]), .Y(n134) );
  INVX1 U518 ( .A(pos_dacis[12]), .Y(n459) );
  INVX1 U519 ( .A(n293), .Y(n478) );
  NAND21X1 U520 ( .B(pos_dacis[13]), .A(n459), .Y(n293) );
  OAI21BBX1 U521 ( .A(N1433), .B(n553), .C(n316), .Y(o_dacv[143]) );
  OAI21BBX1 U522 ( .A(N1334), .B(n544), .C(n309), .Y(o_dacv[71]) );
  OAI21BBX1 U523 ( .A(N1411), .B(n551), .C(n318), .Y(o_dacv[127]) );
  OAI21BBX1 U524 ( .A(N1345), .B(n545), .C(n308), .Y(o_dacv[79]) );
  BUFX3 U525 ( .A(n570), .Y(n82) );
  BUFX3 U526 ( .A(n570), .Y(r_adofs[1]) );
  MUX2AXL U527 ( .D0(r_rpt_v[8]), .D1(n5), .S(n137), .Y(n126) );
  INVX1 U528 ( .A(pos_dacis[13]), .Y(n495) );
  OAI21BBX1 U529 ( .A(N1422), .B(n552), .C(n317), .Y(o_dacv[135]) );
  INVX1 U530 ( .A(n571), .Y(n109) );
  MUX2AXL U531 ( .D0(r_rpt_v[2]), .D1(n225), .S(n137), .Y(n125) );
  BUFX3 U532 ( .A(n569), .Y(n84) );
  BUFX3 U533 ( .A(n569), .Y(r_adofs[2]) );
  AO21X1 U534 ( .B(N1272), .C(n513), .A(n512), .Y(o_dacv[24]) );
  AO21X1 U535 ( .B(N1250), .C(n507), .A(n506), .Y(o_dacv[8]) );
  OAI21BBX1 U536 ( .A(N1431), .B(n553), .C(n316), .Y(o_dacv[141]) );
  OAI21BBX1 U537 ( .A(N1427), .B(n553), .C(n316), .Y(o_dacv[137]) );
  OAI21BBX1 U538 ( .A(N1430), .B(n553), .C(n316), .Y(o_dacv[140]) );
  OAI21BBX1 U539 ( .A(N1429), .B(n553), .C(n316), .Y(o_dacv[139]) );
  OAI21BBX1 U540 ( .A(N1428), .B(n553), .C(n316), .Y(o_dacv[138]) );
  OAI21BBX1 U541 ( .A(N1332), .B(n544), .C(n309), .Y(o_dacv[69]) );
  OAI21BBX1 U542 ( .A(N1328), .B(n544), .C(n309), .Y(o_dacv[65]) );
  OAI21BBX1 U543 ( .A(N1331), .B(n544), .C(n309), .Y(o_dacv[68]) );
  OAI21BBX1 U544 ( .A(N1333), .B(n544), .C(n309), .Y(o_dacv[70]) );
  OAI21BBX1 U545 ( .A(N1327), .B(n544), .C(n309), .Y(o_dacv[64]) );
  OAI21BBX1 U546 ( .A(N1330), .B(n544), .C(n309), .Y(o_dacv[67]) );
  OAI21BBX1 U547 ( .A(N1329), .B(n544), .C(n309), .Y(o_dacv[66]) );
  OAI21BBX1 U548 ( .A(N1343), .B(n545), .C(n308), .Y(o_dacv[77]) );
  OAI21BBX1 U549 ( .A(N1339), .B(n545), .C(n308), .Y(o_dacv[73]) );
  OAI21BBX1 U550 ( .A(N1342), .B(n545), .C(n308), .Y(o_dacv[76]) );
  OAI21BBX1 U551 ( .A(N1344), .B(n545), .C(n308), .Y(o_dacv[78]) );
  OAI21BBX1 U552 ( .A(N1338), .B(n545), .C(n308), .Y(o_dacv[72]) );
  OAI21BBX1 U553 ( .A(N1341), .B(n545), .C(n308), .Y(o_dacv[75]) );
  OAI21BBX1 U554 ( .A(N1340), .B(n545), .C(n308), .Y(o_dacv[74]) );
  OAI21BBX1 U555 ( .A(N1409), .B(n551), .C(n318), .Y(o_dacv[125]) );
  OAI21BBX1 U556 ( .A(N1405), .B(n551), .C(n318), .Y(o_dacv[121]) );
  OAI21BBX1 U557 ( .A(N1408), .B(n551), .C(n318), .Y(o_dacv[124]) );
  OAI21BBX1 U558 ( .A(N1410), .B(n551), .C(n318), .Y(o_dacv[126]) );
  OAI21BBX1 U559 ( .A(N1404), .B(n551), .C(n318), .Y(o_dacv[120]) );
  OAI21BBX1 U560 ( .A(N1407), .B(n551), .C(n318), .Y(o_dacv[123]) );
  OAI21BBX1 U561 ( .A(N1406), .B(n551), .C(n318), .Y(o_dacv[122]) );
  BUFX3 U562 ( .A(n567), .Y(n88) );
  BUFX3 U563 ( .A(n568), .Y(n86) );
  BUFX3 U564 ( .A(n568), .Y(r_adofs[3]) );
  BUFX3 U565 ( .A(n567), .Y(r_adofs[4]) );
  INVX1 U566 ( .A(n508), .Y(n509) );
  NAND21X1 U567 ( .B(r_isofs[7]), .A(N1269), .Y(n508) );
  OAI21BBX1 U568 ( .A(N1426), .B(n553), .C(n316), .Y(o_dacv[136]) );
  OAI21BBX1 U569 ( .A(N1415), .B(n552), .C(n317), .Y(o_dacv[128]) );
  INVX1 U570 ( .A(pos_dacis[14]), .Y(n486) );
  OAI21BBX1 U571 ( .A(N1420), .B(n552), .C(n317), .Y(o_dacv[133]) );
  OAI21BBX1 U572 ( .A(N1416), .B(n552), .C(n317), .Y(o_dacv[129]) );
  OAI21BBX1 U573 ( .A(N1419), .B(n552), .C(n317), .Y(o_dacv[132]) );
  OAI21BBX1 U574 ( .A(N1418), .B(n552), .C(n317), .Y(o_dacv[131]) );
  OAI21BBX1 U575 ( .A(N1417), .B(n552), .C(n317), .Y(o_dacv[130]) );
  OAI21BBX1 U576 ( .A(N1360), .B(n547), .C(n305), .Y(o_dacv[88]) );
  OAI21BBX1 U577 ( .A(N1349), .B(n546), .C(n306), .Y(o_dacv[80]) );
  OAI21BBX1 U578 ( .A(N1393), .B(n550), .C(n319), .Y(o_dacv[112]) );
  OAI21BBX1 U579 ( .A(N1371), .B(n548), .C(n304), .Y(o_dacv[96]) );
  OAI21BBX1 U580 ( .A(N1382), .B(n549), .C(n320), .Y(o_dacv[104]) );
  INVX1 U581 ( .A(pos_dacis[15]), .Y(n484) );
  OAI21BBX1 U582 ( .A(N1421), .B(n552), .C(n317), .Y(o_dacv[134]) );
  OAI21BBX1 U583 ( .A(N1432), .B(n553), .C(n316), .Y(o_dacv[142]) );
  BUFX3 U584 ( .A(n564), .Y(n90) );
  BUFX3 U585 ( .A(n564), .Y(r_adofs[5]) );
  NAND21X1 U586 ( .B(pos_dacis[17]), .A(n487), .Y(n501) );
  BUFX3 U587 ( .A(n563), .Y(n92) );
  BUFX3 U588 ( .A(n563), .Y(r_adofs[6]) );
  INVX1 U589 ( .A(n562), .Y(n115) );
  INVX1 U590 ( .A(pos_dacis[16]), .Y(n487) );
  INVX1 U591 ( .A(n562), .Y(n114) );
  INVX1 U592 ( .A(n115), .Y(r_adofs[7]) );
  NAND21X1 U593 ( .B(cs_ptr[2]), .A(n533), .Y(n203) );
  AO222X1 U594 ( .A(n321), .B(n402), .C(n323), .D(n403), .E(r_dac1v[2]), .F(
        n10), .Y(o_dac1[2]) );
  NAND4X1 U595 ( .A(n408), .B(n409), .C(n410), .D(n411), .Y(n402) );
  NAND4X1 U596 ( .A(n404), .B(n405), .C(n406), .D(n407), .Y(n403) );
  AOI22X1 U597 ( .A(r_dacvs[136]), .B(n53), .C(r_dacvs[8]), .D(n46), .Y(n408)
         );
  AO222X1 U598 ( .A(n321), .B(n392), .C(n323), .D(n393), .E(r_dac1v[3]), .F(
        n11), .Y(o_dac1[3]) );
  NAND4X1 U599 ( .A(n398), .B(n399), .C(n400), .D(n401), .Y(n392) );
  NAND4X1 U600 ( .A(n394), .B(n395), .C(n396), .D(n397), .Y(n393) );
  AOI22X1 U601 ( .A(r_dacvs[137]), .B(n53), .C(r_dacvs[9]), .D(n46), .Y(n398)
         );
  NAND21X1 U602 ( .B(cs_ptr[2]), .A(cs_ptr[3]), .Y(n218) );
  NAND4X1 U603 ( .A(n378), .B(n379), .C(n380), .D(n381), .Y(n372) );
  NAND4X1 U604 ( .A(n374), .B(n375), .C(n376), .D(n377), .Y(n373) );
  AOI22X1 U605 ( .A(r_dacvs[139]), .B(n53), .C(r_dacvs[11]), .D(n46), .Y(n378)
         );
  OA2222XL U606 ( .A(n436), .B(n161), .C(n437), .D(n159), .E(n438), .F(n18), 
        .G(n439), .H(n59), .Y(n435) );
  AOI221XL U607 ( .A(r_sar_en[2]), .B(n528), .C(r_sar_en[14]), .D(n527), .E(
        n443), .Y(n436) );
  AOI221XL U608 ( .A(r_sar_en[1]), .B(n528), .C(r_sar_en[13]), .D(n527), .E(
        n441), .Y(n438) );
  AO222X1 U609 ( .A(n321), .B(n362), .C(n323), .D(n363), .E(r_dac1v[6]), .F(
        n10), .Y(o_dac1[6]) );
  NAND4X1 U610 ( .A(n368), .B(n369), .C(n370), .D(n371), .Y(n362) );
  NAND4X1 U611 ( .A(n364), .B(n365), .C(n366), .D(n367), .Y(n363) );
  AOI22X1 U612 ( .A(r_dacvs[140]), .B(n53), .C(r_dacvs[12]), .D(n46), .Y(n368)
         );
  AO222X1 U613 ( .A(n321), .B(n352), .C(n323), .D(n353), .E(r_dac1v[7]), .F(
        n10), .Y(o_dac1[7]) );
  NAND4X1 U614 ( .A(n358), .B(n359), .C(n360), .D(n361), .Y(n352) );
  NAND4X1 U615 ( .A(n354), .B(n355), .C(n356), .D(n357), .Y(n353) );
  AOI22X1 U616 ( .A(r_dacvs[141]), .B(n53), .C(r_dacvs[13]), .D(n46), .Y(n358)
         );
  AO222X1 U617 ( .A(n321), .B(n322), .C(n323), .D(n324), .E(r_dac1v[9]), .F(
        n11), .Y(o_dac1[9]) );
  NAND4X1 U618 ( .A(n338), .B(n339), .C(n340), .D(n341), .Y(n322) );
  NAND4X1 U619 ( .A(n325), .B(n326), .C(n327), .D(n328), .Y(n324) );
  AOI22X1 U620 ( .A(r_dacvs[143]), .B(n53), .C(r_dacvs[15]), .D(n46), .Y(n338)
         );
  AO222X1 U621 ( .A(n321), .B(n382), .C(n323), .D(n383), .E(r_dac1v[4]), .F(
        n10), .Y(o_dac1[4]) );
  NAND4X1 U622 ( .A(n388), .B(n389), .C(n390), .D(n391), .Y(n382) );
  NAND4X1 U623 ( .A(n384), .B(n385), .C(n386), .D(n387), .Y(n383) );
  AOI22X1 U624 ( .A(r_dacvs[138]), .B(n336), .C(r_dacvs[10]), .D(n337), .Y(
        n388) );
  AO222X1 U625 ( .A(n321), .B(n342), .C(n323), .D(n343), .E(r_dac1v[8]), .F(
        n11), .Y(o_dac1[8]) );
  NAND4X1 U626 ( .A(n348), .B(n349), .C(n350), .D(n351), .Y(n342) );
  NAND4X1 U627 ( .A(n344), .B(n345), .C(n346), .D(n347), .Y(n343) );
  AOI22X1 U628 ( .A(r_dacvs[142]), .B(n53), .C(r_dacvs[14]), .D(n46), .Y(n348)
         );
  AO22X1 U629 ( .A(x_daclsb[0]), .B(n412), .C(r_dac1v[0]), .D(n10), .Y(
        o_dac1[0]) );
  AO22X1 U630 ( .A(x_daclsb[1]), .B(n412), .C(r_dac1v[1]), .D(n11), .Y(
        o_dac1[1]) );
  NAND2X1 U631 ( .A(cs_ptr[2]), .B(n533), .Y(n204) );
  INVX1 U632 ( .A(cs_ptr[2]), .Y(n534) );
  AOI221XL U633 ( .A(r_sar_en[0]), .B(n528), .C(r_sar_en[12]), .D(n527), .E(
        n440), .Y(n439) );
  ENOX1 U634 ( .A(n204), .B(n556), .C(n526), .D(r_sar_en[8]), .Y(n440) );
  AOI221XL U635 ( .A(r_sar_en[3]), .B(n528), .C(r_sar_en[15]), .D(n527), .E(
        n442), .Y(n437) );
  ENOX1 U636 ( .A(n204), .B(n554), .C(n526), .D(r_sar_en[11]), .Y(n442) );
  ENOX1 U637 ( .A(n218), .B(n539), .C(n559), .D(r_sar_en[5]), .Y(n441) );
  INVX1 U638 ( .A(r_sar_en[6]), .Y(n555) );
  AOI222XL U639 ( .A(r_dacvs[112]), .B(n47), .C(r_dacvs[96]), .D(n330), .E(
        r_dacvs[80]), .F(n43), .Y(n407) );
  AOI222XL U640 ( .A(r_dacvs[120]), .B(n47), .C(r_dacvs[104]), .D(n330), .E(
        r_dacvs[88]), .F(n43), .Y(n411) );
  AOI222XL U641 ( .A(r_dacvs[113]), .B(n72), .C(r_dacvs[97]), .D(n39), .E(
        r_dacvs[81]), .F(n71), .Y(n397) );
  AOI222XL U642 ( .A(r_dacvs[121]), .B(n72), .C(r_dacvs[105]), .D(n39), .E(
        r_dacvs[89]), .F(n71), .Y(n401) );
  AOI222XL U643 ( .A(r_dacvs[114]), .B(n72), .C(r_dacvs[98]), .D(n330), .E(
        r_dacvs[82]), .F(n71), .Y(n387) );
  AOI222XL U644 ( .A(r_dacvs[122]), .B(n72), .C(r_dacvs[106]), .D(n330), .E(
        r_dacvs[90]), .F(n71), .Y(n391) );
  AOI222XL U645 ( .A(r_dacvs[115]), .B(n47), .C(r_dacvs[99]), .D(n330), .E(
        r_dacvs[83]), .F(n43), .Y(n377) );
  AOI222XL U646 ( .A(r_dacvs[123]), .B(n47), .C(r_dacvs[107]), .D(n330), .E(
        r_dacvs[91]), .F(n43), .Y(n381) );
  AOI222XL U647 ( .A(r_dacvs[116]), .B(n72), .C(r_dacvs[100]), .D(n39), .E(
        r_dacvs[84]), .F(n71), .Y(n367) );
  AOI222XL U648 ( .A(r_dacvs[124]), .B(n72), .C(r_dacvs[108]), .D(n39), .E(
        r_dacvs[92]), .F(n71), .Y(n371) );
  AOI222XL U649 ( .A(r_dacvs[117]), .B(n47), .C(r_dacvs[101]), .D(n330), .E(
        r_dacvs[85]), .F(n43), .Y(n357) );
  AOI222XL U650 ( .A(r_dacvs[125]), .B(n47), .C(r_dacvs[109]), .D(n330), .E(
        r_dacvs[93]), .F(n43), .Y(n361) );
  AOI222XL U651 ( .A(r_dacvs[118]), .B(n47), .C(r_dacvs[102]), .D(n39), .E(
        r_dacvs[86]), .F(n43), .Y(n347) );
  AOI222XL U652 ( .A(r_dacvs[126]), .B(n47), .C(r_dacvs[110]), .D(n39), .E(
        r_dacvs[94]), .F(n43), .Y(n351) );
  AOI222XL U653 ( .A(r_dacvs[119]), .B(n72), .C(r_dacvs[103]), .D(n39), .E(
        r_dacvs[87]), .F(n71), .Y(n328) );
  AOI222XL U654 ( .A(r_dacvs[127]), .B(n72), .C(r_dacvs[111]), .D(n39), .E(
        r_dacvs[95]), .F(n71), .Y(n341) );
  AOI22X1 U655 ( .A(r_dacvs[16]), .B(n56), .C(r_dacvs[64]), .D(n333), .Y(n406)
         );
  AOI22X1 U656 ( .A(r_dacvs[24]), .B(n56), .C(r_dacvs[72]), .D(n333), .Y(n410)
         );
  AOI22X1 U657 ( .A(r_dacvs[17]), .B(n73), .C(r_dacvs[65]), .D(n61), .Y(n396)
         );
  AOI22X1 U658 ( .A(r_dacvs[25]), .B(n73), .C(r_dacvs[73]), .D(n61), .Y(n400)
         );
  AOI22X1 U659 ( .A(r_dacvs[18]), .B(n73), .C(r_dacvs[66]), .D(n333), .Y(n386)
         );
  AOI22X1 U660 ( .A(r_dacvs[26]), .B(n73), .C(r_dacvs[74]), .D(n333), .Y(n390)
         );
  AOI22X1 U661 ( .A(r_dacvs[19]), .B(n56), .C(r_dacvs[67]), .D(n333), .Y(n376)
         );
  AOI22X1 U662 ( .A(r_dacvs[20]), .B(n73), .C(r_dacvs[68]), .D(n61), .Y(n366)
         );
  AOI22X1 U663 ( .A(r_dacvs[28]), .B(n56), .C(r_dacvs[76]), .D(n333), .Y(n370)
         );
  AOI22X1 U664 ( .A(r_dacvs[21]), .B(n56), .C(r_dacvs[69]), .D(n333), .Y(n356)
         );
  AOI22X1 U665 ( .A(r_dacvs[29]), .B(n56), .C(r_dacvs[77]), .D(n333), .Y(n360)
         );
  AOI22X1 U666 ( .A(r_dacvs[22]), .B(n56), .C(r_dacvs[70]), .D(n61), .Y(n346)
         );
  AOI22X1 U667 ( .A(r_dacvs[30]), .B(n56), .C(r_dacvs[78]), .D(n61), .Y(n350)
         );
  AOI22X1 U668 ( .A(r_dacvs[23]), .B(n73), .C(r_dacvs[71]), .D(n61), .Y(n327)
         );
  AOI22X1 U669 ( .A(r_dacvs[31]), .B(n73), .C(r_dacvs[79]), .D(n61), .Y(n340)
         );
  AOI22X1 U670 ( .A(r_dacvs[48]), .B(n62), .C(r_dacvs[32]), .D(n335), .Y(n405)
         );
  AOI22X1 U671 ( .A(r_dacvs[56]), .B(n62), .C(r_dacvs[40]), .D(n52), .Y(n409)
         );
  AOI22X1 U672 ( .A(r_dacvs[49]), .B(n74), .C(r_dacvs[33]), .D(n335), .Y(n395)
         );
  AOI22X1 U673 ( .A(r_dacvs[57]), .B(n74), .C(r_dacvs[41]), .D(n52), .Y(n399)
         );
  AOI22X1 U674 ( .A(r_dacvs[50]), .B(n74), .C(r_dacvs[34]), .D(n335), .Y(n385)
         );
  AOI22X1 U675 ( .A(r_dacvs[58]), .B(n74), .C(r_dacvs[42]), .D(n335), .Y(n389)
         );
  AOI22X1 U676 ( .A(r_dacvs[51]), .B(n62), .C(r_dacvs[35]), .D(n335), .Y(n375)
         );
  AOI22X1 U677 ( .A(r_dacvs[52]), .B(n74), .C(r_dacvs[36]), .D(n335), .Y(n365)
         );
  AOI22X1 U678 ( .A(r_dacvs[60]), .B(n62), .C(r_dacvs[44]), .D(n52), .Y(n369)
         );
  AOI22X1 U679 ( .A(r_dacvs[53]), .B(n62), .C(r_dacvs[37]), .D(n335), .Y(n355)
         );
  AOI22X1 U680 ( .A(r_dacvs[61]), .B(n62), .C(r_dacvs[45]), .D(n52), .Y(n359)
         );
  AOI22X1 U681 ( .A(r_dacvs[54]), .B(n62), .C(r_dacvs[38]), .D(n335), .Y(n345)
         );
  AOI22X1 U682 ( .A(r_dacvs[62]), .B(n62), .C(r_dacvs[46]), .D(n52), .Y(n349)
         );
  AOI22X1 U683 ( .A(r_dacvs[55]), .B(n74), .C(r_dacvs[39]), .D(n335), .Y(n326)
         );
  AOI22X1 U684 ( .A(r_dacvs[63]), .B(n74), .C(r_dacvs[47]), .D(n52), .Y(n339)
         );
  AOI22X1 U685 ( .A(r_dacvs[128]), .B(n336), .C(r_dacvs[0]), .D(n337), .Y(n404) );
  AOI22X1 U686 ( .A(r_dacvs[129]), .B(n336), .C(r_dacvs[1]), .D(n337), .Y(n394) );
  AOI22X1 U687 ( .A(r_dacvs[130]), .B(n336), .C(r_dacvs[2]), .D(n337), .Y(n384) );
  AOI22X1 U688 ( .A(r_dacvs[131]), .B(n336), .C(r_dacvs[3]), .D(n337), .Y(n374) );
  AOI22X1 U689 ( .A(r_dacvs[132]), .B(n336), .C(r_dacvs[4]), .D(n337), .Y(n364) );
  AOI22X1 U690 ( .A(r_dacvs[133]), .B(n336), .C(r_dacvs[5]), .D(n337), .Y(n354) );
  AOI22X1 U691 ( .A(r_dacvs[134]), .B(n336), .C(r_dacvs[6]), .D(n337), .Y(n344) );
  AOI22X1 U692 ( .A(r_dacvs[135]), .B(n336), .C(r_dacvs[7]), .D(n337), .Y(n325) );
  INVX1 U693 ( .A(r_sar_en[9]), .Y(n539) );
  INVX1 U694 ( .A(r_sar_en[10]), .Y(n540) );
  INVX1 U695 ( .A(r_sar_en[7]), .Y(n554) );
  INVX1 U696 ( .A(r_sar_en[4]), .Y(n556) );
  AOI22X1 U697 ( .A(r_dacvs[27]), .B(n73), .C(r_dacvs[75]), .D(n61), .Y(n380)
         );
  AOI22X1 U698 ( .A(r_dacvs[59]), .B(n74), .C(r_dacvs[43]), .D(n52), .Y(n379)
         );
  INVX1 U699 ( .A(r_sar_en[17]), .Y(n535) );
  INVX1 U700 ( .A(r_sar_en[16]), .Y(n536) );
  BUFX3 U701 ( .A(r_comp_opt[0]), .Y(n97) );
  BUFX3 U702 ( .A(r_comp_opt[0]), .Y(n98) );
  NAND42X1 U703 ( .C(r_dac_en[3]), .D(n124), .A(n123), .B(n122), .Y(n207) );
  NAND21X1 U704 ( .B(r_dac_en[1]), .A(n116), .Y(n124) );
  NOR43XL U705 ( .B(n121), .C(n120), .D(n119), .A(n118), .Y(n122) );
  NOR32XL U706 ( .B(n532), .C(n78), .A(n117), .Y(n123) );
  INVX1 U707 ( .A(r_dac_en[7]), .Y(n557) );
  NAND21X1 U708 ( .B(r_dac_en[0]), .A(n2), .Y(n117) );
  INVX1 U709 ( .A(r_dac_en[15]), .Y(n543) );
  INVX1 U710 ( .A(r_dac_en[17]), .Y(n538) );
  INVX1 U711 ( .A(r_dac_en[8]), .Y(n541) );
  INVX1 U712 ( .A(r_dac_en[9]), .Y(n542) );
  INVX1 U713 ( .A(r_dac_en[16]), .Y(n537) );
  OR4X1 U714 ( .A(r_dac_en[4]), .B(r_dac_en[5]), .C(r_dac_en[11]), .D(
        r_dac_en[10]), .Y(n118) );
  INVX1 U715 ( .A(r_dac_en[6]), .Y(n532) );
  INVX1 U716 ( .A(r_dac_en[2]), .Y(n116) );
  INVX1 U717 ( .A(r_dac_en[12]), .Y(n120) );
  INVX1 U718 ( .A(r_dac_en[14]), .Y(n119) );
  INVX1 U719 ( .A(r_dac_en[13]), .Y(n121) );
  XNOR2XL U720 ( .A(n103), .B(x_daclsb[4]), .Y(n417) );
  NAND4X1 U721 ( .A(o_dactl[6]), .B(n531), .C(n414), .D(n415), .Y(n138) );
  NOR2X1 U722 ( .A(n416), .B(n417), .Y(n415) );
  XNOR2XL U723 ( .A(x_daclsb[3]), .B(n99), .Y(n414) );
  XNOR2XL U724 ( .A(n534), .B(x_daclsb[5]), .Y(n416) );
  NOR42XL U725 ( .C(n196), .D(o_dactl[1]), .A(n558), .B(n140), .Y(n194) );
  XNOR2XL U726 ( .A(syn_comp[1]), .B(n197), .Y(n196) );
  AOI221XL U727 ( .A(n530), .B(n198), .C(n529), .D(n199), .E(n200), .Y(n197)
         );
  OAI22X1 U728 ( .A(n203), .B(n561), .C(n204), .D(n560), .Y(n198) );
  OAI22X1 U729 ( .A(n201), .B(n159), .C(n202), .D(n161), .Y(n200) );
  AOI22X1 U730 ( .A(o_dat[7]), .B(n559), .C(o_dat[3]), .D(n528), .Y(n201) );
  AOI22X1 U731 ( .A(o_dat[6]), .B(n559), .C(o_dat[2]), .D(n528), .Y(n202) );
  INVX1 U732 ( .A(r_sar_en[15]), .Y(n130) );
  AO22X1 U733 ( .A(n528), .B(o_dat[0]), .C(n559), .D(o_dat[4]), .Y(n199) );
  OAI222XL U734 ( .A(n209), .B(n538), .C(n210), .D(n537), .E(cs_ptr[4]), .F(
        n211), .Y(n141) );
  OA2222XL U735 ( .A(n212), .B(n161), .C(n213), .D(n159), .E(n214), .F(n162), 
        .G(n215), .H(n193), .Y(n211) );
  AOI221XL U736 ( .A(r_dac_en[2]), .B(n42), .C(r_dac_en[14]), .D(n527), .E(
        n221), .Y(n212) );
  AOI221XL U737 ( .A(r_dac_en[1]), .B(n528), .C(r_dac_en[13]), .D(n527), .E(
        n219), .Y(n214) );
  AOI221XL U738 ( .A(r_dac_en[0]), .B(n42), .C(r_dac_en[12]), .D(n527), .E(
        n217), .Y(n215) );
  ENOX1 U739 ( .A(n218), .B(n541), .C(n559), .D(r_dac_en[4]), .Y(n217) );
  AOI221XL U740 ( .A(r_dac_en[3]), .B(n528), .C(r_dac_en[15]), .D(n527), .E(
        n220), .Y(n213) );
  ENOX1 U741 ( .A(n204), .B(n557), .C(n526), .D(r_dac_en[11]), .Y(n220) );
  ENOX1 U742 ( .A(n218), .B(n542), .C(n559), .D(r_dac_en[5]), .Y(n219) );
  INVX1 U743 ( .A(o_dat[5]), .Y(n560) );
  INVX1 U744 ( .A(o_dat[1]), .Y(n561) );
  ENOX1 U745 ( .A(n204), .B(n532), .C(n526), .D(r_dac_en[10]), .Y(n221) );
  OAI21X1 U746 ( .B(n143), .C(n444), .A(n445), .Y(datcmp[9]) );
  OAI21X1 U747 ( .B(n162), .C(n143), .A(o_dat[9]), .Y(n445) );
  OAI21X1 U748 ( .B(n156), .C(n444), .A(n451), .Y(datcmp[13]) );
  OAI21X1 U749 ( .B(n162), .C(n156), .A(o_dat[13]), .Y(n451) );
  ENOX1 U750 ( .A(n152), .B(n105), .C(o_dat[17]), .D(n152), .Y(datcmp[17]) );
  NAND2X1 U751 ( .A(syn_comp[1]), .B(n530), .Y(n444) );
  OAI21X1 U752 ( .B(n151), .C(n446), .A(n453), .Y(datcmp[0]) );
  OAI21X1 U753 ( .B(n193), .C(n151), .A(o_dat[0]), .Y(n453) );
  OAI21X1 U754 ( .B(n148), .C(n446), .A(n449), .Y(datcmp[4]) );
  OAI21X1 U755 ( .B(n193), .C(n148), .A(o_dat[4]), .Y(n449) );
  OAI21X1 U756 ( .B(n143), .C(n446), .A(n447), .Y(datcmp[8]) );
  OAI21X1 U757 ( .B(n193), .C(n143), .A(o_dat[8]), .Y(n447) );
  OAI21X1 U758 ( .B(n156), .C(n446), .A(n452), .Y(datcmp[12]) );
  OAI21X1 U759 ( .B(n193), .C(n156), .A(o_dat[12]), .Y(n452) );
  ENOX1 U760 ( .A(n154), .B(n105), .C(o_dat[15]), .D(n154), .Y(datcmp[15]) );
  ENOX1 U761 ( .A(n149), .B(n105), .C(n149), .D(o_dat[3]), .Y(datcmp[3]) );
  ENOX1 U762 ( .A(n146), .B(n105), .C(n146), .D(o_dat[7]), .Y(datcmp[7]) );
  ENOX1 U763 ( .A(n150), .B(n105), .C(n150), .D(o_dat[2]), .Y(datcmp[2]) );
  ENOX1 U764 ( .A(n147), .B(n105), .C(n147), .D(o_dat[6]), .Y(datcmp[6]) );
  ENOX1 U765 ( .A(n153), .B(n105), .C(o_dat[16]), .D(n153), .Y(datcmp[16]) );
  ENOX1 U766 ( .A(n158), .B(n105), .C(o_dat[10]), .D(n158), .Y(datcmp[10]) );
  ENOX1 U767 ( .A(n155), .B(n105), .C(o_dat[14]), .D(n155), .Y(datcmp[14]) );
  ENOX1 U768 ( .A(n157), .B(n105), .C(o_dat[11]), .D(n157), .Y(datcmp[11]) );
  NAND2X1 U769 ( .A(syn_comp[1]), .B(n529), .Y(n446) );
  INVX1 U770 ( .A(syn_comp[1]), .Y(n105) );
  AO222X1 U771 ( .A(n321), .B(n372), .C(n323), .D(n373), .E(r_dac1v[5]), .F(
        n11), .Y(o_dac1[5]) );
  INVXL U772 ( .A(dacv_wr[11]), .Y(n286) );
  AND2XL U773 ( .A(ps_ptr[4]), .B(r_sar_en[16]), .Y(n249) );
  AND2XL U774 ( .A(ps_ptr[4]), .B(r_dac_en[17]), .Y(n259) );
  AND2XL U775 ( .A(ps_ptr[4]), .B(r_dac_en[16]), .Y(n253) );
  AND2XL U776 ( .A(ps_ptr[4]), .B(r_sar_en[17]), .Y(n268) );
  NAND21X1 U777 ( .B(ps_ptr[4]), .A(n262), .Y(n243) );
  NAND32X1 U778 ( .B(pos_dacis[2]), .C(n299), .A(n298), .Y(n464) );
  INVXL U779 ( .A(n299), .Y(n303) );
  XOR2X1 U780 ( .A(n295), .B(pos_dacis[1]), .Y(n299) );
  INVX1 U781 ( .A(dacv_wr[10]), .Y(n287) );
  AND4X1 U782 ( .A(n471), .B(n479), .C(n496), .D(n489), .Y(n472) );
  AO21XL U783 ( .B(n478), .C(n460), .A(n467), .Y(n473) );
  OAI211X1 U784 ( .C(n332), .D(n466), .A(n331), .B(n430), .Y(n418) );
  MUX2XL U785 ( .D0(r_rpt_v[0]), .D1(n50), .S(r_wr[3]), .Y(wdlsb[0]) );
  AND2XL U786 ( .A(r_wr[4]), .B(n51), .Y(clrsta[0]) );
  INVXL U787 ( .A(n51), .Y(n225) );
  NAND6XL U788 ( .A(r_wdat[6]), .B(n51), .C(n226), .D(n3), .E(n223), .F(n7), 
        .Y(n224) );
  MUX2IX4 U789 ( .D0(n272), .D1(n271), .S(ps_ptr[0]), .Y(n273) );
  INVX3 U790 ( .A(n240), .Y(n263) );
  INVXL U791 ( .A(n314), .Y(n315) );
  INVXL U792 ( .A(n491), .Y(n492) );
  AND2X1 U793 ( .A(n491), .B(n484), .Y(n485) );
  NAND21X1 U794 ( .B(n76), .A(pos_dacis[17]), .Y(n491) );
  NAND32XL U795 ( .B(pos_dacis[12]), .C(n462), .A(n461), .Y(n496) );
  NAND21X1 U796 ( .B(n418), .A(n462), .Y(n419) );
  NAND32X1 U797 ( .B(n427), .C(n334), .A(n462), .Y(n413) );
  INVXL U798 ( .A(n95), .Y(n236) );
  INVX2 U799 ( .A(n243), .Y(n260) );
  AO2222X1 U800 ( .A(n264), .B(r_sar_en[12]), .C(n263), .D(r_sar_en[14]), .E(
        n262), .F(r_sar_en[8]), .G(n261), .H(r_sar_en[10]), .Y(n246) );
  AO2222X1 U801 ( .A(n264), .B(r_sar_en[13]), .C(n263), .D(r_sar_en[15]), .E(
        n262), .F(r_sar_en[9]), .G(n261), .H(r_sar_en[11]), .Y(n265) );
  NAND2X2 U802 ( .A(n270), .B(n269), .Y(n271) );
  NAND2X2 U803 ( .A(n255), .B(n254), .Y(n272) );
  AO2222X1 U804 ( .A(n263), .B(r_sar_en[7]), .C(n260), .D(r_sar_en[1]), .E(
        n261), .F(r_sar_en[3]), .G(n264), .H(r_sar_en[5]), .Y(n266) );
  AO2222X1 U805 ( .A(n263), .B(r_dac_en[6]), .C(r_dac_en[0]), .D(n260), .E(
        r_dac_en[2]), .F(n261), .G(r_dac_en[4]), .H(n264), .Y(n251) );
  AO2222X1 U806 ( .A(n263), .B(r_dac_en[7]), .C(r_dac_en[1]), .D(n260), .E(
        r_dac_en[3]), .F(n261), .G(r_dac_en[5]), .H(n264), .Y(n257) );
endmodule


module dacmux_a0_DW01_add_17 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_16 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_15 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_14 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_13 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_12 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_11 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_10 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_9 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_6 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_5 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module glreg_WIDTH2_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n4, n5;

  SDFFRQX1 mem_reg_0_ ( .D(n5), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(n4), .SIN(rdat[0]), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[1]) );
  MUX2XL U2 ( .D0(rdat[1]), .D1(wdat[1]), .S(we), .Y(n4) );
  MUX2XL U3 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n5) );
endmodule


module glreg_WIDTH2_1 ( clk, arstz, we, wdat, rdat, test_si, test_so, test_se
 );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  output test_so;
  wire   n8, n9;

  SDFFRQX1 mem_reg_0_ ( .D(n9), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(n8), .SIN(rdat[0]), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[1]) );
  MUX2XL U2 ( .D0(rdat[1]), .D1(wdat[1]), .S(we), .Y(n8) );
  BUFX3 U3 ( .A(rdat[1]), .Y(test_so) );
  MUX2XL U4 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n9) );
endmodule


module glreg_a0_26 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9734;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_26 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9734), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9734), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9734), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9734), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9734), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9734), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9734), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9734), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9734), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_27 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9752;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_27 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9752), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9752), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9752), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9752), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9752), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9752), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9752), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9752), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9752), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_28 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9770;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_28 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9770), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9770), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9770), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9770), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9770), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9770), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9770), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9770), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9770), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_29 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9788;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_29 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9788), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9788), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9788), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9788), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9788), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9788), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9788), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9788), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9788), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_1 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21;
  wire   [7:0] wd_r;

  glreg_WIDTH8_1 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[5]), .Y(n16) );
  INVX1 U3 ( .A(set2[1]), .Y(n20) );
  NAND21X1 U4 ( .B(set2[5]), .A(n15), .Y(n1) );
  INVX1 U5 ( .A(set2[6]), .Y(n15) );
  INVX1 U6 ( .A(set2[0]), .Y(n21) );
  INVX1 U7 ( .A(set2[2]), .Y(n19) );
  INVX1 U8 ( .A(set2[7]), .Y(n14) );
  INVX1 U9 ( .A(set2[3]), .Y(n18) );
  INVX1 U10 ( .A(set2[4]), .Y(n17) );
  NAND42X1 U11 ( .C(n5), .D(n4), .A(n3), .B(n2), .Y(upd_r) );
  NOR43XL U12 ( .B(n14), .C(n18), .D(n17), .A(n1), .Y(n2) );
  NAND21X1 U13 ( .B(set2[1]), .A(n19), .Y(n4) );
  NAND21X1 U14 ( .B(clr1[0]), .A(n21), .Y(n5) );
  NOR8XL U15 ( .A(clr1[4]), .B(clr1[5]), .C(clr1[6]), .D(clr1[7]), .E(rst0), 
        .F(clr1[1]), .G(clr1[2]), .H(clr1[3]), .Y(n3) );
  AOI211X1 U16 ( .C(n17), .D(n9), .A(clr1[4]), .B(rst0), .Y(wd_r[4]) );
  INVX1 U17 ( .A(rdat[4]), .Y(n9) );
  AOI211X1 U18 ( .C(n19), .D(n11), .A(clr1[2]), .B(rst0), .Y(wd_r[2]) );
  INVX1 U19 ( .A(rdat[2]), .Y(n11) );
  AOI211X1 U20 ( .C(n16), .D(n8), .A(clr1[5]), .B(rst0), .Y(wd_r[5]) );
  INVX1 U21 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U22 ( .C(n21), .D(n13), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U23 ( .A(rdat[0]), .Y(n13) );
  AOI211X1 U24 ( .C(n20), .D(n12), .A(clr1[1]), .B(rst0), .Y(wd_r[1]) );
  INVX1 U25 ( .A(rdat[1]), .Y(n12) );
  AOI211X1 U26 ( .C(n18), .D(n10), .A(clr1[3]), .B(rst0), .Y(wd_r[3]) );
  INVX1 U27 ( .A(rdat[3]), .Y(n10) );
  AOI211X1 U28 ( .C(n15), .D(n7), .A(clr1[6]), .B(rst0), .Y(wd_r[6]) );
  INVX1 U29 ( .A(rdat[6]), .Y(n7) );
  AOI211X1 U30 ( .C(n14), .D(n6), .A(clr1[7]), .B(rst0), .Y(wd_r[7]) );
  INVX1 U31 ( .A(rdat[7]), .Y(n6) );
  NOR2X1 U32 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
  NOR2X1 U33 ( .A(rdat[1]), .B(n20), .Y(irq[1]) );
  NOR2X1 U34 ( .A(rdat[0]), .B(n21), .Y(irq[0]) );
  NOR2X1 U35 ( .A(rdat[4]), .B(n17), .Y(irq[4]) );
  NOR2X1 U36 ( .A(rdat[6]), .B(n15), .Y(irq[6]) );
  NOR2X1 U37 ( .A(rdat[2]), .B(n19), .Y(irq[2]) );
  NOR2X1 U38 ( .A(rdat[7]), .B(n14), .Y(irq[7]) );
  NOR2X1 U39 ( .A(rdat[3]), .B(n18), .Y(irq[3]) );
endmodule


module glreg_WIDTH8_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9806;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9806), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9806), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9806), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9806), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9806), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9806), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9806), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9806), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9806), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_30 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9824;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_30 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9824), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9824), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9824), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9824), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9824), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9824), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9824), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9824), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9824), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_31 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9842;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_31 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9842), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9842), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9842), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9842), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9842), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9842), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9842), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9842), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9842), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_32 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9860;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_32 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9860), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9860), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9860), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9860), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9860), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9860), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9860), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9860), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9860), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_33 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9878;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_33 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9878), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9878), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9878), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9878), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9878), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9878), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9878), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9878), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9878), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_34 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9896;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_34 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9896), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9896), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9896), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9896), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9896), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9896), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9896), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9896), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9896), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_35 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9914;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_35 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9914), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9914), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9914), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9914), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9914), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9914), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9914), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9914), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9914), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_36 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9932;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_36 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9932), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9932), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9932), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9932), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9932), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9932), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9932), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9932), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9932), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_37 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9950;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_37 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9950), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9950), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9950), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9950), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9950), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9950), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9950), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9950), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9950), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_38 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9968;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_38 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9968), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9968), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9968), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9968), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9968), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9968), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9968), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9968), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9968), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_39 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9986;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_39 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9986), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9986), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9986), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9986), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9986), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9986), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9986), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9986), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9986), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_40 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10004;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_40 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10004), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10004), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10004), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10004), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10004), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10004), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10004), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10004), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10004), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_41 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10022;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_41 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10022), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10022), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10022), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10022), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10022), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10022), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10022), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10022), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10022), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_42 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10040;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_42 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10040), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10040), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10040), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10040), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10040), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10040), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10040), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10040), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10040), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_43 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10058;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_43 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10058), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10058), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10058), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10058), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10058), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10058), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10058), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10058), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10058), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_44 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10076;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_44 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10076), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10076), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10076), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10076), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10076), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10076), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10076), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10076), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10076), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_45 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10094;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_45 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10094), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10094), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10094), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10094), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10094), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10094), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10094), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10094), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10094), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_46 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10112;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_46 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10112), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10112), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10112), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10112), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10112), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10112), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10112), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10112), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10112), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_47 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10130;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_47 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10130), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10130), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10130), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10130), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10130), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10130), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10130), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10130), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10130), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10148;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10148), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10148), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10148), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10148), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10148), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10148), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10148), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_48 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10166;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_48 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10166), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10166), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10166), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10166), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10166), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10166), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10166), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10166), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10166), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_49 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10184;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_49 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10184), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10184), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10184), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10184), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10184), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10184), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10184), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10184), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10184), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH7_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10202;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10202), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10202), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10202), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10202), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10202), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10202), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10202), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10202), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module shmux_00000005_00000012_00000012 ( ps_md4ch, r_comp_swtch, r_semi, 
        r_loop, r_dac_en, wr_dacv, busy, sh_hold, stop, semi_start, auto_start, 
        mxcyc_done, sampl_begn, sampl_done, app_dacis, pos_dacis, cs_ptr, 
        ps_ptr, clk, srstz, test_si2, test_si1, test_so1, test_se );
  input [17:0] r_dac_en;
  input [17:0] wr_dacv;
  output [17:0] app_dacis;
  output [17:0] pos_dacis;
  output [4:0] cs_ptr;
  output [4:0] ps_ptr;
  input ps_md4ch, r_comp_swtch, r_semi, r_loop, stop, semi_start, auto_start,
         mxcyc_done, sampl_begn, sampl_done, clk, srstz, test_si2, test_si1,
         test_se;
  output busy, sh_hold, test_so1;
  wire   n772, cs_mux_5_, neg_dacis_16_, neg_dacis_15_, neg_dacis_14_,
         neg_dacis_13_, neg_dacis_12_, neg_dacis_11_, neg_dacis_10_,
         neg_dacis_9_, neg_dacis_8_, neg_dacis_7_, neg_dacis_6_, neg_dacis_5_,
         neg_dacis_4_, neg_dacis_3_, neg_dacis_2_, neg_dacis_1_, neg_dacis_0_,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N971, N972, N973,
         N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984,
         N985, N986, N987, N988, N989, N994, N995, N996, N997, N998, N999,
         N1139, N1148, N1230, N1312, N1394, net10220, net10238, net10243, n671,
         sub_398_S2_I5_aco_carry_4_, sub_398_S2_I4_aco_carry_4_, n62, n63, n64,
         n771, n770, n769, n768, n209, n212, n213, n214, n216, n231, n232,
         n233, n234, n242, n243, n244, n264, n265, n266, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n299, n302,
         n303, n324, n326, n328, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n391, n392, n395, n398, n399, n400, n401,
         n402, n403, n404, n408, n409, n410, n411, n412, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n425, n426, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n439, n441, n444, n445, n446,
         n449, n450, n454, n455, n456, n457, n460, n462, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n479, n482, n483, n484, n485, n486, n487, n488, n489, n490, n492,
         n496, n497, n500, n501, n508, n509, n510, n511, n512, n515, n516,
         n517, n518, n519, n523, n524, n526, n527, n528, n530, n531, n532,
         n533, n534, n535, n536, n540, n541, n542, n546, n547, n548, n549,
         n550, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n579, n582, n583, n584, n585, n587, n588, n589, n590, n591,
         n592, n593, n594, n596, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n43, n44,
         n45, n46, n48, n49, n50, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n210, n211, n215, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n235, n236, n237, n238, n239, n240, n241, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n267, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n300, n301, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n325, n327, n329, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n371, n372, n373, n374, n375, n387, n388, n389, n390,
         n393, n394, n396, n397, n405, n406, n407, n413, n423, n424, n427,
         n437, n438, n440, n442, n443, n447, n448, n451, n452, n453, n458,
         n459, n461, n463, n478, n480, n481, n491, n493, n494, n495, n498,
         n499, n502, n503, n504, n505, n506, n507, n513, n514, n520, n521,
         n522, n525, n529, n537, n538, n539, n543, n544, n545, n551, n564,
         n565, n566, n577, n578, n580, n581, n586, n595, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767;
  wire   [5:4] sub_398_S2_I7_aco_carry;
  wire   [5:4] sub_398_S2_I3_aco_carry;
  wire   [5:4] sub_398_S2_aco_carry;

  FAD1X1 sub_398_S2_I7_aco_U2_4 ( .A(n750), .B(n63), .CI(
        sub_398_S2_I7_aco_carry[4]), .CO(sub_398_S2_I7_aco_carry[5]), .SO(
        N1394) );
  FAD1X1 sub_398_S2_I3_aco_U2_4 ( .A(n764), .B(n64), .CI(
        sub_398_S2_I3_aco_carry[4]), .CO(sub_398_S2_I3_aco_carry[5]), .SO(
        N1230) );
  FAD1X1 sub_398_S2_aco_U2_4 ( .A(N1139), .B(n62), .CI(sub_398_S2_aco_carry[4]), .CO(sub_398_S2_aco_carry[5]), .SO(N1148) );
  SNPS_CLOCK_GATE_LOW_shmux_00000005_00000012_00000012 clk_gate_neg_dacis_reg ( 
        .CLK(clk), .EN(N949), .ENCLK(net10220), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 clk_gate_r_dacis_reg ( 
        .CLK(clk), .EN(N971), .ENCLK(net10238), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 clk_gate_cs_mux_reg ( 
        .CLK(clk), .EN(N994), .ENCLK(net10243), .TE(test_se) );
  SDFFQX1 cs_mux_reg_4_ ( .D(N999), .SIN(n769), .SMC(test_se), .C(net10243), 
        .Q(n768) );
  SDFFQX1 cs_mux_reg_1_ ( .D(N996), .SIN(n44), .SMC(test_se), .C(net10243), 
        .Q(n770) );
  SDFFQX1 cs_mux_reg_0_ ( .D(N995), .SIN(test_si2), .SMC(test_se), .C(net10243), .Q(n771) );
  SDFFQX1 cs_mux_reg_3_ ( .D(N998), .SIN(n7), .SMC(test_se), .C(net10243), .Q(
        n769) );
  SDFFQX1 cs_mux_reg_2_ ( .D(N997), .SIN(n48), .SMC(test_se), .C(net10243), 
        .Q(cs_ptr[2]) );
  SDFFQX1 r_dacis_reg_17_ ( .D(N989), .SIN(pos_dacis[16]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[17]) );
  SDFFQX1 r_dacis_reg_16_ ( .D(N988), .SIN(pos_dacis[15]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[16]) );
  SDFFQX1 r_dacis_reg_15_ ( .D(N987), .SIN(pos_dacis[14]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[15]) );
  SDFFQX1 r_dacis_reg_14_ ( .D(N986), .SIN(pos_dacis[13]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[14]) );
  SDFFQX1 r_dacis_reg_13_ ( .D(N985), .SIN(pos_dacis[12]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[13]) );
  SDFFQX1 r_dacis_reg_12_ ( .D(N984), .SIN(pos_dacis[11]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[12]) );
  SDFFQX1 r_dacis_reg_9_ ( .D(N981), .SIN(pos_dacis[8]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[9]) );
  SDFFQX1 r_dacis_reg_10_ ( .D(N982), .SIN(pos_dacis[9]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[10]) );
  SDFFQX1 r_dacis_reg_8_ ( .D(N980), .SIN(pos_dacis[7]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[8]) );
  SDFFQX1 r_dacis_reg_11_ ( .D(N983), .SIN(pos_dacis[10]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[11]) );
  SDFFQX1 r_dacis_reg_7_ ( .D(N979), .SIN(pos_dacis[6]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[7]) );
  SDFFNQX1 neg_dacis_reg_16_ ( .D(N966), .SIN(neg_dacis_15_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_16_) );
  SDFFNQX1 neg_dacis_reg_15_ ( .D(N965), .SIN(neg_dacis_14_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_15_) );
  SDFFNQX1 neg_dacis_reg_14_ ( .D(N964), .SIN(neg_dacis_13_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_14_) );
  SDFFNQX1 neg_dacis_reg_11_ ( .D(N961), .SIN(neg_dacis_10_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_11_) );
  SDFFNQX1 neg_dacis_reg_10_ ( .D(N960), .SIN(neg_dacis_9_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_10_) );
  SDFFNQX1 neg_dacis_reg_9_ ( .D(N959), .SIN(neg_dacis_8_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_9_) );
  SDFFNQX1 neg_dacis_reg_8_ ( .D(N958), .SIN(neg_dacis_7_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_8_) );
  SDFFNQX1 neg_dacis_reg_7_ ( .D(N957), .SIN(neg_dacis_6_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_7_) );
  SDFFNQX1 neg_dacis_reg_4_ ( .D(N954), .SIN(neg_dacis_3_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_4_) );
  SDFFNQX1 neg_dacis_reg_3_ ( .D(N953), .SIN(neg_dacis_2_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_3_) );
  SDFFNQX1 neg_dacis_reg_2_ ( .D(N952), .SIN(neg_dacis_1_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_2_) );
  SDFFNQX1 neg_dacis_reg_0_ ( .D(N950), .SIN(test_si1), .SMC(test_se), .XC(
        net10220), .Q(neg_dacis_0_) );
  SDFFNQX1 neg_dacis_reg_6_ ( .D(N956), .SIN(neg_dacis_5_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_6_) );
  SDFFNQX1 neg_dacis_reg_1_ ( .D(N951), .SIN(neg_dacis_0_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_1_) );
  SDFFNQX1 neg_dacis_reg_17_ ( .D(N967), .SIN(neg_dacis_16_), .SMC(test_se), 
        .XC(net10220), .Q(test_so1) );
  SDFFNQX1 neg_dacis_reg_5_ ( .D(N955), .SIN(neg_dacis_4_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_5_) );
  SDFFNQX1 neg_dacis_reg_12_ ( .D(N962), .SIN(neg_dacis_11_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_12_) );
  SDFFNQX1 neg_dacis_reg_13_ ( .D(N963), .SIN(neg_dacis_12_), .SMC(test_se), 
        .XC(net10220), .Q(neg_dacis_13_) );
  SDFFQX1 r_dacis_reg_6_ ( .D(N978), .SIN(pos_dacis[5]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[6]) );
  SDFFQX1 r_dacis_reg_5_ ( .D(N977), .SIN(pos_dacis[4]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[5]) );
  SDFFQX1 r_dacis_reg_4_ ( .D(N976), .SIN(pos_dacis[3]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[4]) );
  SDFFQX1 r_dacis_reg_2_ ( .D(N974), .SIN(pos_dacis[1]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[2]) );
  SDFFQX1 cs_mux_reg_5_ ( .D(n671), .SIN(n53), .SMC(test_se), .C(clk), .Q(
        cs_mux_5_) );
  SDFFQX1 r_dacis_reg_0_ ( .D(N972), .SIN(cs_mux_5_), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[0]) );
  SDFFQX1 r_dacis_reg_3_ ( .D(N975), .SIN(pos_dacis[2]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[3]) );
  SDFFQX1 r_dacis_reg_1_ ( .D(N973), .SIN(pos_dacis[0]), .SMC(test_se), .C(
        net10238), .Q(pos_dacis[1]) );
  BUFX3 U3 ( .A(n772), .Y(ps_ptr[2]) );
  BUFX1 U4 ( .A(n606), .Y(n1) );
  INVX1 U5 ( .A(n125), .Y(n91) );
  GEN2XL U6 ( .D(n327), .E(n48), .C(n325), .B(n323), .A(n322), .Y(n342) );
  GEN2XL U7 ( .D(n544), .E(n543), .C(n539), .B(n538), .A(n537), .Y(n354) );
  OAI221X1 U8 ( .A(n320), .B(n504), .C(n10), .D(n505), .E(n319), .Y(n772) );
  NOR21XL U9 ( .B(n315), .A(n314), .Y(n317) );
  OAI221X1 U10 ( .A(n189), .B(n504), .C(n12), .D(n505), .E(n188), .Y(ps_ptr[3]) );
  OA222X1 U11 ( .A(n187), .B(n360), .C(n186), .D(n197), .E(n185), .F(n1), .Y(
        n188) );
  GEN3XL U12 ( .F(n286), .G(n285), .E(n284), .D(n283), .C(n282), .B(n507), .A(
        n281), .Y(ps_ptr[0]) );
  GEN2XL U13 ( .D(n253), .E(n252), .C(n251), .B(n250), .A(n249), .Y(n285) );
  AOI21X1 U14 ( .B(n478), .C(n768), .A(n463), .Y(n3) );
  OA21X1 U15 ( .B(n563), .C(n519), .A(n561), .Y(n4) );
  XNOR2XL U16 ( .A(n50), .B(n44), .Y(n678) );
  INVX1 U17 ( .A(n678), .Y(n5) );
  INVX1 U18 ( .A(n678), .Y(n6) );
  INVX1 U19 ( .A(n601), .Y(n7) );
  INVX1 U20 ( .A(n653), .Y(n8) );
  OR2XL U21 ( .A(n91), .B(n184), .Y(n504) );
  NAND5XL U22 ( .A(n344), .B(n132), .C(n329), .D(n131), .E(n543), .Y(n198) );
  INVXL U23 ( .A(n360), .Y(n564) );
  AND2XL U24 ( .A(n609), .B(ps_ptr[3]), .Y(N998) );
  AND2XL U25 ( .A(n609), .B(ps_ptr[1]), .Y(N996) );
  NAND32XL U26 ( .B(n345), .C(n316), .A(n315), .Y(n197) );
  INVXL U27 ( .A(n505), .Y(n577) );
  INVXL U28 ( .A(n504), .Y(n580) );
  AO21XL U29 ( .B(n564), .C(n551), .A(n545), .Y(n565) );
  MAJ3XL U30 ( .A(n48), .B(n586), .C(n581), .Y(n595) );
  NAND21XL U31 ( .B(n44), .A(ps_ptr[0]), .Y(n581) );
  AND2XL U32 ( .A(n609), .B(ps_ptr[0]), .Y(N995) );
  OAI222XL U33 ( .A(n466), .B(n467), .C(n468), .D(n751), .E(n445), .F(n753), 
        .Y(n369) );
  INVX2 U34 ( .A(n184), .Y(n39) );
  GEN3X1 U35 ( .F(n544), .G(n543), .E(n539), .D(n538), .C(n537), .B(n529), .A(
        n525), .Y(n545) );
  AND2XL U36 ( .A(n507), .B(n506), .Y(n529) );
  NAND21XL U37 ( .B(n769), .A(ps_ptr[3]), .Y(n503) );
  NAND21XL U38 ( .B(n325), .A(n323), .Y(n313) );
  INVXL U39 ( .A(n129), .Y(n253) );
  AOI211XL U40 ( .C(n327), .D(n769), .A(n313), .B(n198), .Y(n186) );
  NAND2X1 U41 ( .A(n9), .B(n611), .Y(n671) );
  MUX2IX1 U42 ( .D0(cs_mux_5_), .D1(n610), .S(n609), .Y(n9) );
  GEN2X1 U43 ( .D(n604), .E(n603), .C(r_loop), .B(n602), .A(cs_mux_5_), .Y(
        n605) );
  NOR3XL U44 ( .A(pos_dacis[1]), .B(pos_dacis[2]), .C(n623), .Y(n624) );
  INVX1 U45 ( .A(wr_dacv[2]), .Y(n254) );
  INVX1 U46 ( .A(n450), .Y(n747) );
  INVX1 U47 ( .A(n94), .Y(n104) );
  INVX1 U48 ( .A(n302), .Y(n296) );
  INVXL U49 ( .A(n1), .Y(n353) );
  INVX1 U50 ( .A(wr_dacv[9]), .Y(n543) );
  NOR2X1 U51 ( .A(n748), .B(n695), .Y(n454) );
  INVX1 U52 ( .A(n341), .Y(n705) );
  INVX1 U53 ( .A(n734), .Y(n706) );
  AOI21X1 U54 ( .B(n748), .C(n695), .A(n454), .Y(n450) );
  NAND21X1 U55 ( .B(n489), .A(n635), .Y(n302) );
  OAI22X1 U56 ( .A(n740), .B(n232), .C(n739), .D(n234), .Y(n326) );
  INVX1 U57 ( .A(n607), .Y(n513) );
  INVX1 U58 ( .A(n77), .Y(n141) );
  INVX1 U59 ( .A(n641), .Y(n401) );
  INVX1 U60 ( .A(n346), .Y(n262) );
  NOR2X1 U61 ( .A(n302), .B(n339), .Y(n485) );
  INVX1 U62 ( .A(n682), .Y(n746) );
  INVX1 U63 ( .A(n466), .Y(n751) );
  OAI22X1 U64 ( .A(n265), .B(n232), .C(n738), .D(n234), .Y(n264) );
  NAND21X1 U65 ( .B(n695), .A(n96), .Y(n94) );
  INVX1 U66 ( .A(n189), .Y(n81) );
  INVX1 U67 ( .A(n511), .Y(n740) );
  INVX1 U68 ( .A(n761), .Y(n383) );
  INVX1 U69 ( .A(n591), .Y(n680) );
  INVX1 U70 ( .A(n672), .Y(n178) );
  INVX1 U71 ( .A(n578), .Y(n357) );
  INVX1 U72 ( .A(n183), .Y(n123) );
  INVXL U73 ( .A(wr_dacv[16]), .Y(n225) );
  INVX1 U74 ( .A(n197), .Y(n217) );
  INVX1 U75 ( .A(wr_dacv[12]), .Y(n240) );
  AND2X1 U76 ( .A(n390), .B(n443), .Y(N984) );
  AND2X1 U77 ( .A(n390), .B(n438), .Y(N986) );
  AND2X1 U78 ( .A(n427), .B(n438), .Y(N978) );
  INVX1 U79 ( .A(n396), .Y(n423) );
  INVX1 U80 ( .A(n437), .Y(n447) );
  AND2X1 U81 ( .A(n438), .B(n447), .Y(N974) );
  INVX1 U82 ( .A(n539), .Y(n315) );
  INVX1 U83 ( .A(n345), .Y(n538) );
  NOR2X1 U84 ( .A(n420), .B(n707), .Y(n421) );
  INVX1 U85 ( .A(n462), .Y(n748) );
  OAI21BX1 U86 ( .C(n766), .B(n216), .A(n420), .Y(n341) );
  AO21X1 U87 ( .B(n420), .C(n707), .A(n421), .Y(n734) );
  INVX1 U88 ( .A(N1148), .Y(n741) );
  AO2222XL U89 ( .A(n206), .B(n694), .C(n513), .D(n205), .E(n204), .F(n680), 
        .G(n262), .H(n22), .Y(n210) );
  INVX1 U90 ( .A(n348), .Y(n206) );
  INVX1 U91 ( .A(n351), .Y(n204) );
  NAND21X1 U92 ( .B(n203), .A(n202), .Y(n205) );
  AOI211X1 U93 ( .C(n764), .D(n765), .A(n477), .B(n213), .Y(n64) );
  AOI21X1 U94 ( .B(n766), .C(n695), .A(n479), .Y(n477) );
  INVX1 U95 ( .A(n764), .Y(n479) );
  INVX1 U96 ( .A(n755), .Y(n695) );
  INVX1 U97 ( .A(n736), .Y(N1312) );
  INVX1 U98 ( .A(n338), .Y(n715) );
  INVX1 U99 ( .A(n337), .Y(n717) );
  INVX1 U100 ( .A(n453), .Y(n708) );
  INVX1 U101 ( .A(n451), .Y(n636) );
  NOR2X1 U102 ( .A(n492), .B(n62), .Y(n489) );
  NOR2X1 U103 ( .A(n756), .B(n755), .Y(n475) );
  INVX1 U104 ( .A(n209), .Y(n681) );
  INVX1 U105 ( .A(n369), .Y(n716) );
  INVX1 U106 ( .A(n277), .Y(n735) );
  INVX1 U107 ( .A(n474), .Y(n756) );
  INVX1 U108 ( .A(n340), .Y(n710) );
  NOR21XL U109 ( .B(n696), .A(n361), .Y(n362) );
  XOR3X1 U110 ( .A(sub_398_S2_I4_aco_carry_4_), .B(n491), .C(n642), .Y(n682)
         );
  NAND21X1 U111 ( .B(n693), .A(n362), .Y(n351) );
  OA2222XL U112 ( .A(n26), .B(n351), .C(n582), .D(n350), .E(n349), .F(n348), 
        .G(n347), .H(n346), .Y(n522) );
  INVX1 U113 ( .A(n324), .Y(n349) );
  NAND2X1 U114 ( .A(n180), .B(n179), .Y(n346) );
  NAND21X1 U115 ( .B(n180), .A(n179), .Y(n607) );
  NAND21X1 U116 ( .B(n404), .A(n579), .Y(n77) );
  NAND21X1 U117 ( .B(n404), .A(n642), .Y(n641) );
  INVX1 U118 ( .A(n177), .Y(n179) );
  NAND32X1 U119 ( .B(n363), .C(n176), .A(n693), .Y(n177) );
  INVX1 U120 ( .A(n362), .Y(n176) );
  INVX1 U121 ( .A(n157), .Y(n158) );
  NAND21X1 U122 ( .B(n196), .A(n308), .Y(n157) );
  NAND3X1 U123 ( .A(n362), .B(n363), .C(n693), .Y(n232) );
  NOR2X1 U124 ( .A(n744), .B(n582), .Y(n572) );
  INVX1 U125 ( .A(n554), .Y(n738) );
  NOR2X1 U126 ( .A(n766), .B(n62), .Y(n339) );
  NAND2X1 U127 ( .A(n562), .B(n557), .Y(n558) );
  INVX1 U128 ( .A(n469), .Y(n757) );
  INVX1 U129 ( .A(n455), .Y(n749) );
  INVX1 U130 ( .A(n275), .Y(n752) );
  INVX1 U131 ( .A(sub_398_S2_I4_aco_carry_4_), .Y(n639) );
  XOR2X1 U132 ( .A(n166), .B(n162), .Y(n672) );
  NAND2X1 U133 ( .A(n361), .B(n696), .Y(n348) );
  NAND21X1 U134 ( .B(n707), .A(n766), .Y(n635) );
  AOI21X1 U135 ( .B(n755), .C(n756), .A(n475), .Y(n466) );
  NAND2X1 U136 ( .A(n196), .B(n308), .Y(n234) );
  OA21X1 U137 ( .B(n692), .C(n518), .A(n515), .Y(n265) );
  NOR2X1 U138 ( .A(n679), .B(n492), .Y(n518) );
  NOR2X1 U139 ( .A(n582), .B(n583), .Y(n573) );
  INVX1 U140 ( .A(n744), .Y(n583) );
  INVX1 U141 ( .A(n754), .Y(n532) );
  INVX1 U142 ( .A(n492), .Y(n172) );
  INVX1 U143 ( .A(n287), .Y(n92) );
  INVX1 U144 ( .A(n634), .Y(n679) );
  INVX1 U145 ( .A(n168), .Y(n163) );
  INVX1 U146 ( .A(n552), .Y(n739) );
  NOR2X1 U147 ( .A(n535), .B(n755), .Y(n528) );
  INVX1 U148 ( .A(n200), .Y(n694) );
  NAND2X1 U149 ( .A(n518), .B(n692), .Y(n515) );
  AO21X1 U150 ( .B(n89), .C(n111), .A(n88), .Y(n125) );
  INVX1 U151 ( .A(n219), .Y(n89) );
  MUX2X1 U152 ( .D0(n87), .D1(n86), .S(n320), .Y(n88) );
  MUX4X1 U153 ( .D0(n102), .D1(n99), .D2(n101), .D3(n98), .S0(n81), .S1(n80), 
        .Y(n87) );
  AO21X1 U154 ( .B(n112), .C(n111), .A(n110), .Y(n183) );
  MUX4X1 U155 ( .D0(n109), .D1(n108), .D2(n107), .D3(n106), .S0(n10), .S1(n105), .Y(n110) );
  XOR2X1 U156 ( .A(n691), .B(n104), .Y(n105) );
  AO21X1 U157 ( .B(n566), .C(n102), .A(n101), .Y(n107) );
  XOR2X1 U158 ( .A(n84), .B(n692), .Y(n189) );
  XNOR2XL U159 ( .A(n766), .B(n679), .Y(n511) );
  NAND21X1 U160 ( .B(n492), .A(n355), .Y(n84) );
  AO21X1 U161 ( .B(n566), .C(n100), .A(n719), .Y(n108) );
  AO21X1 U162 ( .B(n566), .C(n99), .A(n98), .Y(n109) );
  NOR2X1 U163 ( .A(n703), .B(n684), .Y(n596) );
  INVX1 U164 ( .A(n592), .Y(n294) );
  INVX1 U165 ( .A(n566), .Y(n356) );
  AOI21X1 U166 ( .B(n103), .C(n695), .A(n104), .Y(n10) );
  AOI21X1 U167 ( .B(n535), .C(n755), .A(n528), .Y(n11) );
  INVX1 U168 ( .A(n103), .Y(n96) );
  INVX1 U169 ( .A(n218), .Y(n112) );
  INVX1 U170 ( .A(n76), .Y(n195) );
  NAND21X1 U171 ( .B(n294), .A(n75), .Y(n76) );
  NAND21X1 U172 ( .B(n27), .A(n78), .Y(n219) );
  NAND21X1 U173 ( .B(n644), .A(n481), .Y(n761) );
  XOR2X1 U174 ( .A(n678), .B(n78), .Y(n80) );
  INVX1 U175 ( .A(n355), .Y(n78) );
  INVX1 U176 ( .A(n85), .Y(n320) );
  OAI211X1 U177 ( .C(n707), .D(n355), .A(n84), .B(n635), .Y(n85) );
  INVX1 U178 ( .A(n174), .Y(n307) );
  OAI211X1 U179 ( .C(n707), .D(n634), .A(n635), .B(n173), .Y(n174) );
  INVX1 U180 ( .A(n518), .Y(n173) );
  MUX4X1 U181 ( .D0(n726), .D1(n724), .D2(n117), .D3(n720), .S0(n116), .S1(
        n115), .Y(n119) );
  AND2X1 U182 ( .A(n222), .B(n725), .Y(n117) );
  NAND21X1 U183 ( .B(n195), .A(n594), .Y(n591) );
  XNOR2XL U184 ( .A(n592), .B(n596), .Y(n594) );
  NOR2X1 U185 ( .A(n677), .B(n395), .Y(n379) );
  INVX1 U186 ( .A(n645), .Y(n395) );
  INVX1 U187 ( .A(n187), .Y(n116) );
  XOR2X1 U188 ( .A(n355), .B(n678), .Y(n578) );
  XNOR2XL U189 ( .A(n94), .B(n691), .Y(n12) );
  OAI211X1 U190 ( .C(n371), .D(n360), .A(n359), .B(n358), .Y(ps_ptr[1]) );
  INVX1 U191 ( .A(n551), .Y(n371) );
  AOI32X1 U192 ( .A(n507), .B(n506), .C(n354), .D(n353), .E(n352), .Y(n359) );
  MUX2X1 U193 ( .D0(n280), .D1(n267), .S(cs_ptr[0]), .Y(n281) );
  AO21XL U194 ( .B(n353), .C(n263), .A(n564), .Y(n267) );
  NAND43X1 U195 ( .B(n262), .C(n520), .D(n261), .A(n351), .Y(n263) );
  OAI211X1 U196 ( .C(n222), .D(n360), .A(n221), .B(n220), .Y(ps_ptr[4]) );
  AOI32XL U197 ( .A(n217), .B(n312), .C(n215), .D(n353), .E(n211), .Y(n221) );
  NAND21X1 U198 ( .B(n210), .A(n208), .Y(n211) );
  OAI22AX1 U199 ( .D(n599), .C(n595), .A(n52), .B(n597), .Y(n598) );
  AOI221XL U200 ( .A(n580), .B(n578), .C(n577), .D(n566), .E(n565), .Y(n586)
         );
  INVX1 U201 ( .A(n503), .Y(n600) );
  INVX1 U202 ( .A(n198), .Y(n312) );
  INVX1 U203 ( .A(n56), .Y(n609) );
  INVX1 U204 ( .A(n413), .Y(n427) );
  NAND21X1 U205 ( .B(n407), .A(n406), .Y(n413) );
  NAND21X1 U206 ( .B(n394), .A(n407), .Y(n437) );
  NAND21X1 U207 ( .B(n393), .A(n407), .Y(n396) );
  INVX1 U208 ( .A(n388), .Y(n390) );
  NAND21X1 U209 ( .B(n407), .A(n684), .Y(n388) );
  AND2X1 U210 ( .A(n390), .B(n440), .Y(N985) );
  AND2X1 U211 ( .A(n390), .B(n37), .Y(N987) );
  AND2X1 U212 ( .A(n427), .B(n37), .Y(N979) );
  AND2X1 U213 ( .A(n423), .B(n37), .Y(N983) );
  AND2X1 U214 ( .A(n375), .B(n443), .Y(N988) );
  AND2X1 U215 ( .A(n375), .B(n440), .Y(N989) );
  AND2X1 U216 ( .A(n37), .B(n447), .Y(N975) );
  AND2X1 U217 ( .A(n440), .B(n447), .Y(N973) );
  NAND21X1 U218 ( .B(n249), .A(n286), .Y(n345) );
  NAND21X1 U219 ( .B(n251), .A(n250), .Y(n539) );
  INVX1 U220 ( .A(n282), .Y(n506) );
  INVX1 U221 ( .A(n653), .Y(n612) );
  NOR32XL U222 ( .B(n716), .C(n368), .A(n377), .Y(n364) );
  XOR3X1 U223 ( .A(sub_398_S2_I5_aco_carry_4_), .B(n216), .C(n683), .Y(n736)
         );
  NAND21X1 U224 ( .B(n636), .A(n637), .Y(n755) );
  NAND21X1 U225 ( .B(n365), .A(n364), .Y(n243) );
  OR2X1 U226 ( .A(n684), .B(n13), .Y(n750) );
  MUX2IX1 U227 ( .D0(n53), .D1(n638), .S(n637), .Y(n13) );
  NAND21X1 U228 ( .B(n684), .A(n638), .Y(n287) );
  OAI211X1 U229 ( .C(n425), .D(n32), .A(n426), .B(n3), .Y(n216) );
  OAI21X1 U230 ( .B(n707), .C(n766), .A(n683), .Y(n426) );
  OAI221X1 U231 ( .A(n445), .B(n194), .C(n444), .D(n747), .E(n446), .Y(n209)
         );
  GEN2XL U232 ( .D(n688), .E(n686), .C(n749), .B(n449), .A(n450), .Y(n446) );
  INVX1 U233 ( .A(N1394), .Y(n194) );
  AOI22X1 U234 ( .A(n455), .B(n456), .C(n457), .D(n749), .Y(n444) );
  INVX1 U235 ( .A(n5), .Y(n766) );
  NOR2X1 U236 ( .A(n209), .B(n376), .Y(n366) );
  NAND31X1 U237 ( .C(n326), .A(n14), .B(n522), .Y(n352) );
  AOI22X1 U238 ( .A(n328), .B(n513), .C(n520), .D(n514), .Y(n14) );
  INVX1 U239 ( .A(n393), .Y(n684) );
  NOR2X1 U240 ( .A(n5), .B(n63), .Y(n462) );
  NAND2X1 U241 ( .A(n5), .B(n216), .Y(n420) );
  NAND2X1 U242 ( .A(n421), .B(n32), .Y(sub_398_S2_I5_aco_carry_4_) );
  INVX1 U243 ( .A(n519), .Y(n707) );
  INVX1 U244 ( .A(n113), .Y(n677) );
  INVX1 U245 ( .A(n758), .Y(n691) );
  INVX1 U246 ( .A(n632), .Y(n478) );
  INVX1 U247 ( .A(n683), .Y(n425) );
  OAI31XL U248 ( .A(n278), .B(N1394), .C(n460), .D(n690), .Y(n456) );
  AOI211X1 U249 ( .C(n750), .D(n691), .A(n464), .B(n212), .Y(n63) );
  AOI21X1 U250 ( .B(n755), .C(n766), .A(n465), .Y(n464) );
  INVX1 U251 ( .A(n750), .Y(n465) );
  NAND2X1 U252 ( .A(n454), .B(n758), .Y(sub_398_S2_I7_aco_carry[4]) );
  NAND3X1 U253 ( .A(n330), .B(n331), .C(n332), .Y(n328) );
  AOI22X1 U254 ( .A(n704), .B(n341), .C(n209), .D(n749), .Y(n330) );
  AOI22X1 U255 ( .A(n710), .B(n757), .C(n339), .D(n708), .Y(n331) );
  AOI221XL U256 ( .A(n715), .B(n333), .C(n717), .D(n334), .E(n335), .Y(n332)
         );
  OAI21X1 U257 ( .B(n759), .C(n767), .A(n214), .Y(N1139) );
  NAND21X1 U258 ( .B(n519), .A(n5), .Y(n492) );
  OA2222XL U259 ( .A(n242), .B(n746), .C(n383), .D(n338), .E(n453), .F(n741), 
        .G(n736), .H(n458), .Y(n202) );
  OR2X1 U260 ( .A(n684), .B(n15), .Y(n764) );
  MUX2IX1 U261 ( .D0(n53), .D1(n638), .S(n636), .Y(n15) );
  NAND2X1 U262 ( .A(n365), .B(n364), .Y(n453) );
  NAND21X1 U263 ( .B(n44), .A(n643), .Y(n451) );
  OA2222XL U264 ( .A(n24), .B(n346), .C(n304), .D(n351), .E(n301), .F(n607), 
        .G(n11), .H(n348), .Y(n311) );
  INVX1 U265 ( .A(n303), .Y(n304) );
  AND2X1 U266 ( .A(n300), .B(n298), .Y(n301) );
  OA2222XL U267 ( .A(n706), .B(n458), .C(n242), .D(n297), .E(n453), .F(n296), 
        .G(n730), .H(n337), .Y(n300) );
  INVX1 U268 ( .A(N1230), .Y(n753) );
  AOI21X1 U269 ( .B(n472), .C(n757), .A(n473), .Y(n467) );
  AOI22X1 U270 ( .A(n469), .B(n470), .C(n471), .D(n757), .Y(n468) );
  OAI21X1 U271 ( .B(n475), .C(n476), .A(sub_398_S2_I3_aco_carry[4]), .Y(n275)
         );
  OAI21X1 U272 ( .B(n421), .C(n32), .A(sub_398_S2_I5_aco_carry_4_), .Y(n277)
         );
  INVX1 U273 ( .A(n490), .Y(n692) );
  NOR2X1 U274 ( .A(n6), .B(n64), .Y(n474) );
  NAND3X1 U275 ( .A(n716), .B(n377), .C(n368), .Y(n338) );
  NOR3XL U276 ( .A(n692), .B(n492), .C(n214), .Y(n62) );
  NAND2X1 U277 ( .A(n368), .B(n369), .Y(n340) );
  NAND2X1 U278 ( .A(n681), .B(n376), .Y(n337) );
  INVX1 U279 ( .A(n767), .Y(n463) );
  OAI21X1 U280 ( .B(n454), .C(n758), .A(sub_398_S2_I7_aco_carry[4]), .Y(n278)
         );
  INVX1 U281 ( .A(n476), .Y(n765) );
  AO2222XL U282 ( .A(n732), .B(n717), .C(N1394), .D(n209), .E(N1230), .F(n710), 
        .G(n52), .H(n201), .Y(n203) );
  INVX1 U283 ( .A(n244), .Y(n732) );
  INVX1 U284 ( .A(n243), .Y(n201) );
  OAI22X1 U285 ( .A(n242), .B(n649), .C(n243), .D(n648), .Y(n273) );
  INVX1 U286 ( .A(n274), .Y(n649) );
  OAI22X1 U287 ( .A(n709), .B(n752), .C(n689), .D(n275), .Y(n471) );
  OAI31XL U288 ( .A(n275), .B(N1230), .C(n460), .D(n690), .Y(n470) );
  INVX1 U289 ( .A(n458), .Y(n704) );
  INVX1 U290 ( .A(n759), .Y(n452) );
  AND2X1 U291 ( .A(n182), .B(n181), .Y(n185) );
  OA2222XL U292 ( .A(n763), .B(n351), .C(n583), .D(n350), .E(n532), .F(n348), 
        .G(n178), .H(n346), .Y(n182) );
  AOI221XL U293 ( .A(n520), .B(n712), .C(n266), .D(n513), .E(n264), .Y(n181)
         );
  NAND2X1 U294 ( .A(n475), .B(n476), .Y(sub_398_S2_I3_aco_carry[4]) );
  NAND2X1 U295 ( .A(n489), .B(n490), .Y(sub_398_S2_aco_carry[4]) );
  NAND3X1 U296 ( .A(n268), .B(n269), .C(n270), .Y(n266) );
  AOI22X1 U297 ( .A(n704), .B(n277), .C(n209), .D(n278), .Y(n268) );
  AOI22X1 U298 ( .A(n710), .B(n275), .C(n708), .D(n276), .Y(n269) );
  AOI221XL U299 ( .A(n715), .B(n271), .C(n717), .D(n272), .E(n273), .Y(n270)
         );
  OAI21X1 U300 ( .B(n556), .C(n562), .A(n767), .Y(n557) );
  MUX2X1 U301 ( .D0(n630), .D1(n16), .S(n579), .Y(n743) );
  NAND2X1 U302 ( .A(n142), .B(n630), .Y(n16) );
  AO21X1 U303 ( .B(n641), .C(n640), .A(n639), .Y(n274) );
  INVX1 U304 ( .A(n762), .Y(n640) );
  NAND21X1 U305 ( .B(n762), .A(n141), .Y(n142) );
  NOR32XL U306 ( .B(n738), .C(n233), .A(n460), .Y(n555) );
  INVX1 U307 ( .A(n160), .Y(n696) );
  NAND21X1 U308 ( .B(n159), .A(n158), .Y(n160) );
  OAI21BBX1 U309 ( .A(n561), .B(n32), .C(n558), .Y(n554) );
  NAND21X1 U310 ( .B(n193), .A(n192), .Y(n642) );
  NAND21X1 U311 ( .B(n491), .A(n191), .Y(n192) );
  NAND21X1 U312 ( .B(n404), .A(n762), .Y(n191) );
  NAND21X1 U313 ( .B(n584), .A(n585), .Y(n579) );
  INVX1 U314 ( .A(n631), .Y(n584) );
  OAI21X1 U315 ( .B(n762), .C(n404), .A(n697), .Y(n585) );
  INVX1 U316 ( .A(n630), .Y(n697) );
  AOI21X1 U317 ( .B(n6), .C(n64), .A(n474), .Y(n469) );
  AOI21X1 U318 ( .B(n6), .C(n63), .A(n462), .Y(n455) );
  MUX2X1 U319 ( .D0(n556), .D1(n17), .S(n557), .Y(n233) );
  NAND2X1 U320 ( .A(n558), .B(n556), .Y(n17) );
  XOR2X1 U321 ( .A(n433), .B(n48), .Y(n334) );
  NAND21X1 U322 ( .B(n293), .A(cs_ptr[1]), .Y(n404) );
  AO21X1 U323 ( .B(n53), .C(n451), .A(n463), .Y(n213) );
  INVX1 U324 ( .A(n673), .Y(n582) );
  NAND2X1 U325 ( .A(n401), .B(n762), .Y(sub_398_S2_I4_aco_carry_4_) );
  AND3X1 U326 ( .A(n232), .B(n348), .C(n258), .Y(n259) );
  OA21X1 U327 ( .B(n257), .C(n607), .A(n234), .Y(n258) );
  AND4X1 U328 ( .A(n681), .B(n340), .C(n458), .D(n453), .Y(n257) );
  INVX1 U329 ( .A(n167), .Y(n293) );
  NOR3XL U330 ( .A(n32), .B(n707), .C(n766), .Y(n562) );
  OAI22X1 U331 ( .A(n738), .B(n709), .C(n689), .D(n554), .Y(n553) );
  OAI21X1 U332 ( .B(n391), .C(n731), .A(n674), .Y(n430) );
  OAI22X1 U333 ( .A(n738), .B(n688), .C(n686), .D(n554), .Y(n559) );
  OAI21X1 U334 ( .B(n687), .C(n752), .A(n685), .Y(n472) );
  OAI22X1 U335 ( .A(n738), .B(n687), .C(n685), .D(n554), .Y(n560) );
  INVX1 U336 ( .A(n74), .Y(n75) );
  OAI21X1 U337 ( .B(n675), .C(n731), .A(n676), .Y(n435) );
  OAI31XL U338 ( .A(n274), .B(n682), .C(n386), .D(n701), .Y(n402) );
  OAI21X1 U339 ( .B(n233), .C(n445), .A(n147), .Y(n196) );
  MUX2X1 U340 ( .D0(n549), .D1(n550), .S(n4), .Y(n147) );
  AOI22X1 U341 ( .A(n739), .B(n559), .C(n552), .D(n560), .Y(n549) );
  AOI221XL U342 ( .A(n552), .B(n553), .C(n719), .D(n554), .E(n555), .Y(n550)
         );
  AOI21X1 U343 ( .B(n688), .C(n686), .A(n757), .Y(n473) );
  NAND2X1 U344 ( .A(n441), .B(n433), .Y(n432) );
  OAI21BBX1 U345 ( .A(n685), .B(n687), .C(n749), .Y(n449) );
  AO21X1 U346 ( .B(n370), .C(n513), .A(n260), .Y(n261) );
  INVX1 U347 ( .A(n350), .Y(n260) );
  NAND4X1 U348 ( .A(n243), .B(n242), .C(n338), .D(n337), .Y(n370) );
  NAND3X1 U349 ( .A(n557), .B(n519), .C(n6), .Y(n561) );
  INVX1 U350 ( .A(n272), .Y(n731) );
  OA2222XL U351 ( .A(n234), .B(n233), .C(n232), .D(n231), .E(n743), .F(n350), 
        .G(n308), .H(n207), .Y(n208) );
  XOR2X1 U352 ( .A(n476), .B(n528), .Y(n754) );
  NOR21XL U353 ( .B(n393), .A(n190), .Y(n491) );
  MUX2IX1 U354 ( .D0(n52), .D1(n638), .S(n643), .Y(n190) );
  NAND2X1 U355 ( .A(n159), .B(n158), .Y(n350) );
  NAND21X1 U356 ( .B(n6), .A(n531), .Y(n535) );
  OR2X1 U357 ( .A(n52), .B(n18), .Y(n634) );
  AOI21X1 U358 ( .B(n172), .C(n692), .A(n33), .Y(n18) );
  OAI211X1 U359 ( .C(n530), .D(n765), .A(n536), .B(n767), .Y(n531) );
  AO21X1 U360 ( .B(n766), .C(n695), .A(n530), .Y(n536) );
  NAND21X1 U361 ( .B(n167), .A(n163), .Y(n166) );
  XNOR2XL U362 ( .A(n557), .B(n6), .Y(n552) );
  NAND21X1 U363 ( .B(n528), .A(n69), .Y(n200) );
  XNOR2XL U364 ( .A(n531), .B(n530), .Y(n69) );
  NAND21X1 U365 ( .B(n164), .A(cs_ptr[1]), .Y(n168) );
  OAI21X1 U366 ( .B(n445), .C(n200), .A(n70), .Y(n361) );
  MUX2X1 U367 ( .D0(n523), .D1(n524), .S(n11), .Y(n70) );
  AOI22AXL U368 ( .A(n533), .B(n324), .D(n324), .C(n534), .Y(n523) );
  AOI221XL U369 ( .A(n526), .B(n324), .C(n754), .D(n719), .E(n527), .Y(n524)
         );
  XOR2X1 U370 ( .A(n642), .B(cs_ptr[1]), .Y(n336) );
  MUX2X1 U371 ( .D0(n634), .D1(n19), .S(n33), .Y(n231) );
  NAND2X1 U372 ( .A(n515), .B(n634), .Y(n19) );
  AO21X1 U373 ( .B(n22), .C(n718), .A(n171), .Y(n180) );
  MUX2BXL U374 ( .D0(n170), .D1(n169), .S(n24), .Y(n171) );
  MUX2X1 U375 ( .D0(n500), .D1(n501), .S(n347), .Y(n170) );
  AOI221XL U376 ( .A(n496), .B(n165), .C(n672), .D(n720), .E(n497), .Y(n169)
         );
  INVX1 U377 ( .A(n520), .Y(n308) );
  INVX1 U378 ( .A(n733), .Y(n542) );
  OAI21X1 U379 ( .B(n489), .C(n490), .A(sub_398_S2_aco_carry[4]), .Y(n276) );
  INVX1 U380 ( .A(n638), .Y(n703) );
  INVX1 U381 ( .A(n207), .Y(n698) );
  INVX1 U382 ( .A(n161), .Y(n164) );
  OAI22X1 U383 ( .A(n709), .B(n532), .C(n689), .D(n754), .Y(n526) );
  OAI22X1 U384 ( .A(n674), .B(n712), .C(n391), .D(n546), .Y(n540) );
  OAI22X1 U385 ( .A(n676), .B(n712), .C(n675), .D(n546), .Y(n547) );
  OAI22AX1 U386 ( .D(n231), .C(n460), .A(n690), .B(n265), .Y(n510) );
  OAI22X1 U387 ( .A(n687), .B(n532), .C(n685), .D(n754), .Y(n533) );
  OAI22X1 U388 ( .A(n688), .B(n532), .C(n686), .D(n754), .Y(n534) );
  NOR2X1 U389 ( .A(n744), .B(n673), .Y(n571) );
  OAI21X1 U390 ( .B(n178), .C(n700), .A(n699), .Y(n501) );
  OAI21X1 U391 ( .B(n709), .C(n265), .A(n689), .Y(n512) );
  INVX1 U392 ( .A(n633), .Y(n441) );
  OAI21X1 U393 ( .B(n445), .C(n231), .A(n175), .Y(n363) );
  MUX2X1 U394 ( .D0(n508), .D1(n509), .S(n307), .Y(n175) );
  AOI22X1 U395 ( .A(n740), .B(n516), .C(n511), .D(n517), .Y(n508) );
  AOI22X1 U396 ( .A(n740), .B(n510), .C(n511), .D(n512), .Y(n509) );
  NOR3XL U397 ( .A(n754), .B(n460), .C(n694), .Y(n527) );
  NOR3XL U398 ( .A(n672), .B(n386), .C(n22), .Y(n497) );
  NOR3XL U399 ( .A(n698), .B(n386), .C(n712), .Y(n541) );
  INVX1 U400 ( .A(n546), .Y(n712) );
  NOR2X1 U401 ( .A(n673), .B(n583), .Y(n567) );
  OAI21BBX1 U402 ( .A(n77), .B(n762), .C(n142), .Y(n744) );
  NOR2X1 U403 ( .A(n737), .B(n766), .Y(n563) );
  INVX1 U404 ( .A(n557), .Y(n737) );
  OR2X1 U405 ( .A(n463), .B(n20), .Y(n355) );
  AOI21X1 U406 ( .B(n490), .C(n172), .A(n27), .Y(n20) );
  AO21X1 U407 ( .B(n35), .C(n93), .A(n463), .Y(n95) );
  NAND32X1 U408 ( .B(n758), .C(n6), .A(n755), .Y(n93) );
  MUX4X1 U409 ( .D0(n83), .D1(n100), .D2(n82), .D3(n719), .S0(n81), .S1(n80), 
        .Y(n86) );
  INVX1 U410 ( .A(n689), .Y(n83) );
  AND2X1 U411 ( .A(n219), .B(n79), .Y(n82) );
  INVX1 U412 ( .A(n460), .Y(n79) );
  AO21X1 U413 ( .B(n97), .C(n6), .A(n96), .Y(n566) );
  INVX1 U414 ( .A(n95), .Y(n97) );
  OAI21BX1 U415 ( .C(n6), .B(n531), .A(n535), .Y(n324) );
  NAND21X1 U416 ( .B(n644), .A(n643), .Y(n645) );
  NAND21X1 U417 ( .B(n6), .A(n95), .Y(n103) );
  OR2X1 U418 ( .A(n104), .B(n21), .Y(n218) );
  XNOR2XL U419 ( .A(n95), .B(n35), .Y(n21) );
  XOR2X1 U420 ( .A(n733), .B(cs_ptr[1]), .Y(n514) );
  INVX1 U421 ( .A(n279), .Y(n763) );
  INVX1 U422 ( .A(n114), .Y(n162) );
  INVX1 U423 ( .A(n394), .Y(n406) );
  INVX1 U424 ( .A(n165), .Y(n347) );
  XOR2X1 U425 ( .A(n161), .B(n72), .Y(n22) );
  INVX1 U426 ( .A(n760), .Y(n271) );
  OAI21X1 U427 ( .B(n178), .C(n391), .A(n674), .Y(n496) );
  OAI21X1 U428 ( .B(n760), .C(n675), .A(n676), .Y(n392) );
  OAI21X1 U429 ( .B(n178), .C(n675), .A(n676), .Y(n500) );
  OAI22X1 U430 ( .A(n689), .B(n356), .C(n460), .D(n112), .Y(n106) );
  OAI22X1 U431 ( .A(n674), .B(n271), .C(n760), .D(n391), .Y(n384) );
  OAI21X1 U432 ( .B(n688), .C(n265), .A(n686), .Y(n516) );
  OAI21X1 U433 ( .B(n687), .C(n265), .A(n685), .Y(n517) );
  INVX1 U434 ( .A(n646), .Y(n644) );
  INVX1 U435 ( .A(n139), .Y(n693) );
  OAI211X1 U436 ( .C(n587), .D(n26), .A(n588), .B(n589), .Y(n139) );
  AOI32X1 U437 ( .A(n725), .B(n591), .C(n763), .D(n720), .E(n279), .Y(n588) );
  AOI22X1 U438 ( .A(n724), .B(n279), .C(n763), .D(n726), .Y(n587) );
  NOR2X1 U439 ( .A(n125), .B(n124), .Y(n23) );
  NAND2X1 U440 ( .A(n709), .B(n689), .Y(n457) );
  AO21X1 U441 ( .B(n74), .C(n73), .A(n463), .Y(n592) );
  INVX1 U442 ( .A(n596), .Y(n73) );
  AOI21AX1 U443 ( .B(n168), .C(n167), .A(n166), .Y(n24) );
  OR2X1 U444 ( .A(n141), .B(n25), .Y(n305) );
  AOI21X1 U445 ( .B(n579), .C(n48), .A(n167), .Y(n25) );
  INVX1 U446 ( .A(n701), .Y(n720) );
  INVX1 U447 ( .A(n700), .Y(n722) );
  INVX1 U448 ( .A(n386), .Y(n725) );
  INVX1 U449 ( .A(n193), .Y(n481) );
  XNOR2XL U450 ( .A(n592), .B(cs_ptr[1]), .Y(n26) );
  AOI21X1 U451 ( .B(n684), .C(n452), .A(n53), .Y(n27) );
  OAI21X1 U452 ( .B(n386), .C(n761), .A(n701), .Y(n385) );
  NAND2X1 U453 ( .A(n674), .B(n391), .Y(n403) );
  XNOR2XL U454 ( .A(n114), .B(n28), .Y(n187) );
  NAND2X1 U455 ( .A(n321), .B(n293), .Y(n28) );
  INVX1 U456 ( .A(n647), .Y(n333) );
  NAND21X1 U457 ( .B(n48), .A(n646), .Y(n647) );
  INVX1 U458 ( .A(n690), .Y(n719) );
  NAND21X1 U459 ( .B(n113), .A(n684), .Y(n222) );
  INVX1 U460 ( .A(n382), .Y(n718) );
  INVX1 U461 ( .A(n709), .Y(n100) );
  INVX1 U462 ( .A(n674), .Y(n726) );
  INVX1 U463 ( .A(n685), .Y(n102) );
  INVX1 U464 ( .A(n687), .Y(n99) );
  INVX1 U465 ( .A(n686), .Y(n101) );
  INVX1 U466 ( .A(n688), .Y(n98) );
  INVX1 U467 ( .A(n391), .Y(n724) );
  OAI222XL U468 ( .A(n681), .B(n495), .C(n242), .D(n494), .E(n340), .F(n493), 
        .Y(n498) );
  OAI211X1 U469 ( .C(n491), .D(n642), .A(n639), .B(n481), .Y(n494) );
  XOR2X1 U470 ( .A(n213), .B(sub_398_S2_I3_aco_carry[5]), .Y(n493) );
  XOR2X1 U471 ( .A(n212), .B(sub_398_S2_I7_aco_carry[5]), .Y(n495) );
  XNOR2XL U472 ( .A(n118), .B(n293), .Y(n29) );
  INVX1 U473 ( .A(n742), .Y(n297) );
  INVX1 U474 ( .A(n118), .Y(n321) );
  OA21X1 U475 ( .B(n52), .C(n48), .A(n118), .Y(n115) );
  INVX1 U476 ( .A(n445), .Y(n111) );
  XOR2X1 U477 ( .A(n480), .B(n3), .Y(n499) );
  OAI22X1 U478 ( .A(n216), .B(n461), .C(n459), .D(n425), .Y(n480) );
  AND2X1 U479 ( .A(n216), .B(n461), .Y(n459) );
  INVX1 U480 ( .A(sub_398_S2_I5_aco_carry_4_), .Y(n461) );
  XNOR2XL U481 ( .A(sub_398_S2_aco_carry[5]), .B(n214), .Y(n502) );
  INVX1 U482 ( .A(n405), .Y(n443) );
  INVX1 U483 ( .A(n397), .Y(n438) );
  AND2X1 U484 ( .A(n255), .B(n254), .Y(n283) );
  NAND21X1 U485 ( .B(wr_dacv[3]), .A(n714), .Y(n284) );
  NAND2X1 U486 ( .A(n30), .B(n503), .Y(n599) );
  OAI22XL U487 ( .A(ps_ptr[2]), .B(n601), .C(ps_ptr[3]), .D(n648), .Y(n30) );
  AND2X1 U488 ( .A(n311), .B(n310), .Y(n318) );
  NAND32XL U489 ( .B(wr_dacv[15]), .C(n236), .A(n228), .Y(n325) );
  INVX1 U490 ( .A(n199), .Y(n327) );
  AND2X1 U491 ( .A(n344), .B(n343), .Y(n544) );
  AOI221XL U492 ( .A(n520), .B(n514), .C(n328), .D(n513), .E(n326), .Y(n521)
         );
  NAND32XL U493 ( .B(wr_dacv[9]), .C(n248), .A(n247), .Y(n252) );
  AND3X1 U494 ( .A(n246), .B(n329), .C(n245), .Y(n248) );
  AND3X1 U495 ( .A(n240), .B(n239), .C(n238), .Y(n241) );
  NAND21XL U496 ( .B(wr_dacv[8]), .A(n128), .Y(n129) );
  OAI211X1 U497 ( .C(n237), .D(n236), .A(n235), .B(n230), .Y(n238) );
  INVX1 U498 ( .A(wr_dacv[13]), .Y(n235) );
  AND3X1 U499 ( .A(n229), .B(n228), .C(n227), .Y(n237) );
  INVXL U500 ( .A(wr_dacv[15]), .Y(n229) );
  AOI21BBXL U501 ( .B(n52), .C(n199), .A(n313), .Y(n215) );
  INVX1 U502 ( .A(n387), .Y(n407) );
  AND2X1 U503 ( .A(n440), .B(n424), .Y(N981) );
  AND2X1 U504 ( .A(n443), .B(n424), .Y(N980) );
  AND3X1 U505 ( .A(n427), .B(n443), .C(n442), .Y(N976) );
  AND3X1 U506 ( .A(n427), .B(n440), .C(n442), .Y(N977) );
  OAI32X1 U507 ( .A(n405), .B(n437), .C(n442), .D(n397), .E(n396), .Y(N982) );
  INVX1 U508 ( .A(n58), .Y(n611) );
  AND3X1 U509 ( .A(n447), .B(n443), .C(n442), .Y(N972) );
  INVX1 U510 ( .A(n372), .Y(n375) );
  NAND21X1 U511 ( .B(n387), .A(n703), .Y(n372) );
  OR3XL U512 ( .A(sampl_done), .B(n58), .C(sampl_begn), .Y(N971) );
  NAND21X1 U513 ( .B(wr_dacv[5]), .A(n133), .Y(n249) );
  INVX1 U514 ( .A(n134), .Y(n286) );
  NAND21X1 U515 ( .B(wr_dacv[4]), .A(n713), .Y(n134) );
  NAND21X1 U516 ( .B(wr_dacv[1]), .A(n136), .Y(n282) );
  NAND21X1 U517 ( .B(wr_dacv[7]), .A(n729), .Y(n251) );
  INVX1 U518 ( .A(n138), .Y(n250) );
  NAND21X1 U519 ( .B(wr_dacv[6]), .A(n137), .Y(n138) );
  INVX1 U520 ( .A(n50), .Y(cs_ptr[1]) );
  INVX1 U521 ( .A(n45), .Y(cs_ptr[0]) );
  INVX1 U522 ( .A(n55), .Y(cs_ptr[4]) );
  NAND2X1 U523 ( .A(sampl_done), .B(n654), .Y(n653) );
  NAND2X1 U524 ( .A(n654), .B(n653), .Y(N949) );
  NOR32XL U525 ( .B(n366), .C(n367), .A(n378), .Y(n368) );
  MUX2X1 U526 ( .D0(n287), .D1(n54), .S(n478), .Y(n683) );
  XOR2X1 U527 ( .A(n448), .B(n41), .Y(n758) );
  OR2X1 U528 ( .A(n68), .B(n31), .Y(n519) );
  MUX2IX1 U529 ( .D0(n601), .D1(n289), .S(n44), .Y(n31) );
  NAND21X1 U530 ( .B(n52), .A(cs_ptr[3]), .Y(n393) );
  NAND21X1 U531 ( .B(n601), .A(cs_ptr[1]), .Y(n113) );
  AO21X1 U532 ( .B(n46), .C(n601), .A(n643), .Y(n632) );
  NAND3X1 U533 ( .A(n366), .B(n378), .C(n367), .Y(n242) );
  AO21X1 U534 ( .B(n53), .C(n448), .A(n463), .Y(n212) );
  INVX1 U535 ( .A(n295), .Y(n643) );
  INVX1 U536 ( .A(n448), .Y(n637) );
  INVX1 U537 ( .A(n54), .Y(n52) );
  XNOR2XL U538 ( .A(n632), .B(n41), .Y(n32) );
  INVX1 U539 ( .A(n45), .Y(n44) );
  OAI22X1 U540 ( .A(n336), .B(n242), .C(n243), .D(n49), .Y(n335) );
  NAND21X1 U541 ( .B(n41), .A(n52), .Y(n638) );
  XOR2X1 U542 ( .A(n451), .B(n41), .Y(n476) );
  XOR2X1 U543 ( .A(n759), .B(n41), .Y(n490) );
  NAND21X1 U544 ( .B(n55), .A(n41), .Y(n767) );
  NAND21X1 U545 ( .B(n367), .A(n366), .Y(n458) );
  AO21X1 U546 ( .B(n41), .C(n452), .A(n53), .Y(n214) );
  NAND21X1 U547 ( .B(n45), .A(n677), .Y(n759) );
  OA2222XL U548 ( .A(n340), .B(n466), .C(n243), .D(n601), .E(n681), .F(n450), 
        .G(n379), .H(n338), .Y(n298) );
  OAI211X1 U549 ( .C(n741), .D(n445), .A(n61), .B(n709), .Y(n365) );
  MUX2X1 U550 ( .D0(n60), .D1(n59), .S(n43), .Y(n61) );
  NOR2X1 U551 ( .A(n482), .B(n483), .Y(n60) );
  NOR2X1 U552 ( .A(n486), .B(n487), .Y(n59) );
  INVX1 U553 ( .A(n439), .Y(n68) );
  INVX1 U554 ( .A(n54), .Y(n53) );
  INVX1 U555 ( .A(n50), .Y(n48) );
  AO21X1 U556 ( .B(n295), .C(n648), .A(n75), .Y(n762) );
  AO21X1 U557 ( .B(n288), .C(n633), .A(n53), .Y(n433) );
  XOR2X1 U558 ( .A(n50), .B(n579), .Y(n673) );
  NAND21X1 U559 ( .B(n68), .A(n289), .Y(n167) );
  NAND21X1 U560 ( .B(n146), .A(n145), .Y(n159) );
  AOI22X1 U561 ( .A(n305), .B(n144), .C(n143), .D(n718), .Y(n145) );
  AO21X1 U562 ( .B(n567), .C(n720), .A(n140), .Y(n146) );
  INVX1 U563 ( .A(n743), .Y(n143) );
  NAND21X1 U564 ( .B(n295), .A(n41), .Y(n74) );
  OAI221X1 U565 ( .A(n398), .B(n742), .C(n382), .D(n746), .E(n399), .Y(n378)
         );
  OAI31XL U566 ( .A(n400), .B(n728), .C(n722), .D(n742), .Y(n399) );
  AOI22AXL U567 ( .A(n336), .B(n402), .D(n336), .C(n403), .Y(n398) );
  AOI21X1 U568 ( .B(n676), .C(n675), .A(n336), .Y(n400) );
  OA2222XL U569 ( .A(n309), .B(n308), .C(n232), .D(n307), .E(n306), .F(n350), 
        .G(n234), .H(n4), .Y(n310) );
  INVX1 U570 ( .A(n305), .Y(n306) );
  OAI21BBX1 U571 ( .A(n439), .B(n702), .C(n432), .Y(n272) );
  MUX2X1 U572 ( .D0(n569), .D1(n575), .S(cs_ptr[0]), .Y(n140) );
  OAI21X1 U573 ( .B(n246), .C(n745), .A(n570), .Y(n569) );
  OAI21X1 U574 ( .B(n723), .C(n745), .A(n576), .Y(n575) );
  INVX1 U575 ( .A(n573), .Y(n745) );
  OAI222XL U576 ( .A(n730), .B(n428), .C(n429), .D(n299), .E(n382), .F(n244), 
        .Y(n376) );
  AOI22AXL U577 ( .A(n334), .B(n435), .D(n334), .C(n436), .Y(n428) );
  AOI222XL U578 ( .A(n334), .B(n430), .C(n244), .D(n725), .E(n272), .F(n720), 
        .Y(n429) );
  NAND2X1 U579 ( .A(n699), .B(n700), .Y(n436) );
  NAND2X1 U580 ( .A(n431), .B(n432), .Y(n244) );
  XNOR2XL U581 ( .A(n433), .B(n434), .Y(n431) );
  INVX1 U582 ( .A(n288), .Y(n434) );
  MUX2IX1 U583 ( .D0(n151), .D1(n150), .S(n542), .Y(n207) );
  AND2X1 U584 ( .A(n149), .B(n148), .Y(n151) );
  INVX1 U585 ( .A(n150), .Y(n148) );
  XOR2X1 U586 ( .A(n601), .B(n41), .Y(n702) );
  AO21X1 U587 ( .B(n698), .C(n718), .A(n156), .Y(n520) );
  MUX2BXL U588 ( .D0(n155), .D1(n154), .S(n309), .Y(n156) );
  AOI221XL U589 ( .A(n540), .B(n514), .C(n720), .D(n712), .E(n541), .Y(n154)
         );
  AO21X1 U590 ( .B(n547), .C(n514), .A(n152), .Y(n155) );
  AO21X1 U591 ( .B(n149), .C(n150), .A(n463), .Y(n733) );
  AO21X1 U592 ( .B(n72), .C(n71), .A(n53), .Y(n161) );
  NAND32X1 U593 ( .B(n50), .C(n167), .A(n162), .Y(n71) );
  NAND21X1 U594 ( .B(n41), .A(n54), .Y(n394) );
  AO21X1 U595 ( .B(n53), .C(n295), .A(n463), .Y(n193) );
  AO21X1 U596 ( .B(n677), .C(n55), .A(n287), .Y(n72) );
  NAND21X1 U597 ( .B(n767), .A(n295), .Y(n631) );
  OR2X1 U598 ( .A(n439), .B(n702), .Y(n633) );
  OAI21BBX1 U599 ( .A(n733), .B(n441), .C(n548), .Y(n546) );
  OAI21X1 U600 ( .B(n542), .C(n439), .A(n702), .Y(n548) );
  OAI211X1 U601 ( .C(n52), .D(n295), .A(n631), .B(n394), .Y(n630) );
  MUX2X1 U602 ( .D0(n92), .D1(n54), .S(n636), .Y(n530) );
  MUX2X1 U603 ( .D0(n55), .D1(n92), .S(n478), .Y(n556) );
  MUX2X1 U604 ( .D0(n722), .D1(n728), .S(n546), .Y(n152) );
  NAND21X1 U605 ( .B(n439), .A(n702), .Y(n149) );
  AOI21X1 U606 ( .B(n452), .C(n55), .A(n287), .Y(n33) );
  INVX1 U607 ( .A(n299), .Y(n730) );
  INVX1 U608 ( .A(cs_ptr[3]), .Y(n648) );
  OR2X1 U609 ( .A(n195), .B(n34), .Y(n279) );
  AOI21X1 U610 ( .B(n643), .C(n592), .A(n769), .Y(n34) );
  MUX2X1 U611 ( .D0(n136), .D1(n135), .S(cs_ptr[0]), .Y(n460) );
  MUX2X1 U612 ( .D0(n714), .D1(n255), .S(cs_ptr[0]), .Y(n689) );
  MUX2X1 U613 ( .D0(n723), .D1(n246), .S(n44), .Y(n709) );
  MUX2X1 U614 ( .D0(n255), .D1(n714), .S(n43), .Y(n674) );
  AO21X1 U615 ( .B(n246), .C(n46), .A(n132), .Y(n391) );
  MUX2X1 U616 ( .D0(n239), .D1(n230), .S(n43), .Y(n700) );
  NAND21X1 U617 ( .B(n295), .A(n406), .Y(n646) );
  AO21X1 U618 ( .B(n293), .C(n49), .A(n401), .Y(n742) );
  XOR2X1 U619 ( .A(n645), .B(cs_ptr[3]), .Y(n760) );
  XOR2X1 U620 ( .A(n113), .B(cs_ptr[3]), .Y(n114) );
  AO21X1 U621 ( .B(n164), .C(n49), .A(n163), .Y(n165) );
  OAI222XL U622 ( .A(n379), .B(n380), .C(n381), .D(n711), .E(n382), .F(n383), 
        .Y(n377) );
  INVX1 U623 ( .A(n379), .Y(n711) );
  AOI211X1 U624 ( .C(n333), .D(n392), .A(n728), .B(n722), .Y(n380) );
  AOI22AXL U625 ( .A(n333), .B(n384), .D(n333), .C(n385), .Y(n381) );
  INVX1 U626 ( .A(n45), .Y(n43) );
  AOI22X1 U627 ( .A(n590), .B(n303), .C(n680), .D(n718), .Y(n589) );
  OAI222XL U628 ( .A(n699), .B(n279), .C(n763), .D(n700), .E(n593), .F(n26), 
        .Y(n590) );
  AOI22X1 U629 ( .A(n721), .B(n279), .C(n763), .D(n727), .Y(n593) );
  INVX1 U630 ( .A(n322), .Y(n132) );
  MUX2X1 U631 ( .D0(n223), .D1(n67), .S(cs_ptr[0]), .Y(n445) );
  MUX2X1 U632 ( .D0(n729), .D1(n137), .S(n43), .Y(n685) );
  MUX2X1 U633 ( .D0(n228), .D1(n126), .S(n43), .Y(n687) );
  MUX2X1 U634 ( .D0(n133), .D1(n713), .S(n43), .Y(n686) );
  MUX2X1 U635 ( .D0(n230), .D1(n239), .S(n43), .Y(n688) );
  MUX2X1 U636 ( .D0(n135), .D1(n136), .S(cs_ptr[0]), .Y(n386) );
  MUX2X1 U637 ( .D0(n247), .D1(n128), .S(n43), .Y(n690) );
  MUX2X1 U638 ( .D0(n67), .D1(n223), .S(n43), .Y(n382) );
  MUX2X1 U639 ( .D0(n128), .D1(n247), .S(n43), .Y(n701) );
  INVX1 U640 ( .A(n728), .Y(n699) );
  INVX1 U641 ( .A(n727), .Y(n676) );
  INVX1 U642 ( .A(n721), .Y(n675) );
  MUX2IX1 U643 ( .D0(n92), .D1(n54), .S(n637), .Y(n35) );
  AO21X1 U644 ( .B(n122), .C(n718), .A(n121), .Y(n124) );
  INVX1 U645 ( .A(n222), .Y(n122) );
  MUX2X1 U646 ( .D0(n120), .D1(n119), .S(n29), .Y(n121) );
  MUX4X1 U647 ( .D0(n727), .D1(n721), .D2(n728), .D3(n722), .S0(n116), .S1(
        n115), .Y(n120) );
  OR2X1 U648 ( .A(n677), .B(n36), .Y(n303) );
  MUX2IX1 U649 ( .D0(n295), .D1(n601), .S(n294), .Y(n36) );
  NAND21X1 U650 ( .B(n55), .A(cs_ptr[1]), .Y(n118) );
  AO21X1 U651 ( .B(n49), .C(n55), .A(n321), .Y(n551) );
  NAND32X1 U652 ( .B(n50), .C(n389), .A(n46), .Y(n397) );
  NAND32X1 U653 ( .B(n48), .C(n389), .A(n46), .Y(n405) );
  NOR3XL U654 ( .A(n49), .B(n46), .C(n389), .Y(n37) );
  INVX1 U655 ( .A(n374), .Y(n440) );
  NAND32X1 U656 ( .B(n46), .C(n389), .A(n49), .Y(n374) );
  NAND3X1 U657 ( .A(n651), .B(n650), .C(n652), .Y(n659) );
  NAND3X1 U658 ( .A(n665), .B(n664), .C(n666), .Y(n660) );
  NAND3X1 U659 ( .A(n668), .B(n667), .C(n669), .Y(n661) );
  NAND43X1 U660 ( .B(r_dac_en[17]), .C(r_dac_en[16]), .D(wr_dacv[17]), .A(n225), .Y(n199) );
  INVX1 U661 ( .A(r_semi), .Y(n602) );
  AOI221XL U662 ( .A(n708), .B(n502), .C(n704), .D(n499), .E(n498), .Y(n608)
         );
  GEN2XL U663 ( .D(n327), .E(n7), .C(n313), .B(n312), .A(n345), .Y(n314) );
  NAND32X1 U664 ( .B(r_dac_en[16]), .C(n226), .A(n225), .Y(n227) );
  AND3X1 U665 ( .A(n224), .B(n45), .C(n223), .Y(n226) );
  INVXL U666 ( .A(wr_dacv[17]), .Y(n224) );
  INVX1 U667 ( .A(n127), .Y(n323) );
  NAND43X1 U668 ( .B(r_dac_en[13]), .C(r_dac_en[12]), .D(wr_dacv[13]), .A(n240), .Y(n127) );
  INVX1 U669 ( .A(n130), .Y(n344) );
  NAND21X1 U670 ( .B(r_dac_en[9]), .A(n253), .Y(n130) );
  NAND21X1 U671 ( .B(pos_dacis[10]), .A(n663), .Y(app_dacis[10]) );
  NAND21X1 U672 ( .B(pos_dacis[7]), .A(n666), .Y(app_dacis[7]) );
  NAND21X1 U673 ( .B(pos_dacis[8]), .A(n665), .Y(app_dacis[8]) );
  NAND21X1 U674 ( .B(pos_dacis[11]), .A(n662), .Y(app_dacis[11]) );
  NAND21X1 U675 ( .B(pos_dacis[16]), .A(n650), .Y(app_dacis[16]) );
  NAND21X1 U676 ( .B(pos_dacis[3]), .A(n668), .Y(app_dacis[3]) );
  NAND21X1 U677 ( .B(pos_dacis[4]), .A(n667), .Y(app_dacis[4]) );
  NAND21X1 U678 ( .B(pos_dacis[6]), .A(n615), .Y(app_dacis[6]) );
  INVX1 U679 ( .A(neg_dacis_6_), .Y(n615) );
  NAND21X1 U680 ( .B(pos_dacis[5]), .A(n614), .Y(app_dacis[5]) );
  INVX1 U681 ( .A(neg_dacis_5_), .Y(n614) );
  NAND21X1 U682 ( .B(pos_dacis[2]), .A(n669), .Y(app_dacis[2]) );
  NAND21XL U683 ( .B(pos_dacis[0]), .A(n670), .Y(app_dacis[0]) );
  NAND21XL U684 ( .B(pos_dacis[1]), .A(n613), .Y(app_dacis[1]) );
  INVX1 U685 ( .A(neg_dacis_1_), .Y(n613) );
  NAND21X1 U686 ( .B(pos_dacis[17]), .A(n618), .Y(app_dacis[17]) );
  INVX1 U687 ( .A(test_so1), .Y(n618) );
  NAND21X1 U688 ( .B(pos_dacis[14]), .A(n652), .Y(app_dacis[14]) );
  NAND21X1 U689 ( .B(pos_dacis[15]), .A(n651), .Y(app_dacis[15]) );
  NAND21X1 U690 ( .B(pos_dacis[9]), .A(n664), .Y(app_dacis[9]) );
  INVX1 U691 ( .A(neg_dacis_11_), .Y(n662) );
  INVX1 U692 ( .A(neg_dacis_10_), .Y(n663) );
  INVX1 U693 ( .A(neg_dacis_0_), .Y(n670) );
  INVX1 U694 ( .A(neg_dacis_15_), .Y(n651) );
  INVX1 U695 ( .A(neg_dacis_8_), .Y(n665) );
  INVX1 U696 ( .A(neg_dacis_3_), .Y(n668) );
  INVX1 U697 ( .A(neg_dacis_16_), .Y(n650) );
  INVX1 U698 ( .A(neg_dacis_9_), .Y(n664) );
  INVX1 U699 ( .A(neg_dacis_4_), .Y(n667) );
  INVX1 U700 ( .A(neg_dacis_14_), .Y(n652) );
  INVX1 U701 ( .A(neg_dacis_7_), .Y(n666) );
  INVX1 U702 ( .A(neg_dacis_2_), .Y(n669) );
  NAND21X1 U703 ( .B(pos_dacis[13]), .A(n617), .Y(app_dacis[13]) );
  INVX1 U704 ( .A(neg_dacis_13_), .Y(n617) );
  NAND21X1 U705 ( .B(pos_dacis[12]), .A(n616), .Y(app_dacis[12]) );
  INVX1 U706 ( .A(neg_dacis_12_), .Y(n616) );
  AO21X1 U707 ( .B(ps_md4ch), .C(n406), .A(n7), .Y(n387) );
  AO21X1 U708 ( .B(r_comp_swtch), .C(n427), .A(n423), .Y(n424) );
  AO21X1 U709 ( .B(n57), .C(n373), .A(n609), .Y(N994) );
  INVXL U710 ( .A(stop), .Y(n57) );
  NAND21XL U711 ( .B(stop), .A(srstz), .Y(n58) );
  NAND43X1 U712 ( .B(wr_dacv[2]), .C(wr_dacv[3]), .D(r_dac_en[2]), .A(n714), 
        .Y(n537) );
  BUFX3 U713 ( .A(n769), .Y(cs_ptr[3]) );
  INVX1 U714 ( .A(n770), .Y(n50) );
  INVX1 U715 ( .A(n771), .Y(n45) );
  INVX1 U716 ( .A(cs_mux_5_), .Y(busy) );
  AND3X1 U717 ( .A(n655), .B(n656), .C(n657), .Y(n654) );
  NOR3XL U718 ( .A(n661), .B(neg_dacis_1_), .C(test_so1), .Y(n655) );
  NOR3XL U719 ( .A(n660), .B(neg_dacis_6_), .C(neg_dacis_5_), .Y(n656) );
  NOR4XL U720 ( .A(n658), .B(n659), .C(neg_dacis_13_), .D(neg_dacis_12_), .Y(
        n657) );
  INVX1 U721 ( .A(n768), .Y(n55) );
  AND2X1 U722 ( .A(pos_dacis[6]), .B(n612), .Y(N956) );
  AND2X1 U723 ( .A(pos_dacis[2]), .B(n612), .Y(N952) );
  AND2X1 U724 ( .A(pos_dacis[7]), .B(n612), .Y(N957) );
  AND2X1 U725 ( .A(pos_dacis[4]), .B(n612), .Y(N954) );
  AND2X1 U726 ( .A(pos_dacis[11]), .B(n612), .Y(N961) );
  AND2X1 U727 ( .A(pos_dacis[12]), .B(n612), .Y(N962) );
  AND2X1 U728 ( .A(pos_dacis[3]), .B(n612), .Y(N953) );
  AND2X1 U729 ( .A(pos_dacis[8]), .B(n612), .Y(N958) );
  AND2X1 U730 ( .A(pos_dacis[17]), .B(n8), .Y(N967) );
  AND2X1 U731 ( .A(pos_dacis[15]), .B(n8), .Y(N965) );
  AND2X1 U732 ( .A(pos_dacis[16]), .B(n8), .Y(N966) );
  AND2X1 U733 ( .A(pos_dacis[14]), .B(n8), .Y(N964) );
  AND2X1 U734 ( .A(pos_dacis[13]), .B(n8), .Y(N963) );
  AND2XL U735 ( .A(pos_dacis[0]), .B(n612), .Y(N950) );
  AND2XL U736 ( .A(pos_dacis[1]), .B(n612), .Y(N951) );
  AND2X1 U737 ( .A(pos_dacis[5]), .B(n8), .Y(N955) );
  AND2X1 U738 ( .A(pos_dacis[10]), .B(n8), .Y(N960) );
  AND2X1 U739 ( .A(pos_dacis[9]), .B(n8), .Y(N959) );
  NAND4X1 U740 ( .A(srstz), .B(n670), .C(n663), .D(n662), .Y(n658) );
  NAND31X1 U741 ( .C(pos_dacis[5]), .A(n622), .B(n621), .Y(n623) );
  NOR32XL U742 ( .B(n629), .C(n628), .A(n627), .Y(sh_hold) );
  INVX1 U743 ( .A(pos_dacis[8]), .Y(n629) );
  NOR21XL U744 ( .B(n620), .A(n619), .Y(n628) );
  NAND31X1 U745 ( .C(n626), .A(n625), .B(n624), .Y(n627) );
  OR3XL U746 ( .A(pos_dacis[10]), .B(pos_dacis[12]), .C(pos_dacis[11]), .Y(
        n626) );
  OR2X1 U747 ( .A(pos_dacis[9]), .B(pos_dacis[6]), .Y(n619) );
  NOR6XL U748 ( .A(pos_dacis[15]), .B(pos_dacis[13]), .C(pos_dacis[16]), .D(
        pos_dacis[14]), .E(pos_dacis[17]), .F(pos_dacis[0]), .Y(n625) );
  INVX1 U749 ( .A(pos_dacis[4]), .Y(n622) );
  INVX1 U750 ( .A(pos_dacis[3]), .Y(n621) );
  INVX1 U751 ( .A(pos_dacis[7]), .Y(n620) );
  NAND21X1 U752 ( .B(cs_ptr[2]), .A(n49), .Y(n295) );
  NAND21X1 U753 ( .B(cs_ptr[2]), .A(cs_ptr[1]), .Y(n289) );
  AO21X1 U754 ( .B(n44), .C(cs_ptr[2]), .A(n677), .Y(n448) );
  MUX2BXL U755 ( .D0(n66), .D1(n409), .S(n44), .Y(n367) );
  AOI21X1 U756 ( .B(n65), .C(n706), .A(n408), .Y(n66) );
  OAI21BBX1 U757 ( .A(r_dac_en[16]), .B(N1312), .C(n410), .Y(n409) );
  OAI21BBX1 U758 ( .A(r_dac_en[17]), .B(N1312), .C(n417), .Y(n408) );
  INVX1 U759 ( .A(cs_ptr[2]), .Y(n601) );
  OAI32X1 U760 ( .A(n411), .B(r_dac_en[8]), .C(n735), .D(n277), .E(n412), .Y(
        n410) );
  OAI22X1 U761 ( .A(n706), .B(n416), .C(n705), .D(n246), .Y(n411) );
  OAI22X1 U762 ( .A(n706), .B(n414), .C(n415), .D(n734), .Y(n412) );
  AOI21X1 U763 ( .B(r_dac_en[14]), .C(n341), .A(r_dac_en[12]), .Y(n416) );
  INVX1 U764 ( .A(n768), .Y(n54) );
  INVX1 U765 ( .A(n770), .Y(n49) );
  AOI32X1 U766 ( .A(r_dac_en[0]), .B(n736), .C(n705), .D(r_dac_en[2]), .E(n341), .Y(n415) );
  NAND21X1 U767 ( .B(n48), .A(cs_ptr[2]), .Y(n439) );
  GEN2XL U768 ( .D(n228), .E(n729), .C(n705), .B(n418), .A(n706), .Y(n417) );
  OAI21X1 U769 ( .B(r_dac_en[5]), .C(r_dac_en[13]), .A(n705), .Y(n418) );
  BUFX3 U770 ( .A(n769), .Y(n41) );
  AOI21X1 U771 ( .B(r_dac_en[6]), .C(n341), .A(r_dac_en[4]), .Y(n414) );
  AOI31X1 U772 ( .A(n713), .B(n137), .C(n488), .D(n276), .Y(n487) );
  AOI31X1 U773 ( .A(r_dac_en[0]), .B(n741), .C(n485), .D(r_dac_en[2]), .Y(n488) );
  AOI31X1 U774 ( .A(n133), .B(n729), .C(n484), .D(n276), .Y(n483) );
  AOI31X1 U775 ( .A(r_dac_en[1]), .B(n741), .C(n485), .D(r_dac_en[3]), .Y(n484) );
  OAI21AX1 U776 ( .B(n422), .C(n341), .A(n419), .Y(n65) );
  AOI21X1 U777 ( .B(n723), .C(n714), .A(n705), .Y(n419) );
  AOI31X1 U778 ( .A(n735), .B(n736), .C(r_dac_en[1]), .D(r_dac_en[9]), .Y(n422) );
  INVX1 U779 ( .A(n771), .Y(n46) );
  MUX2X1 U780 ( .D0(n287), .D1(n54), .S(n7), .Y(n288) );
  AOI32X1 U781 ( .A(n743), .B(r_dac_en[1]), .C(n571), .D(n572), .E(r_dac_en[3]), .Y(n576) );
  OR2X1 U782 ( .A(n703), .B(n38), .Y(n150) );
  MUX2IX1 U783 ( .D0(n55), .D1(n393), .S(cs_ptr[2]), .Y(n38) );
  NAND21X1 U784 ( .B(n292), .A(n291), .Y(n299) );
  INVX1 U785 ( .A(n289), .Y(n292) );
  MUX2X1 U786 ( .D0(n439), .D1(n7), .S(n290), .Y(n291) );
  INVX1 U787 ( .A(n433), .Y(n290) );
  MUX2X1 U788 ( .D0(n568), .D1(n574), .S(cs_ptr[0]), .Y(n144) );
  AO2222XL U789 ( .A(n567), .B(r_dac_en[12]), .C(n571), .D(r_dac_en[4]), .E(
        n573), .F(r_dac_en[14]), .G(n572), .H(r_dac_en[6]), .Y(n568) );
  AO2222XL U790 ( .A(n567), .B(r_dac_en[13]), .C(n571), .D(r_dac_en[5]), .E(
        n573), .F(r_dac_en[15]), .G(n572), .H(r_dac_en[7]), .Y(n574) );
  AOI32X1 U791 ( .A(n743), .B(r_dac_en[0]), .C(n571), .D(n572), .E(r_dac_en[2]), .Y(n570) );
  NOR21XL U792 ( .B(n289), .A(n153), .Y(n309) );
  MUX2IX1 U793 ( .D0(n439), .D1(n7), .S(n542), .Y(n153) );
  NAND21X1 U794 ( .B(r_dac_en[11]), .A(n246), .Y(n322) );
  INVX1 U795 ( .A(r_dac_en[10]), .Y(n246) );
  INVX1 U796 ( .A(r_dac_en[1]), .Y(n136) );
  INVX1 U797 ( .A(r_dac_en[0]), .Y(n135) );
  AO21X1 U798 ( .B(r_dac_en[5]), .C(n44), .A(r_dac_en[4]), .Y(n728) );
  AO21X1 U799 ( .B(r_dac_en[15]), .C(n771), .A(r_dac_en[14]), .Y(n721) );
  AO21X1 U800 ( .B(n44), .C(r_dac_en[7]), .A(r_dac_en[6]), .Y(n727) );
  INVX1 U801 ( .A(r_dac_en[15]), .Y(n228) );
  INVX1 U802 ( .A(r_dac_en[6]), .Y(n137) );
  INVX1 U803 ( .A(r_dac_en[8]), .Y(n128) );
  INVX1 U804 ( .A(r_dac_en[9]), .Y(n247) );
  INVX1 U805 ( .A(r_dac_en[3]), .Y(n714) );
  INVX1 U806 ( .A(r_dac_en[5]), .Y(n133) );
  INVX1 U807 ( .A(r_dac_en[12]), .Y(n239) );
  INVX1 U808 ( .A(r_dac_en[11]), .Y(n723) );
  INVX1 U809 ( .A(r_dac_en[7]), .Y(n729) );
  INVX1 U810 ( .A(r_dac_en[13]), .Y(n230) );
  INVX1 U811 ( .A(r_dac_en[2]), .Y(n255) );
  INVX1 U812 ( .A(r_dac_en[14]), .Y(n126) );
  INVX1 U813 ( .A(r_dac_en[4]), .Y(n713) );
  NAND32X1 U814 ( .B(r_dac_en[13]), .C(r_dac_en[9]), .A(n228), .Y(n482) );
  OR3XL U815 ( .A(r_dac_en[14]), .B(r_dac_en[8]), .C(r_dac_en[12]), .Y(n486)
         );
  INVX1 U816 ( .A(r_dac_en[17]), .Y(n223) );
  INVX1 U817 ( .A(r_dac_en[16]), .Y(n67) );
  NAND21X1 U818 ( .B(n373), .A(sampl_begn), .Y(n389) );
  INVX1 U819 ( .A(r_comp_swtch), .Y(n442) );
  NAND32XL U820 ( .B(wr_dacv[11]), .C(n342), .A(n329), .Y(n343) );
  NAND32XL U821 ( .B(wr_dacv[11]), .C(n241), .A(n723), .Y(n245) );
  INVXL U822 ( .A(wr_dacv[11]), .Y(n131) );
  AND2XL U823 ( .A(n609), .B(ps_ptr[4]), .Y(N999) );
  NAND21XL U824 ( .B(ps_ptr[4]), .A(n52), .Y(n604) );
  INVX1 U825 ( .A(wr_dacv[10]), .Y(n329) );
  INVXL U826 ( .A(n256), .Y(n507) );
  NAND32X1 U827 ( .B(n39), .C(wr_dacv[0]), .A(n135), .Y(n256) );
  NAND32X1 U828 ( .B(n256), .C(n537), .A(n506), .Y(n316) );
  AND2XL U829 ( .A(n609), .B(ps_ptr[2]), .Y(N997) );
  GEN2XL U830 ( .D(ps_ptr[2]), .E(n601), .C(n600), .B(n599), .A(n598), .Y(n603) );
  INVXL U831 ( .A(ps_ptr[4]), .Y(n597) );
  NAND32XL U832 ( .B(n184), .C(n183), .A(n23), .Y(n606) );
  NAND32XL U833 ( .B(n123), .C(n184), .A(n23), .Y(n505) );
  NAND32XL U834 ( .B(n125), .C(n184), .A(n124), .Y(n360) );
  OA22X1 U835 ( .A(n357), .B(n504), .C(n356), .D(n505), .Y(n358) );
  OAI211XL U836 ( .C(n259), .D(n1), .A(n505), .B(n504), .Y(n280) );
  OA22XL U837 ( .A(n219), .B(n504), .C(n218), .D(n505), .Y(n220) );
  OAI31XL U838 ( .A(n608), .B(n607), .C(n1), .D(n605), .Y(n610) );
  AOI21XL U839 ( .B(n522), .C(n521), .A(n1), .Y(n525) );
  INVX3 U840 ( .A(auto_start), .Y(n90) );
  OAI31XL U841 ( .A(semi_start), .B(mxcyc_done), .C(auto_start), .D(n611), .Y(
        n56) );
  NAND21XL U842 ( .B(wr_dacv[14]), .A(n126), .Y(n236) );
  OA222X1 U843 ( .A(n29), .B(n360), .C(n318), .D(n1), .E(n317), .F(n316), .Y(
        n319) );
  INVX8 U844 ( .A(srstz), .Y(n373) );
  NAND21X4 U845 ( .B(r_semi), .A(n90), .Y(n184) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_LOW_shmux_00000005_00000012_00000012 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLNXL latch ( .CKN(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dac2sar_a0 ( r_dac_t, r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, 
        auto_sar, busy, stop, sync_i, sampl_begn, sampl_done, sh_rst, 
        dacyc_done, sacyc_done, ps_sample, dac_v, rpt_v, clk, srstz, test_si2, 
        test_si1, test_so1, test_se );
  input [1:0] r_dac_t;
  output [9:0] dac_v;
  output [9:0] rpt_v;
  input r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, auto_sar, busy, stop,
         sync_i, clk, srstz, test_si2, test_si1, test_se;
  output sampl_begn, sampl_done, sh_rst, dacyc_done, sacyc_done, ps_sample,
         test_so1;
  wire   N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N71, N72, N73, N74, N75, N79, updlo, updup, upd1v, r_lt_up_8_,
         r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, r_lt_up_3_,
         r_lt_up_2_, r_lt_up_1_, r_lt_up_0_, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102,
         net10260, net10266, n128, n21, n22, n23, n24, n11, n17, n18, n19, n20,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n58, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n104,
         n105, n106, n1, n2, n4, n5, n6, n10, n12, n13, n14, n15, n16, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3;
  wire   [3:0] sarcyc;
  wire   [6:0] dacnt;
  wire   [9:0] r_lt_lo;
  wire   [9:0] r_avg00;
  wire   [9:0] r_avgup;
  wire   [9:0] r_dacvo;

  INVX1 U29 ( .A(n24), .Y(n22) );
  INVX1 U30 ( .A(n24), .Y(n23) );
  INVX1 U31 ( .A(srstz), .Y(n24) );
  INVX1 U32 ( .A(n24), .Y(n21) );
  glreg_WIDTH10_2 u0_dac1v ( .clk(clk), .arstz(n23), .we(upd1v), .wdat(r_dacvo), .rdat({dac_v[9:1], n128}), .test_si(sarcyc[3]), .test_se(test_se) );
  glreg_WIDTH10_1 u0_lt_lo ( .clk(clk), .arstz(n22), .we(updlo), .wdat({n1, 
        n117, n12, n14, n116, n13, n16, n15, n10, n40}), .rdat(r_lt_lo), 
        .test_si(dac_v[9]), .test_se(test_se) );
  glreg_WIDTH10_0 u0_lt_up ( .clk(clk), .arstz(n21), .we(updup), .wdat(r_avgup), .rdat({test_so1, r_lt_up_8_, r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, 
        r_lt_up_3_, r_lt_up_2_, r_lt_up_1_, r_lt_up_0_}), .test_si(r_lt_lo[9]), 
        .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 clk_gate_dacnt_reg ( .CLK(clk), .EN(N54), 
        .ENCLK(net10260), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 clk_gate_sarcyc_reg ( .CLK(clk), .EN(N71), 
        .ENCLK(net10266), .TE(test_se) );
  dac2sar_a0_DW01_add_0 add_312 ( .A({1'b0, n11, n19, n20, n27, n29, n31, n33, 
        n35, n37, n39}), .B({1'b0, n17, n18, n25, n26, n28, n30, n32, n34, n36, 
        n38}), .CI(1'b0), .SUM({N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, SYNOPSYS_UNCONNECTED_1}), .CO() );
  dac2sar_a0_DW01_add_2 add_305 ( .A({1'b0, r_lt_lo}), .B({1'b0, test_so1, 
        r_lt_up_8_, r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, r_lt_up_3_, 
        r_lt_up_2_, r_lt_up_1_, r_lt_up_0_}), .CI(1'b0), .SUM({r_avg00, 
        SYNOPSYS_UNCONNECTED_2}), .CO() );
  dac2sar_a0_DW01_inc_0 add_285 ( .A(dacnt), .SUM({N53, N52, N51, N50, N49, 
        N48, N47}) );
  dac2sar_a0_DW01_add_1 add_310 ( .A({1'b0, n1, n117, n12, n14, n48, n13, n16, 
        n15, n10, n40}), .B({1'b0, r_avgup}), .CI(1'b0), .SUM({N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, SYNOPSYS_UNCONNECTED_3}), .CO() );
  SDFFQX1 dacnt_reg_1_ ( .D(N56), .SIN(dacnt[0]), .SMC(test_se), .C(net10260), 
        .Q(dacnt[1]) );
  SDFFQX1 sarcyc_reg_1_ ( .D(N73), .SIN(sarcyc[0]), .SMC(test_se), .C(net10266), .Q(sarcyc[1]) );
  SDFFQX1 sarcyc_reg_0_ ( .D(N72), .SIN(dacnt[6]), .SMC(test_se), .C(net10266), 
        .Q(sarcyc[0]) );
  SDFFQX1 sarcyc_reg_3_ ( .D(N75), .SIN(sarcyc[2]), .SMC(test_se), .C(net10266), .Q(sarcyc[3]) );
  SDFFQX1 dacnt_reg_5_ ( .D(N60), .SIN(dacnt[4]), .SMC(test_se), .C(net10260), 
        .Q(dacnt[5]) );
  SDFFQX1 sarcyc_reg_2_ ( .D(N74), .SIN(sarcyc[1]), .SMC(test_se), .C(net10266), .Q(sarcyc[2]) );
  SDFFQX1 dacnt_reg_4_ ( .D(N59), .SIN(dacnt[3]), .SMC(test_se), .C(net10260), 
        .Q(dacnt[4]) );
  SDFFQX1 dacnt_reg_0_ ( .D(N55), .SIN(test_si2), .SMC(test_se), .C(net10260), 
        .Q(dacnt[0]) );
  SDFFQX1 dacnt_reg_3_ ( .D(N58), .SIN(dacnt[2]), .SMC(test_se), .C(net10260), 
        .Q(dacnt[3]) );
  SDFFQX1 dacnt_reg_6_ ( .D(N61), .SIN(dacnt[5]), .SMC(test_se), .C(net10260), 
        .Q(dacnt[6]) );
  SDFFQX1 dacnt_reg_2_ ( .D(N57), .SIN(dacnt[1]), .SMC(test_se), .C(net10260), 
        .Q(dacnt[2]) );
  SDFFNQX1 sh_rst_n_reg ( .D(N79), .SIN(test_si1), .SMC(test_se), .XC(clk), 
        .Q(sh_rst) );
  NAND21X1 U6 ( .B(n28), .A(n92), .Y(r_avgup[5]) );
  INVX3 U7 ( .A(sar_ini), .Y(n92) );
  NAND2X1 U8 ( .A(n120), .B(n92), .Y(r_avgup[2]) );
  NAND2X1 U9 ( .A(n121), .B(n92), .Y(r_avgup[3]) );
  NAND21X1 U10 ( .B(n26), .A(n92), .Y(r_avgup[6]) );
  MUX2X1 U11 ( .D0(N89), .D1(r_avg00[7]), .S(n5), .Y(r_dacvo[7]) );
  MUX2X1 U12 ( .D0(N91), .D1(r_avg00[9]), .S(semi_nxt), .Y(r_dacvo[9]) );
  NOR2X1 U13 ( .A(n6), .B(n73), .Y(n1) );
  INVXL U14 ( .A(n128), .Y(n2) );
  INVXL U15 ( .A(n2), .Y(dac_v[0]) );
  INVXL U16 ( .A(n2), .Y(n4) );
  BUFX3 U17 ( .A(semi_nxt), .Y(n5) );
  MUX2X1 U18 ( .D0(N88), .D1(r_avg00[6]), .S(semi_nxt), .Y(r_dacvo[6]) );
  MUX2X1 U19 ( .D0(N87), .D1(r_avg00[5]), .S(semi_nxt), .Y(r_dacvo[5]) );
  MUX2X1 U20 ( .D0(N86), .D1(r_avg00[4]), .S(semi_nxt), .Y(r_dacvo[4]) );
  BUFX3 U21 ( .A(sar_ini), .Y(n6) );
  NAND2XL U22 ( .A(n119), .B(n92), .Y(r_avgup[1]) );
  NAND21X1 U23 ( .B(sar_ini), .A(n29), .Y(n99) );
  NAND2X1 U24 ( .A(n122), .B(n92), .Y(r_avgup[4]) );
  NOR2XL U25 ( .A(sar_ini), .B(n79), .Y(n16) );
  NOR2XL U26 ( .A(sar_ini), .B(n76), .Y(n14) );
  MUX2X2 U27 ( .D0(N90), .D1(r_avg00[8]), .S(n5), .Y(r_dacvo[8]) );
  NOR2XL U28 ( .A(sar_ini), .B(n80), .Y(n15) );
  NOR2XL U33 ( .A(sar_ini), .B(n78), .Y(n13) );
  NAND2XL U34 ( .A(n118), .B(n92), .Y(r_avgup[0]) );
  NAND2XL U35 ( .A(n127), .B(n92), .Y(r_avgup[9]) );
  INVXL U36 ( .A(n95), .Y(n117) );
  INVX1 U37 ( .A(n99), .Y(n48) );
  OR3XL U38 ( .A(sar_nxt), .B(n6), .C(semi_nxt), .Y(upd1v) );
  INVX1 U39 ( .A(n85), .Y(n89) );
  INVX1 U40 ( .A(n84), .Y(n69) );
  OR2X1 U41 ( .A(n89), .B(n88), .Y(N71) );
  INVX1 U42 ( .A(n90), .Y(n61) );
  NAND2XL U43 ( .A(n126), .B(n92), .Y(r_avgup[8]) );
  MUX2X1 U44 ( .D0(N83), .D1(r_avg00[1]), .S(semi_nxt), .Y(r_dacvo[1]) );
  MUX2X1 U45 ( .D0(N85), .D1(r_avg00[3]), .S(semi_nxt), .Y(r_dacvo[3]) );
  MUX2X1 U46 ( .D0(N84), .D1(r_avg00[2]), .S(semi_nxt), .Y(r_dacvo[2]) );
  NOR2XL U47 ( .A(sar_ini), .B(n81), .Y(n10) );
  NOR2XL U48 ( .A(n6), .B(n75), .Y(n12) );
  NOR2XL U49 ( .A(sar_ini), .B(n82), .Y(n40) );
  OR2X1 U50 ( .A(sacyc_done), .B(n91), .Y(n88) );
  NAND21X1 U51 ( .B(n71), .A(n89), .Y(n84) );
  NAND32X1 U52 ( .B(n67), .C(n88), .A(auto_sar), .Y(n85) );
  AND2X1 U53 ( .A(n69), .B(n68), .Y(N73) );
  AND2X1 U54 ( .A(n89), .B(n87), .Y(N72) );
  NAND32X1 U55 ( .B(n60), .C(n91), .A(n67), .Y(n90) );
  INVX1 U56 ( .A(busy), .Y(n60) );
  NAND32X1 U57 ( .B(dacyc_done), .C(n91), .A(n90), .Y(N54) );
  AND2X1 U58 ( .A(N50), .B(n61), .Y(N58) );
  AND2X1 U59 ( .A(N52), .B(n61), .Y(N60) );
  AND2X1 U60 ( .A(N51), .B(n61), .Y(N59) );
  AND2X1 U61 ( .A(N49), .B(n61), .Y(N57) );
  AND2X1 U62 ( .A(N48), .B(n61), .Y(N56) );
  NAND21X1 U63 ( .B(n104), .A(n105), .Y(n58) );
  XNOR2XL U64 ( .A(n113), .B(n105), .Y(n41) );
  XOR2X1 U65 ( .A(n54), .B(n106), .Y(n42) );
  AND3X1 U66 ( .A(busy), .B(n44), .C(n115), .Y(N79) );
  INVX1 U67 ( .A(n80), .Y(n35) );
  INVX1 U68 ( .A(n120), .Y(n34) );
  INVX1 U69 ( .A(n79), .Y(n33) );
  INVX1 U70 ( .A(n121), .Y(n32) );
  INVX1 U71 ( .A(n78), .Y(n31) );
  INVX1 U72 ( .A(n122), .Y(n30) );
  INVX1 U73 ( .A(n77), .Y(n29) );
  INVX1 U74 ( .A(n123), .Y(n28) );
  INVX1 U75 ( .A(n76), .Y(n27) );
  INVX1 U76 ( .A(n124), .Y(n26) );
  INVX1 U77 ( .A(n125), .Y(n25) );
  INVX1 U78 ( .A(n75), .Y(n20) );
  INVX1 U79 ( .A(n126), .Y(n18) );
  INVX1 U80 ( .A(n74), .Y(n19) );
  INVX1 U81 ( .A(n119), .Y(n36) );
  INVX1 U82 ( .A(n81), .Y(n37) );
  INVX1 U83 ( .A(n73), .Y(n11) );
  INVX1 U84 ( .A(n127), .Y(n17) );
  INVX1 U85 ( .A(r_avg00[9]), .Y(n93) );
  INVX1 U86 ( .A(r_avg00[8]), .Y(n94) );
  INVX1 U87 ( .A(r_avg00[3]), .Y(n101) );
  INVX1 U88 ( .A(r_avg00[4]), .Y(n100) );
  INVX1 U89 ( .A(r_avg00[5]), .Y(n98) );
  INVX1 U90 ( .A(r_avg00[6]), .Y(n97) );
  INVX1 U91 ( .A(r_avg00[7]), .Y(n96) );
  INVX1 U92 ( .A(r_avg00[2]), .Y(n102) );
  INVX1 U93 ( .A(r_avg00[1]), .Y(n103) );
  INVX1 U94 ( .A(r_avg00[0]), .Y(n107) );
  INVX1 U95 ( .A(n51), .Y(n50) );
  INVX1 U96 ( .A(n51), .Y(n49) );
  INVX1 U97 ( .A(n67), .Y(dacyc_done) );
  INVX1 U98 ( .A(n118), .Y(n38) );
  INVX1 U99 ( .A(n82), .Y(n39) );
  NAND21XL U100 ( .B(stop), .A(n23), .Y(n91) );
  ENOX1 U101 ( .A(dac_v[0]), .B(n125), .C(N100), .D(n4), .Y(rpt_v[7]) );
  ENOX1 U102 ( .A(n4), .B(n122), .C(N97), .D(n4), .Y(rpt_v[4]) );
  ENOX1 U103 ( .A(n4), .B(n123), .C(N98), .D(dac_v[0]), .Y(rpt_v[5]) );
  MUX2X1 U104 ( .D0(n70), .D1(n69), .S(sarcyc[2]), .Y(N74) );
  AND2X1 U105 ( .A(n71), .B(n89), .Y(n70) );
  ENOX1 U106 ( .A(dac_v[0]), .B(n121), .C(N96), .D(n4), .Y(rpt_v[3]) );
  ENOX1 U107 ( .A(n4), .B(n124), .C(N99), .D(n4), .Y(rpt_v[6]) );
  ENOX1 U108 ( .A(n128), .B(n126), .C(N101), .D(dac_v[0]), .Y(rpt_v[8]) );
  ENOX1 U109 ( .A(dac_v[0]), .B(n127), .C(dac_v[0]), .D(N102), .Y(rpt_v[9]) );
  OAI22X1 U110 ( .A(n86), .B(n85), .C(n84), .D(n83), .Y(N75) );
  MUX2BXL U111 ( .D0(n83), .D1(n72), .S(sarcyc[2]), .Y(n86) );
  AND2X1 U112 ( .A(n71), .B(n83), .Y(n72) );
  INVX1 U113 ( .A(sarcyc[3]), .Y(n83) );
  ENOX1 U114 ( .A(dac_v[0]), .B(n120), .C(N95), .D(n4), .Y(rpt_v[2]) );
  ENOX1 U115 ( .A(n4), .B(n119), .C(N94), .D(n4), .Y(rpt_v[1]) );
  AND2X1 U116 ( .A(N47), .B(n61), .Y(N55) );
  AND2X1 U117 ( .A(N53), .B(n61), .Y(N61) );
  ENOX1 U118 ( .A(n128), .B(n118), .C(N93), .D(n128), .Y(rpt_v[0]) );
  AOI21BBXL U119 ( .B(r_dac_t[0]), .C(n104), .A(n106), .Y(n105) );
  AND4X1 U120 ( .A(n111), .B(n115), .C(n110), .D(n109), .Y(sampl_done) );
  XOR2X1 U121 ( .A(n112), .B(n58), .Y(n110) );
  AND4X1 U122 ( .A(dacnt[1]), .B(n42), .C(n108), .D(n41), .Y(n109) );
  XOR2X1 U123 ( .A(n58), .B(dacnt[6]), .Y(n108) );
  NOR2X1 U124 ( .A(r_dac_t[1]), .B(n104), .Y(n106) );
  XOR2X1 U125 ( .A(dacnt[4]), .B(n43), .Y(n111) );
  OA21X1 U126 ( .B(r_dac_t[0]), .C(n104), .A(n58), .Y(n43) );
  NOR2X1 U127 ( .A(r_dac_t[0]), .B(r_dac_t[1]), .Y(n104) );
  INVX1 U128 ( .A(dacnt[3]), .Y(n113) );
  INVX1 U129 ( .A(dacnt[2]), .Y(n54) );
  NAND21X1 U130 ( .B(sarcyc[1]), .A(n87), .Y(n68) );
  NOR4XL U131 ( .A(dacnt[4]), .B(dacnt[2]), .C(dacnt[1]), .D(n45), .Y(n44) );
  NAND4X1 U132 ( .A(n46), .B(n114), .C(n113), .D(n112), .Y(n45) );
  NOR3XL U133 ( .A(sarcyc[3]), .B(n68), .C(sarcyc[2]), .Y(n46) );
  INVX1 U134 ( .A(dacnt[0]), .Y(n115) );
  INVX1 U135 ( .A(sarcyc[0]), .Y(n87) );
  INVX1 U136 ( .A(dacnt[5]), .Y(n112) );
  INVX1 U137 ( .A(dacnt[6]), .Y(n114) );
  MUX2AXL U138 ( .D0(r_lt_lo[1]), .D1(n103), .S(n49), .Y(n81) );
  MUX2BXL U139 ( .D0(n96), .D1(r_lt_up_7_), .S(n50), .Y(n125) );
  MUX2BXL U140 ( .D0(n102), .D1(r_lt_up_2_), .S(n50), .Y(n120) );
  MUX2BXL U141 ( .D0(n101), .D1(r_lt_up_3_), .S(n50), .Y(n121) );
  MUX2BXL U142 ( .D0(n100), .D1(r_lt_up_4_), .S(n50), .Y(n122) );
  MUX2BXL U143 ( .D0(n98), .D1(r_lt_up_5_), .S(n50), .Y(n123) );
  MUX2BXL U144 ( .D0(n97), .D1(r_lt_up_6_), .S(n50), .Y(n124) );
  MUX2BXL U145 ( .D0(n94), .D1(r_lt_up_8_), .S(n50), .Y(n126) );
  MUX2BXL U146 ( .D0(n93), .D1(test_so1), .S(n49), .Y(n127) );
  MUX2BXL U147 ( .D0(n103), .D1(r_lt_up_1_), .S(n50), .Y(n119) );
  MUX2AXL U148 ( .D0(r_lt_lo[2]), .D1(n102), .S(n49), .Y(n80) );
  MUX2AXL U149 ( .D0(r_lt_lo[3]), .D1(n101), .S(n49), .Y(n79) );
  MUX2AXL U150 ( .D0(r_lt_lo[4]), .D1(n100), .S(n49), .Y(n78) );
  MUX2AXL U151 ( .D0(r_lt_lo[5]), .D1(n98), .S(n49), .Y(n77) );
  MUX2AXL U152 ( .D0(r_lt_lo[6]), .D1(n97), .S(n49), .Y(n76) );
  MUX2AXL U153 ( .D0(r_lt_lo[7]), .D1(n96), .S(n49), .Y(n75) );
  MUX2AXL U154 ( .D0(r_lt_lo[8]), .D1(n94), .S(n49), .Y(n74) );
  NOR43XL U155 ( .B(n66), .C(n65), .D(n64), .A(n63), .Y(sacyc_done) );
  XOR2X1 U156 ( .A(sarcyc[3]), .B(r_sar10), .Y(n63) );
  XOR2X1 U157 ( .A(r_sar10), .B(sarcyc[1]), .Y(n66) );
  XOR2X1 U158 ( .A(r_sar10), .B(sarcyc[2]), .Y(n65) );
  MUX2BXL U159 ( .D0(n107), .D1(r_lt_up_0_), .S(n50), .Y(n118) );
  MUX2AXL U160 ( .D0(r_lt_lo[0]), .D1(n107), .S(n50), .Y(n82) );
  MUX2AXL U161 ( .D0(r_lt_lo[9]), .D1(n93), .S(n49), .Y(n73) );
  OAI211X1 U162 ( .C(n114), .D(n112), .A(n59), .B(n57), .Y(n67) );
  AND2X1 U163 ( .A(dacnt[1]), .B(dacnt[0]), .Y(n57) );
  MUX2X1 U164 ( .D0(n56), .D1(n55), .S(n46), .Y(n59) );
  AND4X1 U165 ( .A(n53), .B(n52), .C(n114), .D(n112), .Y(n56) );
  NOR43XL U166 ( .B(n41), .C(n42), .D(n111), .A(n47), .Y(n55) );
  MUX2IX1 U167 ( .D0(dacnt[6]), .D1(dacnt[5]), .S(n58), .Y(n47) );
  AND2X1 U168 ( .A(sarcyc[0]), .B(dacyc_done), .Y(n64) );
  INVX1 U169 ( .A(sync_i), .Y(n51) );
  MUX2X1 U170 ( .D0(n54), .D1(n113), .S(dacnt[4]), .Y(n53) );
  MUX2X1 U171 ( .D0(dacnt[3]), .D1(dacnt[2]), .S(r_dacyc), .Y(n52) );
  AND2X1 U172 ( .A(dacnt[0]), .B(n44), .Y(sampl_begn) );
  INVX1 U173 ( .A(n62), .Y(n71) );
  NAND21X1 U174 ( .B(n87), .A(sarcyc[1]), .Y(n62) );
  NAND21X1 U175 ( .B(n25), .A(n92), .Y(r_avgup[7]) );
  AO21XL U176 ( .B(sar_nxt), .C(sync_i), .A(n6), .Y(updlo) );
  AO21XL U177 ( .B(sar_nxt), .C(n51), .A(n6), .Y(updup) );
  NAND21XL U178 ( .B(n6), .A(n19), .Y(n95) );
  INVXL U179 ( .A(n99), .Y(n116) );
  MUX2X1 U180 ( .D0(N82), .D1(r_avg00[0]), .S(semi_nxt), .Y(r_dacvo[0]) );
endmodule


module dac2sar_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n7, n8, n10, n18, n19, n21, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n37, n38, n39, n40, n41, n42,
         n45, n46, n49, n50, n51, n52, n53, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n68, n69, n70, n71, n72, n73, n74, n113, n114,
         n115, n116, n117, n118, n119, n120, n121;

  OAI21X1 U23 ( .B(n53), .C(n25), .A(n26), .Y(n24) );
  OAI21X1 U27 ( .B(n29), .C(n37), .A(n30), .Y(n28) );
  NOR2X1 U34 ( .A(n41), .B(n34), .Y(n32) );
  OAI21X1 U35 ( .B(n42), .C(n34), .A(n37), .Y(n33) );
  OAI21X1 U49 ( .B(n45), .C(n51), .A(n46), .Y(n40) );
  OAI21X1 U66 ( .B(n56), .C(n60), .A(n57), .Y(n55) );
  XOR2X1 U71 ( .A(n61), .B(n8), .Y(SUM[2]) );
  OAI21X1 U72 ( .B(n61), .C(n59), .A(n60), .Y(n58) );
  NOR2XL U88 ( .A(n34), .B(n29), .Y(n27) );
  NOR2X1 U89 ( .A(A[3]), .B(B[3]), .Y(n56) );
  NOR2X1 U90 ( .A(A[7]), .B(B[7]), .Y(n29) );
  NOR2X1 U91 ( .A(A[6]), .B(B[6]), .Y(n34) );
  NOR2X1 U92 ( .A(A[2]), .B(B[2]), .Y(n59) );
  XNOR2XL U93 ( .A(n115), .B(n119), .Y(SUM[5]) );
  OAI21BBX1 U94 ( .A(n118), .B(n21), .C(n18), .Y(n113) );
  AND2X1 U95 ( .A(n117), .B(n118), .Y(n114) );
  AOI21X1 U96 ( .B(n24), .C(n117), .A(n21), .Y(n19) );
  NAND2X1 U97 ( .A(A[5]), .B(B[5]), .Y(n46) );
  NOR2X1 U98 ( .A(A[5]), .B(B[5]), .Y(n45) );
  NAND2XL U99 ( .A(A[3]), .B(B[3]), .Y(n57) );
  NAND2X1 U100 ( .A(A[2]), .B(B[2]), .Y(n60) );
  AOI21XL U101 ( .B(n27), .C(n40), .A(n28), .Y(n26) );
  INVXL U102 ( .A(n50), .Y(n71) );
  INVXL U103 ( .A(n34), .Y(n69) );
  NAND2X1 U104 ( .A(A[6]), .B(B[6]), .Y(n37) );
  NAND2XL U105 ( .A(A[8]), .B(B[8]), .Y(n23) );
  OR2X2 U106 ( .A(A[9]), .B(B[9]), .Y(n118) );
  NAND2XL U107 ( .A(A[9]), .B(B[9]), .Y(n18) );
  AOI21X1 U108 ( .B(n52), .C(n71), .A(n49), .Y(n115) );
  AOI21BX1 U109 ( .C(n116), .B(n62), .A(n55), .Y(n53) );
  OR2X1 U110 ( .A(n59), .B(n56), .Y(n116) );
  INVX1 U111 ( .A(n23), .Y(n21) );
  INVX1 U112 ( .A(n45), .Y(n70) );
  INVX1 U113 ( .A(n56), .Y(n72) );
  NOR2X1 U114 ( .A(A[4]), .B(B[4]), .Y(n50) );
  OR2X1 U115 ( .A(A[8]), .B(B[8]), .Y(n117) );
  NAND2XL U116 ( .A(A[7]), .B(B[7]), .Y(n30) );
  NOR2X1 U117 ( .A(A[1]), .B(B[1]), .Y(n63) );
  NAND2X1 U118 ( .A(A[4]), .B(B[4]), .Y(n51) );
  NAND2X1 U119 ( .A(A[0]), .B(B[0]), .Y(n65) );
  NAND2XL U120 ( .A(n117), .B(n23), .Y(n2) );
  AND2XL U121 ( .A(n70), .B(n46), .Y(n119) );
  NAND2XL U122 ( .A(n73), .B(n60), .Y(n8) );
  XNOR2XL U123 ( .A(n120), .B(n65), .Y(SUM[1]) );
  AND2X1 U124 ( .A(n74), .B(n121), .Y(n120) );
  XNOR2XL U125 ( .A(n6), .B(n52), .Y(SUM[4]) );
  XNOR2XL U126 ( .A(n7), .B(n58), .Y(SUM[3]) );
  NAND2XL U127 ( .A(n72), .B(n57), .Y(n7) );
  NAND2XL U128 ( .A(n69), .B(n37), .Y(n4) );
  NAND2XL U129 ( .A(n68), .B(n30), .Y(n3) );
  NAND2XL U130 ( .A(n118), .B(n18), .Y(n1) );
  INVX1 U131 ( .A(n53), .Y(n52) );
  NAND2XL U132 ( .A(n71), .B(n51), .Y(n6) );
  INVXL U133 ( .A(n51), .Y(n49) );
  NAND2X1 U134 ( .A(n39), .B(n27), .Y(n25) );
  INVXL U135 ( .A(n29), .Y(n68) );
  INVX1 U136 ( .A(n59), .Y(n73) );
  INVXL U137 ( .A(n40), .Y(n42) );
  XOR2XL U138 ( .A(n31), .B(n3), .Y(SUM[7]) );
  AOI21XL U139 ( .B(n52), .C(n32), .A(n33), .Y(n31) );
  XOR2XL U140 ( .A(n38), .B(n4), .Y(SUM[6]) );
  AOI21XL U141 ( .B(n52), .C(n39), .A(n40), .Y(n38) );
  AOI21XL U142 ( .B(n24), .C(n114), .A(n113), .Y(n10) );
  BUFXL U143 ( .A(n64), .Y(n121) );
  NAND2X1 U144 ( .A(A[1]), .B(B[1]), .Y(n64) );
  INVXL U145 ( .A(n62), .Y(n61) );
  INVX1 U146 ( .A(n63), .Y(n74) );
  INVXL U147 ( .A(n39), .Y(n41) );
  NOR2XL U148 ( .A(n50), .B(n45), .Y(n39) );
  OAI21X1 U149 ( .B(n63), .C(n65), .A(n64), .Y(n62) );
  XOR2XL U150 ( .A(n19), .B(n1), .Y(SUM[9]) );
  INVXL U151 ( .A(n10), .Y(SUM[10]) );
  XNOR2XL U152 ( .A(n2), .B(n24), .Y(SUM[8]) );
endmodule


module dac2sar_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module dac2sar_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module dac2sar_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10283;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10283), .TE(test_se) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10283), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10301;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10301), .TE(test_se) );
  SDFFRQXL mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10301), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10319;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10319), .TE(test_se) );
  SDFFRQXL mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[5]) );
  SDFFRQXL mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[6]) );
  SDFFRQXL mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[4]) );
  SDFFRQXL mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[9]) );
  SDFFRQXL mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[8]) );
  SDFFRQXL mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[3]) );
  SDFFRQXL mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[2]) );
  SDFFRQXL mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[0]) );
  SDFFRQXL mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10319), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_00000012 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [17:0] wdat;
  output [17:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10337, n1, n2, n3;

  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(arstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_glreg_00000012 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10337), .TE(test_se) );
  SDFFRQX1 mem_reg_14_ ( .D(wdat[14]), .SIN(rdat[13]), .SMC(test_se), .C(
        net10337), .XR(n1), .Q(rdat[14]) );
  SDFFRQX1 mem_reg_11_ ( .D(wdat[11]), .SIN(rdat[10]), .SMC(test_se), .C(
        net10337), .XR(n1), .Q(rdat[11]) );
  SDFFRQX1 mem_reg_10_ ( .D(wdat[10]), .SIN(rdat[9]), .SMC(test_se), .C(
        net10337), .XR(n1), .Q(rdat[10]) );
  SDFFRQX1 mem_reg_16_ ( .D(wdat[16]), .SIN(rdat[15]), .SMC(test_se), .C(
        net10337), .XR(n1), .Q(rdat[16]) );
  SDFFRQX1 mem_reg_17_ ( .D(wdat[17]), .SIN(rdat[16]), .SMC(test_se), .C(
        net10337), .XR(n1), .Q(rdat[17]) );
  SDFFRQX1 mem_reg_13_ ( .D(wdat[13]), .SIN(rdat[12]), .SMC(test_se), .C(
        net10337), .XR(n1), .Q(rdat[13]) );
  SDFFRQX1 mem_reg_12_ ( .D(wdat[12]), .SIN(rdat[11]), .SMC(test_se), .C(
        net10337), .XR(n1), .Q(rdat[12]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10337), .XR(n1), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10337), .XR(n1), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10337), .XR(n2), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10337), .XR(n2), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10337), .XR(n2), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10337), .XR(n2), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10337), .XR(n2), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10337), .XR(n2), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10337), .XR(n2), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10337), .XR(n2), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_15_ ( .D(wdat[15]), .SIN(rdat[14]), .SMC(test_se), .C(
        net10337), .XR(n1), .Q(rdat[15]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_00000012 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( i_cc, i_cc_49, i_sqlch, r_sqlch, 
        r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, 
        r_fiforst, r_unlock, r_first, r_last, r_set_cpmsgid, r_rdy, r_wdat, 
        r_rdat, r_txnumk, r_txendk, r_txshrt, r_auto_discard, r_txauto, 
        r_rxords_ena, r_spec, r_dat_spec, r_auto_gdcrc, r_rxdb_opt, r_pshords, 
        r_dat_portrole, r_dat_datarole, r_discard, pid_goidle, pid_gobusy, 
        pff_ack, pff_rdat, pff_rxpart, prx_rcvinf, pff_obsd, pff_ptr, 
        pff_empty, pff_full, ptx_ack, ptx_cc, ptx_oe, prx_setsta, prx_rst, 
        prl_c0set, prl_cany0, prl_cany0r, prl_cany0w, prl_discard, 
        prl_GCTxDone, prl_cany0adr, prl_cpmsgid, prx_fifowdat, ptx_fsm, 
        prl_fsm, prx_fsm, prx_adpn, dbgpo, clk, srstz, test_si, test_so, 
        test_se );
  input [1:0] r_sqlch;
  input [7:0] r_wdat;
  input [7:0] r_rdat;
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [6:0] r_rxords_ena;
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [1:0] r_auto_gdcrc;
  input [1:0] r_rxdb_opt;
  output [1:0] pff_ack;
  output [7:0] pff_rdat;
  output [15:0] pff_rxpart;
  output [4:0] prx_rcvinf;
  output [5:0] pff_ptr;
  output [6:0] prx_setsta;
  output [1:0] prx_rst;
  output [7:0] prl_cany0adr;
  output [2:0] prl_cpmsgid;
  output [7:0] prx_fifowdat;
  output [2:0] ptx_fsm;
  output [3:0] prl_fsm;
  output [3:0] prx_fsm;
  output [5:0] prx_adpn;
  output [31:0] dbgpo;
  input i_cc, i_cc_49, i_sqlch, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4,
         r_fifopsh, r_fifopop, r_fiforst, r_unlock, r_first, r_last,
         r_set_cpmsgid, r_rdy, r_txendk, r_txshrt, r_auto_discard, r_pshords,
         r_dat_portrole, r_dat_datarole, r_discard, clk, srstz, test_si,
         test_se;
  output pid_goidle, pid_gobusy, pff_obsd, pff_empty, pff_full, ptx_ack,
         ptx_cc, ptx_oe, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_discard, prl_GCTxDone, test_so;
  wire   n108, rx_pshords, auto_rx_gdcrc, prx_trans, prx_fiforst, pcc_rxgood,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd, x_trans, ptx_goidle,
         c0_txendk, mux_one, ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4,
         crcstart, crcshfi4, crcshfo4, prl_idle, lockena, fifosrstz,
         fifopop_pff, fifopsh_pff, pff_txreq, pff_one, obsd, prl_last,
         prl_txreq, fifopop_prl, fifopsh_prl, prx_gdmsgrcvd, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, d_sqlch, net10355, n61, n62, n63, n64,
         n55, n56, n57, n58, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n5, n6, n7, n10, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n59, n60, n65, n66, n67, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;
  wire   [1:0] prx_cccnt;
  wire   [3:0] prx_crcsidat;
  wire   [4:0] c0_txnumk;
  wire   [6:0] c0_txauto;
  wire   [7:0] mux_rdat;
  wire   [3:0] ptx_crcsidat;
  wire   [3:0] crc32_3_0;
  wire   [3:0] crcsidat;
  wire   [55:0] pff_dat_7_1;
  wire   [47:16] pff_c0dat;
  wire   [7:0] prl_rdat;
  wire   [4:0] prl_txauto;
  wire   [1:0] d_cc;
  wire   [8:0] cclow_cnt;

  phyrx_a0 u0_phyrx ( .i_cc(i_cc), .ptx_txact(n6), .r_adprx_en(r_adprx_en), 
        .r_adp2nd(r_adp2nd), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), 
        .r_rxdb_opt(r_rxdb_opt), .r_ords_ena(r_rxords_ena), .r_pshords(
        rx_pshords), .r_rgdcrc(auto_rx_gdcrc), .prx_cccnt(prx_cccnt), 
        .prx_rst(prx_rst), .prx_setsta({prx_setsta[6:1], 
        SYNOPSYS_UNCONNECTED_1}), .prx_idle(), .prx_d_cc(dbgpo[17]), .prx_bmc(
        dbgpo[18]), .prx_trans(prx_trans), .prx_fiforst(prx_fiforst), 
        .prx_fifopsh(dbgpo[29]), .prx_fifowdat(prx_fifowdat), .pff_txreq(n10), 
        .pid_gobusy(pid_gobusy), .pid_goidle(pid_goidle), .pid_ccidle(
        prx_rcvinf[4]), .pcc_rxgood(pcc_rxgood), .prx_crcstart(prx_crcstart), 
        .prx_crcshfi4(prx_crcshfi4), .prx_crcsidat(prx_crcsidat), .prx_rxcode(
        dbgpo[28:24]), .prx_adpn(prx_adpn), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_eoprcvd(prx_eoprcvd), .prx_fsm(prx_fsm), .clk(clk), .srstz(n35), 
        .test_si(n63), .test_so(n62), .test_se(test_se) );
  phyidd_a0 u0_phyidd ( .i_trans(x_trans), .i_goidle(ptx_goidle), .o_ccidle(
        prx_rcvinf[4]), .o_goidle(pid_goidle), .o_gobusy(pid_gobusy), .clk(clk), .srstz(srstz), .test_si(pff_ptr[5]), .test_so(n63), .test_se(test_se) );
  phytx_a0 u0_phytx ( .r_txnumk(c0_txnumk), .r_txendk(c0_txendk), .r_txshrt(
        r_txshrt), .r_txauto(c0_txauto), .prx_cccnt(prx_cccnt), .ptx_txact(
        ptx_oe), .ptx_cc(ptx_cc), .ptx_goidle(ptx_goidle), .ptx_fifopop(
        dbgpo[30]), .ptx_pspyld(), .i_rdat(mux_rdat), .i_txreq(n10), .i_one(
        mux_one), .ptx_crcstart(ptx_crcstart), .ptx_crcshfi4(ptx_crcshfi4), 
        .ptx_crcshfo4(ptx_crcshfo4), .ptx_crcsidat(ptx_crcsidat), .ptx_fsm(
        ptx_fsm), .pcc_crc30(crc32_3_0), .clk(clk), .srstz(srstz), .test_si(
        n62), .test_se(test_se) );
  phycrc_a0 u0_phycrc ( .crc32_3_0(crc32_3_0), .rx_good(pcc_rxgood), 
        .i_shfidat(crcsidat), .i_start(crcstart), .i_shfi4(crcshfi4), 
        .i_shfo4(crcshfo4), .clk(clk), .test_si(d_cc[1]), .test_so(n64), 
        .test_se(test_se) );
  phyff_DEPTH_NUM34_DEPTH_NBT6 u0_phyff ( .r_psh(r_fifopsh), .r_pop(r_fifopop), 
        .prx_psh(fifopsh_pff), .ptx_pop(fifopop_pff), .r_last(r_last), 
        .r_unlock(r_unlock), .i_lockena(lockena), .r_fiforst(r_fiforst), 
        .i_ccidle(prx_rcvinf[4]), .r_wdat(r_wdat), .prx_wdat(prx_fifowdat), 
        .txreq(pff_txreq), .ffack(pff_ack), .rdat0(pff_rdat), .full(pff_full), 
        .empty(pff_empty), .one(pff_one), .half(), .obsd(obsd), .dat_7_1(
        pff_dat_7_1), .ptr(pff_ptr), .fifowdat(dbgpo[7:0]), .fifopsh(dbgpo[16]), .clk(clk), .srstz(fifosrstz), .test_si(n64), .test_se(test_se) );
  updprl_a0 u0_updprl ( .r_spec(r_spec), .r_dat_spec(r_dat_spec), 
        .r_auto_txgdcrc(r_auto_gdcrc[0]), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_auto_discard(r_auto_discard), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_dat_cpmsgid(r_wdat[2:0]), .r_rdat(
        r_rdat), .r_rdy(r_rdy), .pid_ccidle(prx_rcvinf[4]), .r_discard(
        r_discard), .ptx_ack(ptx_goidle), .ptx_txact(n6), .ptx_fifopop(
        fifopop_prl), .prx_fifopsh(fifopsh_prl), .prx_gdmsgrcvd(prx_gdmsgrcvd), 
        .prx_eoprcvd(prx_eoprcvd), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_fifowdat(prx_fifowdat), .pff_c0dat({pff_c0dat, pff_rxpart}), 
        .prl_rdat(prl_rdat), .prl_txauto({SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, prl_txauto[4], SYNOPSYS_UNCONNECTED_4, 
        prl_txauto[2:0]}), .prl_last(prl_last), .prl_txreq(prl_txreq), 
        .prl_c0set(prl_c0set), .prl_cany0(n108), .prl_cany0r(prl_cany0r), 
        .prl_cany0w(prl_cany0w), .prl_idle(prl_idle), .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_fsm(prl_fsm), .prl_cpmsgid(prl_cpmsgid), 
        .prl_cany0adr(prl_cany0adr), .clk(clk), .srstz(n35), .test_si(n61), 
        .test_so(test_so), .test_se(test_se) );
  dbnc_WIDTH3 u0_sqlch_db ( .o_dbc(d_sqlch), .o_chg(), .i_org(i_sqlch), .clk(
        clk), .rstz(n35), .test_si(ptx_cc), .test_so(n61), .test_se(test_se)
         );
  SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 clk_gate_cclow_cnt_reg ( 
        .CLK(clk), .EN(N34), .ENCLK(net10355), .TE(test_se) );
  SDFFSQX1 d_cc_reg_0_ ( .D(i_cc_49), .SIN(cclow_cnt[8]), .SMC(test_se), .C(
        clk), .XS(n35), .Q(d_cc[0]) );
  SDFFSQX1 d_cc_reg_1_ ( .D(d_cc[0]), .SIN(d_cc[0]), .SMC(test_se), .C(clk), 
        .XS(n35), .Q(d_cc[1]) );
  SDFFQX1 cclow_cnt_reg_1_ ( .D(N36), .SIN(cclow_cnt[0]), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[1]) );
  SDFFQX1 cclow_cnt_reg_3_ ( .D(N38), .SIN(cclow_cnt[2]), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[3]) );
  SDFFQX1 cclow_cnt_reg_8_ ( .D(n102), .SIN(cclow_cnt[7]), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[8]) );
  SDFFQX1 cclow_cnt_reg_4_ ( .D(N39), .SIN(cclow_cnt[3]), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[4]) );
  SDFFQX1 cclow_cnt_reg_5_ ( .D(N40), .SIN(cclow_cnt[4]), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[5]) );
  SDFFQX1 cclow_cnt_reg_6_ ( .D(N41), .SIN(cclow_cnt[5]), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[6]) );
  SDFFQX1 cclow_cnt_reg_2_ ( .D(N37), .SIN(cclow_cnt[1]), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[2]) );
  SDFFQX1 cclow_cnt_reg_7_ ( .D(N42), .SIN(cclow_cnt[6]), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[7]) );
  SDFFQX1 cclow_cnt_reg_0_ ( .D(N35), .SIN(test_si), .SMC(test_se), .C(
        net10355), .Q(cclow_cnt[0]) );
  INVX1 U3 ( .A(1'b1), .Y(dbgpo[31]) );
  AND2X1 U5 ( .A(r_txnumk[0]), .B(n33), .Y(c0_txnumk[0]) );
  MUX2X1 U6 ( .D0(prl_last), .D1(pff_one), .S(n32), .Y(mux_one) );
  AND2X1 U7 ( .A(n32), .B(n40), .Y(rx_pshords) );
  INVX1 U8 ( .A(n34), .Y(n33) );
  MUX2IX1 U9 ( .D0(n44), .D1(n100), .S(n38), .Y(pff_rxpart[5]) );
  MUX2IX1 U10 ( .D0(n45), .D1(n98), .S(n38), .Y(pff_rxpart[7]) );
  INVX1 U11 ( .A(ptx_oe), .Y(n5) );
  INVX1 U12 ( .A(n5), .Y(n6) );
  INVX1 U13 ( .A(n108), .Y(n7) );
  INVX1 U14 ( .A(n7), .Y(prl_cany0) );
  BUFX3 U15 ( .A(prx_fsm[3]), .Y(dbgpo[23]) );
  BUFX3 U16 ( .A(prx_rcvinf[4]), .Y(dbgpo[19]) );
  BUFX3 U17 ( .A(prx_fsm[0]), .Y(dbgpo[20]) );
  BUFX3 U18 ( .A(prx_fsm[1]), .Y(dbgpo[21]) );
  BUFX3 U19 ( .A(prx_fsm[2]), .Y(dbgpo[22]) );
  BUFX3 U20 ( .A(pff_rdat[0]), .Y(dbgpo[8]) );
  BUFX3 U21 ( .A(pff_rdat[7]), .Y(dbgpo[15]) );
  BUFX3 U22 ( .A(pff_rdat[1]), .Y(dbgpo[9]) );
  BUFX3 U23 ( .A(pff_rdat[2]), .Y(dbgpo[10]) );
  BUFX3 U24 ( .A(pff_rdat[6]), .Y(dbgpo[14]) );
  BUFX3 U25 ( .A(pff_rdat[3]), .Y(dbgpo[11]) );
  BUFX3 U26 ( .A(pff_rdat[4]), .Y(dbgpo[12]) );
  BUFX3 U27 ( .A(pff_rdat[5]), .Y(dbgpo[13]) );
  AND2X1 U28 ( .A(r_txnumk[2]), .B(n33), .Y(c0_txnumk[2]) );
  AND2XL U29 ( .A(r_txnumk[1]), .B(n33), .Y(c0_txnumk[1]) );
  INVXL U30 ( .A(n34), .Y(n32) );
  INVXL U31 ( .A(n34), .Y(n31) );
  AND2X1 U32 ( .A(dbgpo[30]), .B(n34), .Y(fifopop_prl) );
  MUX2XL U33 ( .D0(prl_txreq), .D1(pff_txreq), .S(n31), .Y(n10) );
  AND2XL U34 ( .A(r_txendk), .B(n32), .Y(c0_txendk) );
  MUX2XL U35 ( .D0(prl_rdat[5]), .D1(pff_rdat[5]), .S(n32), .Y(mux_rdat[5]) );
  BUFXL U36 ( .A(dbgpo[17]), .Y(prx_rcvinf[3]) );
  AND2XL U37 ( .A(r_txnumk[3]), .B(n33), .Y(c0_txnumk[3]) );
  MUX2XL U38 ( .D0(prl_rdat[1]), .D1(pff_rdat[1]), .S(n32), .Y(mux_rdat[1]) );
  AND2XL U39 ( .A(r_txauto[6]), .B(n32), .Y(c0_txauto[6]) );
  AO22XL U40 ( .A(ptx_crcsidat[3]), .B(n6), .C(prx_crcsidat[3]), .D(n5), .Y(
        crcsidat[3]) );
  MUX2IXL U41 ( .D0(pff_rdat[1]), .D1(pff_dat_7_1[9]), .S(n37), .Y(n51) );
  MUX2XL U42 ( .D0(pff_rdat[0]), .D1(pff_dat_7_1[8]), .S(n37), .Y(
        pff_rxpart[0]) );
  MUX2XL U43 ( .D0(pff_rdat[3]), .D1(pff_dat_7_1[11]), .S(n38), .Y(
        pff_rxpart[3]) );
  MUX2XL U44 ( .D0(pff_rdat[2]), .D1(pff_dat_7_1[10]), .S(n37), .Y(
        pff_rxpart[2]) );
  MUX2XL U45 ( .D0(pff_rdat[4]), .D1(pff_dat_7_1[12]), .S(n37), .Y(
        pff_rxpart[4]) );
  MUX2XL U46 ( .D0(prl_txauto[0]), .D1(r_txauto[0]), .S(n31), .Y(c0_txauto[0])
         );
  MUX2XL U47 ( .D0(prl_txauto[2]), .D1(r_txauto[2]), .S(n31), .Y(c0_txauto[2])
         );
  MUX2XL U48 ( .D0(prl_txauto[1]), .D1(r_txauto[1]), .S(n31), .Y(c0_txauto[1])
         );
  NAND21XL U49 ( .B(r_txauto[3]), .A(n31), .Y(c0_txauto[3]) );
  MUX2XL U50 ( .D0(prl_txauto[4]), .D1(r_txauto[4]), .S(n31), .Y(c0_txauto[4])
         );
  NAND21XL U51 ( .B(r_txauto[5]), .A(n31), .Y(c0_txauto[5]) );
  INVXL U52 ( .A(pff_rdat[7]), .Y(n45) );
  INVXL U53 ( .A(pff_rdat[5]), .Y(n44) );
  INVX1 U54 ( .A(prl_idle), .Y(n34) );
  NOR21XL U55 ( .B(ptx_crcshfo4), .A(n5), .Y(crcshfo4) );
  AND2X1 U56 ( .A(prx_setsta[3]), .B(n58), .Y(prx_gdmsgrcvd) );
  NOR2X1 U57 ( .A(prx_fiforst), .B(n36), .Y(fifosrstz) );
  AND2XL U58 ( .A(dbgpo[30]), .B(n33), .Y(fifopop_pff) );
  MUX2X1 U59 ( .D0(pff_dat_7_1[18]), .D1(pff_dat_7_1[34]), .S(n39), .Y(
        pff_c0dat[26]) );
  MUX2X1 U60 ( .D0(pff_dat_7_1[17]), .D1(pff_dat_7_1[33]), .S(n39), .Y(
        pff_c0dat[25]) );
  MUX2X1 U61 ( .D0(pff_dat_7_1[15]), .D1(pff_dat_7_1[31]), .S(n39), .Y(
        pff_c0dat[23]) );
  INVX1 U62 ( .A(n36), .Y(n35) );
  INVX1 U63 ( .A(n43), .Y(n40) );
  AO22X1 U64 ( .A(ptx_crcstart), .B(n6), .C(prx_crcstart), .D(n5), .Y(crcstart) );
  AO22X1 U65 ( .A(ptx_crcshfi4), .B(n6), .C(prx_crcshfi4), .D(n5), .Y(crcshfi4) );
  MUX2X1 U66 ( .D0(pff_dat_7_1[11]), .D1(pff_dat_7_1[27]), .S(n38), .Y(
        pff_c0dat[19]) );
  NAND42X1 U67 ( .C(pff_rxpart[14]), .D(pff_rxpart[13]), .A(n54), .B(n53), .Y(
        n58) );
  AND3X1 U68 ( .A(n52), .B(pff_rxpart[0]), .C(n51), .Y(n53) );
  NOR32XL U69 ( .B(n50), .C(n49), .A(n48), .Y(n54) );
  NAND21X1 U70 ( .B(pff_rxpart[4]), .A(n47), .Y(n48) );
  INVX1 U71 ( .A(n43), .Y(n38) );
  INVX1 U72 ( .A(pff_rxpart[12]), .Y(n47) );
  INVX1 U73 ( .A(pff_rxpart[2]), .Y(n49) );
  INVX1 U74 ( .A(pff_rxpart[3]), .Y(n50) );
  MUX2IX1 U75 ( .D0(n97), .D1(n92), .S(n39), .Y(pff_c0dat[24]) );
  MUX2IX1 U76 ( .D0(n100), .D1(n83), .S(n39), .Y(pff_c0dat[21]) );
  INVX1 U77 ( .A(n43), .Y(n39) );
  MUX2X1 U78 ( .D0(pff_dat_7_1[20]), .D1(pff_dat_7_1[36]), .S(n39), .Y(
        pff_c0dat[28]) );
  MUX2X1 U79 ( .D0(pff_dat_7_1[19]), .D1(pff_dat_7_1[35]), .S(n39), .Y(
        pff_c0dat[27]) );
  INVX1 U80 ( .A(n43), .Y(n41) );
  INVX1 U81 ( .A(n43), .Y(n42) );
  INVX1 U82 ( .A(n52), .Y(pff_rxpart[15]) );
  MUX2IX1 U83 ( .D0(n99), .D1(n66), .S(n39), .Y(pff_c0dat[22]) );
  MUX2BXL U84 ( .D0(pff_dat_7_1[12]), .D1(n85), .S(n39), .Y(pff_c0dat[20]) );
  MUX2BXL U85 ( .D0(pff_dat_7_1[21]), .D1(n67), .S(n39), .Y(pff_c0dat[29]) );
  INVX1 U86 ( .A(n51), .Y(pff_rxpart[1]) );
  INVX1 U87 ( .A(srstz), .Y(n36) );
  INVX1 U88 ( .A(n72), .Y(n104) );
  INVX1 U89 ( .A(n76), .Y(n106) );
  INVX1 U90 ( .A(n74), .Y(n105) );
  MUX2X1 U91 ( .D0(prl_rdat[7]), .D1(pff_rdat[7]), .S(n31), .Y(mux_rdat[7]) );
  MUX2X1 U92 ( .D0(prl_rdat[4]), .D1(pff_rdat[4]), .S(n32), .Y(mux_rdat[4]) );
  MUX2X1 U93 ( .D0(prl_rdat[6]), .D1(pff_rdat[6]), .S(n31), .Y(mux_rdat[6]) );
  MUX2X1 U94 ( .D0(prl_rdat[0]), .D1(pff_rdat[0]), .S(n32), .Y(mux_rdat[0]) );
  MUX2X1 U95 ( .D0(prl_rdat[2]), .D1(pff_rdat[2]), .S(n31), .Y(mux_rdat[2]) );
  MUX2X1 U96 ( .D0(prl_rdat[3]), .D1(pff_rdat[3]), .S(n32), .Y(mux_rdat[3]) );
  AND2XL U97 ( .A(r_txnumk[4]), .B(n33), .Y(c0_txnumk[4]) );
  INVX1 U98 ( .A(r_pshords), .Y(n43) );
  AOI21AXL U99 ( .B(n6), .C(n33), .A(r_first), .Y(lockena) );
  AO22X1 U100 ( .A(ptx_crcsidat[1]), .B(n6), .C(prx_crcsidat[1]), .D(n5), .Y(
        crcsidat[1]) );
  AO22X1 U101 ( .A(ptx_crcsidat[0]), .B(n6), .C(prx_crcsidat[0]), .D(n5), .Y(
        crcsidat[0]) );
  MUX2BXL U102 ( .D0(pff_rdat[6]), .D1(n99), .S(n37), .Y(pff_rxpart[6]) );
  INVX1 U103 ( .A(n46), .Y(pff_rxpart[8]) );
  MUX2AXL U104 ( .D0(pff_dat_7_1[0]), .D1(n97), .S(n37), .Y(n46) );
  NOR21XL U105 ( .B(obsd), .A(prx_setsta[6]), .Y(pff_obsd) );
  MUX2X1 U106 ( .D0(pff_dat_7_1[4]), .D1(pff_dat_7_1[20]), .S(n38), .Y(
        pff_rxpart[12]) );
  MUX2IX1 U107 ( .D0(pff_dat_7_1[7]), .D1(pff_dat_7_1[23]), .S(n37), .Y(n52)
         );
  MUX2X1 U108 ( .D0(pff_dat_7_1[5]), .D1(pff_dat_7_1[21]), .S(n38), .Y(
        pff_rxpart[13]) );
  MUX2X1 U109 ( .D0(pff_dat_7_1[6]), .D1(pff_dat_7_1[22]), .S(n38), .Y(
        pff_rxpart[14]) );
  INVX1 U110 ( .A(n43), .Y(n37) );
  NOR21XL U111 ( .B(r_auto_gdcrc[1]), .A(n58), .Y(auto_rx_gdcrc) );
  ENOX1 U112 ( .A(n41), .B(n60), .C(pff_dat_7_1[55]), .D(r_pshords), .Y(
        pff_c0dat[47]) );
  ENOX1 U113 ( .A(n41), .B(n67), .C(pff_dat_7_1[53]), .D(r_pshords), .Y(
        pff_c0dat[45]) );
  ENOX1 U114 ( .A(n40), .B(n91), .C(pff_dat_7_1[41]), .D(n42), .Y(
        pff_c0dat[33]) );
  MUX2X1 U115 ( .D0(pff_dat_7_1[22]), .D1(pff_dat_7_1[38]), .S(n40), .Y(
        pff_c0dat[30]) );
  MUX2X1 U116 ( .D0(pff_dat_7_1[8]), .D1(pff_dat_7_1[24]), .S(n38), .Y(
        pff_c0dat[16]) );
  MUX2X1 U117 ( .D0(pff_dat_7_1[10]), .D1(pff_dat_7_1[26]), .S(n38), .Y(
        pff_c0dat[18]) );
  ENOX1 U118 ( .A(n41), .B(n86), .C(pff_dat_7_1[51]), .D(r_pshords), .Y(
        pff_c0dat[43]) );
  ENOX1 U119 ( .A(n41), .B(n88), .C(pff_dat_7_1[50]), .D(n42), .Y(
        pff_c0dat[42]) );
  ENOX1 U120 ( .A(n41), .B(n84), .C(pff_dat_7_1[52]), .D(r_pshords), .Y(
        pff_c0dat[44]) );
  ENOX1 U121 ( .A(n40), .B(n93), .C(pff_dat_7_1[40]), .D(n41), .Y(
        pff_c0dat[32]) );
  ENOX1 U122 ( .A(n40), .B(n83), .C(pff_dat_7_1[45]), .D(n42), .Y(
        pff_c0dat[37]) );
  ENOX1 U123 ( .A(n40), .B(n87), .C(pff_dat_7_1[43]), .D(n42), .Y(
        pff_c0dat[35]) );
  MUX2BXL U124 ( .D0(pff_dat_7_1[9]), .D1(n91), .S(n38), .Y(pff_c0dat[17]) );
  MUX2BXL U125 ( .D0(pff_dat_7_1[23]), .D1(n60), .S(n40), .Y(pff_c0dat[31]) );
  ENOX1 U126 ( .A(n41), .B(n90), .C(pff_dat_7_1[49]), .D(n42), .Y(
        pff_c0dat[41]) );
  ENOX1 U127 ( .A(n41), .B(n65), .C(pff_dat_7_1[47]), .D(n42), .Y(
        pff_c0dat[39]) );
  ENOX1 U128 ( .A(n40), .B(n66), .C(pff_dat_7_1[46]), .D(n42), .Y(
        pff_c0dat[38]) );
  ENOX1 U129 ( .A(n40), .B(n85), .C(pff_dat_7_1[44]), .D(n42), .Y(
        pff_c0dat[36]) );
  INVX1 U130 ( .A(pff_dat_7_1[26]), .Y(n89) );
  INVX1 U131 ( .A(pff_dat_7_1[24]), .Y(n93) );
  INVX1 U132 ( .A(pff_dat_7_1[29]), .Y(n83) );
  INVX1 U133 ( .A(pff_dat_7_1[32]), .Y(n92) );
  INVX1 U134 ( .A(pff_dat_7_1[38]), .Y(n101) );
  INVX1 U135 ( .A(pff_dat_7_1[35]), .Y(n86) );
  INVX1 U136 ( .A(pff_dat_7_1[36]), .Y(n84) );
  INVX1 U137 ( .A(pff_dat_7_1[34]), .Y(n88) );
  INVX1 U138 ( .A(pff_dat_7_1[25]), .Y(n91) );
  INVX1 U139 ( .A(pff_dat_7_1[37]), .Y(n67) );
  INVX1 U140 ( .A(pff_dat_7_1[39]), .Y(n60) );
  INVX1 U141 ( .A(pff_dat_7_1[31]), .Y(n65) );
  INVX1 U142 ( .A(pff_dat_7_1[33]), .Y(n90) );
  INVX1 U143 ( .A(pff_dat_7_1[30]), .Y(n66) );
  INVX1 U144 ( .A(pff_dat_7_1[16]), .Y(n97) );
  INVX1 U145 ( .A(pff_dat_7_1[19]), .Y(n94) );
  INVX1 U146 ( .A(pff_dat_7_1[17]), .Y(n96) );
  INVX1 U147 ( .A(pff_dat_7_1[18]), .Y(n95) );
  ENOX1 U148 ( .A(n40), .B(n89), .C(pff_dat_7_1[42]), .D(n42), .Y(
        pff_c0dat[34]) );
  INVX1 U149 ( .A(pff_dat_7_1[15]), .Y(n98) );
  INVX1 U150 ( .A(pff_dat_7_1[13]), .Y(n100) );
  ENOX1 U151 ( .A(n41), .B(n101), .C(pff_dat_7_1[54]), .D(r_pshords), .Y(
        pff_c0dat[46]) );
  ENOX1 U152 ( .A(n41), .B(n92), .C(pff_dat_7_1[48]), .D(n42), .Y(
        pff_c0dat[40]) );
  INVX1 U153 ( .A(pff_dat_7_1[27]), .Y(n87) );
  INVX1 U154 ( .A(pff_dat_7_1[28]), .Y(n85) );
  INVX1 U155 ( .A(pff_dat_7_1[14]), .Y(n99) );
  AOI31X1 U156 ( .A(d_sqlch), .B(n55), .C(r_sqlch[0]), .D(n59), .Y(x_trans) );
  OAI21X1 U157 ( .B(n6), .C(prx_fsm[3]), .A(r_sqlch[1]), .Y(n55) );
  INVX1 U158 ( .A(prx_trans), .Y(n59) );
  NOR21XL U159 ( .B(ptx_goidle), .A(prl_cany0), .Y(ptx_ack) );
  NOR4XL U160 ( .A(n56), .B(n57), .C(cclow_cnt[5]), .D(cclow_cnt[4]), .Y(
        prx_setsta[0]) );
  OR3XL U161 ( .A(cclow_cnt[7]), .B(cclow_cnt[6]), .C(cclow_cnt[8]), .Y(n57)
         );
  NAND43X1 U162 ( .B(cclow_cnt[3]), .C(cclow_cnt[1]), .D(cclow_cnt[2]), .A(
        cclow_cnt[0]), .Y(n56) );
  OAI211X1 U163 ( .C(cclow_cnt[8]), .D(n69), .A(n35), .B(n82), .Y(n72) );
  XNOR2XL U164 ( .A(d_cc[1]), .B(d_cc[0]), .Y(n82) );
  GEN2XL U165 ( .D(cclow_cnt[1]), .E(cclow_cnt[0]), .C(n80), .B(n104), .A(n70), 
        .Y(N36) );
  GEN2XL U166 ( .D(cclow_cnt[4]), .E(n75), .C(n76), .B(n104), .A(n70), .Y(N39)
         );
  GEN2XL U167 ( .D(cclow_cnt[6]), .E(n105), .C(n73), .B(n104), .A(n70), .Y(N41) );
  GEN2XL U168 ( .D(cclow_cnt[5]), .E(n106), .C(n74), .B(n104), .A(n70), .Y(N40) );
  NAND21X1 U169 ( .B(cclow_cnt[2]), .A(n80), .Y(n78) );
  NAND21X1 U170 ( .B(cclow_cnt[7]), .A(n73), .Y(n69) );
  NOR2X1 U171 ( .A(n75), .B(cclow_cnt[4]), .Y(n76) );
  NOR2X1 U172 ( .A(n106), .B(cclow_cnt[5]), .Y(n74) );
  NOR2X1 U173 ( .A(n105), .B(cclow_cnt[6]), .Y(n73) );
  NOR2X1 U174 ( .A(cclow_cnt[1]), .B(cclow_cnt[0]), .Y(n80) );
  AOI21X1 U175 ( .B(n69), .C(n71), .A(n72), .Y(N42) );
  NAND21X1 U176 ( .B(n73), .A(cclow_cnt[7]), .Y(n71) );
  AOI21X1 U178 ( .B(n78), .C(n79), .A(n72), .Y(N37) );
  NAND21X1 U179 ( .B(n80), .A(cclow_cnt[2]), .Y(n79) );
  AOI21X1 U180 ( .B(n75), .C(n77), .A(n72), .Y(N38) );
  NAND2X1 U181 ( .A(cclow_cnt[3]), .B(n78), .Y(n77) );
  OR2X1 U182 ( .A(n78), .B(cclow_cnt[3]), .Y(n75) );
  NOR2X1 U183 ( .A(cclow_cnt[0]), .B(n72), .Y(N35) );
  INVX1 U184 ( .A(n68), .Y(n102) );
  AOI31X1 U185 ( .A(n104), .B(n69), .C(cclow_cnt[8]), .D(n70), .Y(n68) );
  NAND31X1 U186 ( .C(n70), .A(n72), .B(n81), .Y(N34) );
  AOI21X1 U187 ( .B(d_cc[0]), .C(n103), .A(n36), .Y(n81) );
  NOR3XL U188 ( .A(n36), .B(d_cc[0]), .C(n103), .Y(n70) );
  MUX2BXL U189 ( .D0(pff_dat_7_1[3]), .D1(n94), .S(n37), .Y(pff_rxpart[11]) );
  MUX2BXL U190 ( .D0(pff_dat_7_1[2]), .D1(n95), .S(n37), .Y(pff_rxpart[10]) );
  MUX2BXL U191 ( .D0(pff_dat_7_1[1]), .D1(n96), .S(n37), .Y(pff_rxpart[9]) );
  INVX1 U192 ( .A(d_cc[1]), .Y(n103) );
  AND2XL U193 ( .A(dbgpo[29]), .B(n32), .Y(fifopsh_pff) );
  AO22XL U194 ( .A(ptx_crcsidat[2]), .B(n6), .C(prx_crcsidat[2]), .D(n5), .Y(
        crcsidat[2]) );
  AND2X2 U195 ( .A(dbgpo[29]), .B(n34), .Y(fifopsh_prl) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_1_, db_cnt_0_, N14, N15, N16, N17, net10373, n8, n1,
         n2, n3, n4, n5;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N14), 
        .ENCLK(net10373), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N17), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net10373), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N16), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net10373), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N15), .SIN(o_dbc), .SMC(test_se), .C(net10373), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n8), .SIN(d_org_0_), .SMC(test_se), .C(net10373), 
        .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n2), .A(n1), .Y(n4) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U5 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n8) );
  NOR2X1 U6 ( .A(n1), .B(n2), .Y(o_chg) );
  NAND3X1 U7 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(test_so), .Y(n1) );
  NOR2X1 U8 ( .A(n5), .B(n4), .Y(N16) );
  XNOR2XL U9 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n5) );
  NOR2X1 U10 ( .A(db_cnt_0_), .B(n4), .Y(N15) );
  NOR2X1 U11 ( .A(n3), .B(n4), .Y(N17) );
  AOI21X1 U12 ( .B(db_cnt_1_), .C(db_cnt_0_), .A(test_so), .Y(n3) );
  NAND43X1 U13 ( .B(test_so), .C(db_cnt_0_), .D(db_cnt_1_), .A(n2), .Y(N14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updprl_a0 ( r_spec, r_dat_spec, r_auto_txgdcrc, r_dat_portrole, 
        r_dat_datarole, r_auto_discard, r_set_cpmsgid, r_dat_cpmsgid, r_rdat, 
        r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact, ptx_fifopop, 
        prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, prx_rcvdords, prx_fifowdat, 
        pff_c0dat, prl_rdat, prl_txauto, prl_last, prl_txreq, prl_c0set, 
        prl_cany0, prl_cany0r, prl_cany0w, prl_idle, prl_discard, prl_GCTxDone, 
        prl_fsm, prl_cpmsgid, prl_cany0adr, clk, srstz, test_si, test_so, 
        test_se );
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [2:0] r_dat_cpmsgid;
  input [7:0] r_rdat;
  input [2:0] prx_rcvdords;
  input [7:0] prx_fifowdat;
  input [47:0] pff_c0dat;
  output [7:0] prl_rdat;
  output [6:0] prl_txauto;
  output [3:0] prl_fsm;
  output [2:0] prl_cpmsgid;
  output [7:0] prl_cany0adr;
  input r_auto_txgdcrc, r_dat_portrole, r_dat_datarole, r_auto_discard,
         r_set_cpmsgid, r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact,
         ptx_fifopop, prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, clk, srstz,
         test_si, test_se;
  output prl_last, prl_txreq, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_idle, prl_discard, prl_GCTxDone, test_so;
  wire   sendgdcrc, stoptimer, N41, c0_iop, N113, N114, N115, N116, N117, N118,
         N119, N120, N151, N152, N153, N154, N155, N156, N157, N158, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N189, N190, N191,
         N192, N193, N194, N196, N203, N204, N205, N206, net10396, net10402,
         net10407, net10412, net10417, n99, n100, n37, n39, n51, n57, n67, n68,
         n72, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n101, n7, n8, n9, n10, n11, n12, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n52, n53, n54, n55, n56, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n69, n70, n71, n73, n74, n75, n76, n77, n78, n79, n80, n97, n98,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147;
  wire   [1:0] PrlTo;
  wire   [8:0] c0_cnt;
  wire   [7:0] txbuf;

  PrlTimer_1112a0 u0_PrlTimer ( .to(PrlTo), .restart(sendgdcrc), .stop(
        stoptimer), .clk(clk), .srstz(n16), .test_si(txbuf[7]), .test_so(
        test_so), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_0 clk_gate_txbuf_reg ( .CLK(clk), .EN(N41), 
        .ENCLK(net10396), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_4 clk_gate_c0_adr_reg ( .CLK(clk), .EN(N194), 
        .ENCLK(net10402), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_3 clk_gate_cs_prcl_reg ( .CLK(clk), .EN(N189), 
        .ENCLK(net10407), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_2 clk_gate_c0_cnt_reg ( .CLK(clk), .EN(N196), 
        .ENCLK(net10412), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_1 clk_gate_CpMsgId_reg ( .CLK(clk), .EN(N203), 
        .ENCLK(net10417), .TE(test_se) );
  updprl_a0_DW01_inc_0 r328 ( .A(prl_cany0adr), .SUM({N120, N119, N118, N117, 
        N116, N115, N114, N113}) );
  SDFFQXL txbuf_reg_3_ ( .D(r_rdat[3]), .SIN(txbuf[2]), .SMC(test_se), .C(
        net10396), .Q(txbuf[3]) );
  SDFFQX1 c0_iop_reg ( .D(n99), .SIN(c0_cnt[8]), .SMC(test_se), .C(net10407), 
        .Q(c0_iop) );
  SDFFQX1 canyon_m0_reg ( .D(n100), .SIN(c0_iop), .SMC(test_se), .C(clk), .Q(
        prl_cany0) );
  SDFFQX1 c0_adr_reg_6_ ( .D(N157), .SIN(prl_cany0adr[5]), .SMC(test_se), .C(
        net10402), .Q(prl_cany0adr[6]) );
  SDFFQX1 c0_adr_reg_2_ ( .D(N153), .SIN(prl_cany0adr[1]), .SMC(test_se), .C(
        net10402), .Q(prl_cany0adr[2]) );
  SDFFQX1 c0_adr_reg_4_ ( .D(N155), .SIN(prl_cany0adr[3]), .SMC(test_se), .C(
        net10402), .Q(prl_cany0adr[4]) );
  SDFFQX1 c0_adr_reg_1_ ( .D(N152), .SIN(prl_cany0adr[0]), .SMC(test_se), .C(
        net10402), .Q(prl_cany0adr[1]) );
  SDFFQX1 c0_adr_reg_3_ ( .D(N154), .SIN(prl_cany0adr[2]), .SMC(test_se), .C(
        net10402), .Q(prl_cany0adr[3]) );
  SDFFQX1 c0_adr_reg_5_ ( .D(N156), .SIN(prl_cany0adr[4]), .SMC(test_se), .C(
        net10402), .Q(prl_cany0adr[5]) );
  SDFFQX1 c0_adr_reg_7_ ( .D(N158), .SIN(prl_cany0adr[6]), .SMC(test_se), .C(
        net10402), .Q(prl_cany0adr[7]) );
  SDFFQX1 c0_adr_reg_0_ ( .D(N151), .SIN(prl_cpmsgid[2]), .SMC(test_se), .C(
        net10402), .Q(prl_cany0adr[0]) );
  SDFFQX1 txbuf_reg_2_ ( .D(r_rdat[2]), .SIN(txbuf[1]), .SMC(test_se), .C(
        net10396), .Q(txbuf[2]) );
  SDFFQX1 txbuf_reg_1_ ( .D(r_rdat[1]), .SIN(txbuf[0]), .SMC(test_se), .C(
        net10396), .Q(txbuf[1]) );
  SDFFQX1 txbuf_reg_6_ ( .D(r_rdat[6]), .SIN(txbuf[5]), .SMC(test_se), .C(
        net10396), .Q(txbuf[6]) );
  SDFFQX1 txbuf_reg_7_ ( .D(r_rdat[7]), .SIN(txbuf[6]), .SMC(test_se), .C(
        net10396), .Q(txbuf[7]) );
  SDFFQX1 CpMsgId_reg_1_ ( .D(N205), .SIN(prl_cpmsgid[0]), .SMC(test_se), .C(
        net10417), .Q(prl_cpmsgid[1]) );
  SDFFQX1 c0_cnt_reg_8_ ( .D(N173), .SIN(c0_cnt[7]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[8]) );
  SDFFQX1 c0_cnt_reg_7_ ( .D(N172), .SIN(c0_cnt[6]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[7]) );
  SDFFQX1 txbuf_reg_0_ ( .D(r_rdat[0]), .SIN(prl_fsm[3]), .SMC(test_se), .C(
        net10396), .Q(txbuf[0]) );
  SDFFQX1 c0_cnt_reg_3_ ( .D(N168), .SIN(c0_cnt[2]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[3]) );
  SDFFQX1 c0_cnt_reg_2_ ( .D(N167), .SIN(c0_cnt[1]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[2]) );
  SDFFQX1 c0_cnt_reg_6_ ( .D(N171), .SIN(c0_cnt[5]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[6]) );
  SDFFQX1 c0_cnt_reg_5_ ( .D(N170), .SIN(c0_cnt[4]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[5]) );
  SDFFQX1 c0_cnt_reg_4_ ( .D(N169), .SIN(c0_cnt[3]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[4]) );
  SDFFQX1 txbuf_reg_5_ ( .D(r_rdat[5]), .SIN(txbuf[4]), .SMC(test_se), .C(
        net10396), .Q(txbuf[5]) );
  SDFFQXL CpMsgId_reg_0_ ( .D(N204), .SIN(test_si), .SMC(test_se), .C(net10417), .Q(prl_cpmsgid[0]) );
  SDFFQXL CpMsgId_reg_2_ ( .D(N206), .SIN(prl_cpmsgid[1]), .SMC(test_se), .C(
        net10417), .Q(prl_cpmsgid[2]) );
  SDFFQX1 txbuf_reg_4_ ( .D(r_rdat[4]), .SIN(txbuf[3]), .SMC(test_se), .C(
        net10396), .Q(txbuf[4]) );
  SDFFQX1 cs_prcl_reg_1_ ( .D(N191), .SIN(prl_fsm[0]), .SMC(test_se), .C(
        net10407), .Q(prl_fsm[1]) );
  SDFFQX1 cs_prcl_reg_0_ ( .D(N190), .SIN(prl_cany0), .SMC(test_se), .C(
        net10407), .Q(prl_fsm[0]) );
  SDFFQX1 cs_prcl_reg_3_ ( .D(N193), .SIN(prl_fsm[2]), .SMC(test_se), .C(
        net10407), .Q(prl_fsm[3]) );
  SDFFQX1 cs_prcl_reg_2_ ( .D(N192), .SIN(prl_fsm[1]), .SMC(test_se), .C(
        net10407), .Q(prl_fsm[2]) );
  SDFFQX1 c0_cnt_reg_0_ ( .D(N165), .SIN(prl_cany0adr[7]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[0]) );
  SDFFQX1 c0_cnt_reg_1_ ( .D(N166), .SIN(c0_cnt[0]), .SMC(test_se), .C(
        net10412), .Q(c0_cnt[1]) );
  INVX1 U3 ( .A(1'b0), .Y(prl_txauto[3]) );
  INVX1 U5 ( .A(1'b0), .Y(prl_txauto[5]) );
  INVX1 U7 ( .A(1'b1), .Y(prl_txauto[6]) );
  INVX1 U9 ( .A(n22), .Y(n24) );
  INVX1 U10 ( .A(prl_fsm[1]), .Y(n61) );
  NAND21X1 U11 ( .B(n79), .A(n128), .Y(n142) );
  OR2X1 U12 ( .A(prl_fsm[2]), .B(n25), .Y(n143) );
  NAND21X1 U13 ( .B(c0_cnt[3]), .A(n35), .Y(n42) );
  INVX1 U14 ( .A(n45), .Y(n43) );
  NAND21X1 U15 ( .B(c0_cnt[4]), .A(n40), .Y(n45) );
  INVX1 U16 ( .A(n48), .Y(n46) );
  NAND21X1 U17 ( .B(c0_cnt[5]), .A(n43), .Y(n48) );
  INVX1 U18 ( .A(n52), .Y(n49) );
  INVX1 U19 ( .A(c0_cnt[0]), .Y(n30) );
  INVX1 U20 ( .A(n38), .Y(n35) );
  NAND21X1 U21 ( .B(c0_cnt[2]), .A(n32), .Y(n38) );
  INVX1 U22 ( .A(n42), .Y(n40) );
  NAND21X1 U23 ( .B(c0_cnt[6]), .A(n46), .Y(n52) );
  INVX1 U24 ( .A(n55), .Y(n53) );
  NAND21X1 U25 ( .B(c0_cnt[7]), .A(n49), .Y(n55) );
  INVX1 U26 ( .A(n54), .Y(n122) );
  NAND21X1 U27 ( .B(c0_cnt[8]), .A(n53), .Y(n54) );
  INVX1 U28 ( .A(prl_fsm[0]), .Y(n106) );
  INVX1 U29 ( .A(n108), .Y(n7) );
  OAI21X1 U30 ( .B(prx_eoprcvd), .C(pid_ccidle), .A(n56), .Y(n20) );
  NAND32X1 U31 ( .B(prl_fsm[2]), .C(n18), .A(n61), .Y(n108) );
  NAND32XL U32 ( .B(prl_fsm[2]), .C(prl_fsm[1]), .A(n24), .Y(n80) );
  INVX2 U33 ( .A(n118), .Y(prl_cany0w) );
  INVX3 U34 ( .A(prx_fifopsh), .Y(n107) );
  INVXL U35 ( .A(prl_txauto[4]), .Y(n121) );
  OAI211XL U36 ( .C(n128), .D(n17), .A(n60), .B(n112), .Y(N192) );
  NAND21XL U37 ( .B(n56), .A(n97), .Y(n29) );
  INVXL U38 ( .A(n128), .Y(n120) );
  OAI22AXL U39 ( .D(prl_cpmsgid[1]), .C(n128), .A(n142), .B(n126), .Y(
        prl_rdat[2]) );
  NAND21X1 U40 ( .B(c0_cnt[1]), .A(n30), .Y(n34) );
  NAND42XL U41 ( .C(n143), .D(r_dat_datarole), .A(n132), .B(n131), .Y(n133) );
  NAND21XL U42 ( .B(prl_fsm[3]), .A(prl_fsm[0]), .Y(n62) );
  INVXL U43 ( .A(prl_fsm[2]), .Y(n58) );
  OAI22XL U44 ( .A(n142), .B(n125), .C(n128), .D(n124), .Y(prl_rdat[1]) );
  INVXL U45 ( .A(txbuf[1]), .Y(n125) );
  INVXL U46 ( .A(prl_cpmsgid[0]), .Y(n124) );
  INVXL U47 ( .A(r_spec[0]), .Y(n136) );
  INVXL U48 ( .A(prl_cpmsgid[2]), .Y(n127) );
  NAND21XL U49 ( .B(n61), .A(prl_fsm[2]), .Y(n21) );
  OAI211XL U50 ( .C(prl_fsm[0]), .D(n20), .A(n16), .B(n19), .Y(n109) );
  NAND4XL U51 ( .A(n105), .B(n27), .C(n106), .D(n69), .Y(n11) );
  BUFXL U52 ( .A(prx_rcvdords[0]), .Y(prl_txauto[0]) );
  BUFXL U53 ( .A(prx_rcvdords[2]), .Y(prl_txauto[2]) );
  BUFXL U54 ( .A(prx_rcvdords[1]), .Y(prl_txauto[1]) );
  NAND32XL U55 ( .B(prl_fsm[2]), .C(n62), .A(n61), .Y(n77) );
  NAND21XL U56 ( .B(n25), .A(prl_fsm[2]), .Y(n74) );
  INVX1 U57 ( .A(r_discard), .Y(n145) );
  INVX1 U58 ( .A(n17), .Y(n16) );
  NOR21XL U59 ( .B(prx_gdmsgrcvd), .A(r_set_cpmsgid), .Y(n57) );
  NAND32X1 U60 ( .B(r_set_cpmsgid), .C(prx_gdmsgrcvd), .A(n16), .Y(N203) );
  INVX1 U61 ( .A(srstz), .Y(n17) );
  NAND21X1 U62 ( .B(prl_txauto[4]), .A(ptx_fifopop), .Y(n110) );
  INVX1 U63 ( .A(n51), .Y(prl_c0set) );
  OR3XL U64 ( .A(pff_c0dat[26]), .B(pff_c0dat[25]), .C(pff_c0dat[23]), .Y(n89)
         );
  INVX1 U65 ( .A(n97), .Y(n73) );
  INVX1 U66 ( .A(n75), .Y(n59) );
  NAND32X1 U67 ( .B(n62), .C(n61), .A(n58), .Y(n128) );
  NAND21X1 U68 ( .B(n106), .A(n7), .Y(prl_txauto[4]) );
  NAND32X1 U69 ( .B(n108), .C(n107), .A(n106), .Y(n118) );
  AO21X1 U70 ( .B(n122), .C(n121), .A(n120), .Y(prl_last) );
  INVX1 U71 ( .A(n108), .Y(n56) );
  OAI22X1 U72 ( .A(n107), .B(n97), .C(n122), .D(n110), .Y(prl_cany0r) );
  INVX1 U73 ( .A(n80), .Y(prl_idle) );
  INVX1 U74 ( .A(n34), .Y(n32) );
  INVX1 U75 ( .A(n143), .Y(n79) );
  NAND21X1 U76 ( .B(n62), .A(n27), .Y(n97) );
  OAI21X1 U77 ( .B(ptx_txact), .C(prl_txauto[4]), .A(n119), .Y(prl_txreq) );
  NAND21X1 U78 ( .B(n66), .A(n112), .Y(N191) );
  GEN2XL U79 ( .D(n67), .E(n65), .C(n79), .B(n16), .A(n64), .Y(n66) );
  INVX1 U80 ( .A(n119), .Y(n65) );
  INVX1 U81 ( .A(n63), .Y(n64) );
  NOR2X1 U82 ( .A(r_discard), .B(n68), .Y(n67) );
  NAND4X1 U83 ( .A(n81), .B(n82), .C(n83), .D(n84), .Y(n51) );
  NOR4XL U84 ( .A(n88), .B(n89), .C(pff_c0dat[22]), .D(pff_c0dat[20]), .Y(n83)
         );
  NOR4XL U85 ( .A(n85), .B(n86), .C(pff_c0dat[36]), .D(pff_c0dat[34]), .Y(n84)
         );
  NOR42XL U86 ( .C(pff_c0dat[46]), .D(pff_c0dat[40]), .A(n94), .B(n95), .Y(n81) );
  NAND5XL U87 ( .A(n105), .B(n119), .C(n146), .D(n104), .E(n103), .Y(N189) );
  AOI221XL U88 ( .A(n117), .B(ptx_ack), .C(ptx_fifopop), .D(n142), .E(n102), 
        .Y(n103) );
  OA21X1 U89 ( .B(n77), .C(n145), .A(n76), .Y(n104) );
  AO21XL U90 ( .B(sendgdcrc), .C(prl_idle), .A(n98), .Y(n102) );
  NOR42XL U91 ( .C(pff_c0dat[1]), .D(pff_c0dat[19]), .A(n91), .B(n92), .Y(n82)
         );
  NAND3X1 U92 ( .A(pff_c0dat[12]), .B(pff_c0dat[0]), .C(pff_c0dat[17]), .Y(n92) );
  NAND42X1 U93 ( .C(pff_c0dat[14]), .D(pff_c0dat[13]), .A(prx_gdmsgrcvd), .B(
        n93), .Y(n91) );
  OAI21BBX1 U94 ( .A(r_dat_cpmsgid[1]), .B(r_set_cpmsgid), .C(n8), .Y(N205) );
  AOI21X1 U95 ( .B(pff_c0dat[10]), .C(n57), .A(n17), .Y(n8) );
  OAI21BBX1 U96 ( .A(r_dat_cpmsgid[2]), .B(r_set_cpmsgid), .C(n9), .Y(N206) );
  AOI21X1 U97 ( .B(pff_c0dat[11]), .C(n57), .A(n17), .Y(n9) );
  OAI21BBX1 U98 ( .A(r_dat_cpmsgid[0]), .B(r_set_cpmsgid), .C(n10), .Y(N204)
         );
  AOI21X1 U99 ( .B(pff_c0dat[9]), .C(n57), .A(n17), .Y(n10) );
  INVX1 U100 ( .A(n109), .Y(n105) );
  OAI211X1 U101 ( .C(n97), .D(n109), .A(n60), .B(n26), .Y(N190) );
  AO21X1 U102 ( .B(n80), .C(n143), .A(n17), .Y(n26) );
  INVX1 U103 ( .A(n23), .Y(n60) );
  OAI31XL U104 ( .A(n78), .B(n147), .C(n17), .D(n63), .Y(n23) );
  NAND21X1 U105 ( .B(n109), .A(n59), .Y(n112) );
  AO21XL U106 ( .B(n75), .C(n74), .A(n107), .Y(n76) );
  INVX1 U107 ( .A(n72), .Y(n69) );
  AO22X1 U108 ( .A(N117), .B(n29), .C(n59), .D(prx_fifowdat[4]), .Y(N155) );
  NAND32X1 U109 ( .B(pff_c0dat[28]), .C(pff_c0dat[27]), .A(n90), .Y(n88) );
  NOR3XL U110 ( .A(pff_c0dat[29]), .B(pff_c0dat[32]), .C(pff_c0dat[31]), .Y(
        n90) );
  AO22XL U111 ( .A(N118), .B(n29), .C(prx_fifowdat[5]), .D(n59), .Y(N156) );
  OR2X1 U112 ( .A(n39), .B(n77), .Y(n119) );
  NAND21X1 U113 ( .B(n77), .A(n68), .Y(n146) );
  INVX1 U114 ( .A(n78), .Y(n117) );
  INVX1 U115 ( .A(n74), .Y(n70) );
  INVX1 U116 ( .A(n111), .Y(n98) );
  NAND32X1 U117 ( .B(n62), .C(n58), .A(n61), .Y(n75) );
  AO22X1 U118 ( .A(N116), .B(n29), .C(n59), .D(prx_fifowdat[3]), .Y(N154) );
  OAI22X1 U119 ( .A(n144), .B(n143), .C(n142), .D(n141), .Y(prl_rdat[7]) );
  INVX1 U120 ( .A(txbuf[7]), .Y(n141) );
  MUX2BXL U121 ( .D0(n140), .D1(r_dat_spec[1]), .S(n139), .Y(n144) );
  AND2X1 U122 ( .A(txbuf[4]), .B(n130), .Y(prl_rdat[4]) );
  INVX1 U123 ( .A(n142), .Y(n130) );
  OAI22X1 U124 ( .A(n138), .B(n143), .C(n142), .D(n137), .Y(prl_rdat[6]) );
  INVX1 U125 ( .A(txbuf[6]), .Y(n137) );
  MUX2BXL U126 ( .D0(n136), .D1(r_dat_spec[0]), .S(n139), .Y(n138) );
  OAI221X1 U127 ( .A(n142), .B(n123), .C(r_dat_portrole), .D(n128), .E(n143), 
        .Y(prl_rdat[0]) );
  INVX1 U128 ( .A(txbuf[0]), .Y(n123) );
  INVX1 U129 ( .A(txbuf[2]), .Y(n126) );
  NAND32X1 U130 ( .B(prl_fsm[0]), .C(n61), .A(n18), .Y(n25) );
  OAI22X1 U131 ( .A(n142), .B(n129), .C(n128), .D(n127), .Y(prl_rdat[3]) );
  INVX1 U132 ( .A(txbuf[3]), .Y(n129) );
  NAND21X1 U133 ( .B(prl_fsm[3]), .A(n106), .Y(n22) );
  INVX1 U134 ( .A(n135), .Y(n139) );
  NAND21X1 U135 ( .B(n140), .A(r_spec[0]), .Y(n135) );
  INVXL U136 ( .A(prl_fsm[3]), .Y(n18) );
  INVX1 U137 ( .A(r_spec[1]), .Y(n140) );
  NAND21X1 U138 ( .B(n134), .A(n133), .Y(prl_rdat[5]) );
  NOR21XL U139 ( .B(txbuf[5]), .A(n142), .Y(n134) );
  NOR21XL U140 ( .B(prx_rcvdords[0]), .A(prx_rcvdords[1]), .Y(n132) );
  INVX1 U141 ( .A(prx_rcvdords[2]), .Y(n131) );
  INVX1 U142 ( .A(n21), .Y(n27) );
  OAI21BX1 U143 ( .C(PrlTo[0]), .B(r_auto_discard), .A(n37), .Y(stoptimer) );
  AND3X1 U144 ( .A(n39), .B(n146), .C(n145), .Y(n37) );
  NAND21X1 U145 ( .B(r_rdy), .A(n116), .Y(N41) );
  NAND43X1 U146 ( .B(prx_fifowdat[0]), .C(n72), .D(n74), .A(n105), .Y(n63) );
  OAI21BBX1 U147 ( .A(r_auto_txgdcrc), .B(prx_gdmsgrcvd), .C(n51), .Y(
        sendgdcrc) );
  MUX2X1 U148 ( .D0(prx_fifowdat[1]), .D1(c0_iop), .S(n11), .Y(n99) );
  OA21X1 U149 ( .B(prl_cany0), .C(prl_c0set), .A(n105), .Y(n100) );
  INVX1 U150 ( .A(c0_iop), .Y(n114) );
  INVX1 U151 ( .A(n112), .Y(n113) );
  OA21X1 U152 ( .B(n73), .C(n71), .A(n105), .Y(N193) );
  AND3X1 U153 ( .A(prx_fifowdat[0]), .B(n70), .C(n69), .Y(n71) );
  NAND43X1 U154 ( .B(prx_fifowdat[3]), .C(prx_fifowdat[4]), .D(prx_fifowdat[2]), .A(n101), .Y(n72) );
  GEN2XL U155 ( .D(c0_cnt[7]), .E(n52), .C(n53), .B(n56), .A(n50), .Y(N172) );
  AND2X1 U156 ( .A(prx_fifowdat[7]), .B(n73), .Y(n50) );
  NAND42X1 U157 ( .C(pff_c0dat[47]), .D(pff_c0dat[45]), .A(n147), .B(n87), .Y(
        n85) );
  NOR3XL U158 ( .A(pff_c0dat[42]), .B(pff_c0dat[44]), .C(pff_c0dat[43]), .Y(
        n87) );
  GEN2XL U159 ( .D(c0_cnt[4]), .E(n42), .C(n43), .B(n56), .A(n41), .Y(N169) );
  AND2X1 U160 ( .A(n73), .B(prx_fifowdat[4]), .Y(n41) );
  AO22X1 U161 ( .A(N120), .B(n29), .C(prx_fifowdat[7]), .D(n59), .Y(N158) );
  NAND4X1 U162 ( .A(pff_c0dat[33]), .B(pff_c0dat[30]), .C(n96), .D(
        pff_c0dat[2]), .Y(n94) );
  AND2X1 U163 ( .A(pff_c0dat[24]), .B(pff_c0dat[21]), .Y(n96) );
  NOR3XL U164 ( .A(pff_c0dat[15]), .B(pff_c0dat[18]), .C(pff_c0dat[16]), .Y(
        n93) );
  NAND3X1 U168 ( .A(pff_c0dat[37]), .B(pff_c0dat[35]), .C(pff_c0dat[3]), .Y(
        n95) );
  GEN2XL U169 ( .D(c0_cnt[5]), .E(n45), .C(n46), .B(n56), .A(n44), .Y(N170) );
  AND2XL U170 ( .A(prx_fifowdat[5]), .B(n73), .Y(n44) );
  GEN2XL U171 ( .D(c0_cnt[6]), .E(n48), .C(n49), .B(n56), .A(n47), .Y(N171) );
  OR3XL U172 ( .A(pff_c0dat[41]), .B(pff_c0dat[39]), .C(pff_c0dat[38]), .Y(n86) );
  INVX1 U173 ( .A(prl_cany0), .Y(n147) );
  NAND2X1 U174 ( .A(pid_ccidle), .B(PrlTo[0]), .Y(n39) );
  AND3X1 U175 ( .A(ptx_ack), .B(n147), .C(n117), .Y(prl_GCTxDone) );
  AND2X1 U176 ( .A(r_auto_discard), .B(PrlTo[1]), .Y(n68) );
  INVX1 U177 ( .A(n146), .Y(prl_discard) );
  NAND21X1 U178 ( .B(n97), .A(pid_ccidle), .Y(n111) );
  NAND32XL U179 ( .B(prl_fsm[1]), .C(n58), .A(n24), .Y(n78) );
  AND2X1 U180 ( .A(n73), .B(prx_fifowdat[2]), .Y(n33) );
  AND2X1 U181 ( .A(n73), .B(prx_fifowdat[3]), .Y(n36) );
  NOR21XL U182 ( .B(n56), .A(n12), .Y(N173) );
  AOI21XL U183 ( .B(c0_cnt[8]), .C(n55), .A(n122), .Y(n12) );
  GEN2XL U184 ( .D(c0_cnt[1]), .E(c0_cnt[0]), .C(n32), .B(n56), .A(n31), .Y(
        N166) );
  AND2X1 U185 ( .A(prx_fifowdat[1]), .B(n73), .Y(n31) );
  AO22X1 U186 ( .A(N113), .B(n29), .C(prx_fifowdat[0]), .D(n59), .Y(N151) );
  AO22X1 U187 ( .A(N114), .B(n29), .C(prx_fifowdat[1]), .D(n59), .Y(N152) );
  AO22X1 U188 ( .A(N115), .B(n29), .C(n59), .D(prx_fifowdat[2]), .Y(N153) );
  OAI22XL U189 ( .A(n97), .B(n28), .C(c0_cnt[0]), .D(n108), .Y(N165) );
  INVX1 U190 ( .A(prx_fifowdat[0]), .Y(n28) );
  AO22XL U191 ( .A(n115), .B(n114), .C(n113), .D(prx_fifopsh), .Y(N194) );
  AOI32XL U192 ( .A(n72), .B(prx_fifopsh), .C(n70), .D(ptx_ack), .E(n121), .Y(
        n19) );
  AO22XL U193 ( .A(N119), .B(n29), .C(prx_fifowdat[6]), .D(n59), .Y(N157) );
  AND2XL U194 ( .A(prx_fifowdat[6]), .B(n73), .Y(n47) );
  NOR3XL U195 ( .A(prx_fifowdat[5]), .B(prx_fifowdat[7]), .C(prx_fifowdat[6]), 
        .Y(n101) );
  INVXL U196 ( .A(prl_cany0r), .Y(n116) );
  AND2XL U197 ( .A(n105), .B(prl_cany0r), .Y(N196) );
  GEN2XL U198 ( .D(c0_cnt[3]), .E(n38), .C(n40), .B(n56), .A(n36), .Y(N168) );
  GEN2XL U199 ( .D(c0_cnt[2]), .E(n34), .C(n35), .B(n56), .A(n33), .Y(N167) );
  AOI31XL U200 ( .A(n111), .B(n118), .C(n110), .D(n109), .Y(n115) );
endmodule


module updprl_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module PrlTimer_1112a0 ( to, restart, stop, clk, srstz, test_si, test_so, 
        test_se );
  output [1:0] to;
  input restart, stop, clk, srstz, test_si, test_se;
  output test_so;
  wire   timer_10_, timer_9_, timer_8_, timer_7_, timer_6_, timer_5_, timer_4_,
         timer_3_, timer_2_, timer_1_, timer_0_, ena, N4, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, net10434, n7, n8, n9, n10, n11, n12, n13, n1,
         n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 clk_gate_timer_reg ( .CLK(clk), .EN(N18), .ENCLK(net10434), .TE(test_se) );
  PrlTimer_1112a0_DW01_inc_0 add_25 ( .A({test_so, timer_10_, timer_9_, 
        timer_8_, timer_7_, timer_6_, timer_5_, timer_4_, timer_3_, timer_2_, 
        timer_1_, timer_0_}), .SUM({N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, N4}) );
  SDFFQX1 ena_reg ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .Q(ena) );
  SDFFQX1 timer_reg_1_ ( .D(N20), .SIN(timer_0_), .SMC(test_se), .C(net10434), 
        .Q(timer_1_) );
  SDFFQX1 timer_reg_2_ ( .D(N21), .SIN(timer_1_), .SMC(test_se), .C(net10434), 
        .Q(timer_2_) );
  SDFFQX1 timer_reg_0_ ( .D(N19), .SIN(ena), .SMC(test_se), .C(net10434), .Q(
        timer_0_) );
  SDFFQX1 timer_reg_11_ ( .D(N30), .SIN(timer_10_), .SMC(test_se), .C(net10434), .Q(test_so) );
  SDFFQX1 timer_reg_9_ ( .D(N28), .SIN(timer_8_), .SMC(test_se), .C(net10434), 
        .Q(timer_9_) );
  SDFFQX1 timer_reg_10_ ( .D(N29), .SIN(timer_9_), .SMC(test_se), .C(net10434), 
        .Q(timer_10_) );
  SDFFQX1 timer_reg_7_ ( .D(N26), .SIN(timer_6_), .SMC(test_se), .C(net10434), 
        .Q(timer_7_) );
  SDFFQX1 timer_reg_6_ ( .D(N25), .SIN(timer_5_), .SMC(test_se), .C(net10434), 
        .Q(timer_6_) );
  SDFFQX1 timer_reg_8_ ( .D(N27), .SIN(timer_7_), .SMC(test_se), .C(net10434), 
        .Q(timer_8_) );
  SDFFQX1 timer_reg_3_ ( .D(N22), .SIN(timer_2_), .SMC(test_se), .C(net10434), 
        .Q(timer_3_) );
  SDFFQX1 timer_reg_4_ ( .D(N23), .SIN(timer_3_), .SMC(test_se), .C(net10434), 
        .Q(timer_4_) );
  SDFFQX1 timer_reg_5_ ( .D(N24), .SIN(timer_4_), .SMC(test_se), .C(net10434), 
        .Q(timer_5_) );
  BUFX3 U3 ( .A(n11), .Y(n1) );
  NOR21XL U4 ( .B(N9), .A(n11), .Y(N24) );
  NOR21XL U5 ( .B(N7), .A(n11), .Y(N22) );
  NOR21XL U6 ( .B(N8), .A(n11), .Y(N23) );
  NOR21XL U7 ( .B(N14), .A(n11), .Y(N29) );
  NOR21XL U8 ( .B(N13), .A(n11), .Y(N28) );
  NOR21XL U9 ( .B(N12), .A(n11), .Y(N27) );
  NOR21XL U10 ( .B(N11), .A(n11), .Y(N26) );
  NOR21XL U11 ( .B(N10), .A(n11), .Y(N25) );
  NOR21XL U12 ( .B(N6), .A(n11), .Y(N21) );
  NOR21XL U13 ( .B(N5), .A(n1), .Y(N20) );
  NAND31X1 U14 ( .C(restart), .A(n1), .B(srstz), .Y(N18) );
  NAND3X1 U15 ( .A(srstz), .B(ena), .C(n12), .Y(n11) );
  NOR3XL U16 ( .A(to[1]), .B(stop), .C(restart), .Y(n12) );
  NOR21XL U17 ( .B(N15), .A(n1), .Y(N30) );
  NOR21XL U18 ( .B(N4), .A(n1), .Y(N19) );
  INVX1 U19 ( .A(n10), .Y(n2) );
  AOI31X1 U20 ( .A(srstz), .B(n3), .C(ena), .D(restart), .Y(n10) );
  INVX1 U21 ( .A(stop), .Y(n3) );
  INVX1 U22 ( .A(n7), .Y(to[0]) );
  AOI211X1 U23 ( .C(n4), .D(timer_9_), .A(timer_10_), .B(test_so), .Y(n7) );
  INVX1 U24 ( .A(n8), .Y(n4) );
  AOI211X1 U25 ( .C(timer_6_), .D(n9), .A(timer_8_), .B(timer_7_), .Y(n8) );
  AO21X1 U26 ( .B(timer_4_), .C(timer_3_), .A(timer_5_), .Y(n9) );
  OAI31XL U27 ( .A(timer_10_), .B(timer_9_), .C(timer_8_), .D(test_so), .Y(n13) );
  INVX1 U28 ( .A(n13), .Y(to[1]) );
endmodule


module PrlTimer_1112a0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyff_DEPTH_NUM34_DEPTH_NBT6 ( r_psh, r_pop, prx_psh, ptx_pop, r_last, 
        r_unlock, i_lockena, r_fiforst, i_ccidle, r_wdat, prx_wdat, txreq, 
        ffack, rdat0, full, empty, one, half, obsd, dat_7_1, ptr, fifowdat, 
        fifopsh, clk, srstz, test_si, test_se );
  input [7:0] r_wdat;
  input [7:0] prx_wdat;
  output [1:0] ffack;
  output [7:0] rdat0;
  output [55:0] dat_7_1;
  output [5:0] ptr;
  output [7:0] fifowdat;
  input r_psh, r_pop, prx_psh, ptx_pop, r_last, r_unlock, i_lockena, r_fiforst,
         i_ccidle, clk, srstz, test_si, test_se;
  output txreq, full, empty, one, half, obsd, fifopsh;
  wire   ps_locked, locked, mem_8__7_, mem_8__6_, mem_8__5_, mem_8__4_,
         mem_8__3_, mem_8__2_, mem_8__1_, mem_8__0_, mem_9__7_, mem_9__6_,
         mem_9__5_, mem_9__4_, mem_9__3_, mem_9__2_, mem_9__1_, mem_9__0_,
         mem_10__7_, mem_10__6_, mem_10__5_, mem_10__4_, mem_10__3_,
         mem_10__2_, mem_10__1_, mem_10__0_, mem_11__7_, mem_11__6_,
         mem_11__5_, mem_11__4_, mem_11__3_, mem_11__2_, mem_11__1_,
         mem_11__0_, mem_12__7_, mem_12__6_, mem_12__5_, mem_12__4_,
         mem_12__3_, mem_12__2_, mem_12__1_, mem_12__0_, mem_13__7_,
         mem_13__6_, mem_13__5_, mem_13__4_, mem_13__3_, mem_13__2_,
         mem_13__1_, mem_13__0_, mem_14__7_, mem_14__6_, mem_14__5_,
         mem_14__4_, mem_14__3_, mem_14__2_, mem_14__1_, mem_14__0_,
         mem_15__7_, mem_15__6_, mem_15__5_, mem_15__4_, mem_15__3_,
         mem_15__2_, mem_15__1_, mem_15__0_, mem_16__7_, mem_16__6_,
         mem_16__5_, mem_16__4_, mem_16__3_, mem_16__2_, mem_16__1_,
         mem_16__0_, mem_17__7_, mem_17__6_, mem_17__5_, mem_17__4_,
         mem_17__3_, mem_17__2_, mem_17__1_, mem_17__0_, mem_18__7_,
         mem_18__6_, mem_18__5_, mem_18__4_, mem_18__3_, mem_18__2_,
         mem_18__1_, mem_18__0_, mem_19__7_, mem_19__6_, mem_19__5_,
         mem_19__4_, mem_19__3_, mem_19__2_, mem_19__1_, mem_19__0_,
         mem_20__7_, mem_20__6_, mem_20__5_, mem_20__4_, mem_20__3_,
         mem_20__2_, mem_20__1_, mem_20__0_, mem_21__7_, mem_21__6_,
         mem_21__5_, mem_21__4_, mem_21__3_, mem_21__2_, mem_21__1_,
         mem_21__0_, mem_22__7_, mem_22__6_, mem_22__5_, mem_22__4_,
         mem_22__3_, mem_22__2_, mem_22__1_, mem_22__0_, mem_23__7_,
         mem_23__6_, mem_23__5_, mem_23__4_, mem_23__3_, mem_23__2_,
         mem_23__1_, mem_23__0_, mem_24__7_, mem_24__6_, mem_24__5_,
         mem_24__4_, mem_24__3_, mem_24__2_, mem_24__1_, mem_24__0_,
         mem_25__7_, mem_25__6_, mem_25__5_, mem_25__4_, mem_25__3_,
         mem_25__2_, mem_25__1_, mem_25__0_, mem_26__7_, mem_26__6_,
         mem_26__5_, mem_26__4_, mem_26__3_, mem_26__2_, mem_26__1_,
         mem_26__0_, mem_27__7_, mem_27__6_, mem_27__5_, mem_27__4_,
         mem_27__3_, mem_27__2_, mem_27__1_, mem_27__0_, mem_28__7_,
         mem_28__6_, mem_28__5_, mem_28__4_, mem_28__3_, mem_28__2_,
         mem_28__1_, mem_28__0_, mem_29__7_, mem_29__6_, mem_29__5_,
         mem_29__4_, mem_29__3_, mem_29__2_, mem_29__1_, mem_29__0_,
         mem_30__7_, mem_30__6_, mem_30__5_, mem_30__4_, mem_30__3_,
         mem_30__2_, mem_30__1_, mem_30__0_, mem_31__7_, mem_31__6_,
         mem_31__5_, mem_31__4_, mem_31__3_, mem_31__2_, mem_31__1_,
         mem_31__0_, mem_32__7_, mem_32__6_, mem_32__5_, mem_32__4_,
         mem_32__3_, mem_32__2_, mem_32__1_, mem_32__0_, mem_33__7_,
         mem_33__6_, mem_33__5_, mem_33__4_, mem_33__3_, mem_33__2_,
         mem_33__1_, mem_33__0_, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1053, N1054, N1055,
         N1056, N1057, N1058, N1059, net10452, net10458, net10463, net10468,
         net10473, net10478, net10483, net10488, net10493, net10498, net10503,
         net10508, net10513, net10518, net10523, net10528, net10533, net10538,
         net10543, net10548, net10553, net10558, net10563, net10568, net10573,
         net10578, net10583, net10588, net10593, net10598, net10603, net10608,
         net10613, net10618, net10623, n48, n50, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n436, n442,
         n443, n444, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38,
         n39, n40, n42, n43, n44, n45, n46, n47, n49, n66, n92, n105, n141,
         n142, n154, n165, n176, n187, n199, n211, n223, n245, n246, n257,
         n268, n280, n291, n335, n348, n349, n383, n384, n419, n420, n421,
         n422, n423, n424, n425, n427, n428, n429, n430, n431, n432, n433,
         n435, n437, n438, n439, n440, n441, n445, n446, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555;

  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 clk_gate_mem_reg_0_ ( 
        .CLK(clk), .EN(N1022), .ENCLK(net10452), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 clk_gate_mem_reg_1_ ( 
        .CLK(clk), .EN(N1013), .ENCLK(net10458), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 clk_gate_mem_reg_2_ ( 
        .CLK(clk), .EN(N1004), .ENCLK(net10463), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 clk_gate_mem_reg_3_ ( 
        .CLK(clk), .EN(N995), .ENCLK(net10468), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 clk_gate_mem_reg_4_ ( 
        .CLK(clk), .EN(N986), .ENCLK(net10473), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 clk_gate_mem_reg_5_ ( 
        .CLK(clk), .EN(N977), .ENCLK(net10478), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 clk_gate_mem_reg_6_ ( 
        .CLK(clk), .EN(N968), .ENCLK(net10483), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 clk_gate_mem_reg_7_ ( 
        .CLK(clk), .EN(N959), .ENCLK(net10488), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 clk_gate_mem_reg_8_ ( 
        .CLK(clk), .EN(N950), .ENCLK(net10493), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 clk_gate_mem_reg_9_ ( 
        .CLK(clk), .EN(N941), .ENCLK(net10498), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 clk_gate_mem_reg_10_ ( 
        .CLK(clk), .EN(N932), .ENCLK(net10503), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 clk_gate_mem_reg_11_ ( 
        .CLK(clk), .EN(N923), .ENCLK(net10508), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 clk_gate_mem_reg_12_ ( 
        .CLK(clk), .EN(N914), .ENCLK(net10513), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 clk_gate_mem_reg_13_ ( 
        .CLK(clk), .EN(N905), .ENCLK(net10518), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 clk_gate_mem_reg_14_ ( 
        .CLK(clk), .EN(N896), .ENCLK(net10523), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 clk_gate_mem_reg_15_ ( 
        .CLK(clk), .EN(N887), .ENCLK(net10528), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 clk_gate_mem_reg_16_ ( 
        .CLK(clk), .EN(N878), .ENCLK(net10533), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 clk_gate_mem_reg_17_ ( 
        .CLK(clk), .EN(N869), .ENCLK(net10538), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 clk_gate_mem_reg_18_ ( 
        .CLK(clk), .EN(N860), .ENCLK(net10543), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 clk_gate_mem_reg_19_ ( 
        .CLK(clk), .EN(N851), .ENCLK(net10548), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 clk_gate_mem_reg_20_ ( 
        .CLK(clk), .EN(N842), .ENCLK(net10553), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 clk_gate_mem_reg_21_ ( 
        .CLK(clk), .EN(N833), .ENCLK(net10558), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 clk_gate_mem_reg_22_ ( 
        .CLK(clk), .EN(N824), .ENCLK(net10563), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 clk_gate_mem_reg_23_ ( 
        .CLK(clk), .EN(N815), .ENCLK(net10568), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 clk_gate_mem_reg_24_ ( 
        .CLK(clk), .EN(N806), .ENCLK(net10573), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 clk_gate_mem_reg_25_ ( 
        .CLK(clk), .EN(N797), .ENCLK(net10578), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 clk_gate_mem_reg_26_ ( 
        .CLK(clk), .EN(N788), .ENCLK(net10583), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 clk_gate_mem_reg_27_ ( 
        .CLK(clk), .EN(N779), .ENCLK(net10588), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 clk_gate_mem_reg_28_ ( 
        .CLK(clk), .EN(N770), .ENCLK(net10593), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 clk_gate_mem_reg_29_ ( 
        .CLK(clk), .EN(N761), .ENCLK(net10598), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 clk_gate_mem_reg_30_ ( 
        .CLK(clk), .EN(N752), .ENCLK(net10603), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 clk_gate_mem_reg_31_ ( 
        .CLK(clk), .EN(N743), .ENCLK(net10608), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 clk_gate_mem_reg_32_ ( 
        .CLK(clk), .EN(N734), .ENCLK(net10613), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 clk_gate_mem_reg_33_ ( 
        .CLK(clk), .EN(N733), .ENCLK(net10618), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 clk_gate_pshptr_reg ( 
        .CLK(clk), .EN(N1053), .ENCLK(net10623), .TE(test_se) );
  SDFFQX1 mem_reg_33__7_ ( .D(fifowdat[7]), .SIN(mem_33__6_), .SMC(test_se), 
        .C(net10618), .Q(mem_33__7_) );
  SDFFQX1 mem_reg_32__7_ ( .D(N742), .SIN(mem_32__6_), .SMC(test_se), .C(
        net10613), .Q(mem_32__7_) );
  SDFFQX1 mem_reg_31__7_ ( .D(N751), .SIN(mem_31__6_), .SMC(test_se), .C(
        net10608), .Q(mem_31__7_) );
  SDFFQX1 mem_reg_30__7_ ( .D(N760), .SIN(mem_30__6_), .SMC(test_se), .C(
        net10603), .Q(mem_30__7_) );
  SDFFQX1 mem_reg_29__7_ ( .D(N769), .SIN(mem_29__6_), .SMC(test_se), .C(
        net10598), .Q(mem_29__7_) );
  SDFFQX1 mem_reg_28__7_ ( .D(N778), .SIN(mem_28__6_), .SMC(test_se), .C(
        net10593), .Q(mem_28__7_) );
  SDFFQX1 mem_reg_33__6_ ( .D(fifowdat[6]), .SIN(mem_33__5_), .SMC(test_se), 
        .C(net10618), .Q(mem_33__6_) );
  SDFFQX1 mem_reg_32__6_ ( .D(N741), .SIN(mem_32__5_), .SMC(test_se), .C(
        net10613), .Q(mem_32__6_) );
  SDFFQX1 mem_reg_31__6_ ( .D(N750), .SIN(mem_31__5_), .SMC(test_se), .C(
        net10608), .Q(mem_31__6_) );
  SDFFQX1 mem_reg_30__6_ ( .D(N759), .SIN(mem_30__5_), .SMC(test_se), .C(
        net10603), .Q(mem_30__6_) );
  SDFFQX1 mem_reg_29__6_ ( .D(N768), .SIN(mem_29__5_), .SMC(test_se), .C(
        net10598), .Q(mem_29__6_) );
  SDFFQX1 mem_reg_28__6_ ( .D(N777), .SIN(mem_28__5_), .SMC(test_se), .C(
        net10593), .Q(mem_28__6_) );
  SDFFQX1 mem_reg_33__5_ ( .D(fifowdat[5]), .SIN(mem_33__4_), .SMC(test_se), 
        .C(net10618), .Q(mem_33__5_) );
  SDFFQX1 mem_reg_32__5_ ( .D(N740), .SIN(mem_32__4_), .SMC(test_se), .C(
        net10613), .Q(mem_32__5_) );
  SDFFQX1 mem_reg_31__5_ ( .D(N749), .SIN(mem_31__4_), .SMC(test_se), .C(
        net10608), .Q(mem_31__5_) );
  SDFFQX1 mem_reg_30__5_ ( .D(N758), .SIN(mem_30__4_), .SMC(test_se), .C(
        net10603), .Q(mem_30__5_) );
  SDFFQX1 mem_reg_29__5_ ( .D(N767), .SIN(mem_29__4_), .SMC(test_se), .C(
        net10598), .Q(mem_29__5_) );
  SDFFQX1 mem_reg_28__5_ ( .D(N776), .SIN(mem_28__4_), .SMC(test_se), .C(
        net10593), .Q(mem_28__5_) );
  SDFFQX1 mem_reg_33__4_ ( .D(fifowdat[4]), .SIN(mem_33__3_), .SMC(test_se), 
        .C(net10618), .Q(mem_33__4_) );
  SDFFQX1 mem_reg_32__4_ ( .D(N739), .SIN(mem_32__3_), .SMC(test_se), .C(
        net10613), .Q(mem_32__4_) );
  SDFFQX1 mem_reg_31__4_ ( .D(N748), .SIN(mem_31__3_), .SMC(test_se), .C(
        net10608), .Q(mem_31__4_) );
  SDFFQX1 mem_reg_30__4_ ( .D(N757), .SIN(mem_30__3_), .SMC(test_se), .C(
        net10603), .Q(mem_30__4_) );
  SDFFQX1 mem_reg_29__4_ ( .D(N766), .SIN(mem_29__3_), .SMC(test_se), .C(
        net10598), .Q(mem_29__4_) );
  SDFFQX1 mem_reg_28__4_ ( .D(N775), .SIN(mem_28__3_), .SMC(test_se), .C(
        net10593), .Q(mem_28__4_) );
  SDFFQX1 mem_reg_33__3_ ( .D(fifowdat[3]), .SIN(mem_33__2_), .SMC(test_se), 
        .C(net10618), .Q(mem_33__3_) );
  SDFFQX1 mem_reg_32__3_ ( .D(N738), .SIN(mem_32__2_), .SMC(test_se), .C(
        net10613), .Q(mem_32__3_) );
  SDFFQX1 mem_reg_31__3_ ( .D(N747), .SIN(mem_31__2_), .SMC(test_se), .C(
        net10608), .Q(mem_31__3_) );
  SDFFQX1 mem_reg_30__3_ ( .D(N756), .SIN(mem_30__2_), .SMC(test_se), .C(
        net10603), .Q(mem_30__3_) );
  SDFFQX1 mem_reg_29__3_ ( .D(N765), .SIN(mem_29__2_), .SMC(test_se), .C(
        net10598), .Q(mem_29__3_) );
  SDFFQX1 mem_reg_28__3_ ( .D(N774), .SIN(mem_28__2_), .SMC(test_se), .C(
        net10593), .Q(mem_28__3_) );
  SDFFQX1 mem_reg_33__2_ ( .D(fifowdat[2]), .SIN(mem_33__1_), .SMC(test_se), 
        .C(net10618), .Q(mem_33__2_) );
  SDFFQX1 mem_reg_32__2_ ( .D(N737), .SIN(mem_32__1_), .SMC(test_se), .C(
        net10613), .Q(mem_32__2_) );
  SDFFQX1 mem_reg_31__2_ ( .D(N746), .SIN(mem_31__1_), .SMC(test_se), .C(
        net10608), .Q(mem_31__2_) );
  SDFFQX1 mem_reg_30__2_ ( .D(N755), .SIN(mem_30__1_), .SMC(test_se), .C(
        net10603), .Q(mem_30__2_) );
  SDFFQX1 mem_reg_29__2_ ( .D(N764), .SIN(mem_29__1_), .SMC(test_se), .C(
        net10598), .Q(mem_29__2_) );
  SDFFQX1 mem_reg_28__2_ ( .D(N773), .SIN(mem_28__1_), .SMC(test_se), .C(
        net10593), .Q(mem_28__2_) );
  SDFFQX1 mem_reg_33__1_ ( .D(fifowdat[1]), .SIN(mem_33__0_), .SMC(test_se), 
        .C(net10618), .Q(mem_33__1_) );
  SDFFQX1 mem_reg_32__1_ ( .D(N736), .SIN(mem_32__0_), .SMC(test_se), .C(
        net10613), .Q(mem_32__1_) );
  SDFFQX1 mem_reg_31__1_ ( .D(N745), .SIN(mem_31__0_), .SMC(test_se), .C(
        net10608), .Q(mem_31__1_) );
  SDFFQX1 mem_reg_30__1_ ( .D(N754), .SIN(mem_30__0_), .SMC(test_se), .C(
        net10603), .Q(mem_30__1_) );
  SDFFQX1 mem_reg_29__1_ ( .D(N763), .SIN(mem_29__0_), .SMC(test_se), .C(
        net10598), .Q(mem_29__1_) );
  SDFFQX1 mem_reg_28__1_ ( .D(N772), .SIN(mem_28__0_), .SMC(test_se), .C(
        net10593), .Q(mem_28__1_) );
  SDFFQX1 mem_reg_33__0_ ( .D(fifowdat[0]), .SIN(mem_32__7_), .SMC(test_se), 
        .C(net10618), .Q(mem_33__0_) );
  SDFFQX1 mem_reg_32__0_ ( .D(N735), .SIN(mem_31__7_), .SMC(test_se), .C(
        net10613), .Q(mem_32__0_) );
  SDFFQX1 mem_reg_31__0_ ( .D(N744), .SIN(mem_30__7_), .SMC(test_se), .C(
        net10608), .Q(mem_31__0_) );
  SDFFQX1 mem_reg_30__0_ ( .D(N753), .SIN(mem_29__7_), .SMC(test_se), .C(
        net10603), .Q(mem_30__0_) );
  SDFFQX1 mem_reg_29__0_ ( .D(N762), .SIN(mem_28__7_), .SMC(test_se), .C(
        net10598), .Q(mem_29__0_) );
  SDFFQX1 mem_reg_28__0_ ( .D(N771), .SIN(mem_27__7_), .SMC(test_se), .C(
        net10593), .Q(mem_28__0_) );
  SDFFQX1 mem_reg_27__7_ ( .D(N787), .SIN(mem_27__6_), .SMC(test_se), .C(
        net10588), .Q(mem_27__7_) );
  SDFFQX1 mem_reg_26__7_ ( .D(N796), .SIN(mem_26__6_), .SMC(test_se), .C(
        net10583), .Q(mem_26__7_) );
  SDFFQX1 mem_reg_25__7_ ( .D(N805), .SIN(mem_25__6_), .SMC(test_se), .C(
        net10578), .Q(mem_25__7_) );
  SDFFQX1 mem_reg_24__7_ ( .D(N814), .SIN(mem_24__6_), .SMC(test_se), .C(
        net10573), .Q(mem_24__7_) );
  SDFFQX1 mem_reg_23__7_ ( .D(N823), .SIN(mem_23__6_), .SMC(test_se), .C(
        net10568), .Q(mem_23__7_) );
  SDFFQX1 mem_reg_22__7_ ( .D(N832), .SIN(mem_22__6_), .SMC(test_se), .C(
        net10563), .Q(mem_22__7_) );
  SDFFQX1 mem_reg_21__7_ ( .D(N841), .SIN(mem_21__6_), .SMC(test_se), .C(
        net10558), .Q(mem_21__7_) );
  SDFFQX1 mem_reg_20__7_ ( .D(N850), .SIN(mem_20__6_), .SMC(test_se), .C(
        net10553), .Q(mem_20__7_) );
  SDFFQX1 mem_reg_19__7_ ( .D(N859), .SIN(mem_19__6_), .SMC(test_se), .C(
        net10548), .Q(mem_19__7_) );
  SDFFQX1 mem_reg_18__7_ ( .D(N868), .SIN(mem_18__6_), .SMC(test_se), .C(
        net10543), .Q(mem_18__7_) );
  SDFFQX1 mem_reg_17__7_ ( .D(N877), .SIN(mem_17__6_), .SMC(test_se), .C(
        net10538), .Q(mem_17__7_) );
  SDFFQX1 mem_reg_16__7_ ( .D(N886), .SIN(mem_16__6_), .SMC(test_se), .C(
        net10533), .Q(mem_16__7_) );
  SDFFQX1 mem_reg_15__7_ ( .D(N895), .SIN(mem_15__6_), .SMC(test_se), .C(
        net10528), .Q(mem_15__7_) );
  SDFFQX1 mem_reg_14__7_ ( .D(N904), .SIN(mem_14__6_), .SMC(test_se), .C(
        net10523), .Q(mem_14__7_) );
  SDFFQX1 mem_reg_13__7_ ( .D(N913), .SIN(mem_13__6_), .SMC(test_se), .C(
        net10518), .Q(mem_13__7_) );
  SDFFQX1 mem_reg_12__7_ ( .D(N922), .SIN(mem_12__6_), .SMC(test_se), .C(
        net10513), .Q(mem_12__7_) );
  SDFFQX1 mem_reg_11__7_ ( .D(N931), .SIN(mem_11__6_), .SMC(test_se), .C(
        net10508), .Q(mem_11__7_) );
  SDFFQX1 mem_reg_10__7_ ( .D(N940), .SIN(mem_10__6_), .SMC(test_se), .C(
        net10503), .Q(mem_10__7_) );
  SDFFQX1 mem_reg_9__7_ ( .D(N949), .SIN(mem_9__6_), .SMC(test_se), .C(
        net10498), .Q(mem_9__7_) );
  SDFFQX1 mem_reg_8__7_ ( .D(N958), .SIN(mem_8__6_), .SMC(test_se), .C(
        net10493), .Q(mem_8__7_) );
  SDFFQX1 mem_reg_27__6_ ( .D(N786), .SIN(mem_27__5_), .SMC(test_se), .C(
        net10588), .Q(mem_27__6_) );
  SDFFQX1 mem_reg_26__6_ ( .D(N795), .SIN(mem_26__5_), .SMC(test_se), .C(
        net10583), .Q(mem_26__6_) );
  SDFFQX1 mem_reg_25__6_ ( .D(N804), .SIN(mem_25__5_), .SMC(test_se), .C(
        net10578), .Q(mem_25__6_) );
  SDFFQX1 mem_reg_24__6_ ( .D(N813), .SIN(mem_24__5_), .SMC(test_se), .C(
        net10573), .Q(mem_24__6_) );
  SDFFQX1 mem_reg_23__6_ ( .D(N822), .SIN(mem_23__5_), .SMC(test_se), .C(
        net10568), .Q(mem_23__6_) );
  SDFFQX1 mem_reg_22__6_ ( .D(N831), .SIN(mem_22__5_), .SMC(test_se), .C(
        net10563), .Q(mem_22__6_) );
  SDFFQX1 mem_reg_21__6_ ( .D(N840), .SIN(mem_21__5_), .SMC(test_se), .C(
        net10558), .Q(mem_21__6_) );
  SDFFQX1 mem_reg_20__6_ ( .D(N849), .SIN(mem_20__5_), .SMC(test_se), .C(
        net10553), .Q(mem_20__6_) );
  SDFFQX1 mem_reg_19__6_ ( .D(N858), .SIN(mem_19__5_), .SMC(test_se), .C(
        net10548), .Q(mem_19__6_) );
  SDFFQX1 mem_reg_18__6_ ( .D(N867), .SIN(mem_18__5_), .SMC(test_se), .C(
        net10543), .Q(mem_18__6_) );
  SDFFQX1 mem_reg_17__6_ ( .D(N876), .SIN(mem_17__5_), .SMC(test_se), .C(
        net10538), .Q(mem_17__6_) );
  SDFFQX1 mem_reg_16__6_ ( .D(N885), .SIN(mem_16__5_), .SMC(test_se), .C(
        net10533), .Q(mem_16__6_) );
  SDFFQX1 mem_reg_15__6_ ( .D(N894), .SIN(mem_15__5_), .SMC(test_se), .C(
        net10528), .Q(mem_15__6_) );
  SDFFQX1 mem_reg_14__6_ ( .D(N903), .SIN(mem_14__5_), .SMC(test_se), .C(
        net10523), .Q(mem_14__6_) );
  SDFFQX1 mem_reg_13__6_ ( .D(N912), .SIN(mem_13__5_), .SMC(test_se), .C(
        net10518), .Q(mem_13__6_) );
  SDFFQX1 mem_reg_12__6_ ( .D(N921), .SIN(mem_12__5_), .SMC(test_se), .C(
        net10513), .Q(mem_12__6_) );
  SDFFQX1 mem_reg_11__6_ ( .D(N930), .SIN(mem_11__5_), .SMC(test_se), .C(
        net10508), .Q(mem_11__6_) );
  SDFFQX1 mem_reg_10__6_ ( .D(N939), .SIN(mem_10__5_), .SMC(test_se), .C(
        net10503), .Q(mem_10__6_) );
  SDFFQX1 mem_reg_9__6_ ( .D(N948), .SIN(mem_9__5_), .SMC(test_se), .C(
        net10498), .Q(mem_9__6_) );
  SDFFQX1 mem_reg_8__6_ ( .D(N957), .SIN(mem_8__5_), .SMC(test_se), .C(
        net10493), .Q(mem_8__6_) );
  SDFFQX1 mem_reg_27__5_ ( .D(N785), .SIN(mem_27__4_), .SMC(test_se), .C(
        net10588), .Q(mem_27__5_) );
  SDFFQX1 mem_reg_26__5_ ( .D(N794), .SIN(mem_26__4_), .SMC(test_se), .C(
        net10583), .Q(mem_26__5_) );
  SDFFQX1 mem_reg_25__5_ ( .D(N803), .SIN(mem_25__4_), .SMC(test_se), .C(
        net10578), .Q(mem_25__5_) );
  SDFFQX1 mem_reg_24__5_ ( .D(N812), .SIN(mem_24__4_), .SMC(test_se), .C(
        net10573), .Q(mem_24__5_) );
  SDFFQX1 mem_reg_23__5_ ( .D(N821), .SIN(mem_23__4_), .SMC(test_se), .C(
        net10568), .Q(mem_23__5_) );
  SDFFQX1 mem_reg_22__5_ ( .D(N830), .SIN(mem_22__4_), .SMC(test_se), .C(
        net10563), .Q(mem_22__5_) );
  SDFFQX1 mem_reg_21__5_ ( .D(N839), .SIN(mem_21__4_), .SMC(test_se), .C(
        net10558), .Q(mem_21__5_) );
  SDFFQX1 mem_reg_20__5_ ( .D(N848), .SIN(mem_20__4_), .SMC(test_se), .C(
        net10553), .Q(mem_20__5_) );
  SDFFQX1 mem_reg_19__5_ ( .D(N857), .SIN(mem_19__4_), .SMC(test_se), .C(
        net10548), .Q(mem_19__5_) );
  SDFFQX1 mem_reg_18__5_ ( .D(N866), .SIN(mem_18__4_), .SMC(test_se), .C(
        net10543), .Q(mem_18__5_) );
  SDFFQX1 mem_reg_17__5_ ( .D(N875), .SIN(mem_17__4_), .SMC(test_se), .C(
        net10538), .Q(mem_17__5_) );
  SDFFQX1 mem_reg_16__5_ ( .D(N884), .SIN(mem_16__4_), .SMC(test_se), .C(
        net10533), .Q(mem_16__5_) );
  SDFFQX1 mem_reg_15__5_ ( .D(N893), .SIN(mem_15__4_), .SMC(test_se), .C(
        net10528), .Q(mem_15__5_) );
  SDFFQX1 mem_reg_14__5_ ( .D(N902), .SIN(mem_14__4_), .SMC(test_se), .C(
        net10523), .Q(mem_14__5_) );
  SDFFQX1 mem_reg_13__5_ ( .D(N911), .SIN(mem_13__4_), .SMC(test_se), .C(
        net10518), .Q(mem_13__5_) );
  SDFFQX1 mem_reg_12__5_ ( .D(N920), .SIN(mem_12__4_), .SMC(test_se), .C(
        net10513), .Q(mem_12__5_) );
  SDFFQX1 mem_reg_11__5_ ( .D(N929), .SIN(mem_11__4_), .SMC(test_se), .C(
        net10508), .Q(mem_11__5_) );
  SDFFQX1 mem_reg_10__5_ ( .D(N938), .SIN(mem_10__4_), .SMC(test_se), .C(
        net10503), .Q(mem_10__5_) );
  SDFFQX1 mem_reg_9__5_ ( .D(N947), .SIN(mem_9__4_), .SMC(test_se), .C(
        net10498), .Q(mem_9__5_) );
  SDFFQX1 mem_reg_8__5_ ( .D(N956), .SIN(mem_8__4_), .SMC(test_se), .C(
        net10493), .Q(mem_8__5_) );
  SDFFQX1 mem_reg_27__4_ ( .D(N784), .SIN(mem_27__3_), .SMC(test_se), .C(
        net10588), .Q(mem_27__4_) );
  SDFFQX1 mem_reg_26__4_ ( .D(N793), .SIN(mem_26__3_), .SMC(test_se), .C(
        net10583), .Q(mem_26__4_) );
  SDFFQX1 mem_reg_25__4_ ( .D(N802), .SIN(mem_25__3_), .SMC(test_se), .C(
        net10578), .Q(mem_25__4_) );
  SDFFQX1 mem_reg_24__4_ ( .D(N811), .SIN(mem_24__3_), .SMC(test_se), .C(
        net10573), .Q(mem_24__4_) );
  SDFFQX1 mem_reg_23__4_ ( .D(N820), .SIN(mem_23__3_), .SMC(test_se), .C(
        net10568), .Q(mem_23__4_) );
  SDFFQX1 mem_reg_22__4_ ( .D(N829), .SIN(mem_22__3_), .SMC(test_se), .C(
        net10563), .Q(mem_22__4_) );
  SDFFQX1 mem_reg_21__4_ ( .D(N838), .SIN(mem_21__3_), .SMC(test_se), .C(
        net10558), .Q(mem_21__4_) );
  SDFFQX1 mem_reg_20__4_ ( .D(N847), .SIN(mem_20__3_), .SMC(test_se), .C(
        net10553), .Q(mem_20__4_) );
  SDFFQX1 mem_reg_19__4_ ( .D(N856), .SIN(mem_19__3_), .SMC(test_se), .C(
        net10548), .Q(mem_19__4_) );
  SDFFQX1 mem_reg_18__4_ ( .D(N865), .SIN(mem_18__3_), .SMC(test_se), .C(
        net10543), .Q(mem_18__4_) );
  SDFFQX1 mem_reg_17__4_ ( .D(N874), .SIN(mem_17__3_), .SMC(test_se), .C(
        net10538), .Q(mem_17__4_) );
  SDFFQX1 mem_reg_16__4_ ( .D(N883), .SIN(mem_16__3_), .SMC(test_se), .C(
        net10533), .Q(mem_16__4_) );
  SDFFQX1 mem_reg_15__4_ ( .D(N892), .SIN(mem_15__3_), .SMC(test_se), .C(
        net10528), .Q(mem_15__4_) );
  SDFFQX1 mem_reg_14__4_ ( .D(N901), .SIN(mem_14__3_), .SMC(test_se), .C(
        net10523), .Q(mem_14__4_) );
  SDFFQX1 mem_reg_13__4_ ( .D(N910), .SIN(mem_13__3_), .SMC(test_se), .C(
        net10518), .Q(mem_13__4_) );
  SDFFQX1 mem_reg_12__4_ ( .D(N919), .SIN(mem_12__3_), .SMC(test_se), .C(
        net10513), .Q(mem_12__4_) );
  SDFFQX1 mem_reg_11__4_ ( .D(N928), .SIN(mem_11__3_), .SMC(test_se), .C(
        net10508), .Q(mem_11__4_) );
  SDFFQX1 mem_reg_10__4_ ( .D(N937), .SIN(mem_10__3_), .SMC(test_se), .C(
        net10503), .Q(mem_10__4_) );
  SDFFQX1 mem_reg_9__4_ ( .D(N946), .SIN(mem_9__3_), .SMC(test_se), .C(
        net10498), .Q(mem_9__4_) );
  SDFFQX1 mem_reg_8__4_ ( .D(N955), .SIN(mem_8__3_), .SMC(test_se), .C(
        net10493), .Q(mem_8__4_) );
  SDFFQX1 mem_reg_27__3_ ( .D(N783), .SIN(mem_27__2_), .SMC(test_se), .C(
        net10588), .Q(mem_27__3_) );
  SDFFQX1 mem_reg_26__3_ ( .D(N792), .SIN(mem_26__2_), .SMC(test_se), .C(
        net10583), .Q(mem_26__3_) );
  SDFFQX1 mem_reg_25__3_ ( .D(N801), .SIN(mem_25__2_), .SMC(test_se), .C(
        net10578), .Q(mem_25__3_) );
  SDFFQX1 mem_reg_24__3_ ( .D(N810), .SIN(mem_24__2_), .SMC(test_se), .C(
        net10573), .Q(mem_24__3_) );
  SDFFQX1 mem_reg_23__3_ ( .D(N819), .SIN(mem_23__2_), .SMC(test_se), .C(
        net10568), .Q(mem_23__3_) );
  SDFFQX1 mem_reg_22__3_ ( .D(N828), .SIN(mem_22__2_), .SMC(test_se), .C(
        net10563), .Q(mem_22__3_) );
  SDFFQX1 mem_reg_21__3_ ( .D(N837), .SIN(mem_21__2_), .SMC(test_se), .C(
        net10558), .Q(mem_21__3_) );
  SDFFQX1 mem_reg_20__3_ ( .D(N846), .SIN(mem_20__2_), .SMC(test_se), .C(
        net10553), .Q(mem_20__3_) );
  SDFFQX1 mem_reg_19__3_ ( .D(N855), .SIN(mem_19__2_), .SMC(test_se), .C(
        net10548), .Q(mem_19__3_) );
  SDFFQX1 mem_reg_18__3_ ( .D(N864), .SIN(mem_18__2_), .SMC(test_se), .C(
        net10543), .Q(mem_18__3_) );
  SDFFQX1 mem_reg_17__3_ ( .D(N873), .SIN(mem_17__2_), .SMC(test_se), .C(
        net10538), .Q(mem_17__3_) );
  SDFFQX1 mem_reg_16__3_ ( .D(N882), .SIN(mem_16__2_), .SMC(test_se), .C(
        net10533), .Q(mem_16__3_) );
  SDFFQX1 mem_reg_15__3_ ( .D(N891), .SIN(mem_15__2_), .SMC(test_se), .C(
        net10528), .Q(mem_15__3_) );
  SDFFQX1 mem_reg_14__3_ ( .D(N900), .SIN(mem_14__2_), .SMC(test_se), .C(
        net10523), .Q(mem_14__3_) );
  SDFFQX1 mem_reg_13__3_ ( .D(N909), .SIN(mem_13__2_), .SMC(test_se), .C(
        net10518), .Q(mem_13__3_) );
  SDFFQX1 mem_reg_12__3_ ( .D(N918), .SIN(mem_12__2_), .SMC(test_se), .C(
        net10513), .Q(mem_12__3_) );
  SDFFQX1 mem_reg_11__3_ ( .D(N927), .SIN(mem_11__2_), .SMC(test_se), .C(
        net10508), .Q(mem_11__3_) );
  SDFFQX1 mem_reg_10__3_ ( .D(N936), .SIN(mem_10__2_), .SMC(test_se), .C(
        net10503), .Q(mem_10__3_) );
  SDFFQX1 mem_reg_9__3_ ( .D(N945), .SIN(mem_9__2_), .SMC(test_se), .C(
        net10498), .Q(mem_9__3_) );
  SDFFQX1 mem_reg_8__3_ ( .D(N954), .SIN(mem_8__2_), .SMC(test_se), .C(
        net10493), .Q(mem_8__3_) );
  SDFFQX1 mem_reg_27__2_ ( .D(N782), .SIN(mem_27__1_), .SMC(test_se), .C(
        net10588), .Q(mem_27__2_) );
  SDFFQX1 mem_reg_26__2_ ( .D(N791), .SIN(mem_26__1_), .SMC(test_se), .C(
        net10583), .Q(mem_26__2_) );
  SDFFQX1 mem_reg_25__2_ ( .D(N800), .SIN(mem_25__1_), .SMC(test_se), .C(
        net10578), .Q(mem_25__2_) );
  SDFFQX1 mem_reg_24__2_ ( .D(N809), .SIN(mem_24__1_), .SMC(test_se), .C(
        net10573), .Q(mem_24__2_) );
  SDFFQX1 mem_reg_23__2_ ( .D(N818), .SIN(mem_23__1_), .SMC(test_se), .C(
        net10568), .Q(mem_23__2_) );
  SDFFQX1 mem_reg_22__2_ ( .D(N827), .SIN(mem_22__1_), .SMC(test_se), .C(
        net10563), .Q(mem_22__2_) );
  SDFFQX1 mem_reg_21__2_ ( .D(N836), .SIN(mem_21__1_), .SMC(test_se), .C(
        net10558), .Q(mem_21__2_) );
  SDFFQX1 mem_reg_20__2_ ( .D(N845), .SIN(mem_20__1_), .SMC(test_se), .C(
        net10553), .Q(mem_20__2_) );
  SDFFQX1 mem_reg_19__2_ ( .D(N854), .SIN(mem_19__1_), .SMC(test_se), .C(
        net10548), .Q(mem_19__2_) );
  SDFFQX1 mem_reg_18__2_ ( .D(N863), .SIN(mem_18__1_), .SMC(test_se), .C(
        net10543), .Q(mem_18__2_) );
  SDFFQX1 mem_reg_17__2_ ( .D(N872), .SIN(mem_17__1_), .SMC(test_se), .C(
        net10538), .Q(mem_17__2_) );
  SDFFQX1 mem_reg_16__2_ ( .D(N881), .SIN(mem_16__1_), .SMC(test_se), .C(
        net10533), .Q(mem_16__2_) );
  SDFFQX1 mem_reg_15__2_ ( .D(N890), .SIN(mem_15__1_), .SMC(test_se), .C(
        net10528), .Q(mem_15__2_) );
  SDFFQX1 mem_reg_14__2_ ( .D(N899), .SIN(mem_14__1_), .SMC(test_se), .C(
        net10523), .Q(mem_14__2_) );
  SDFFQX1 mem_reg_13__2_ ( .D(N908), .SIN(mem_13__1_), .SMC(test_se), .C(
        net10518), .Q(mem_13__2_) );
  SDFFQX1 mem_reg_12__2_ ( .D(N917), .SIN(mem_12__1_), .SMC(test_se), .C(
        net10513), .Q(mem_12__2_) );
  SDFFQX1 mem_reg_11__2_ ( .D(N926), .SIN(mem_11__1_), .SMC(test_se), .C(
        net10508), .Q(mem_11__2_) );
  SDFFQX1 mem_reg_10__2_ ( .D(N935), .SIN(mem_10__1_), .SMC(test_se), .C(
        net10503), .Q(mem_10__2_) );
  SDFFQX1 mem_reg_9__2_ ( .D(N944), .SIN(mem_9__1_), .SMC(test_se), .C(
        net10498), .Q(mem_9__2_) );
  SDFFQX1 mem_reg_8__2_ ( .D(N953), .SIN(mem_8__1_), .SMC(test_se), .C(
        net10493), .Q(mem_8__2_) );
  SDFFQX1 mem_reg_27__1_ ( .D(N781), .SIN(mem_27__0_), .SMC(test_se), .C(
        net10588), .Q(mem_27__1_) );
  SDFFQX1 mem_reg_26__1_ ( .D(N790), .SIN(mem_26__0_), .SMC(test_se), .C(
        net10583), .Q(mem_26__1_) );
  SDFFQX1 mem_reg_25__1_ ( .D(N799), .SIN(mem_25__0_), .SMC(test_se), .C(
        net10578), .Q(mem_25__1_) );
  SDFFQX1 mem_reg_24__1_ ( .D(N808), .SIN(mem_24__0_), .SMC(test_se), .C(
        net10573), .Q(mem_24__1_) );
  SDFFQX1 mem_reg_23__1_ ( .D(N817), .SIN(mem_23__0_), .SMC(test_se), .C(
        net10568), .Q(mem_23__1_) );
  SDFFQX1 mem_reg_22__1_ ( .D(N826), .SIN(mem_22__0_), .SMC(test_se), .C(
        net10563), .Q(mem_22__1_) );
  SDFFQX1 mem_reg_21__1_ ( .D(N835), .SIN(mem_21__0_), .SMC(test_se), .C(
        net10558), .Q(mem_21__1_) );
  SDFFQX1 mem_reg_20__1_ ( .D(N844), .SIN(mem_20__0_), .SMC(test_se), .C(
        net10553), .Q(mem_20__1_) );
  SDFFQX1 mem_reg_19__1_ ( .D(N853), .SIN(mem_19__0_), .SMC(test_se), .C(
        net10548), .Q(mem_19__1_) );
  SDFFQX1 mem_reg_18__1_ ( .D(N862), .SIN(mem_18__0_), .SMC(test_se), .C(
        net10543), .Q(mem_18__1_) );
  SDFFQX1 mem_reg_17__1_ ( .D(N871), .SIN(mem_17__0_), .SMC(test_se), .C(
        net10538), .Q(mem_17__1_) );
  SDFFQX1 mem_reg_16__1_ ( .D(N880), .SIN(mem_16__0_), .SMC(test_se), .C(
        net10533), .Q(mem_16__1_) );
  SDFFQX1 mem_reg_15__1_ ( .D(N889), .SIN(mem_15__0_), .SMC(test_se), .C(
        net10528), .Q(mem_15__1_) );
  SDFFQX1 mem_reg_14__1_ ( .D(N898), .SIN(mem_14__0_), .SMC(test_se), .C(
        net10523), .Q(mem_14__1_) );
  SDFFQX1 mem_reg_13__1_ ( .D(N907), .SIN(mem_13__0_), .SMC(test_se), .C(
        net10518), .Q(mem_13__1_) );
  SDFFQX1 mem_reg_12__1_ ( .D(N916), .SIN(mem_12__0_), .SMC(test_se), .C(
        net10513), .Q(mem_12__1_) );
  SDFFQX1 mem_reg_11__1_ ( .D(N925), .SIN(mem_11__0_), .SMC(test_se), .C(
        net10508), .Q(mem_11__1_) );
  SDFFQX1 mem_reg_10__1_ ( .D(N934), .SIN(mem_10__0_), .SMC(test_se), .C(
        net10503), .Q(mem_10__1_) );
  SDFFQX1 mem_reg_9__1_ ( .D(N943), .SIN(mem_9__0_), .SMC(test_se), .C(
        net10498), .Q(mem_9__1_) );
  SDFFQX1 mem_reg_8__1_ ( .D(N952), .SIN(mem_8__0_), .SMC(test_se), .C(
        net10493), .Q(mem_8__1_) );
  SDFFQX1 mem_reg_27__0_ ( .D(N780), .SIN(mem_26__7_), .SMC(test_se), .C(
        net10588), .Q(mem_27__0_) );
  SDFFQX1 mem_reg_26__0_ ( .D(N789), .SIN(mem_25__7_), .SMC(test_se), .C(
        net10583), .Q(mem_26__0_) );
  SDFFQX1 mem_reg_25__0_ ( .D(N798), .SIN(mem_24__7_), .SMC(test_se), .C(
        net10578), .Q(mem_25__0_) );
  SDFFQX1 mem_reg_24__0_ ( .D(N807), .SIN(mem_23__7_), .SMC(test_se), .C(
        net10573), .Q(mem_24__0_) );
  SDFFQX1 mem_reg_23__0_ ( .D(N816), .SIN(mem_22__7_), .SMC(test_se), .C(
        net10568), .Q(mem_23__0_) );
  SDFFQX1 mem_reg_22__0_ ( .D(N825), .SIN(mem_21__7_), .SMC(test_se), .C(
        net10563), .Q(mem_22__0_) );
  SDFFQX1 mem_reg_21__0_ ( .D(N834), .SIN(mem_20__7_), .SMC(test_se), .C(
        net10558), .Q(mem_21__0_) );
  SDFFQX1 mem_reg_20__0_ ( .D(N843), .SIN(mem_19__7_), .SMC(test_se), .C(
        net10553), .Q(mem_20__0_) );
  SDFFQX1 mem_reg_19__0_ ( .D(N852), .SIN(mem_18__7_), .SMC(test_se), .C(
        net10548), .Q(mem_19__0_) );
  SDFFQX1 mem_reg_18__0_ ( .D(N861), .SIN(mem_17__7_), .SMC(test_se), .C(
        net10543), .Q(mem_18__0_) );
  SDFFQX1 mem_reg_17__0_ ( .D(N870), .SIN(mem_16__7_), .SMC(test_se), .C(
        net10538), .Q(mem_17__0_) );
  SDFFQX1 mem_reg_16__0_ ( .D(N879), .SIN(mem_15__7_), .SMC(test_se), .C(
        net10533), .Q(mem_16__0_) );
  SDFFQX1 mem_reg_15__0_ ( .D(N888), .SIN(mem_14__7_), .SMC(test_se), .C(
        net10528), .Q(mem_15__0_) );
  SDFFQX1 mem_reg_14__0_ ( .D(N897), .SIN(mem_13__7_), .SMC(test_se), .C(
        net10523), .Q(mem_14__0_) );
  SDFFQX1 mem_reg_13__0_ ( .D(N906), .SIN(mem_12__7_), .SMC(test_se), .C(
        net10518), .Q(mem_13__0_) );
  SDFFQX1 mem_reg_12__0_ ( .D(N915), .SIN(mem_11__7_), .SMC(test_se), .C(
        net10513), .Q(mem_12__0_) );
  SDFFQX1 mem_reg_11__0_ ( .D(N924), .SIN(mem_10__7_), .SMC(test_se), .C(
        net10508), .Q(mem_11__0_) );
  SDFFQX1 mem_reg_10__0_ ( .D(N933), .SIN(mem_9__7_), .SMC(test_se), .C(
        net10503), .Q(mem_10__0_) );
  SDFFQX1 mem_reg_9__0_ ( .D(N942), .SIN(mem_8__7_), .SMC(test_se), .C(
        net10498), .Q(mem_9__0_) );
  SDFFQX1 mem_reg_8__0_ ( .D(N951), .SIN(dat_7_1[55]), .SMC(test_se), .C(
        net10493), .Q(mem_8__0_) );
  SDFFQX1 mem_reg_1__0_ ( .D(N1014), .SIN(rdat0[7]), .SMC(test_se), .C(
        net10458), .Q(dat_7_1[0]) );
  SDFFQX1 mem_reg_1__3_ ( .D(N1017), .SIN(dat_7_1[2]), .SMC(test_se), .C(
        net10458), .Q(dat_7_1[3]) );
  SDFFQX1 mem_reg_1__2_ ( .D(N1016), .SIN(dat_7_1[1]), .SMC(test_se), .C(
        net10458), .Q(dat_7_1[2]) );
  SDFFQX1 mem_reg_1__1_ ( .D(N1015), .SIN(dat_7_1[0]), .SMC(test_se), .C(
        net10458), .Q(dat_7_1[1]) );
  SDFFQX1 locked_reg ( .D(ps_locked), .SIN(test_si), .SMC(test_se), .C(clk), 
        .Q(locked) );
  SDFFQX1 mem_reg_6__7_ ( .D(N976), .SIN(dat_7_1[46]), .SMC(test_se), .C(
        net10483), .Q(dat_7_1[47]) );
  SDFFQX1 mem_reg_7__6_ ( .D(N966), .SIN(dat_7_1[53]), .SMC(test_se), .C(
        net10488), .Q(dat_7_1[54]) );
  SDFFQX1 mem_reg_6__4_ ( .D(N973), .SIN(dat_7_1[43]), .SMC(test_se), .C(
        net10483), .Q(dat_7_1[44]) );
  SDFFQX1 mem_reg_6__2_ ( .D(N971), .SIN(dat_7_1[41]), .SMC(test_se), .C(
        net10483), .Q(dat_7_1[42]) );
  SDFFQX1 mem_reg_7__1_ ( .D(N961), .SIN(dat_7_1[48]), .SMC(test_se), .C(
        net10488), .Q(dat_7_1[49]) );
  SDFFQX1 mem_reg_6__1_ ( .D(N970), .SIN(dat_7_1[40]), .SMC(test_se), .C(
        net10483), .Q(dat_7_1[41]) );
  SDFFQX1 mem_reg_7__0_ ( .D(N960), .SIN(dat_7_1[47]), .SMC(test_se), .C(
        net10488), .Q(dat_7_1[48]) );
  SDFFQX1 mem_reg_4__4_ ( .D(N991), .SIN(dat_7_1[27]), .SMC(test_se), .C(
        net10473), .Q(dat_7_1[28]) );
  SDFFQX1 mem_reg_4__3_ ( .D(N990), .SIN(dat_7_1[26]), .SMC(test_se), .C(
        net10473), .Q(dat_7_1[27]) );
  SDFFQX1 mem_reg_2__6_ ( .D(N1011), .SIN(dat_7_1[13]), .SMC(test_se), .C(
        net10463), .Q(dat_7_1[14]) );
  SDFFQX1 mem_reg_7__7_ ( .D(N967), .SIN(dat_7_1[54]), .SMC(test_se), .C(
        net10488), .Q(dat_7_1[55]) );
  SDFFQX1 mem_reg_6__6_ ( .D(N975), .SIN(dat_7_1[45]), .SMC(test_se), .C(
        net10483), .Q(dat_7_1[46]) );
  SDFFQX1 mem_reg_7__5_ ( .D(N965), .SIN(dat_7_1[52]), .SMC(test_se), .C(
        net10488), .Q(dat_7_1[53]) );
  SDFFQX1 mem_reg_6__5_ ( .D(N974), .SIN(dat_7_1[44]), .SMC(test_se), .C(
        net10483), .Q(dat_7_1[45]) );
  SDFFQX1 mem_reg_7__4_ ( .D(N964), .SIN(dat_7_1[51]), .SMC(test_se), .C(
        net10488), .Q(dat_7_1[52]) );
  SDFFQX1 mem_reg_7__3_ ( .D(N963), .SIN(dat_7_1[50]), .SMC(test_se), .C(
        net10488), .Q(dat_7_1[51]) );
  SDFFQX1 mem_reg_6__3_ ( .D(N972), .SIN(dat_7_1[42]), .SMC(test_se), .C(
        net10483), .Q(dat_7_1[43]) );
  SDFFQX1 mem_reg_7__2_ ( .D(N962), .SIN(dat_7_1[49]), .SMC(test_se), .C(
        net10488), .Q(dat_7_1[50]) );
  SDFFQX1 mem_reg_6__0_ ( .D(N969), .SIN(dat_7_1[39]), .SMC(test_se), .C(
        net10483), .Q(dat_7_1[40]) );
  SDFFQX1 mem_reg_5__7_ ( .D(N985), .SIN(dat_7_1[38]), .SMC(test_se), .C(
        net10478), .Q(dat_7_1[39]) );
  SDFFQX1 mem_reg_4__7_ ( .D(N994), .SIN(dat_7_1[30]), .SMC(test_se), .C(
        net10473), .Q(dat_7_1[31]) );
  SDFFQX1 mem_reg_4__6_ ( .D(N993), .SIN(dat_7_1[29]), .SMC(test_se), .C(
        net10473), .Q(dat_7_1[30]) );
  SDFFQX1 mem_reg_5__5_ ( .D(N983), .SIN(dat_7_1[36]), .SMC(test_se), .C(
        net10478), .Q(dat_7_1[37]) );
  SDFFQX1 mem_reg_4__5_ ( .D(N992), .SIN(dat_7_1[28]), .SMC(test_se), .C(
        net10473), .Q(dat_7_1[29]) );
  SDFFQX1 mem_reg_5__4_ ( .D(N982), .SIN(dat_7_1[35]), .SMC(test_se), .C(
        net10478), .Q(dat_7_1[36]) );
  SDFFQX1 mem_reg_5__3_ ( .D(N981), .SIN(dat_7_1[34]), .SMC(test_se), .C(
        net10478), .Q(dat_7_1[35]) );
  SDFFQX1 mem_reg_5__2_ ( .D(N980), .SIN(dat_7_1[33]), .SMC(test_se), .C(
        net10478), .Q(dat_7_1[34]) );
  SDFFQX1 mem_reg_4__2_ ( .D(N989), .SIN(dat_7_1[25]), .SMC(test_se), .C(
        net10473), .Q(dat_7_1[26]) );
  SDFFQX1 mem_reg_5__1_ ( .D(N979), .SIN(dat_7_1[32]), .SMC(test_se), .C(
        net10478), .Q(dat_7_1[33]) );
  SDFFQX1 mem_reg_4__1_ ( .D(N988), .SIN(dat_7_1[24]), .SMC(test_se), .C(
        net10473), .Q(dat_7_1[25]) );
  SDFFQX1 mem_reg_5__0_ ( .D(N978), .SIN(dat_7_1[31]), .SMC(test_se), .C(
        net10478), .Q(dat_7_1[32]) );
  SDFFQX1 mem_reg_4__0_ ( .D(N987), .SIN(dat_7_1[23]), .SMC(test_se), .C(
        net10473), .Q(dat_7_1[24]) );
  SDFFQX1 mem_reg_3__3_ ( .D(N999), .SIN(dat_7_1[18]), .SMC(test_se), .C(
        net10468), .Q(dat_7_1[19]) );
  SDFFQX1 mem_reg_3__2_ ( .D(N998), .SIN(dat_7_1[17]), .SMC(test_se), .C(
        net10468), .Q(dat_7_1[18]) );
  SDFFQX1 mem_reg_3__1_ ( .D(N997), .SIN(dat_7_1[16]), .SMC(test_se), .C(
        net10468), .Q(dat_7_1[17]) );
  SDFFQX1 mem_reg_3__0_ ( .D(N996), .SIN(dat_7_1[15]), .SMC(test_se), .C(
        net10468), .Q(dat_7_1[16]) );
  SDFFQX1 mem_reg_2__7_ ( .D(N1012), .SIN(dat_7_1[14]), .SMC(test_se), .C(
        net10463), .Q(dat_7_1[15]) );
  SDFFQX1 mem_reg_2__5_ ( .D(N1010), .SIN(dat_7_1[12]), .SMC(test_se), .C(
        net10463), .Q(dat_7_1[13]) );
  SDFFQX1 mem_reg_5__6_ ( .D(N984), .SIN(dat_7_1[37]), .SMC(test_se), .C(
        net10478), .Q(dat_7_1[38]) );
  SDFFQX1 mem_reg_1__7_ ( .D(N1021), .SIN(dat_7_1[6]), .SMC(test_se), .C(
        net10458), .Q(dat_7_1[7]) );
  SDFFQX1 mem_reg_1__6_ ( .D(N1020), .SIN(dat_7_1[5]), .SMC(test_se), .C(
        net10458), .Q(dat_7_1[6]) );
  SDFFQX1 mem_reg_1__5_ ( .D(N1019), .SIN(dat_7_1[4]), .SMC(test_se), .C(
        net10458), .Q(dat_7_1[5]) );
  SDFFQX1 mem_reg_1__4_ ( .D(N1018), .SIN(dat_7_1[3]), .SMC(test_se), .C(
        net10458), .Q(dat_7_1[4]) );
  SDFFQX1 mem_reg_3__6_ ( .D(N1002), .SIN(dat_7_1[21]), .SMC(test_se), .C(
        net10468), .Q(dat_7_1[22]) );
  SDFFQX1 mem_reg_3__5_ ( .D(N1001), .SIN(dat_7_1[20]), .SMC(test_se), .C(
        net10468), .Q(dat_7_1[21]) );
  SDFFQX1 mem_reg_3__4_ ( .D(N1000), .SIN(dat_7_1[19]), .SMC(test_se), .C(
        net10468), .Q(dat_7_1[20]) );
  SDFFQX1 mem_reg_2__4_ ( .D(N1009), .SIN(dat_7_1[11]), .SMC(test_se), .C(
        net10463), .Q(dat_7_1[12]) );
  SDFFQX1 mem_reg_2__3_ ( .D(N1008), .SIN(dat_7_1[10]), .SMC(test_se), .C(
        net10463), .Q(dat_7_1[11]) );
  SDFFQX1 mem_reg_2__2_ ( .D(N1007), .SIN(dat_7_1[9]), .SMC(test_se), .C(
        net10463), .Q(dat_7_1[10]) );
  SDFFQX1 mem_reg_3__7_ ( .D(N1003), .SIN(dat_7_1[22]), .SMC(test_se), .C(
        net10468), .Q(dat_7_1[23]) );
  SDFFQX1 mem_reg_2__1_ ( .D(N1006), .SIN(dat_7_1[8]), .SMC(test_se), .C(
        net10463), .Q(dat_7_1[9]) );
  SDFFQX1 mem_reg_2__0_ ( .D(N1005), .SIN(dat_7_1[7]), .SMC(test_se), .C(
        net10463), .Q(dat_7_1[8]) );
  SDFFQX1 mem_reg_0__1_ ( .D(N1024), .SIN(rdat0[0]), .SMC(test_se), .C(
        net10452), .Q(rdat0[1]) );
  SDFFQX1 mem_reg_0__5_ ( .D(N1028), .SIN(rdat0[4]), .SMC(test_se), .C(
        net10452), .Q(rdat0[5]) );
  SDFFQX1 mem_reg_0__2_ ( .D(N1025), .SIN(rdat0[1]), .SMC(test_se), .C(
        net10452), .Q(rdat0[2]) );
  SDFFQX1 mem_reg_0__4_ ( .D(N1027), .SIN(rdat0[3]), .SMC(test_se), .C(
        net10452), .Q(rdat0[4]) );
  SDFFQX1 mem_reg_0__6_ ( .D(N1029), .SIN(rdat0[5]), .SMC(test_se), .C(
        net10452), .Q(rdat0[6]) );
  SDFFQX1 mem_reg_0__7_ ( .D(N1030), .SIN(rdat0[6]), .SMC(test_se), .C(
        net10452), .Q(rdat0[7]) );
  SDFFQX1 pshptr_reg_3_ ( .D(N1057), .SIN(ptr[2]), .SMC(test_se), .C(net10623), 
        .Q(ptr[3]) );
  SDFFQX1 pshptr_reg_2_ ( .D(N1056), .SIN(ptr[1]), .SMC(test_se), .C(net10623), 
        .Q(ptr[2]) );
  SDFFQX1 pshptr_reg_4_ ( .D(N1058), .SIN(ptr[3]), .SMC(test_se), .C(net10623), 
        .Q(ptr[4]) );
  SDFFQX1 mem_reg_0__3_ ( .D(N1026), .SIN(rdat0[2]), .SMC(test_se), .C(
        net10452), .Q(rdat0[3]) );
  SDFFQX1 mem_reg_0__0_ ( .D(N1023), .SIN(locked), .SMC(test_se), .C(net10452), 
        .Q(rdat0[0]) );
  SDFFQX1 pshptr_reg_1_ ( .D(N1055), .SIN(ptr[0]), .SMC(test_se), .C(net10623), 
        .Q(ptr[1]) );
  SDFFQX1 pshptr_reg_5_ ( .D(N1059), .SIN(ptr[4]), .SMC(test_se), .C(net10623), 
        .Q(ptr[5]) );
  SDFFQX1 pshptr_reg_0_ ( .D(N1054), .SIN(mem_33__7_), .SMC(test_se), .C(
        net10623), .Q(ptr[0]) );
  BUFX3 U3 ( .A(n68), .Y(n1) );
  BUFX3 U4 ( .A(n222), .Y(n2) );
  BUFX3 U5 ( .A(n128), .Y(n3) );
  INVX1 U6 ( .A(n521), .Y(n4) );
  BUFX3 U7 ( .A(n313), .Y(n5) );
  INVX1 U8 ( .A(ptr[4]), .Y(n502) );
  INVXL U9 ( .A(n503), .Y(n501) );
  INVXL U10 ( .A(n505), .Y(one) );
  NAND32XL U11 ( .B(ptr[0]), .C(n503), .A(n502), .Y(n500) );
  INVXL U12 ( .A(ptr[5]), .Y(n438) );
  NAND32XL U13 ( .B(ptr[3]), .C(ptr[2]), .A(n435), .Y(n437) );
  AND2XL U14 ( .A(n441), .B(n502), .Y(n435) );
  NAND21XL U15 ( .B(n498), .A(ptr[5]), .Y(n524) );
  NAND21XL U16 ( .B(n498), .A(ptr[3]), .Y(n527) );
  NAND21XL U17 ( .B(n498), .A(ptr[4]), .Y(n518) );
  OR4X1 U18 ( .A(ptx_pop), .B(n498), .C(prx_psh), .D(n6), .Y(n506) );
  AOI21X1 U19 ( .B(i_lockena), .C(n50), .A(locked), .Y(n6) );
  NAND21XL U20 ( .B(n498), .A(ptr[2]), .Y(n531) );
  NAND21XL U21 ( .B(n498), .A(ptr[0]), .Y(n514) );
  NAND21XL U22 ( .B(n498), .A(ptr[1]), .Y(n510) );
  AND2XL U23 ( .A(one), .B(r_pop), .Y(n507) );
  INVX1 U24 ( .A(n430), .Y(n428) );
  INVX1 U25 ( .A(n21), .Y(n20) );
  INVX1 U26 ( .A(n21), .Y(n19) );
  INVX1 U27 ( .A(n430), .Y(n429) );
  INVX1 U28 ( .A(n430), .Y(n427) );
  INVX1 U29 ( .A(n21), .Y(n18) );
  INVX1 U30 ( .A(n83), .Y(n21) );
  INVX1 U31 ( .A(n29), .Y(n28) );
  INVX1 U32 ( .A(n29), .Y(n27) );
  INVX1 U33 ( .A(n37), .Y(n36) );
  INVX1 U34 ( .A(n37), .Y(n35) );
  INVX1 U35 ( .A(n45), .Y(n44) );
  INVX1 U36 ( .A(n45), .Y(n43) );
  INVX1 U37 ( .A(n54), .Y(n430) );
  INVX1 U38 ( .A(n444), .Y(n498) );
  NOR21XL U39 ( .B(n70), .A(n66), .Y(n74) );
  NOR21XL U40 ( .B(n361), .A(n105), .Y(n363) );
  NOR21XL U41 ( .B(n106), .A(n66), .Y(n108) );
  NOR21XL U42 ( .B(n385), .A(n105), .Y(n387) );
  NAND21X1 U43 ( .B(n442), .A(n550), .Y(n490) );
  INVX1 U44 ( .A(n245), .Y(n211) );
  INVX1 U45 ( .A(n348), .Y(n291) );
  INVX1 U46 ( .A(n422), .Y(n420) );
  INVX1 U47 ( .A(n245), .Y(n223) );
  INVX1 U48 ( .A(n348), .Y(n335) );
  INVX1 U49 ( .A(n422), .Y(n421) );
  NAND2X1 U50 ( .A(fifowdat[3]), .B(n141), .Y(n54) );
  NAND2X1 U51 ( .A(fifowdat[4]), .B(n141), .Y(n83) );
  INVX1 U52 ( .A(r_psh), .Y(n552) );
  INVX1 U53 ( .A(n29), .Y(n26) );
  INVX1 U54 ( .A(n80), .Y(n29) );
  INVX1 U55 ( .A(n37), .Y(n34) );
  INVX1 U56 ( .A(n77), .Y(n37) );
  INVX1 U57 ( .A(n45), .Y(n42) );
  INVX1 U58 ( .A(n73), .Y(n45) );
  NAND2X1 U59 ( .A(n442), .B(n444), .Y(N1053) );
  INVX1 U60 ( .A(fifowdat[3]), .Y(n431) );
  INVX1 U61 ( .A(fifowdat[3]), .Y(n432) );
  INVX1 U62 ( .A(fifowdat[4]), .Y(n22) );
  INVX1 U63 ( .A(fifowdat[4]), .Y(n23) );
  INVX1 U64 ( .A(fifowdat[3]), .Y(n433) );
  INVX1 U65 ( .A(fifowdat[4]), .Y(n24) );
  NOR21XL U66 ( .B(srstz), .A(r_fiforst), .Y(n444) );
  NOR21XL U67 ( .B(n407), .A(n141), .Y(n409) );
  NOR21XL U68 ( .B(n458), .A(n105), .Y(n460) );
  NOR21XL U69 ( .B(n52), .A(n141), .Y(n56) );
  NOR21XL U70 ( .B(n93), .A(n66), .Y(n95) );
  NOR21XL U71 ( .B(n118), .A(n66), .Y(n120) );
  NOR21XL U72 ( .B(n448), .A(n105), .Y(n450) );
  NOR21XL U73 ( .B(n130), .A(n66), .Y(n132) );
  NOR21XL U74 ( .B(n143), .A(n66), .Y(n145) );
  NOR21XL U75 ( .B(n155), .A(n66), .Y(n157) );
  NOR21XL U76 ( .B(n166), .A(n66), .Y(n168) );
  NOR21XL U77 ( .B(n177), .A(n66), .Y(n179) );
  NOR21XL U78 ( .B(n189), .A(n66), .Y(n191) );
  NOR21XL U79 ( .B(n212), .A(n92), .Y(n214) );
  NOR21XL U80 ( .B(n224), .A(n92), .Y(n226) );
  NOR21XL U81 ( .B(n235), .A(n92), .Y(n237) );
  NOR21XL U82 ( .B(n247), .A(n92), .Y(n249) );
  NOR21XL U83 ( .B(n258), .A(n92), .Y(n260) );
  NOR21XL U84 ( .B(n269), .A(n92), .Y(n271) );
  NOR21XL U85 ( .B(n281), .A(n92), .Y(n283) );
  NOR21XL U86 ( .B(n303), .A(n92), .Y(n305) );
  NOR21XL U87 ( .B(n314), .A(n92), .Y(n316) );
  NOR21XL U88 ( .B(n325), .A(n105), .Y(n327) );
  NOR21XL U89 ( .B(n337), .A(n105), .Y(n339) );
  NOR21XL U90 ( .B(n350), .A(n105), .Y(n352) );
  NOR21XL U91 ( .B(n373), .A(n105), .Y(n375) );
  NOR21XL U92 ( .B(n200), .A(n92), .Y(n202) );
  NOR21XL U93 ( .B(n292), .A(n105), .Y(n294) );
  AOI21BBXL U94 ( .B(n88), .C(n313), .A(n371), .Y(n361) );
  AOI21BBXL U95 ( .B(n68), .C(n88), .A(n89), .Y(n70) );
  NAND21X1 U96 ( .B(n442), .A(n443), .Y(n491) );
  XNOR2XL U97 ( .A(n7), .B(n550), .Y(n442) );
  AND2X1 U98 ( .A(n395), .B(n313), .Y(n385) );
  AND2X1 U99 ( .A(n116), .B(n68), .Y(n106) );
  INVX1 U100 ( .A(n176), .Y(n141) );
  INVX1 U101 ( .A(n104), .Y(n545) );
  INVX1 U102 ( .A(n534), .Y(n537) );
  INVX1 U103 ( .A(n348), .Y(n280) );
  INVX1 U104 ( .A(n422), .Y(n419) );
  INVX1 U105 ( .A(n245), .Y(n199) );
  INVX1 U106 ( .A(n64), .Y(n245) );
  INVX1 U107 ( .A(n443), .Y(n550) );
  INVX1 U108 ( .A(n494), .Y(n475) );
  INVX1 U109 ( .A(n495), .Y(n476) );
  INVX1 U110 ( .A(n61), .Y(n348) );
  INVX1 U111 ( .A(n58), .Y(n422) );
  NAND2X1 U112 ( .A(fifowdat[5]), .B(n141), .Y(n80) );
  NAND2X1 U113 ( .A(fifowdat[6]), .B(n141), .Y(n77) );
  NAND2X1 U114 ( .A(fifowdat[7]), .B(n141), .Y(n73) );
  NAND2X1 U115 ( .A(n552), .B(n554), .Y(n50) );
  INVX1 U116 ( .A(n187), .Y(n66) );
  INVX1 U117 ( .A(n187), .Y(n92) );
  INVX1 U118 ( .A(n176), .Y(n105) );
  AOI21X1 U119 ( .B(n549), .C(n548), .A(n336), .Y(n347) );
  INVX1 U120 ( .A(n520), .Y(n541) );
  INVX1 U121 ( .A(n522), .Y(n538) );
  INVX1 U122 ( .A(n519), .Y(n539) );
  NOR2X1 U123 ( .A(n104), .B(n546), .Y(n91) );
  INVX1 U124 ( .A(n176), .Y(n142) );
  INVX1 U125 ( .A(n187), .Y(n154) );
  INVX1 U126 ( .A(n187), .Y(n165) );
  INVX1 U127 ( .A(n511), .Y(n543) );
  OAI22X1 U128 ( .A(n1), .B(n88), .C(n91), .D(n165), .Y(N977) );
  INVX1 U129 ( .A(fifowdat[6]), .Y(n38) );
  INVX1 U130 ( .A(fifowdat[6]), .Y(n39) );
  INVX1 U131 ( .A(fifowdat[6]), .Y(n40) );
  INVX1 U132 ( .A(n53), .Y(fifowdat[3]) );
  INVX1 U133 ( .A(n81), .Y(fifowdat[4]) );
  INVX1 U134 ( .A(fifowdat[5]), .Y(n30) );
  INVX1 U135 ( .A(fifowdat[5]), .Y(n31) );
  INVX1 U136 ( .A(fifowdat[7]), .Y(n46) );
  INVX1 U137 ( .A(fifowdat[7]), .Y(n47) );
  INVX1 U138 ( .A(fifowdat[5]), .Y(n32) );
  INVX1 U139 ( .A(fifowdat[7]), .Y(n49) );
  NOR21XL U140 ( .B(n17), .A(n105), .Y(n398) );
  NOR21XL U141 ( .B(n417), .A(n418), .Y(n407) );
  NAND21X1 U142 ( .B(n526), .A(n548), .Y(n313) );
  AOI21BBXL U143 ( .B(n128), .C(n129), .A(n545), .Y(n118) );
  AOI21BBXL U144 ( .B(n129), .C(n313), .A(n541), .Y(n303) );
  AOI21BBXL U145 ( .B(n140), .C(n313), .A(n324), .Y(n314) );
  AOI21BBXL U146 ( .B(n153), .C(n313), .A(n16), .Y(n325) );
  AOI21BBXL U147 ( .B(n69), .C(n313), .A(n347), .Y(n337) );
  AOI21BBXL U148 ( .B(n90), .C(n313), .A(n360), .Y(n350) );
  AOI21BBXL U149 ( .B(n103), .C(n313), .A(n372), .Y(n373) );
  AOI21BBXL U150 ( .B(n69), .C(n128), .A(n9), .Y(n155) );
  AOI21BBXL U151 ( .B(n90), .C(n128), .A(n551), .Y(n166) );
  AOI21BBXL U152 ( .B(n88), .C(n128), .A(n10), .Y(n177) );
  AOI21BBXL U153 ( .B(n103), .C(n128), .A(n188), .Y(n189) );
  AOI21BBXL U154 ( .B(n129), .C(n222), .A(n547), .Y(n212) );
  AOI21BBXL U155 ( .B(n140), .C(n222), .A(n234), .Y(n224) );
  AOI21BBXL U156 ( .B(n153), .C(n222), .A(n14), .Y(n235) );
  AOI21BBXL U157 ( .B(n69), .C(n222), .A(n11), .Y(n247) );
  AOI21BBXL U158 ( .B(n90), .C(n222), .A(n538), .Y(n258) );
  AOI21BBXL U159 ( .B(n88), .C(n222), .A(n15), .Y(n269) );
  AOI21BBXL U160 ( .B(n103), .C(n222), .A(n539), .Y(n281) );
  AOI21BBXL U161 ( .B(n90), .C(n68), .A(n544), .Y(n52) );
  AOI21BBXL U162 ( .B(n68), .C(n69), .A(n468), .Y(n458) );
  AOI21BBXL U163 ( .B(n68), .C(n103), .A(n91), .Y(n93) );
  AOI21BBXL U164 ( .B(n128), .C(n153), .A(n537), .Y(n143) );
  AOI21BBXL U165 ( .B(n68), .C(n153), .A(n543), .Y(n448) );
  AOI21BBXL U166 ( .B(n128), .C(n140), .A(n8), .Y(n130) );
  NAND21X1 U167 ( .B(n526), .A(n545), .Y(n68) );
  AO21X1 U168 ( .B(n547), .C(n530), .A(n545), .Y(n188) );
  OR2X1 U169 ( .A(n477), .B(n491), .Y(n494) );
  NAND21X1 U170 ( .B(n536), .A(n547), .Y(n104) );
  AO21X1 U171 ( .B(n536), .C(n533), .A(n532), .Y(n534) );
  OR2X1 U172 ( .A(n440), .B(n490), .Y(n495) );
  OAI21AX1 U173 ( .B(n542), .C(n554), .A(ptx_pop), .Y(n443) );
  AOI21BBXL U174 ( .B(n542), .C(n552), .A(prx_psh), .Y(n7) );
  INVX1 U175 ( .A(n7), .Y(fifopsh) );
  AND2X1 U176 ( .A(n210), .B(n128), .Y(n200) );
  AND2X1 U177 ( .A(n302), .B(n222), .Y(n292) );
  NAND21X1 U178 ( .B(n526), .A(n516), .Y(n417) );
  INVX1 U179 ( .A(n528), .Y(n547) );
  MUX2X1 U180 ( .D0(n481), .D1(n480), .S(n523), .Y(N1058) );
  OAI22X1 U181 ( .A(n492), .B(n491), .C(n479), .D(n490), .Y(n480) );
  AO21X1 U182 ( .B(n476), .C(n536), .A(n475), .Y(n481) );
  AND2X1 U183 ( .A(n478), .B(n536), .Y(n479) );
  AOI21X1 U184 ( .B(n536), .C(n535), .A(n534), .Y(n8) );
  AOI21X1 U185 ( .B(n536), .C(n549), .A(n532), .Y(n9) );
  AOI21AX1 U186 ( .B(n540), .C(n536), .A(n188), .Y(n10) );
  INVX1 U187 ( .A(n551), .Y(n532) );
  INVX1 U188 ( .A(n67), .Y(n176) );
  NAND2X1 U189 ( .A(fifowdat[0]), .B(n141), .Y(n64) );
  NAND2X1 U190 ( .A(fifowdat[1]), .B(n141), .Y(n61) );
  NAND2X1 U191 ( .A(fifowdat[2]), .B(n141), .Y(n58) );
  INVX1 U192 ( .A(r_pop), .Y(n554) );
  NOR21XL U193 ( .B(n91), .A(n540), .Y(n89) );
  NAND21X1 U194 ( .B(n516), .A(n513), .Y(n520) );
  AO21X1 U195 ( .B(n523), .C(n521), .A(n520), .Y(n522) );
  AO21X1 U196 ( .B(n523), .C(n546), .A(n520), .Y(n519) );
  AOI21X1 U197 ( .B(n523), .C(n549), .A(n522), .Y(n11) );
  NAND21X1 U198 ( .B(n533), .A(n544), .Y(n511) );
  NAND21X1 U199 ( .B(n533), .A(n540), .Y(n88) );
  AO21X1 U200 ( .B(n548), .C(n529), .A(n516), .Y(n395) );
  AO21X1 U201 ( .B(n523), .C(n529), .A(n520), .Y(n302) );
  AO21X1 U202 ( .B(n536), .C(n529), .A(n528), .Y(n210) );
  AO21X1 U203 ( .B(n548), .C(n521), .A(n516), .Y(n336) );
  AOI21AX1 U204 ( .B(n540), .C(n548), .A(n372), .Y(n371) );
  INVX1 U205 ( .A(n129), .Y(n517) );
  AND2X1 U206 ( .A(n544), .B(n436), .Y(n468) );
  NOR2X1 U207 ( .A(n142), .B(n13), .Y(n12) );
  AOI21X1 U208 ( .B(n535), .C(n526), .A(n511), .Y(n13) );
  INVX1 U209 ( .A(n513), .Y(n548) );
  AOI21X1 U210 ( .B(n523), .C(n533), .A(n522), .Y(n14) );
  AOI21X1 U211 ( .B(n523), .C(n540), .A(n519), .Y(n15) );
  AOI21X1 U212 ( .B(n548), .C(n533), .A(n336), .Y(n16) );
  INVX1 U213 ( .A(n530), .Y(n546) );
  OAI32X1 U214 ( .A(n535), .B(empty), .C(n491), .D(n482), .E(n490), .Y(N1054)
         );
  XOR2X1 U215 ( .A(n535), .B(full), .Y(n482) );
  INVX1 U216 ( .A(n117), .Y(n529) );
  INVX1 U217 ( .A(n436), .Y(n549) );
  OAI22X1 U218 ( .A(n547), .B(n165), .C(n3), .D(n117), .Y(N887) );
  OAI22X1 U219 ( .A(n541), .B(n165), .C(n117), .D(n222), .Y(N815) );
  OAI22X1 U220 ( .A(n90), .B(n5), .C(n371), .D(n154), .Y(N770) );
  OAI22X1 U221 ( .A(n153), .B(n5), .C(n347), .D(n154), .Y(N788) );
  OAI22X1 U222 ( .A(n140), .B(n5), .C(n16), .D(n154), .Y(N797) );
  OAI22X1 U223 ( .A(n88), .B(n2), .C(n539), .D(n154), .Y(N833) );
  OAI22X1 U224 ( .A(n90), .B(n2), .C(n15), .D(n154), .Y(N842) );
  OAI22X1 U225 ( .A(n69), .B(n2), .C(n538), .D(n154), .Y(N851) );
  OAI22X1 U226 ( .A(n153), .B(n2), .C(n11), .D(n165), .Y(N860) );
  OAI22X1 U227 ( .A(n140), .B(n2), .C(n14), .D(n154), .Y(N869) );
  OAI22X1 U228 ( .A(n90), .B(n128), .C(n10), .D(n154), .Y(N914) );
  OAI22X1 U229 ( .A(n3), .B(n153), .C(n9), .D(n154), .Y(N932) );
  OAI22X1 U230 ( .A(n3), .B(n140), .C(n537), .D(n165), .Y(N941) );
  OAI22X1 U231 ( .A(n3), .B(n129), .C(n8), .D(n165), .Y(N950) );
  OAI22X1 U232 ( .A(n90), .B(n68), .C(n89), .D(n165), .Y(N986) );
  OAI22X1 U233 ( .A(n1), .B(n129), .C(n447), .D(n154), .Y(N1022) );
  AND2X1 U234 ( .A(n545), .B(n517), .Y(n447) );
  OAI22X1 U235 ( .A(n88), .B(n3), .C(n142), .D(n188), .Y(N905) );
  OAI22X1 U236 ( .A(n69), .B(n3), .C(n142), .D(n551), .Y(N923) );
  OAI22X1 U237 ( .A(n69), .B(n5), .C(n142), .D(n360), .Y(N779) );
  OAI22X1 U238 ( .A(n129), .B(n5), .C(n142), .D(n324), .Y(N806) );
  OAI22X1 U239 ( .A(n129), .B(n2), .C(n142), .D(n234), .Y(N878) );
  INVX1 U240 ( .A(n67), .Y(n187) );
  NAND2X1 U241 ( .A(n545), .B(n117), .Y(n116) );
  INVX1 U242 ( .A(n486), .Y(n445) );
  INVX1 U243 ( .A(n477), .Y(n492) );
  OAI22X1 U244 ( .A(n545), .B(n67), .C(n1), .D(n117), .Y(N959) );
  OAI22X1 U245 ( .A(n544), .B(n165), .C(n68), .D(n69), .Y(N995) );
  OAI22X1 U246 ( .A(n468), .B(n165), .C(n68), .D(n153), .Y(N1004) );
  OAI22X1 U247 ( .A(n543), .B(n165), .C(n1), .D(n140), .Y(N1013) );
  OAI22X1 U248 ( .A(n142), .B(n372), .C(n88), .D(n313), .Y(N761) );
  OAI21X1 U249 ( .B(n142), .C(n418), .A(n406), .Y(N734) );
  NAND21X1 U250 ( .B(n417), .A(n517), .Y(n406) );
  INVX1 U251 ( .A(n440), .Y(n478) );
  ENOX1 U252 ( .A(n103), .B(n5), .C(n395), .D(n187), .Y(N752) );
  ENOX1 U253 ( .A(n103), .B(n2), .C(n302), .D(n187), .Y(N824) );
  ENOX1 U254 ( .A(n103), .B(n3), .C(n210), .D(n187), .Y(N896) );
  ENOX1 U255 ( .A(n1), .B(n103), .C(n116), .D(n187), .Y(N968) );
  MUX2IX1 U256 ( .D0(r_wdat[3]), .D1(prx_wdat[3]), .S(prx_psh), .Y(n53) );
  MUX2IX1 U257 ( .D0(r_wdat[4]), .D1(prx_wdat[4]), .S(prx_psh), .Y(n81) );
  INVX1 U258 ( .A(n75), .Y(fifowdat[6]) );
  INVX1 U259 ( .A(n71), .Y(fifowdat[7]) );
  INVX1 U260 ( .A(fifowdat[0]), .Y(n246) );
  INVX1 U261 ( .A(fifowdat[0]), .Y(n257) );
  INVX1 U262 ( .A(fifowdat[1]), .Y(n349) );
  INVX1 U263 ( .A(fifowdat[1]), .Y(n383) );
  INVX1 U264 ( .A(fifowdat[2]), .Y(n423) );
  INVX1 U265 ( .A(fifowdat[2]), .Y(n424) );
  INVX1 U266 ( .A(fifowdat[0]), .Y(n268) );
  INVX1 U267 ( .A(fifowdat[1]), .Y(n384) );
  INVX1 U268 ( .A(fifowdat[2]), .Y(n425) );
  INVX1 U269 ( .A(n78), .Y(fifowdat[5]) );
  AND3X1 U270 ( .A(ptr[0]), .B(ptr[4]), .C(n501), .Y(half) );
  NOR3XL U271 ( .A(n555), .B(n542), .C(n48), .Y(txreq) );
  INVX1 U272 ( .A(n496), .Y(full) );
  INVX1 U273 ( .A(n500), .Y(empty) );
  INVX1 U274 ( .A(n509), .Y(n542) );
  NAND32X1 U275 ( .B(n527), .C(n526), .A(n547), .Y(n128) );
  NAND32X1 U276 ( .B(n526), .C(n518), .A(n527), .Y(n222) );
  NAND21X1 U277 ( .B(n7), .A(n496), .Y(n526) );
  AO21X1 U278 ( .B(n547), .C(n531), .A(n545), .Y(n551) );
  NAND21X1 U279 ( .B(n523), .A(n524), .Y(n528) );
  OAI221X1 U280 ( .A(n513), .B(n495), .C(n528), .D(n494), .E(n493), .Y(N1059)
         );
  GEN2XL U281 ( .D(n492), .E(n518), .C(n491), .B(n490), .A(n524), .Y(n493) );
  NAND21X1 U282 ( .B(n550), .A(n500), .Y(n67) );
  INVX1 U283 ( .A(n527), .Y(n536) );
  NAND21X1 U284 ( .B(n474), .A(n494), .Y(N1057) );
  MUX2X1 U285 ( .D0(n476), .D1(n473), .S(n536), .Y(n474) );
  OAI22X1 U286 ( .A(n478), .B(n490), .C(n446), .D(n491), .Y(n473) );
  AND2X1 U287 ( .A(n445), .B(n531), .Y(n446) );
  INVX1 U288 ( .A(n518), .Y(n523) );
  AOI21BX1 U289 ( .C(n526), .B(n517), .A(n524), .Y(n17) );
  NAND32X1 U290 ( .B(n521), .C(n533), .A(n514), .Y(n129) );
  NAND21X1 U291 ( .B(n514), .A(n546), .Y(n117) );
  NAND21X1 U292 ( .B(n514), .A(n533), .Y(n436) );
  NAND21X1 U293 ( .B(n527), .A(n523), .Y(n513) );
  NAND21X1 U294 ( .B(n4), .A(n533), .Y(n530) );
  NAND21X1 U295 ( .B(n531), .A(n487), .Y(n440) );
  NAND21X1 U296 ( .B(n530), .A(n514), .Y(n103) );
  NAND32X1 U297 ( .B(n521), .C(n510), .A(n514), .Y(n153) );
  NAND21X1 U298 ( .B(n436), .A(n531), .Y(n69) );
  INVX1 U299 ( .A(n515), .Y(n540) );
  NAND21X1 U300 ( .B(n514), .A(n521), .Y(n515) );
  NAND32X1 U301 ( .B(n521), .C(n514), .A(n510), .Y(n140) );
  AO21X1 U302 ( .B(n530), .C(n524), .A(n541), .Y(n372) );
  AO21X1 U303 ( .B(n524), .C(n517), .A(n541), .Y(n324) );
  AO21X1 U304 ( .B(n525), .C(n524), .A(n547), .Y(n234) );
  AO21X1 U305 ( .B(n524), .C(n531), .A(n541), .Y(n360) );
  AO21X1 U306 ( .B(n525), .C(n518), .A(n524), .Y(n418) );
  INVX1 U307 ( .A(n531), .Y(n521) );
  INVX1 U308 ( .A(n510), .Y(n533) );
  INVX1 U309 ( .A(n524), .Y(n516) );
  INVX1 U310 ( .A(n497), .Y(n544) );
  NAND21X1 U311 ( .B(n104), .A(n531), .Y(n497) );
  OAI32X1 U312 ( .A(n496), .B(n7), .C(n142), .D(n417), .E(n140), .Y(N733) );
  INVX1 U313 ( .A(n439), .Y(n487) );
  NAND21X1 U314 ( .B(n436), .A(n496), .Y(n439) );
  OAI22X1 U315 ( .A(n489), .B(n491), .C(n488), .D(n490), .Y(N1056) );
  XOR2X1 U316 ( .A(n486), .B(n521), .Y(n489) );
  OA22X1 U317 ( .A(n487), .B(n531), .C(n69), .D(full), .Y(n488) );
  OAI22X1 U318 ( .A(n485), .B(n491), .C(n484), .D(n490), .Y(N1055) );
  AND2X1 U319 ( .A(n486), .B(n436), .Y(n485) );
  XOR2X1 U320 ( .A(n510), .B(n483), .Y(n484) );
  AND2X1 U321 ( .A(n535), .B(n496), .Y(n483) );
  INVX1 U322 ( .A(n512), .Y(n525) );
  NAND21X1 U323 ( .B(n129), .A(n527), .Y(n512) );
  NAND32X1 U324 ( .B(n533), .C(empty), .A(n514), .Y(n486) );
  NAND32X1 U325 ( .B(n533), .C(n531), .A(n514), .Y(n90) );
  NAND32X1 U326 ( .B(n536), .C(n486), .A(n531), .Y(n477) );
  INVX1 U327 ( .A(n514), .Y(n535) );
  OAI22X1 U328 ( .A(n142), .B(n524), .C(n5), .D(n117), .Y(N743) );
  INVX1 U329 ( .A(n48), .Y(n553) );
  INVX1 U330 ( .A(n506), .Y(ps_locked) );
  MUX2IX1 U331 ( .D0(r_wdat[7]), .D1(prx_wdat[7]), .S(prx_psh), .Y(n71) );
  INVX1 U332 ( .A(n63), .Y(fifowdat[0]) );
  INVX1 U333 ( .A(n60), .Y(fifowdat[1]) );
  INVX1 U334 ( .A(n57), .Y(fifowdat[2]) );
  MUX2IXL U335 ( .D0(r_wdat[5]), .D1(prx_wdat[5]), .S(prx_psh), .Y(n78) );
  NAND43X1 U336 ( .B(ptr[2]), .C(ptr[3]), .D(ptr[5]), .A(n441), .Y(n503) );
  INVX1 U337 ( .A(ptr[1]), .Y(n441) );
  NAND32X1 U338 ( .B(n504), .C(n503), .A(n502), .Y(n505) );
  INVX1 U339 ( .A(ptr[0]), .Y(n504) );
  NAND21X1 U340 ( .B(n438), .A(n437), .Y(n496) );
  NAND21X1 U341 ( .B(r_unlock), .A(n506), .Y(n509) );
  AO2222XL U342 ( .A(r_pop), .B(empty), .C(r_psh), .D(full), .E(n555), .F(n553), .G(n542), .H(n50), .Y(ffack[1]) );
  NOR21XL U343 ( .B(n509), .A(n508), .Y(ffack[0]) );
  NOR21XL U344 ( .B(n48), .A(n507), .Y(n508) );
  OAI211X1 U345 ( .C(n448), .D(n22), .A(n18), .B(n453), .Y(N1018) );
  NAND2X1 U346 ( .A(dat_7_1[12]), .B(n450), .Y(n453) );
  OAI211X1 U347 ( .C(n448), .D(n30), .A(n26), .B(n452), .Y(N1019) );
  NAND2X1 U348 ( .A(dat_7_1[13]), .B(n450), .Y(n452) );
  OAI211X1 U349 ( .C(n448), .D(n38), .A(n34), .B(n451), .Y(N1020) );
  NAND2X1 U350 ( .A(dat_7_1[14]), .B(n450), .Y(n451) );
  OAI211X1 U351 ( .C(n93), .D(n38), .A(n96), .B(n77), .Y(N984) );
  NAND2X1 U352 ( .A(dat_7_1[46]), .B(n95), .Y(n96) );
  OAI211X1 U353 ( .C(n448), .D(n46), .A(n42), .B(n449), .Y(N1021) );
  NAND2X1 U354 ( .A(dat_7_1[15]), .B(n450), .Y(n449) );
  OAI211X1 U355 ( .C(n52), .D(n246), .A(n199), .B(n65), .Y(N996) );
  NAND2X1 U356 ( .A(dat_7_1[24]), .B(n56), .Y(n65) );
  OAI211X1 U357 ( .C(n52), .D(n349), .A(n280), .B(n62), .Y(N997) );
  NAND2X1 U358 ( .A(dat_7_1[25]), .B(n56), .Y(n62) );
  OAI211X1 U359 ( .C(n52), .D(n423), .A(n419), .B(n59), .Y(N998) );
  NAND2X1 U360 ( .A(dat_7_1[26]), .B(n56), .Y(n59) );
  OAI211X1 U361 ( .C(n52), .D(n431), .A(n427), .B(n55), .Y(N999) );
  NAND2X1 U362 ( .A(dat_7_1[27]), .B(n56), .Y(n55) );
  OAI211X1 U363 ( .C(n70), .D(n246), .A(n87), .B(n199), .Y(N987) );
  NAND2X1 U364 ( .A(dat_7_1[32]), .B(n74), .Y(n87) );
  OAI211X1 U365 ( .C(n93), .D(n246), .A(n102), .B(n199), .Y(N978) );
  NAND2X1 U366 ( .A(dat_7_1[40]), .B(n95), .Y(n102) );
  OAI211X1 U367 ( .C(n70), .D(n349), .A(n86), .B(n280), .Y(N988) );
  NAND2X1 U368 ( .A(dat_7_1[33]), .B(n74), .Y(n86) );
  OAI211X1 U369 ( .C(n93), .D(n349), .A(n101), .B(n280), .Y(N979) );
  NAND2X1 U370 ( .A(dat_7_1[41]), .B(n95), .Y(n101) );
  OAI211X1 U371 ( .C(n70), .D(n423), .A(n85), .B(n419), .Y(N989) );
  NAND2X1 U372 ( .A(dat_7_1[34]), .B(n74), .Y(n85) );
  OAI211X1 U373 ( .C(n93), .D(n423), .A(n100), .B(n419), .Y(N980) );
  NAND2X1 U374 ( .A(dat_7_1[42]), .B(n95), .Y(n100) );
  OAI211X1 U375 ( .C(n70), .D(n431), .A(n84), .B(n427), .Y(N990) );
  NAND2X1 U376 ( .A(dat_7_1[35]), .B(n74), .Y(n84) );
  OAI211X1 U377 ( .C(n93), .D(n431), .A(n99), .B(n427), .Y(N981) );
  NAND2X1 U378 ( .A(dat_7_1[43]), .B(n95), .Y(n99) );
  OAI211X1 U379 ( .C(n70), .D(n22), .A(n82), .B(n83), .Y(N991) );
  NAND2X1 U380 ( .A(dat_7_1[36]), .B(n74), .Y(n82) );
  OAI211X1 U381 ( .C(n93), .D(n22), .A(n98), .B(n83), .Y(N982) );
  NAND2X1 U382 ( .A(dat_7_1[44]), .B(n95), .Y(n98) );
  OAI211X1 U383 ( .C(n70), .D(n30), .A(n79), .B(n80), .Y(N992) );
  NAND2X1 U384 ( .A(dat_7_1[37]), .B(n74), .Y(n79) );
  OAI211X1 U385 ( .C(n93), .D(n30), .A(n97), .B(n80), .Y(N983) );
  NAND2X1 U386 ( .A(dat_7_1[45]), .B(n95), .Y(n97) );
  OAI211X1 U387 ( .C(n70), .D(n38), .A(n76), .B(n77), .Y(N993) );
  NAND2X1 U388 ( .A(dat_7_1[38]), .B(n74), .Y(n76) );
  OAI211X1 U389 ( .C(n70), .D(n46), .A(n72), .B(n73), .Y(N994) );
  NAND2X1 U390 ( .A(dat_7_1[39]), .B(n74), .Y(n72) );
  OAI211X1 U391 ( .C(n93), .D(n46), .A(n94), .B(n73), .Y(N985) );
  NAND2X1 U392 ( .A(dat_7_1[47]), .B(n95), .Y(n94) );
  OAI211X1 U393 ( .C(n106), .D(n246), .A(n115), .B(n199), .Y(N969) );
  NAND2X1 U394 ( .A(dat_7_1[48]), .B(n108), .Y(n115) );
  OAI211X1 U395 ( .C(n118), .D(n246), .A(n127), .B(n199), .Y(N960) );
  NAND2X1 U396 ( .A(mem_8__0_), .B(n120), .Y(n127) );
  OAI211X1 U397 ( .C(n106), .D(n349), .A(n114), .B(n280), .Y(N970) );
  NAND2X1 U398 ( .A(dat_7_1[49]), .B(n108), .Y(n114) );
  OAI211X1 U399 ( .C(n118), .D(n349), .A(n126), .B(n280), .Y(N961) );
  NAND2X1 U400 ( .A(mem_8__1_), .B(n120), .Y(n126) );
  OAI211X1 U401 ( .C(n106), .D(n423), .A(n113), .B(n419), .Y(N971) );
  NAND2X1 U402 ( .A(dat_7_1[50]), .B(n108), .Y(n113) );
  OAI211X1 U403 ( .C(n118), .D(n423), .A(n125), .B(n419), .Y(N962) );
  NAND2X1 U404 ( .A(mem_8__2_), .B(n120), .Y(n125) );
  OAI211X1 U405 ( .C(n106), .D(n431), .A(n112), .B(n427), .Y(N972) );
  NAND2X1 U406 ( .A(dat_7_1[51]), .B(n108), .Y(n112) );
  OAI211X1 U407 ( .C(n118), .D(n431), .A(n124), .B(n427), .Y(N963) );
  NAND2X1 U408 ( .A(mem_8__3_), .B(n120), .Y(n124) );
  OAI211X1 U409 ( .C(n106), .D(n22), .A(n111), .B(n20), .Y(N973) );
  NAND2X1 U410 ( .A(dat_7_1[52]), .B(n108), .Y(n111) );
  OAI211X1 U411 ( .C(n118), .D(n22), .A(n123), .B(n20), .Y(N964) );
  NAND2X1 U412 ( .A(mem_8__4_), .B(n120), .Y(n123) );
  OAI211X1 U413 ( .C(n106), .D(n30), .A(n110), .B(n28), .Y(N974) );
  NAND2X1 U414 ( .A(dat_7_1[53]), .B(n108), .Y(n110) );
  OAI211X1 U415 ( .C(n118), .D(n30), .A(n122), .B(n28), .Y(N965) );
  NAND2X1 U416 ( .A(mem_8__5_), .B(n120), .Y(n122) );
  OAI211X1 U417 ( .C(n106), .D(n38), .A(n109), .B(n36), .Y(N975) );
  NAND2X1 U418 ( .A(dat_7_1[54]), .B(n108), .Y(n109) );
  OAI211X1 U419 ( .C(n118), .D(n38), .A(n121), .B(n36), .Y(N966) );
  NAND2X1 U420 ( .A(mem_8__6_), .B(n120), .Y(n121) );
  OAI211X1 U421 ( .C(n106), .D(n46), .A(n107), .B(n44), .Y(N976) );
  NAND2X1 U422 ( .A(dat_7_1[55]), .B(n108), .Y(n107) );
  OAI211X1 U423 ( .C(n118), .D(n46), .A(n119), .B(n44), .Y(N967) );
  NAND2X1 U424 ( .A(mem_8__7_), .B(n120), .Y(n119) );
  OAI211X1 U425 ( .C(n448), .D(n349), .A(n280), .B(n456), .Y(N1015) );
  NAND2X1 U426 ( .A(dat_7_1[9]), .B(n450), .Y(n456) );
  OAI211X1 U427 ( .C(n448), .D(n423), .A(n419), .B(n455), .Y(N1016) );
  NAND2X1 U428 ( .A(dat_7_1[10]), .B(n450), .Y(n455) );
  OAI211X1 U429 ( .C(n448), .D(n431), .A(n427), .B(n454), .Y(N1017) );
  NAND2X1 U430 ( .A(dat_7_1[11]), .B(n450), .Y(n454) );
  OAI211X1 U431 ( .C(n448), .D(n246), .A(n199), .B(n457), .Y(N1014) );
  NAND2X1 U432 ( .A(dat_7_1[8]), .B(n450), .Y(n457) );
  OAI211X1 U433 ( .C(n130), .D(n246), .A(n139), .B(n199), .Y(N951) );
  NAND2X1 U434 ( .A(mem_9__0_), .B(n132), .Y(n139) );
  OAI211X1 U435 ( .C(n143), .D(n246), .A(n152), .B(n199), .Y(N942) );
  NAND2X1 U436 ( .A(mem_10__0_), .B(n145), .Y(n152) );
  OAI211X1 U437 ( .C(n155), .D(n246), .A(n164), .B(n199), .Y(N933) );
  NAND2X1 U438 ( .A(mem_11__0_), .B(n157), .Y(n164) );
  OAI211X1 U439 ( .C(n166), .D(n246), .A(n175), .B(n211), .Y(N924) );
  NAND2X1 U440 ( .A(mem_12__0_), .B(n168), .Y(n175) );
  OAI211X1 U441 ( .C(n177), .D(n257), .A(n186), .B(n211), .Y(N915) );
  NAND2X1 U442 ( .A(mem_13__0_), .B(n179), .Y(n186) );
  OAI211X1 U443 ( .C(n189), .D(n257), .A(n198), .B(n211), .Y(N906) );
  NAND2X1 U444 ( .A(mem_14__0_), .B(n191), .Y(n198) );
  OAI211X1 U445 ( .C(n200), .D(n257), .A(n209), .B(n211), .Y(N897) );
  NAND2X1 U446 ( .A(mem_15__0_), .B(n202), .Y(n209) );
  OAI211X1 U447 ( .C(n212), .D(n257), .A(n221), .B(n211), .Y(N888) );
  NAND2X1 U448 ( .A(mem_16__0_), .B(n214), .Y(n221) );
  OAI211X1 U449 ( .C(n224), .D(n257), .A(n233), .B(n211), .Y(N879) );
  NAND2X1 U450 ( .A(mem_17__0_), .B(n226), .Y(n233) );
  OAI211X1 U451 ( .C(n235), .D(n257), .A(n244), .B(n211), .Y(N870) );
  NAND2X1 U452 ( .A(mem_18__0_), .B(n237), .Y(n244) );
  OAI211X1 U453 ( .C(n247), .D(n257), .A(n256), .B(n211), .Y(N861) );
  NAND2X1 U454 ( .A(mem_19__0_), .B(n249), .Y(n256) );
  OAI211X1 U455 ( .C(n258), .D(n257), .A(n267), .B(n211), .Y(N852) );
  NAND2X1 U456 ( .A(mem_20__0_), .B(n260), .Y(n267) );
  OAI211X1 U457 ( .C(n269), .D(n257), .A(n278), .B(n211), .Y(N843) );
  NAND2X1 U458 ( .A(mem_21__0_), .B(n271), .Y(n278) );
  OAI211X1 U459 ( .C(n281), .D(n257), .A(n290), .B(n223), .Y(N834) );
  NAND2X1 U460 ( .A(mem_22__0_), .B(n283), .Y(n290) );
  OAI211X1 U461 ( .C(n292), .D(n268), .A(n301), .B(n223), .Y(N825) );
  NAND2X1 U462 ( .A(mem_23__0_), .B(n294), .Y(n301) );
  OAI211X1 U463 ( .C(n303), .D(n268), .A(n312), .B(n223), .Y(N816) );
  NAND2X1 U464 ( .A(mem_24__0_), .B(n305), .Y(n312) );
  OAI211X1 U465 ( .C(n314), .D(n268), .A(n323), .B(n223), .Y(N807) );
  NAND2X1 U466 ( .A(mem_25__0_), .B(n316), .Y(n323) );
  OAI211X1 U467 ( .C(n325), .D(n268), .A(n334), .B(n223), .Y(N798) );
  NAND2X1 U468 ( .A(mem_26__0_), .B(n327), .Y(n334) );
  OAI211X1 U469 ( .C(n337), .D(n268), .A(n346), .B(n223), .Y(N789) );
  NAND2X1 U470 ( .A(mem_27__0_), .B(n339), .Y(n346) );
  OAI211X1 U471 ( .C(n350), .D(n268), .A(n359), .B(n223), .Y(N780) );
  NAND2X1 U472 ( .A(mem_28__0_), .B(n352), .Y(n359) );
  OAI211X1 U473 ( .C(n130), .D(n349), .A(n138), .B(n291), .Y(N952) );
  NAND2X1 U474 ( .A(mem_9__1_), .B(n132), .Y(n138) );
  OAI211X1 U475 ( .C(n143), .D(n349), .A(n151), .B(n280), .Y(N943) );
  NAND2X1 U476 ( .A(mem_10__1_), .B(n145), .Y(n151) );
  OAI211X1 U477 ( .C(n155), .D(n349), .A(n163), .B(n280), .Y(N934) );
  NAND2X1 U478 ( .A(mem_11__1_), .B(n157), .Y(n163) );
  OAI211X1 U479 ( .C(n166), .D(n349), .A(n174), .B(n291), .Y(N925) );
  NAND2X1 U480 ( .A(mem_12__1_), .B(n168), .Y(n174) );
  OAI211X1 U481 ( .C(n177), .D(n383), .A(n185), .B(n291), .Y(N916) );
  NAND2X1 U482 ( .A(mem_13__1_), .B(n179), .Y(n185) );
  OAI211X1 U483 ( .C(n189), .D(n383), .A(n197), .B(n291), .Y(N907) );
  NAND2X1 U484 ( .A(mem_14__1_), .B(n191), .Y(n197) );
  OAI211X1 U485 ( .C(n200), .D(n383), .A(n208), .B(n291), .Y(N898) );
  NAND2X1 U486 ( .A(mem_15__1_), .B(n202), .Y(n208) );
  OAI211X1 U487 ( .C(n212), .D(n383), .A(n220), .B(n291), .Y(N889) );
  NAND2X1 U488 ( .A(mem_16__1_), .B(n214), .Y(n220) );
  OAI211X1 U489 ( .C(n224), .D(n383), .A(n232), .B(n291), .Y(N880) );
  NAND2X1 U490 ( .A(mem_17__1_), .B(n226), .Y(n232) );
  OAI211X1 U491 ( .C(n235), .D(n383), .A(n243), .B(n291), .Y(N871) );
  NAND2X1 U492 ( .A(mem_18__1_), .B(n237), .Y(n243) );
  OAI211X1 U493 ( .C(n247), .D(n383), .A(n255), .B(n291), .Y(N862) );
  NAND2X1 U494 ( .A(mem_19__1_), .B(n249), .Y(n255) );
  OAI211X1 U495 ( .C(n258), .D(n383), .A(n266), .B(n291), .Y(N853) );
  NAND2X1 U496 ( .A(mem_20__1_), .B(n260), .Y(n266) );
  OAI211X1 U497 ( .C(n269), .D(n383), .A(n277), .B(n335), .Y(N844) );
  NAND2X1 U498 ( .A(mem_21__1_), .B(n271), .Y(n277) );
  OAI211X1 U499 ( .C(n281), .D(n383), .A(n289), .B(n335), .Y(N835) );
  NAND2X1 U500 ( .A(mem_22__1_), .B(n283), .Y(n289) );
  OAI211X1 U501 ( .C(n292), .D(n384), .A(n300), .B(n335), .Y(N826) );
  NAND2X1 U502 ( .A(mem_23__1_), .B(n294), .Y(n300) );
  OAI211X1 U503 ( .C(n303), .D(n384), .A(n311), .B(n335), .Y(N817) );
  NAND2X1 U504 ( .A(mem_24__1_), .B(n305), .Y(n311) );
  OAI211X1 U505 ( .C(n314), .D(n384), .A(n322), .B(n335), .Y(N808) );
  NAND2X1 U506 ( .A(mem_25__1_), .B(n316), .Y(n322) );
  OAI211X1 U507 ( .C(n325), .D(n384), .A(n333), .B(n335), .Y(N799) );
  NAND2X1 U508 ( .A(mem_26__1_), .B(n327), .Y(n333) );
  OAI211X1 U509 ( .C(n337), .D(n384), .A(n345), .B(n335), .Y(N790) );
  NAND2X1 U510 ( .A(mem_27__1_), .B(n339), .Y(n345) );
  OAI211X1 U511 ( .C(n350), .D(n384), .A(n358), .B(n335), .Y(N781) );
  NAND2X1 U512 ( .A(mem_28__1_), .B(n352), .Y(n358) );
  OAI211X1 U513 ( .C(n130), .D(n423), .A(n137), .B(n420), .Y(N953) );
  NAND2X1 U514 ( .A(mem_9__2_), .B(n132), .Y(n137) );
  OAI211X1 U515 ( .C(n143), .D(n423), .A(n150), .B(n419), .Y(N944) );
  NAND2X1 U516 ( .A(mem_10__2_), .B(n145), .Y(n150) );
  OAI211X1 U517 ( .C(n155), .D(n423), .A(n162), .B(n419), .Y(N935) );
  NAND2X1 U518 ( .A(mem_11__2_), .B(n157), .Y(n162) );
  OAI211X1 U519 ( .C(n166), .D(n423), .A(n173), .B(n420), .Y(N926) );
  NAND2X1 U520 ( .A(mem_12__2_), .B(n168), .Y(n173) );
  OAI211X1 U521 ( .C(n177), .D(n424), .A(n184), .B(n420), .Y(N917) );
  NAND2X1 U522 ( .A(mem_13__2_), .B(n179), .Y(n184) );
  OAI211X1 U523 ( .C(n189), .D(n424), .A(n196), .B(n420), .Y(N908) );
  NAND2X1 U524 ( .A(mem_14__2_), .B(n191), .Y(n196) );
  OAI211X1 U525 ( .C(n200), .D(n424), .A(n207), .B(n420), .Y(N899) );
  NAND2X1 U526 ( .A(mem_15__2_), .B(n202), .Y(n207) );
  OAI211X1 U527 ( .C(n212), .D(n424), .A(n219), .B(n420), .Y(N890) );
  NAND2X1 U528 ( .A(mem_16__2_), .B(n214), .Y(n219) );
  OAI211X1 U529 ( .C(n224), .D(n424), .A(n231), .B(n420), .Y(N881) );
  NAND2X1 U530 ( .A(mem_17__2_), .B(n226), .Y(n231) );
  OAI211X1 U531 ( .C(n235), .D(n424), .A(n242), .B(n420), .Y(N872) );
  NAND2X1 U532 ( .A(mem_18__2_), .B(n237), .Y(n242) );
  OAI211X1 U533 ( .C(n247), .D(n424), .A(n254), .B(n420), .Y(N863) );
  NAND2X1 U534 ( .A(mem_19__2_), .B(n249), .Y(n254) );
  OAI211X1 U535 ( .C(n258), .D(n424), .A(n265), .B(n420), .Y(N854) );
  NAND2X1 U536 ( .A(mem_20__2_), .B(n260), .Y(n265) );
  OAI211X1 U537 ( .C(n269), .D(n424), .A(n276), .B(n421), .Y(N845) );
  NAND2X1 U538 ( .A(mem_21__2_), .B(n271), .Y(n276) );
  OAI211X1 U539 ( .C(n281), .D(n424), .A(n288), .B(n421), .Y(N836) );
  NAND2X1 U540 ( .A(mem_22__2_), .B(n283), .Y(n288) );
  OAI211X1 U541 ( .C(n292), .D(n425), .A(n299), .B(n421), .Y(N827) );
  NAND2X1 U542 ( .A(mem_23__2_), .B(n294), .Y(n299) );
  OAI211X1 U543 ( .C(n303), .D(n425), .A(n310), .B(n421), .Y(N818) );
  NAND2X1 U544 ( .A(mem_24__2_), .B(n305), .Y(n310) );
  OAI211X1 U545 ( .C(n314), .D(n425), .A(n321), .B(n421), .Y(N809) );
  NAND2X1 U546 ( .A(mem_25__2_), .B(n316), .Y(n321) );
  OAI211X1 U547 ( .C(n325), .D(n425), .A(n332), .B(n421), .Y(N800) );
  NAND2X1 U548 ( .A(mem_26__2_), .B(n327), .Y(n332) );
  OAI211X1 U549 ( .C(n337), .D(n425), .A(n344), .B(n421), .Y(N791) );
  NAND2X1 U550 ( .A(mem_27__2_), .B(n339), .Y(n344) );
  OAI211X1 U551 ( .C(n350), .D(n425), .A(n357), .B(n421), .Y(N782) );
  NAND2X1 U552 ( .A(mem_28__2_), .B(n352), .Y(n357) );
  OAI211X1 U553 ( .C(n130), .D(n431), .A(n136), .B(n428), .Y(N954) );
  NAND2X1 U554 ( .A(mem_9__3_), .B(n132), .Y(n136) );
  OAI211X1 U555 ( .C(n143), .D(n431), .A(n149), .B(n427), .Y(N945) );
  NAND2X1 U556 ( .A(mem_10__3_), .B(n145), .Y(n149) );
  OAI211X1 U557 ( .C(n155), .D(n431), .A(n161), .B(n427), .Y(N936) );
  NAND2X1 U558 ( .A(mem_11__3_), .B(n157), .Y(n161) );
  OAI211X1 U559 ( .C(n166), .D(n431), .A(n172), .B(n428), .Y(N927) );
  NAND2X1 U560 ( .A(mem_12__3_), .B(n168), .Y(n172) );
  OAI211X1 U561 ( .C(n177), .D(n432), .A(n183), .B(n428), .Y(N918) );
  NAND2X1 U562 ( .A(mem_13__3_), .B(n179), .Y(n183) );
  OAI211X1 U563 ( .C(n189), .D(n432), .A(n195), .B(n428), .Y(N909) );
  NAND2X1 U564 ( .A(mem_14__3_), .B(n191), .Y(n195) );
  OAI211X1 U565 ( .C(n200), .D(n432), .A(n206), .B(n428), .Y(N900) );
  NAND2X1 U566 ( .A(mem_15__3_), .B(n202), .Y(n206) );
  OAI211X1 U567 ( .C(n212), .D(n432), .A(n218), .B(n428), .Y(N891) );
  NAND2X1 U568 ( .A(mem_16__3_), .B(n214), .Y(n218) );
  OAI211X1 U569 ( .C(n224), .D(n432), .A(n230), .B(n428), .Y(N882) );
  NAND2X1 U570 ( .A(mem_17__3_), .B(n226), .Y(n230) );
  OAI211X1 U571 ( .C(n235), .D(n432), .A(n241), .B(n428), .Y(N873) );
  NAND2X1 U572 ( .A(mem_18__3_), .B(n237), .Y(n241) );
  OAI211X1 U573 ( .C(n247), .D(n432), .A(n253), .B(n428), .Y(N864) );
  NAND2X1 U574 ( .A(mem_19__3_), .B(n249), .Y(n253) );
  OAI211X1 U575 ( .C(n258), .D(n432), .A(n264), .B(n428), .Y(N855) );
  NAND2X1 U576 ( .A(mem_20__3_), .B(n260), .Y(n264) );
  OAI211X1 U577 ( .C(n269), .D(n432), .A(n275), .B(n429), .Y(N846) );
  NAND2X1 U578 ( .A(mem_21__3_), .B(n271), .Y(n275) );
  OAI211X1 U579 ( .C(n281), .D(n432), .A(n287), .B(n429), .Y(N837) );
  NAND2X1 U580 ( .A(mem_22__3_), .B(n283), .Y(n287) );
  OAI211X1 U581 ( .C(n292), .D(n433), .A(n298), .B(n429), .Y(N828) );
  NAND2X1 U582 ( .A(mem_23__3_), .B(n294), .Y(n298) );
  OAI211X1 U583 ( .C(n303), .D(n433), .A(n309), .B(n429), .Y(N819) );
  NAND2X1 U584 ( .A(mem_24__3_), .B(n305), .Y(n309) );
  OAI211X1 U585 ( .C(n314), .D(n433), .A(n320), .B(n429), .Y(N810) );
  NAND2X1 U586 ( .A(mem_25__3_), .B(n316), .Y(n320) );
  OAI211X1 U587 ( .C(n325), .D(n433), .A(n331), .B(n429), .Y(N801) );
  NAND2X1 U588 ( .A(mem_26__3_), .B(n327), .Y(n331) );
  OAI211X1 U589 ( .C(n337), .D(n433), .A(n343), .B(n429), .Y(N792) );
  NAND2X1 U590 ( .A(mem_27__3_), .B(n339), .Y(n343) );
  OAI211X1 U591 ( .C(n350), .D(n433), .A(n356), .B(n429), .Y(N783) );
  NAND2X1 U592 ( .A(mem_28__3_), .B(n352), .Y(n356) );
  OAI211X1 U593 ( .C(n130), .D(n22), .A(n135), .B(n20), .Y(N955) );
  NAND2X1 U594 ( .A(mem_9__4_), .B(n132), .Y(n135) );
  OAI211X1 U595 ( .C(n143), .D(n22), .A(n148), .B(n20), .Y(N946) );
  NAND2X1 U596 ( .A(mem_10__4_), .B(n145), .Y(n148) );
  OAI211X1 U597 ( .C(n155), .D(n22), .A(n160), .B(n20), .Y(N937) );
  NAND2X1 U598 ( .A(mem_11__4_), .B(n157), .Y(n160) );
  OAI211X1 U599 ( .C(n166), .D(n22), .A(n171), .B(n20), .Y(N928) );
  NAND2X1 U600 ( .A(mem_12__4_), .B(n168), .Y(n171) );
  OAI211X1 U601 ( .C(n177), .D(n22), .A(n182), .B(n20), .Y(N919) );
  NAND2X1 U602 ( .A(mem_13__4_), .B(n179), .Y(n182) );
  OAI211X1 U603 ( .C(n189), .D(n23), .A(n194), .B(n20), .Y(N910) );
  NAND2X1 U604 ( .A(mem_14__4_), .B(n191), .Y(n194) );
  OAI211X1 U605 ( .C(n200), .D(n23), .A(n205), .B(n20), .Y(N901) );
  NAND2X1 U606 ( .A(mem_15__4_), .B(n202), .Y(n205) );
  OAI211X1 U607 ( .C(n212), .D(n23), .A(n217), .B(n20), .Y(N892) );
  NAND2X1 U608 ( .A(mem_16__4_), .B(n214), .Y(n217) );
  OAI211X1 U609 ( .C(n224), .D(n23), .A(n229), .B(n19), .Y(N883) );
  NAND2X1 U610 ( .A(mem_17__4_), .B(n226), .Y(n229) );
  OAI211X1 U611 ( .C(n235), .D(n23), .A(n240), .B(n19), .Y(N874) );
  NAND2X1 U612 ( .A(mem_18__4_), .B(n237), .Y(n240) );
  OAI211X1 U613 ( .C(n247), .D(n23), .A(n252), .B(n19), .Y(N865) );
  NAND2X1 U614 ( .A(mem_19__4_), .B(n249), .Y(n252) );
  OAI211X1 U615 ( .C(n258), .D(n23), .A(n263), .B(n19), .Y(N856) );
  NAND2X1 U616 ( .A(mem_20__4_), .B(n260), .Y(n263) );
  OAI211X1 U617 ( .C(n269), .D(n23), .A(n274), .B(n19), .Y(N847) );
  NAND2X1 U618 ( .A(mem_21__4_), .B(n271), .Y(n274) );
  OAI211X1 U619 ( .C(n281), .D(n23), .A(n286), .B(n19), .Y(N838) );
  NAND2X1 U620 ( .A(mem_22__4_), .B(n283), .Y(n286) );
  OAI211X1 U621 ( .C(n292), .D(n23), .A(n297), .B(n19), .Y(N829) );
  NAND2X1 U622 ( .A(mem_23__4_), .B(n294), .Y(n297) );
  OAI211X1 U623 ( .C(n303), .D(n24), .A(n308), .B(n19), .Y(N820) );
  NAND2X1 U624 ( .A(mem_24__4_), .B(n305), .Y(n308) );
  OAI211X1 U625 ( .C(n314), .D(n24), .A(n319), .B(n19), .Y(N811) );
  NAND2X1 U626 ( .A(mem_25__4_), .B(n316), .Y(n319) );
  OAI211X1 U627 ( .C(n325), .D(n24), .A(n330), .B(n19), .Y(N802) );
  NAND2X1 U628 ( .A(mem_26__4_), .B(n327), .Y(n330) );
  OAI211X1 U629 ( .C(n337), .D(n24), .A(n342), .B(n18), .Y(N793) );
  NAND2X1 U630 ( .A(mem_27__4_), .B(n339), .Y(n342) );
  OAI211X1 U631 ( .C(n350), .D(n24), .A(n355), .B(n18), .Y(N784) );
  NAND2X1 U632 ( .A(mem_28__4_), .B(n352), .Y(n355) );
  OAI211X1 U633 ( .C(n130), .D(n30), .A(n134), .B(n28), .Y(N956) );
  NAND2X1 U634 ( .A(mem_9__5_), .B(n132), .Y(n134) );
  OAI211X1 U635 ( .C(n143), .D(n30), .A(n147), .B(n28), .Y(N947) );
  NAND2X1 U636 ( .A(mem_10__5_), .B(n145), .Y(n147) );
  OAI211X1 U637 ( .C(n155), .D(n30), .A(n159), .B(n28), .Y(N938) );
  NAND2X1 U638 ( .A(mem_11__5_), .B(n157), .Y(n159) );
  OAI211X1 U639 ( .C(n166), .D(n30), .A(n170), .B(n28), .Y(N929) );
  NAND2X1 U640 ( .A(mem_12__5_), .B(n168), .Y(n170) );
  OAI211X1 U641 ( .C(n177), .D(n30), .A(n181), .B(n28), .Y(N920) );
  NAND2X1 U642 ( .A(mem_13__5_), .B(n179), .Y(n181) );
  OAI211X1 U643 ( .C(n189), .D(n31), .A(n193), .B(n28), .Y(N911) );
  NAND2X1 U644 ( .A(mem_14__5_), .B(n191), .Y(n193) );
  OAI211X1 U645 ( .C(n200), .D(n31), .A(n204), .B(n28), .Y(N902) );
  NAND2X1 U646 ( .A(mem_15__5_), .B(n202), .Y(n204) );
  OAI211X1 U647 ( .C(n212), .D(n31), .A(n216), .B(n28), .Y(N893) );
  NAND2X1 U648 ( .A(mem_16__5_), .B(n214), .Y(n216) );
  OAI211X1 U649 ( .C(n224), .D(n31), .A(n228), .B(n27), .Y(N884) );
  NAND2X1 U650 ( .A(mem_17__5_), .B(n226), .Y(n228) );
  OAI211X1 U651 ( .C(n235), .D(n31), .A(n239), .B(n27), .Y(N875) );
  NAND2X1 U652 ( .A(mem_18__5_), .B(n237), .Y(n239) );
  OAI211X1 U653 ( .C(n247), .D(n31), .A(n251), .B(n27), .Y(N866) );
  NAND2X1 U654 ( .A(mem_19__5_), .B(n249), .Y(n251) );
  OAI211X1 U655 ( .C(n258), .D(n31), .A(n262), .B(n27), .Y(N857) );
  NAND2X1 U656 ( .A(mem_20__5_), .B(n260), .Y(n262) );
  OAI211X1 U657 ( .C(n269), .D(n31), .A(n273), .B(n27), .Y(N848) );
  NAND2X1 U658 ( .A(mem_21__5_), .B(n271), .Y(n273) );
  OAI211X1 U659 ( .C(n281), .D(n31), .A(n285), .B(n27), .Y(N839) );
  NAND2X1 U660 ( .A(mem_22__5_), .B(n283), .Y(n285) );
  OAI211X1 U661 ( .C(n292), .D(n31), .A(n296), .B(n27), .Y(N830) );
  NAND2X1 U662 ( .A(mem_23__5_), .B(n294), .Y(n296) );
  OAI211X1 U663 ( .C(n303), .D(n32), .A(n307), .B(n27), .Y(N821) );
  NAND2X1 U664 ( .A(mem_24__5_), .B(n305), .Y(n307) );
  OAI211X1 U665 ( .C(n314), .D(n32), .A(n318), .B(n27), .Y(N812) );
  NAND2X1 U666 ( .A(mem_25__5_), .B(n316), .Y(n318) );
  OAI211X1 U667 ( .C(n325), .D(n32), .A(n329), .B(n27), .Y(N803) );
  NAND2X1 U668 ( .A(mem_26__5_), .B(n327), .Y(n329) );
  OAI211X1 U669 ( .C(n337), .D(n32), .A(n341), .B(n26), .Y(N794) );
  NAND2X1 U670 ( .A(mem_27__5_), .B(n339), .Y(n341) );
  OAI211X1 U671 ( .C(n350), .D(n32), .A(n354), .B(n26), .Y(N785) );
  NAND2X1 U672 ( .A(mem_28__5_), .B(n352), .Y(n354) );
  OAI211X1 U673 ( .C(n130), .D(n38), .A(n133), .B(n36), .Y(N957) );
  NAND2X1 U674 ( .A(mem_9__6_), .B(n132), .Y(n133) );
  OAI211X1 U675 ( .C(n143), .D(n38), .A(n146), .B(n36), .Y(N948) );
  NAND2X1 U676 ( .A(mem_10__6_), .B(n145), .Y(n146) );
  OAI211X1 U677 ( .C(n155), .D(n38), .A(n158), .B(n36), .Y(N939) );
  NAND2X1 U678 ( .A(mem_11__6_), .B(n157), .Y(n158) );
  OAI211X1 U679 ( .C(n166), .D(n38), .A(n169), .B(n36), .Y(N930) );
  NAND2X1 U680 ( .A(mem_12__6_), .B(n168), .Y(n169) );
  OAI211X1 U681 ( .C(n177), .D(n38), .A(n180), .B(n36), .Y(N921) );
  NAND2X1 U682 ( .A(mem_13__6_), .B(n179), .Y(n180) );
  OAI211X1 U683 ( .C(n189), .D(n39), .A(n192), .B(n36), .Y(N912) );
  NAND2X1 U684 ( .A(mem_14__6_), .B(n191), .Y(n192) );
  OAI211X1 U685 ( .C(n200), .D(n39), .A(n203), .B(n36), .Y(N903) );
  NAND2X1 U686 ( .A(mem_15__6_), .B(n202), .Y(n203) );
  OAI211X1 U687 ( .C(n212), .D(n39), .A(n215), .B(n36), .Y(N894) );
  NAND2X1 U688 ( .A(mem_16__6_), .B(n214), .Y(n215) );
  OAI211X1 U689 ( .C(n224), .D(n39), .A(n227), .B(n35), .Y(N885) );
  NAND2X1 U690 ( .A(mem_17__6_), .B(n226), .Y(n227) );
  OAI211X1 U691 ( .C(n235), .D(n39), .A(n238), .B(n35), .Y(N876) );
  NAND2X1 U692 ( .A(mem_18__6_), .B(n237), .Y(n238) );
  OAI211X1 U693 ( .C(n247), .D(n39), .A(n250), .B(n35), .Y(N867) );
  NAND2X1 U694 ( .A(mem_19__6_), .B(n249), .Y(n250) );
  OAI211X1 U695 ( .C(n258), .D(n39), .A(n261), .B(n35), .Y(N858) );
  NAND2X1 U696 ( .A(mem_20__6_), .B(n260), .Y(n261) );
  OAI211X1 U697 ( .C(n269), .D(n39), .A(n272), .B(n35), .Y(N849) );
  NAND2X1 U698 ( .A(mem_21__6_), .B(n271), .Y(n272) );
  OAI211X1 U699 ( .C(n281), .D(n39), .A(n284), .B(n35), .Y(N840) );
  NAND2X1 U700 ( .A(mem_22__6_), .B(n283), .Y(n284) );
  OAI211X1 U701 ( .C(n292), .D(n39), .A(n295), .B(n35), .Y(N831) );
  NAND2X1 U702 ( .A(mem_23__6_), .B(n294), .Y(n295) );
  OAI211X1 U703 ( .C(n303), .D(n40), .A(n306), .B(n35), .Y(N822) );
  NAND2X1 U704 ( .A(mem_24__6_), .B(n305), .Y(n306) );
  OAI211X1 U705 ( .C(n314), .D(n40), .A(n317), .B(n35), .Y(N813) );
  NAND2X1 U706 ( .A(mem_25__6_), .B(n316), .Y(n317) );
  OAI211X1 U707 ( .C(n325), .D(n40), .A(n328), .B(n35), .Y(N804) );
  NAND2X1 U708 ( .A(mem_26__6_), .B(n327), .Y(n328) );
  OAI211X1 U709 ( .C(n337), .D(n40), .A(n340), .B(n34), .Y(N795) );
  NAND2X1 U710 ( .A(mem_27__6_), .B(n339), .Y(n340) );
  OAI211X1 U711 ( .C(n350), .D(n40), .A(n353), .B(n34), .Y(N786) );
  NAND2X1 U712 ( .A(mem_28__6_), .B(n352), .Y(n353) );
  OAI211X1 U713 ( .C(n130), .D(n46), .A(n131), .B(n44), .Y(N958) );
  NAND2X1 U714 ( .A(mem_9__7_), .B(n132), .Y(n131) );
  OAI211X1 U715 ( .C(n143), .D(n46), .A(n144), .B(n44), .Y(N949) );
  NAND2X1 U716 ( .A(mem_10__7_), .B(n145), .Y(n144) );
  OAI211X1 U717 ( .C(n155), .D(n46), .A(n156), .B(n44), .Y(N940) );
  NAND2X1 U718 ( .A(mem_11__7_), .B(n157), .Y(n156) );
  OAI211X1 U719 ( .C(n166), .D(n46), .A(n167), .B(n44), .Y(N931) );
  NAND2X1 U720 ( .A(mem_12__7_), .B(n168), .Y(n167) );
  OAI211X1 U721 ( .C(n177), .D(n46), .A(n178), .B(n44), .Y(N922) );
  NAND2X1 U722 ( .A(mem_13__7_), .B(n179), .Y(n178) );
  OAI211X1 U723 ( .C(n189), .D(n47), .A(n190), .B(n44), .Y(N913) );
  NAND2X1 U724 ( .A(mem_14__7_), .B(n191), .Y(n190) );
  OAI211X1 U725 ( .C(n200), .D(n47), .A(n201), .B(n44), .Y(N904) );
  NAND2X1 U726 ( .A(mem_15__7_), .B(n202), .Y(n201) );
  OAI211X1 U727 ( .C(n212), .D(n47), .A(n213), .B(n44), .Y(N895) );
  NAND2X1 U728 ( .A(mem_16__7_), .B(n214), .Y(n213) );
  OAI211X1 U729 ( .C(n224), .D(n47), .A(n225), .B(n43), .Y(N886) );
  NAND2X1 U730 ( .A(mem_17__7_), .B(n226), .Y(n225) );
  OAI211X1 U731 ( .C(n235), .D(n47), .A(n236), .B(n43), .Y(N877) );
  NAND2X1 U732 ( .A(mem_18__7_), .B(n237), .Y(n236) );
  OAI211X1 U733 ( .C(n247), .D(n47), .A(n248), .B(n43), .Y(N868) );
  NAND2X1 U734 ( .A(mem_19__7_), .B(n249), .Y(n248) );
  OAI211X1 U735 ( .C(n258), .D(n47), .A(n259), .B(n43), .Y(N859) );
  NAND2X1 U736 ( .A(mem_20__7_), .B(n260), .Y(n259) );
  OAI211X1 U737 ( .C(n269), .D(n47), .A(n270), .B(n43), .Y(N850) );
  NAND2X1 U738 ( .A(mem_21__7_), .B(n271), .Y(n270) );
  OAI211X1 U739 ( .C(n281), .D(n47), .A(n282), .B(n43), .Y(N841) );
  NAND2X1 U740 ( .A(mem_22__7_), .B(n283), .Y(n282) );
  OAI211X1 U741 ( .C(n292), .D(n47), .A(n293), .B(n43), .Y(N832) );
  NAND2X1 U742 ( .A(mem_23__7_), .B(n294), .Y(n293) );
  OAI211X1 U743 ( .C(n303), .D(n49), .A(n304), .B(n43), .Y(N823) );
  NAND2X1 U744 ( .A(mem_24__7_), .B(n305), .Y(n304) );
  OAI211X1 U745 ( .C(n314), .D(n49), .A(n315), .B(n43), .Y(N814) );
  NAND2X1 U746 ( .A(mem_25__7_), .B(n316), .Y(n315) );
  OAI211X1 U747 ( .C(n325), .D(n49), .A(n326), .B(n43), .Y(N805) );
  NAND2X1 U748 ( .A(mem_26__7_), .B(n327), .Y(n326) );
  OAI211X1 U749 ( .C(n337), .D(n49), .A(n338), .B(n42), .Y(N796) );
  NAND2X1 U750 ( .A(mem_27__7_), .B(n339), .Y(n338) );
  OAI211X1 U751 ( .C(n350), .D(n49), .A(n351), .B(n42), .Y(N787) );
  NAND2X1 U752 ( .A(mem_28__7_), .B(n352), .Y(n351) );
  OAI211X1 U753 ( .C(n361), .D(n268), .A(n370), .B(n223), .Y(N771) );
  NAND2X1 U754 ( .A(mem_29__0_), .B(n363), .Y(n370) );
  OAI211X1 U755 ( .C(n373), .D(n268), .A(n382), .B(n223), .Y(N762) );
  NAND2X1 U756 ( .A(mem_30__0_), .B(n375), .Y(n382) );
  OAI211X1 U757 ( .C(n385), .D(n268), .A(n394), .B(n223), .Y(N753) );
  NAND2X1 U758 ( .A(mem_31__0_), .B(n387), .Y(n394) );
  OAI211X1 U759 ( .C(n17), .D(n268), .A(n405), .B(n64), .Y(N744) );
  NAND2X1 U760 ( .A(mem_32__0_), .B(n398), .Y(n405) );
  OAI211X1 U761 ( .C(n361), .D(n384), .A(n369), .B(n335), .Y(N772) );
  NAND2X1 U762 ( .A(mem_29__1_), .B(n363), .Y(n369) );
  OAI211X1 U763 ( .C(n373), .D(n384), .A(n381), .B(n335), .Y(N763) );
  NAND2X1 U764 ( .A(mem_30__1_), .B(n375), .Y(n381) );
  OAI211X1 U765 ( .C(n385), .D(n384), .A(n393), .B(n61), .Y(N754) );
  NAND2X1 U766 ( .A(mem_31__1_), .B(n387), .Y(n393) );
  OAI211X1 U767 ( .C(n17), .D(n384), .A(n404), .B(n61), .Y(N745) );
  NAND2X1 U768 ( .A(mem_32__1_), .B(n398), .Y(n404) );
  OAI211X1 U769 ( .C(n361), .D(n425), .A(n368), .B(n421), .Y(N773) );
  NAND2X1 U770 ( .A(mem_29__2_), .B(n363), .Y(n368) );
  OAI211X1 U771 ( .C(n373), .D(n425), .A(n380), .B(n421), .Y(N764) );
  NAND2X1 U772 ( .A(mem_30__2_), .B(n375), .Y(n380) );
  OAI211X1 U773 ( .C(n385), .D(n425), .A(n392), .B(n58), .Y(N755) );
  NAND2X1 U774 ( .A(mem_31__2_), .B(n387), .Y(n392) );
  OAI211X1 U775 ( .C(n17), .D(n425), .A(n403), .B(n58), .Y(N746) );
  NAND2X1 U776 ( .A(mem_32__2_), .B(n398), .Y(n403) );
  OAI211X1 U777 ( .C(n361), .D(n433), .A(n367), .B(n429), .Y(N774) );
  NAND2X1 U778 ( .A(mem_29__3_), .B(n363), .Y(n367) );
  OAI211X1 U779 ( .C(n373), .D(n433), .A(n379), .B(n429), .Y(N765) );
  NAND2X1 U780 ( .A(mem_30__3_), .B(n375), .Y(n379) );
  OAI211X1 U781 ( .C(n385), .D(n433), .A(n391), .B(n54), .Y(N756) );
  NAND2X1 U782 ( .A(mem_31__3_), .B(n387), .Y(n391) );
  OAI211X1 U783 ( .C(n17), .D(n433), .A(n402), .B(n54), .Y(N747) );
  NAND2X1 U784 ( .A(mem_32__3_), .B(n398), .Y(n402) );
  OAI211X1 U785 ( .C(n361), .D(n24), .A(n366), .B(n18), .Y(N775) );
  NAND2X1 U786 ( .A(mem_29__4_), .B(n363), .Y(n366) );
  OAI211X1 U787 ( .C(n373), .D(n24), .A(n378), .B(n18), .Y(N766) );
  NAND2X1 U788 ( .A(mem_30__4_), .B(n375), .Y(n378) );
  OAI211X1 U789 ( .C(n385), .D(n24), .A(n390), .B(n18), .Y(N757) );
  NAND2X1 U790 ( .A(mem_31__4_), .B(n387), .Y(n390) );
  OAI211X1 U791 ( .C(n17), .D(n24), .A(n401), .B(n18), .Y(N748) );
  NAND2X1 U792 ( .A(mem_32__4_), .B(n398), .Y(n401) );
  OAI211X1 U793 ( .C(n407), .D(n24), .A(n412), .B(n18), .Y(N739) );
  NAND2X1 U794 ( .A(mem_33__4_), .B(n409), .Y(n412) );
  OAI211X1 U795 ( .C(n361), .D(n32), .A(n365), .B(n26), .Y(N776) );
  NAND2X1 U796 ( .A(mem_29__5_), .B(n363), .Y(n365) );
  OAI211X1 U797 ( .C(n373), .D(n32), .A(n377), .B(n26), .Y(N767) );
  NAND2X1 U798 ( .A(mem_30__5_), .B(n375), .Y(n377) );
  OAI211X1 U799 ( .C(n385), .D(n32), .A(n389), .B(n26), .Y(N758) );
  NAND2X1 U800 ( .A(mem_31__5_), .B(n387), .Y(n389) );
  OAI211X1 U801 ( .C(n17), .D(n32), .A(n400), .B(n26), .Y(N749) );
  NAND2X1 U802 ( .A(mem_32__5_), .B(n398), .Y(n400) );
  OAI211X1 U803 ( .C(n407), .D(n32), .A(n411), .B(n26), .Y(N740) );
  NAND2X1 U804 ( .A(mem_33__5_), .B(n409), .Y(n411) );
  OAI211X1 U805 ( .C(n361), .D(n40), .A(n364), .B(n34), .Y(N777) );
  NAND2X1 U806 ( .A(mem_29__6_), .B(n363), .Y(n364) );
  OAI211X1 U807 ( .C(n373), .D(n40), .A(n376), .B(n34), .Y(N768) );
  NAND2X1 U808 ( .A(mem_30__6_), .B(n375), .Y(n376) );
  OAI211X1 U809 ( .C(n385), .D(n40), .A(n388), .B(n34), .Y(N759) );
  NAND2X1 U810 ( .A(mem_31__6_), .B(n387), .Y(n388) );
  OAI211X1 U811 ( .C(n17), .D(n40), .A(n399), .B(n34), .Y(N750) );
  NAND2X1 U812 ( .A(mem_32__6_), .B(n398), .Y(n399) );
  OAI211X1 U813 ( .C(n407), .D(n40), .A(n410), .B(n34), .Y(N741) );
  NAND2X1 U814 ( .A(mem_33__6_), .B(n409), .Y(n410) );
  OAI211X1 U815 ( .C(n361), .D(n49), .A(n362), .B(n42), .Y(N778) );
  NAND2X1 U816 ( .A(mem_29__7_), .B(n363), .Y(n362) );
  OAI211X1 U817 ( .C(n373), .D(n49), .A(n374), .B(n42), .Y(N769) );
  NAND2X1 U818 ( .A(mem_30__7_), .B(n375), .Y(n374) );
  OAI211X1 U819 ( .C(n385), .D(n49), .A(n386), .B(n42), .Y(N760) );
  NAND2X1 U820 ( .A(mem_31__7_), .B(n387), .Y(n386) );
  OAI211X1 U821 ( .C(n17), .D(n49), .A(n397), .B(n42), .Y(N751) );
  NAND2X1 U822 ( .A(mem_32__7_), .B(n398), .Y(n397) );
  OAI211X1 U823 ( .C(n407), .D(n49), .A(n408), .B(n42), .Y(N742) );
  NAND2X1 U824 ( .A(mem_33__7_), .B(n409), .Y(n408) );
  OAI211X1 U825 ( .C(n458), .D(n63), .A(n467), .B(n199), .Y(N1005) );
  NAND2X1 U826 ( .A(dat_7_1[16]), .B(n460), .Y(n467) );
  OAI211X1 U827 ( .C(n458), .D(n60), .A(n280), .B(n466), .Y(N1006) );
  NAND2X1 U828 ( .A(dat_7_1[17]), .B(n460), .Y(n466) );
  OAI211X1 U829 ( .C(n458), .D(n57), .A(n419), .B(n465), .Y(N1007) );
  NAND2X1 U830 ( .A(dat_7_1[18]), .B(n460), .Y(n465) );
  OAI211X1 U831 ( .C(n458), .D(n53), .A(n427), .B(n464), .Y(N1008) );
  NAND2X1 U832 ( .A(dat_7_1[19]), .B(n460), .Y(n464) );
  OAI211X1 U833 ( .C(n458), .D(n81), .A(n463), .B(n18), .Y(N1009) );
  NAND2X1 U834 ( .A(dat_7_1[20]), .B(n460), .Y(n463) );
  OAI211X1 U835 ( .C(n52), .D(n81), .A(n472), .B(n18), .Y(N1000) );
  NAND2X1 U836 ( .A(dat_7_1[28]), .B(n56), .Y(n472) );
  OAI211X1 U837 ( .C(n52), .D(n78), .A(n26), .B(n471), .Y(N1001) );
  NAND2X1 U838 ( .A(dat_7_1[29]), .B(n56), .Y(n471) );
  OAI211X1 U839 ( .C(n52), .D(n75), .A(n34), .B(n470), .Y(N1002) );
  NAND2X1 U840 ( .A(dat_7_1[30]), .B(n56), .Y(n470) );
  OAI211X1 U841 ( .C(n52), .D(n71), .A(n42), .B(n469), .Y(N1003) );
  NAND2X1 U842 ( .A(dat_7_1[31]), .B(n56), .Y(n469) );
  OAI211X1 U843 ( .C(n458), .D(n78), .A(n462), .B(n26), .Y(N1010) );
  NAND2X1 U844 ( .A(dat_7_1[21]), .B(n460), .Y(n462) );
  OAI211X1 U845 ( .C(n458), .D(n75), .A(n461), .B(n34), .Y(N1011) );
  NAND2X1 U846 ( .A(dat_7_1[22]), .B(n460), .Y(n461) );
  OAI211X1 U847 ( .C(n458), .D(n71), .A(n459), .B(n42), .Y(N1012) );
  NAND2X1 U848 ( .A(dat_7_1[23]), .B(n460), .Y(n459) );
  OAI211X1 U849 ( .C(n407), .D(n63), .A(n416), .B(n64), .Y(N735) );
  NAND2X1 U850 ( .A(mem_33__0_), .B(n409), .Y(n416) );
  OAI211X1 U851 ( .C(n407), .D(n60), .A(n415), .B(n280), .Y(N736) );
  NAND2X1 U852 ( .A(mem_33__1_), .B(n409), .Y(n415) );
  OAI211X1 U853 ( .C(n407), .D(n57), .A(n414), .B(n419), .Y(N737) );
  NAND2X1 U854 ( .A(mem_33__2_), .B(n409), .Y(n414) );
  OAI211X1 U855 ( .C(n407), .D(n53), .A(n413), .B(n427), .Y(N738) );
  NAND2X1 U856 ( .A(mem_33__3_), .B(n409), .Y(n413) );
  MUX2X1 U857 ( .D0(fifowdat[7]), .D1(dat_7_1[7]), .S(n12), .Y(N1030) );
  MUX2X1 U858 ( .D0(fifowdat[2]), .D1(dat_7_1[2]), .S(n12), .Y(N1025) );
  MUX2X1 U859 ( .D0(fifowdat[4]), .D1(dat_7_1[4]), .S(n12), .Y(N1027) );
  MUX2X1 U860 ( .D0(fifowdat[3]), .D1(dat_7_1[3]), .S(n12), .Y(N1026) );
  MUX2X1 U861 ( .D0(fifowdat[0]), .D1(dat_7_1[0]), .S(n12), .Y(N1023) );
  MUX2X1 U862 ( .D0(fifowdat[6]), .D1(dat_7_1[6]), .S(n12), .Y(N1029) );
  MUX2X1 U863 ( .D0(fifowdat[1]), .D1(dat_7_1[1]), .S(n12), .Y(N1024) );
  MUX2X1 U864 ( .D0(fifowdat[5]), .D1(dat_7_1[5]), .S(n12), .Y(N1028) );
  NAND2X1 U865 ( .A(r_psh), .B(r_last), .Y(n48) );
  MUX2IX1 U866 ( .D0(r_wdat[0]), .D1(prx_wdat[0]), .S(prx_psh), .Y(n63) );
  MUX2IX1 U867 ( .D0(r_wdat[1]), .D1(prx_wdat[1]), .S(prx_psh), .Y(n60) );
  MUX2IX1 U868 ( .D0(r_wdat[2]), .D1(prx_wdat[2]), .S(prx_psh), .Y(n57) );
  AND2X1 U869 ( .A(n500), .B(n499), .Y(obsd) );
  INVX1 U870 ( .A(srstz), .Y(n499) );
  INVX1 U871 ( .A(i_ccidle), .Y(n555) );
  MUX2IXL U872 ( .D0(r_wdat[6]), .D1(prx_wdat[6]), .S(prx_psh), .Y(n75) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phycrc_a0 ( crc32_3_0, rx_good, i_shfidat, i_start, i_shfi4, i_shfo4, 
        clk, test_si, test_so, test_se );
  output [3:0] crc32_3_0;
  input [3:0] i_shfidat;
  input i_start, i_shfi4, i_shfo4, clk, test_si, test_se;
  output rx_good, test_so;
  wire   crc32_r_30_, crc32_r_29_, crc32_r_28_, crc32_r_27_, crc32_r_26_,
         crc32_r_25_, crc32_r_24_, crc32_r_23_, crc32_r_22_, crc32_r_21_,
         crc32_r_20_, crc32_r_19_, crc32_r_18_, crc32_r_17_, crc32_r_16_,
         crc32_r_15_, crc32_r_14_, crc32_r_13_, crc32_r_12_, crc32_r_11_,
         crc32_r_10_, crc32_r_9_, crc32_r_8_, crc32_r_7_, crc32_r_6_,
         crc32_r_5_, crc32_r_4_, crc32_r_3_, crc32_r_2_, crc32_r_1_,
         crc32_r_0_, N188, N189, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, net10640, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n58, n121, n122, n123, n124, n127, n128, n129;

  SNPS_CLOCK_GATE_HIGH_phycrc_a0 clk_gate_crc32_r_reg ( .CLK(clk), .EN(N188), 
        .ENCLK(net10640), .TE(test_se) );
  SDFFQX1 crc32_r_reg_26_ ( .D(N215), .SIN(crc32_r_25_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_26_) );
  SDFFQX1 crc32_r_reg_16_ ( .D(N205), .SIN(crc32_r_15_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_16_) );
  SDFFQX1 crc32_r_reg_4_ ( .D(N193), .SIN(crc32_r_3_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_4_) );
  SDFFQX1 crc32_r_reg_25_ ( .D(N214), .SIN(crc32_r_24_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_25_) );
  SDFFQX1 crc32_r_reg_24_ ( .D(N213), .SIN(crc32_r_23_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_24_) );
  SDFFQX1 crc32_r_reg_27_ ( .D(N216), .SIN(crc32_r_26_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_27_) );
  SDFFQX1 crc32_r_reg_17_ ( .D(N206), .SIN(crc32_r_16_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_17_) );
  SDFFQX1 crc32_r_reg_8_ ( .D(N197), .SIN(crc32_r_7_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_8_) );
  SDFFQX1 crc32_r_reg_5_ ( .D(N194), .SIN(crc32_r_4_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_5_) );
  SDFFQX1 crc32_r_reg_0_ ( .D(N189), .SIN(test_si), .SMC(test_se), .C(net10640), .Q(crc32_r_0_) );
  SDFFQX1 crc32_r_reg_1_ ( .D(N190), .SIN(crc32_r_0_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_1_) );
  SDFFQX1 crc32_r_reg_10_ ( .D(N199), .SIN(crc32_r_9_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_10_) );
  SDFFQX1 crc32_r_reg_6_ ( .D(N195), .SIN(crc32_r_5_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_6_) );
  SDFFQX1 crc32_r_reg_11_ ( .D(N200), .SIN(crc32_r_10_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_11_) );
  SDFFQX1 crc32_r_reg_15_ ( .D(N204), .SIN(crc32_r_14_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_15_) );
  SDFFQX1 crc32_r_reg_12_ ( .D(N201), .SIN(crc32_r_11_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_12_) );
  SDFFQX1 crc32_r_reg_14_ ( .D(N203), .SIN(crc32_r_13_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_14_) );
  SDFFQX1 crc32_r_reg_18_ ( .D(N207), .SIN(crc32_r_17_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_18_) );
  SDFFQX1 crc32_r_reg_3_ ( .D(N192), .SIN(crc32_r_2_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_3_) );
  SDFFQX1 crc32_r_reg_20_ ( .D(N209), .SIN(crc32_r_19_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_20_) );
  SDFFQX1 crc32_r_reg_9_ ( .D(N198), .SIN(crc32_r_8_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_9_) );
  SDFFQX1 crc32_r_reg_21_ ( .D(N210), .SIN(crc32_r_20_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_21_) );
  SDFFQX1 crc32_r_reg_7_ ( .D(N196), .SIN(crc32_r_6_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_7_) );
  SDFFQX1 crc32_r_reg_22_ ( .D(N211), .SIN(crc32_r_21_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_22_) );
  SDFFQX1 crc32_r_reg_2_ ( .D(N191), .SIN(crc32_r_1_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_2_) );
  SDFFQX1 crc32_r_reg_13_ ( .D(N202), .SIN(crc32_r_12_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_13_) );
  SDFFQX1 crc32_r_reg_23_ ( .D(N212), .SIN(crc32_r_22_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_23_) );
  SDFFQX1 crc32_r_reg_28_ ( .D(N217), .SIN(crc32_r_27_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_28_) );
  SDFFQX1 crc32_r_reg_29_ ( .D(N218), .SIN(crc32_r_28_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_29_) );
  SDFFQX1 crc32_r_reg_19_ ( .D(N208), .SIN(crc32_r_18_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_19_) );
  SDFFQX1 crc32_r_reg_31_ ( .D(N220), .SIN(crc32_r_30_), .SMC(test_se), .C(
        net10640), .Q(test_so) );
  SDFFQX1 crc32_r_reg_30_ ( .D(N219), .SIN(crc32_r_29_), .SMC(test_se), .C(
        net10640), .Q(crc32_r_30_) );
  INVX1 U3 ( .A(n18), .Y(n1) );
  XNOR2XL U4 ( .A(i_shfidat[2]), .B(n119), .Y(n56) );
  INVX1 U5 ( .A(n17), .Y(n2) );
  XNOR2XL U6 ( .A(i_shfidat[3]), .B(n120), .Y(n71) );
  INVX1 U7 ( .A(n19), .Y(n3) );
  XNOR2XL U8 ( .A(i_shfidat[1]), .B(n117), .Y(n51) );
  INVX1 U9 ( .A(n16), .Y(n4) );
  XNOR2XL U10 ( .A(i_shfidat[0]), .B(n114), .Y(n62) );
  INVX1 U11 ( .A(n62), .Y(n5) );
  INVX1 U12 ( .A(n62), .Y(n6) );
  AND2X1 U13 ( .A(i_shfo4), .B(n12), .Y(n60) );
  INVX1 U14 ( .A(n60), .Y(n7) );
  INVX1 U15 ( .A(n60), .Y(n8) );
  INVX1 U16 ( .A(n78), .Y(n9) );
  INVX1 U17 ( .A(n78), .Y(n10) );
  INVX1 U18 ( .A(n11), .Y(n12) );
  NAND2X1 U19 ( .A(n12), .B(n7), .Y(N188) );
  INVX1 U20 ( .A(n11), .Y(n14) );
  INVX1 U21 ( .A(n78), .Y(n15) );
  INVX1 U22 ( .A(n11), .Y(n13) );
  NAND21X1 U23 ( .B(n81), .A(n80), .Y(n63) );
  NAND2X1 U24 ( .A(i_start), .B(n19), .Y(n49) );
  OAI21X1 U25 ( .B(n14), .C(n115), .A(n9), .Y(N191) );
  XNOR2XL U26 ( .A(n17), .B(n116), .Y(n115) );
  XNOR2XL U27 ( .A(n18), .B(n19), .Y(n116) );
  INVX1 U28 ( .A(i_start), .Y(n16) );
  OR2X1 U29 ( .A(i_start), .B(i_shfi4), .Y(n11) );
  NAND21X1 U30 ( .B(n12), .A(n81), .Y(n46) );
  OAI21X1 U31 ( .B(n14), .C(n118), .A(n10), .Y(N190) );
  XNOR2XL U32 ( .A(n17), .B(n18), .Y(n118) );
  AOI21X1 U33 ( .B(n18), .C(n4), .A(n78), .Y(n55) );
  AOI21X1 U34 ( .B(n17), .C(n4), .A(n78), .Y(n74) );
  NOR2X1 U35 ( .A(i_shfi4), .B(n12), .Y(n78) );
  AND2X1 U36 ( .A(n80), .B(n15), .Y(n48) );
  NOR2X1 U37 ( .A(n12), .B(n4), .Y(n52) );
  OAI21X1 U38 ( .B(n14), .C(n17), .A(n15), .Y(N189) );
  INVX1 U39 ( .A(n51), .Y(n19) );
  AOI21AX1 U40 ( .B(n16), .C(n51), .A(n49), .Y(n68) );
  NOR2X1 U41 ( .A(n5), .B(i_start), .Y(n81) );
  NAND2X1 U42 ( .A(i_start), .B(n5), .Y(n80) );
  OAI21X1 U43 ( .B(n14), .C(n112), .A(n9), .Y(N192) );
  XNOR2XL U44 ( .A(n18), .B(n113), .Y(n112) );
  XNOR2XL U45 ( .A(n19), .B(n6), .Y(n113) );
  INVX1 U46 ( .A(n56), .Y(n18) );
  INVX1 U47 ( .A(n71), .Y(n17) );
  OAI21BX1 U48 ( .C(n7), .B(n6), .A(N188), .Y(n47) );
  OAI21X1 U49 ( .B(n14), .C(n3), .A(n7), .Y(n53) );
  OAI21X1 U50 ( .B(n14), .C(n56), .A(n7), .Y(n57) );
  OAI21X1 U51 ( .B(n14), .C(n71), .A(n7), .Y(n75) );
  NOR4XL U52 ( .A(n22), .B(n27), .C(n20), .D(n30), .Y(n41) );
  NOR4XL U53 ( .A(n31), .B(n21), .C(n32), .D(n26), .Y(n40) );
  NOR4XL U54 ( .A(n23), .B(n25), .C(n29), .D(n24), .Y(n38) );
  NOR2X1 U55 ( .A(crc32_r_30_), .B(i_start), .Y(n117) );
  NOR2X1 U56 ( .A(test_so), .B(i_start), .Y(n114) );
  OAI221X1 U57 ( .A(n13), .B(n106), .C(n26), .D(n7), .E(n9), .Y(N194) );
  XNOR2XL U58 ( .A(n107), .B(n71), .Y(n106) );
  XNOR2XL U59 ( .A(n56), .B(n108), .Y(n107) );
  OAI22X1 U60 ( .A(n26), .B(n6), .C(crc32_r_1_), .D(n63), .Y(n108) );
  OAI221X1 U61 ( .A(n13), .B(n98), .C(n23), .D(n7), .E(n10), .Y(N197) );
  XNOR2XL U62 ( .A(n99), .B(n71), .Y(n98) );
  XNOR2XL U63 ( .A(n56), .B(n100), .Y(n99) );
  OAI22X1 U64 ( .A(n23), .B(n6), .C(crc32_r_4_), .D(n63), .Y(n100) );
  OAI221X1 U65 ( .A(n13), .B(n90), .C(n8), .D(n122), .E(n15), .Y(N200) );
  XNOR2XL U66 ( .A(n91), .B(n71), .Y(n90) );
  XNOR2XL U67 ( .A(n56), .B(n92), .Y(n91) );
  OAI22X1 U68 ( .A(n6), .B(n122), .C(crc32_r_7_), .D(n63), .Y(n92) );
  OAI221X1 U69 ( .A(n12), .B(n84), .C(n8), .D(n35), .E(n9), .Y(N202) );
  XNOR2XL U70 ( .A(n85), .B(n56), .Y(n84) );
  XNOR2XL U71 ( .A(n51), .B(n86), .Y(n85) );
  OAI22X1 U72 ( .A(n6), .B(n35), .C(crc32_r_9_), .D(n63), .Y(n86) );
  OAI221X1 U73 ( .A(n13), .B(n101), .C(n28), .D(n7), .E(n10), .Y(N196) );
  XNOR2XL U74 ( .A(n102), .B(n71), .Y(n101) );
  XNOR2XL U75 ( .A(n51), .B(n103), .Y(n102) );
  OAI22X1 U76 ( .A(n28), .B(n5), .C(crc32_r_3_), .D(n63), .Y(n103) );
  OAI221X1 U77 ( .A(n13), .B(n93), .C(n29), .D(n7), .E(n15), .Y(N199) );
  XNOR2XL U78 ( .A(n94), .B(n71), .Y(n93) );
  XNOR2XL U79 ( .A(n51), .B(n95), .Y(n94) );
  OAI22X1 U80 ( .A(n29), .B(n5), .C(crc32_r_6_), .D(n63), .Y(n95) );
  OAI221X1 U81 ( .A(n13), .B(n109), .C(n22), .D(n7), .E(n9), .Y(N193) );
  XNOR2XL U82 ( .A(n110), .B(n71), .Y(n109) );
  XNOR2XL U83 ( .A(n51), .B(n111), .Y(n110) );
  OAI22X1 U84 ( .A(n22), .B(n6), .C(crc32_r_0_), .D(n63), .Y(n111) );
  OAI221X1 U85 ( .A(n12), .B(n64), .C(n8), .D(n58), .E(n10), .Y(N214) );
  XNOR2XL U86 ( .A(n19), .B(n65), .Y(n64) );
  OAI22X1 U87 ( .A(n6), .B(n58), .C(crc32_r_21_), .D(n63), .Y(n65) );
  INVX1 U88 ( .A(crc32_r_21_), .Y(n58) );
  OAI221X1 U89 ( .A(n13), .B(n59), .C(n127), .D(n8), .E(n15), .Y(N215) );
  XNOR2XL U90 ( .A(n17), .B(n61), .Y(n59) );
  OAI22X1 U91 ( .A(n6), .B(n127), .C(crc32_r_22_), .D(n63), .Y(n61) );
  INVX1 U92 ( .A(crc32_r_22_), .Y(n127) );
  OAI221X1 U93 ( .A(n12), .B(n82), .C(n27), .D(n8), .E(n9), .Y(N203) );
  XNOR2XL U94 ( .A(n19), .B(n83), .Y(n82) );
  OAI22X1 U95 ( .A(n27), .B(n6), .C(crc32_r_10_), .D(n63), .Y(n83) );
  OAI221X1 U96 ( .A(n13), .B(n96), .C(n25), .D(n8), .E(n10), .Y(N198) );
  XNOR2XL U97 ( .A(n97), .B(n56), .Y(n96) );
  AOI22X1 U98 ( .A(n68), .B(n25), .C(n51), .D(crc32_r_5_), .Y(n97) );
  OAI221X1 U99 ( .A(n13), .B(n87), .C(n24), .D(n8), .E(n15), .Y(N201) );
  XNOR2XL U100 ( .A(n88), .B(n71), .Y(n87) );
  XNOR2XL U101 ( .A(n89), .B(n18), .Y(n88) );
  AOI22X1 U102 ( .A(n68), .B(n24), .C(n51), .D(crc32_r_8_), .Y(n89) );
  OAI221X1 U103 ( .A(n12), .B(n66), .C(n8), .D(n121), .E(n9), .Y(N213) );
  XNOR2XL U104 ( .A(n67), .B(n56), .Y(n66) );
  AOI22X1 U105 ( .A(n68), .B(n121), .C(crc32_r_20_), .D(n51), .Y(n67) );
  INVX1 U106 ( .A(crc32_r_20_), .Y(n121) );
  OAI221X1 U107 ( .A(n13), .B(n104), .C(n8), .D(n128), .E(n10), .Y(N195) );
  XNOR2XL U108 ( .A(n105), .B(n56), .Y(n104) );
  AOI22X1 U109 ( .A(n68), .B(n128), .C(crc32_r_2_), .D(n51), .Y(n105) );
  INVX1 U110 ( .A(crc32_r_2_), .Y(n128) );
  NOR2X1 U111 ( .A(crc32_r_29_), .B(i_start), .Y(n119) );
  NAND2X1 U112 ( .A(n73), .B(n74), .Y(N211) );
  AOI32X1 U113 ( .A(n52), .B(n32), .C(n2), .D(crc32_r_18_), .E(n75), .Y(n73)
         );
  NAND2X1 U114 ( .A(n77), .B(n55), .Y(N206) );
  AOI32X1 U115 ( .A(n52), .B(n123), .C(n1), .D(crc32_r_13_), .E(n57), .Y(n77)
         );
  INVX1 U116 ( .A(crc32_r_13_), .Y(n123) );
  NAND2X1 U117 ( .A(n54), .B(n55), .Y(N216) );
  AOI32X1 U118 ( .A(n52), .B(n129), .C(n1), .D(crc32_r_23_), .E(n57), .Y(n54)
         );
  INVX1 U119 ( .A(crc32_r_23_), .Y(n129) );
  NAND2X1 U120 ( .A(n79), .B(n74), .Y(N205) );
  AOI32X1 U121 ( .A(n52), .B(n30), .C(n2), .D(crc32_r_12_), .E(n75), .Y(n79)
         );
  OAI221X1 U122 ( .A(crc32_r_25_), .B(n46), .C(n33), .D(n47), .E(n48), .Y(N218) );
  INVX1 U123 ( .A(crc32_r_25_), .Y(n33) );
  OAI221X1 U124 ( .A(crc32_r_15_), .B(n46), .C(n21), .D(n47), .E(n48), .Y(N208) );
  OAI221X1 U125 ( .A(crc32_r_11_), .B(n46), .C(n20), .D(n47), .E(n48), .Y(N204) );
  OAI221X1 U126 ( .A(n12), .B(n69), .C(n8), .D(n124), .E(n15), .Y(N212) );
  INVX1 U127 ( .A(crc32_r_19_), .Y(n124) );
  XNOR2XL U128 ( .A(n70), .B(n71), .Y(n69) );
  XNOR2XL U129 ( .A(n72), .B(n56), .Y(n70) );
  NOR2X1 U130 ( .A(crc32_r_28_), .B(i_start), .Y(n120) );
  NAND3X1 U131 ( .A(n49), .B(n10), .C(n50), .Y(N217) );
  AOI32X1 U132 ( .A(n3), .B(n34), .C(n52), .D(crc32_r_24_), .E(n53), .Y(n50)
         );
  INVX1 U133 ( .A(crc32_r_24_), .Y(n34) );
  NAND3X1 U134 ( .A(n49), .B(n15), .C(n76), .Y(N207) );
  AOI32X1 U135 ( .A(n3), .B(n31), .C(n52), .D(crc32_r_14_), .E(n53), .Y(n76)
         );
  OAI21BBX1 U136 ( .A(N188), .B(crc32_r_26_), .C(n16), .Y(N219) );
  OAI21BBX1 U137 ( .A(N188), .B(crc32_r_27_), .C(n16), .Y(N220) );
  OAI21BBX1 U138 ( .A(N188), .B(crc32_r_16_), .C(n16), .Y(N209) );
  OAI21BBX1 U139 ( .A(N188), .B(crc32_r_17_), .C(n16), .Y(N210) );
  NOR2X1 U140 ( .A(crc32_r_19_), .B(i_start), .Y(n72) );
  INVX1 U141 ( .A(crc32_r_28_), .Y(crc32_3_0[3]) );
  INVX1 U142 ( .A(crc32_r_29_), .Y(crc32_3_0[2]) );
  AND4X1 U143 ( .A(crc32_r_24_), .B(crc32_r_25_), .C(crc32_r_26_), .D(
        crc32_r_3_), .Y(n39) );
  NOR2X1 U144 ( .A(n36), .B(n37), .Y(rx_good) );
  NAND4X1 U145 ( .A(n42), .B(n43), .C(n44), .D(n45), .Y(n36) );
  NAND4X1 U146 ( .A(n38), .B(n39), .C(n40), .D(n41), .Y(n37) );
  NOR4XL U147 ( .A(crc32_r_21_), .B(crc32_r_20_), .C(crc32_r_19_), .D(
        crc32_r_17_), .Y(n43) );
  NOR4XL U148 ( .A(crc32_r_9_), .B(crc32_r_7_), .C(crc32_r_2_), .D(crc32_r_29_), .Y(n45) );
  NOR4XL U149 ( .A(crc32_r_28_), .B(crc32_r_27_), .C(crc32_r_23_), .D(
        crc32_r_22_), .Y(n44) );
  NOR4XL U150 ( .A(crc32_r_16_), .B(crc32_r_13_), .C(crc32_3_0[1]), .D(
        crc32_3_0[0]), .Y(n42) );
  INVX1 U151 ( .A(crc32_r_30_), .Y(crc32_3_0[1]) );
  INVX1 U152 ( .A(test_so), .Y(crc32_3_0[0]) );
  INVX1 U153 ( .A(crc32_r_6_), .Y(n29) );
  INVX1 U154 ( .A(crc32_r_1_), .Y(n26) );
  INVX1 U155 ( .A(crc32_r_10_), .Y(n27) );
  INVX1 U156 ( .A(crc32_r_0_), .Y(n22) );
  INVX1 U157 ( .A(crc32_r_8_), .Y(n24) );
  INVX1 U158 ( .A(crc32_r_5_), .Y(n25) );
  INVX1 U159 ( .A(crc32_r_18_), .Y(n32) );
  INVX1 U160 ( .A(crc32_r_12_), .Y(n30) );
  INVX1 U161 ( .A(crc32_r_14_), .Y(n31) );
  INVX1 U162 ( .A(crc32_r_11_), .Y(n20) );
  INVX1 U163 ( .A(crc32_r_15_), .Y(n21) );
  INVX1 U164 ( .A(crc32_r_4_), .Y(n23) );
  INVX1 U165 ( .A(crc32_r_7_), .Y(n122) );
  INVX1 U166 ( .A(crc32_r_9_), .Y(n35) );
  INVX1 U167 ( .A(crc32_r_3_), .Y(n28) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phycrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phytx_a0 ( r_txnumk, r_txendk, r_txshrt, r_txauto, prx_cccnt, ptx_txact, 
        ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, i_rdat, i_txreq, i_one, 
        ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4, ptx_crcsidat, ptx_fsm, 
        pcc_crc30, clk, srstz, test_si, test_se );
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [1:0] prx_cccnt;
  input [7:0] i_rdat;
  output [3:0] ptx_crcsidat;
  output [2:0] ptx_fsm;
  input [3:0] pcc_crc30;
  input r_txendk, r_txshrt, i_txreq, i_one, clk, srstz, test_si, test_se;
  output ptx_txact, ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, ptx_crcstart,
         ptx_crcshfi4, ptx_crcshfo4;
  wire   hinib, N251, N254, N255, N268, N270, N271, N272, N273, N297, N298,
         N299, net10662, net10668, n237, n238, n122, n133, n134, n135, n152,
         n154, n155, n156, n170, n189, n190, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n153, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272;
  wire   [4:0] bytcnt;
  wire   [3:0] bitcnt;

  SNPS_CLOCK_GATE_HIGH_phytx_a0_0 clk_gate_bitcnt_reg ( .CLK(clk), .EN(N251), 
        .ENCLK(net10662), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phytx_a0_1 clk_gate_bytcnt_reg ( .CLK(clk), .EN(N268), 
        .ENCLK(net10668), .TE(test_se) );
  SDFFQX1 ptx_cc_reg ( .D(n238), .SIN(n4), .SMC(test_se), .C(clk), .Q(ptx_cc)
         );
  SDFFQX1 bitcnt_reg_3_ ( .D(N255), .SIN(bitcnt[2]), .SMC(test_se), .C(
        net10662), .Q(bitcnt[3]) );
  SDFFQX1 bitcnt_reg_1_ ( .D(n266), .SIN(bitcnt[0]), .SMC(test_se), .C(
        net10662), .Q(bitcnt[1]) );
  SDFFQX1 bitcnt_reg_2_ ( .D(N254), .SIN(bitcnt[1]), .SMC(test_se), .C(
        net10662), .Q(bitcnt[2]) );
  SDFFQX1 bitcnt_reg_0_ ( .D(n263), .SIN(test_si), .SMC(test_se), .C(net10662), 
        .Q(bitcnt[0]) );
  SDFFQX1 cs_txph_reg_0_ ( .D(N297), .SIN(bytcnt[4]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[0]) );
  SDFFQX1 cs_txph_reg_2_ ( .D(N299), .SIN(ptx_fsm[1]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[2]) );
  SDFFQX1 bytcnt_reg_3_ ( .D(N272), .SIN(bytcnt[2]), .SMC(test_se), .C(
        net10668), .Q(bytcnt[3]) );
  SDFFQX1 bytcnt_reg_4_ ( .D(N273), .SIN(bytcnt[3]), .SMC(test_se), .C(
        net10668), .Q(bytcnt[4]) );
  SDFFQX1 bytcnt_reg_1_ ( .D(N270), .SIN(bytcnt[0]), .SMC(test_se), .C(
        net10668), .Q(bytcnt[1]) );
  SDFFQX1 cs_txph_reg_1_ ( .D(N298), .SIN(ptx_fsm[0]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[1]) );
  SDFFQX1 hinib_reg ( .D(n237), .SIN(ptx_fsm[2]), .SMC(test_se), .C(net10662), 
        .Q(hinib) );
  SDFFQX1 bytcnt_reg_2_ ( .D(N271), .SIN(bytcnt[1]), .SMC(test_se), .C(
        net10668), .Q(bytcnt[2]) );
  SDFFQX1 bytcnt_reg_0_ ( .D(n264), .SIN(bitcnt[3]), .SMC(test_se), .C(
        net10668), .Q(bytcnt[0]) );
  BUFX1 U3 ( .A(n163), .Y(n1) );
  BUFXL U4 ( .A(n163), .Y(n2) );
  INVX1 U5 ( .A(r_txnumk[0]), .Y(n14) );
  NAND5XL U6 ( .A(bytcnt[0]), .B(n245), .C(n39), .D(n98), .E(n86), .Y(n49) );
  NAND21X1 U7 ( .B(n5), .A(n262), .Y(ptx_fifopop) );
  MUX2X1 U8 ( .D0(n25), .D1(n126), .S(ptx_crcsidat[3]), .Y(n27) );
  NAND31X1 U9 ( .C(n225), .A(bitcnt[3]), .B(n112), .Y(n102) );
  AND3X1 U10 ( .A(n271), .B(n269), .C(r_txauto[0]), .Y(n3) );
  INVX1 U11 ( .A(n149), .Y(n4) );
  MUX2X1 U12 ( .D0(n53), .D1(n24), .S(hinib), .Y(n126) );
  MUX2X1 U13 ( .D0(n51), .D1(n23), .S(hinib), .Y(n130) );
  MUX2BXL U14 ( .D0(n144), .D1(i_rdat[7]), .S(hinib), .Y(n164) );
  NOR2X1 U15 ( .A(n101), .B(n258), .Y(n5) );
  AND3XL U16 ( .A(n248), .B(n250), .C(n247), .Y(ptx_crcshfi4) );
  OAI22XL U17 ( .A(n145), .B(n144), .C(n212), .D(n177), .Y(n171) );
  INVX1 U18 ( .A(ptx_fsm[2]), .Y(n59) );
  INVX1 U19 ( .A(bytcnt[3]), .Y(n98) );
  INVX1 U20 ( .A(ptx_fsm[1]), .Y(n124) );
  GEN2X1 U21 ( .D(n27), .E(n123), .C(n115), .B(n207), .A(n166), .Y(n163) );
  OAI31XL U22 ( .A(n30), .B(n250), .C(n253), .D(n38), .Y(n57) );
  AOI31XL U23 ( .A(n26), .B(n23), .C(n52), .D(n115), .Y(n30) );
  OAI221XL U24 ( .A(n5), .B(n87), .C(n86), .D(n95), .E(n265), .Y(n170) );
  AOI31XL U25 ( .A(n158), .B(n68), .C(n71), .D(n38), .Y(n87) );
  AOI32XL U26 ( .A(n267), .B(i_txreq), .C(n75), .D(n166), .E(n62), .Y(n66) );
  INVXL U27 ( .A(n262), .Y(n64) );
  AO21XL U28 ( .B(n46), .C(n166), .A(n61), .Y(n69) );
  AOI211XL U29 ( .C(i_rdat[0]), .D(n222), .A(n142), .B(n141), .Y(n173) );
  AND2XL U30 ( .A(i_rdat[6]), .B(n194), .Y(n196) );
  NAND32XL U31 ( .B(n130), .C(n115), .A(n125), .Y(n165) );
  AO21XL U32 ( .B(i_rdat[4]), .C(n222), .A(n204), .Y(n215) );
  INVXL U33 ( .A(n103), .Y(n104) );
  XOR2X1 U34 ( .A(n1), .B(bitcnt[1]), .Y(n29) );
  GEN2X1 U35 ( .D(bytcnt[4]), .E(n22), .C(n21), .B(n20), .A(n258), .Y(n250) );
  INVXL U36 ( .A(r_txnumk[4]), .Y(n21) );
  AOI32XL U37 ( .A(n252), .B(n16), .C(n249), .D(r_txnumk[2]), .E(n39), .Y(n17)
         );
  NAND21X1 U38 ( .B(r_txnumk[1]), .A(bytcnt[1]), .Y(n249) );
  NAND21XL U39 ( .B(r_txnumk[2]), .A(bytcnt[2]), .Y(n252) );
  OR2XL U40 ( .A(ptx_fsm[2]), .B(n188), .Y(ptx_txact) );
  INVXL U41 ( .A(ptx_fsm[0]), .Y(n37) );
  NAND21XL U42 ( .B(ptx_fsm[1]), .A(n37), .Y(n188) );
  NAND32XL U43 ( .B(ptx_fsm[1]), .C(n37), .A(n59), .Y(n68) );
  XOR2XL U44 ( .A(ptx_fsm[0]), .B(n261), .Y(n82) );
  NOR2XL U45 ( .A(n68), .B(n268), .Y(n81) );
  AND2XL U46 ( .A(n69), .B(ptx_fsm[0]), .Y(n80) );
  NAND21XL U47 ( .B(bytcnt[0]), .A(n96), .Y(n90) );
  MUX2IXL U48 ( .D0(n91), .D1(bytcnt[1]), .S(bytcnt[2]), .Y(n92) );
  OA21XL U49 ( .B(bytcnt[4]), .C(n97), .A(n96), .Y(N273) );
  MUX2XL U50 ( .D0(n109), .D1(n4), .S(n108), .Y(n237) );
  AOI211XL U51 ( .C(n10), .D(n107), .A(i_txreq), .B(n106), .Y(n108) );
  INVXL U52 ( .A(n102), .Y(n107) );
  INVXL U53 ( .A(n123), .Y(ptx_crcsidat[1]) );
  INVXL U54 ( .A(n130), .Y(ptx_crcsidat[0]) );
  OAI21BBXL U55 ( .A(r_txshrt), .B(n245), .C(n72), .Y(n62) );
  OAI21BBX1 U56 ( .A(n224), .B(n149), .C(n6), .Y(n213) );
  MUX2IXL U57 ( .D0(n113), .D1(n121), .S(n112), .Y(n6) );
  NAND21XL U58 ( .B(n110), .A(n4), .Y(n111) );
  AND2XL U59 ( .A(n135), .B(hinib), .Y(n148) );
  MUX2XL U60 ( .D0(ptx_crcsidat[3]), .D1(pcc_crc30[3]), .S(n246), .Y(n201) );
  OAI211XL U61 ( .C(hinib), .D(bytcnt[0]), .A(n156), .B(n157), .Y(n137) );
  INVXL U62 ( .A(bytcnt[0]), .Y(n251) );
  INVXL U63 ( .A(hinib), .Y(n149) );
  NAND21XL U64 ( .B(n251), .A(hinib), .Y(n157) );
  INVXL U65 ( .A(bytcnt[1]), .Y(n89) );
  NAND21XL U66 ( .B(n89), .A(bytcnt[0]), .Y(n91) );
  NAND21XL U67 ( .B(n91), .A(bytcnt[2]), .Y(n99) );
  INVX1 U68 ( .A(n32), .Y(n244) );
  NAND21X1 U69 ( .B(n233), .A(n243), .Y(n32) );
  NAND21X1 U70 ( .B(n244), .A(n243), .Y(N251) );
  INVX1 U71 ( .A(n129), .Y(n146) );
  INVX1 U72 ( .A(n177), .Y(n180) );
  INVX1 U73 ( .A(n210), .Y(n183) );
  INVX1 U74 ( .A(n189), .Y(n268) );
  INVX1 U75 ( .A(n133), .Y(n116) );
  INVX1 U76 ( .A(srstz), .Y(n11) );
  INVX1 U77 ( .A(n38), .Y(n245) );
  INVX1 U78 ( .A(n57), .Y(n101) );
  NAND21X1 U79 ( .B(n75), .A(prx_cccnt[0]), .Y(n233) );
  INVX1 U80 ( .A(n170), .Y(n96) );
  INVX1 U81 ( .A(n31), .Y(n243) );
  NAND32X1 U82 ( .B(i_txreq), .C(n57), .A(n55), .Y(n31) );
  AND2X1 U83 ( .A(srstz), .B(n259), .Y(N298) );
  INVX1 U84 ( .A(i_txreq), .Y(n234) );
  AND2X1 U85 ( .A(n246), .B(n247), .Y(ptx_crcshfo4) );
  INVX1 U86 ( .A(n56), .Y(n77) );
  NAND21X1 U87 ( .B(n64), .A(n55), .Y(n56) );
  NAND21X1 U88 ( .B(n127), .A(n176), .Y(n129) );
  NAND21X1 U89 ( .B(n207), .A(n200), .Y(n210) );
  NAND21X1 U90 ( .B(n129), .A(n211), .Y(n177) );
  INVX1 U91 ( .A(n114), .Y(n125) );
  INVX1 U92 ( .A(n127), .Y(n200) );
  MUX2AXL U93 ( .D0(n7), .D1(n8), .S(n178), .Y(n141) );
  NAND2X1 U94 ( .A(n203), .B(n146), .Y(n7) );
  NAND2X1 U95 ( .A(n177), .B(n210), .Y(n8) );
  NAND21X1 U96 ( .B(n245), .A(n253), .Y(n247) );
  INVX1 U97 ( .A(n253), .Y(n100) );
  INVX1 U98 ( .A(n165), .Y(n219) );
  AND2X1 U99 ( .A(n178), .B(n208), .Y(n179) );
  INVX1 U100 ( .A(n128), .Y(n208) );
  NAND21X1 U101 ( .B(n211), .A(n146), .Y(n128) );
  INVX1 U102 ( .A(n168), .Y(n185) );
  NAND21X1 U103 ( .B(n217), .A(n216), .Y(n168) );
  INVX1 U104 ( .A(n167), .Y(n216) );
  INVX1 U105 ( .A(n145), .Y(n222) );
  AND2X1 U106 ( .A(srstz), .B(n257), .Y(N299) );
  NOR3XL U107 ( .A(n269), .B(n271), .C(n272), .Y(n135) );
  INVX1 U108 ( .A(n143), .Y(n212) );
  NAND21X1 U109 ( .B(n175), .A(n178), .Y(n143) );
  OAI21BBX1 U110 ( .A(n272), .B(n134), .C(n155), .Y(n154) );
  AND2X1 U111 ( .A(n178), .B(n176), .Y(n174) );
  INVX1 U112 ( .A(n155), .Y(n270) );
  INVX1 U113 ( .A(n71), .Y(n246) );
  NOR2X1 U114 ( .A(n135), .B(n156), .Y(n133) );
  NAND3X1 U115 ( .A(n133), .B(n155), .C(n190), .Y(n189) );
  NOR3XL U116 ( .A(n3), .B(n122), .C(n134), .Y(n190) );
  INVX1 U117 ( .A(n158), .Y(n197) );
  INVX1 U118 ( .A(n95), .Y(n97) );
  INVX1 U119 ( .A(n257), .Y(n260) );
  AND2X1 U120 ( .A(n130), .B(ptx_crcsidat[2]), .Y(n25) );
  NAND43X1 U121 ( .B(n29), .C(n103), .D(n233), .A(n105), .Y(n253) );
  NAND32X1 U122 ( .B(n233), .C(n102), .A(n10), .Y(n38) );
  INVX1 U123 ( .A(n250), .Y(n207) );
  INVX1 U124 ( .A(i_one), .Y(n58) );
  INVX1 U125 ( .A(n29), .Y(n112) );
  INVX1 U126 ( .A(i_rdat[6]), .Y(n24) );
  INVX1 U127 ( .A(n164), .Y(ptx_crcsidat[3]) );
  OAI22X1 U128 ( .A(r_txnumk[4]), .B(n86), .C(r_txnumk[3]), .D(n98), .Y(n254)
         );
  INVX1 U129 ( .A(i_rdat[4]), .Y(n23) );
  INVX1 U130 ( .A(i_rdat[0]), .Y(n51) );
  INVX1 U131 ( .A(i_rdat[2]), .Y(n53) );
  INVX1 U132 ( .A(n126), .Y(ptx_crcsidat[2]) );
  INVX1 U133 ( .A(r_txnumk[1]), .Y(n15) );
  INVX1 U134 ( .A(r_txnumk[2]), .Y(n13) );
  INVX1 U135 ( .A(i_rdat[5]), .Y(n26) );
  INVX1 U136 ( .A(i_rdat[1]), .Y(n54) );
  INVX1 U137 ( .A(r_txauto[6]), .Y(n115) );
  INVX1 U138 ( .A(n68), .Y(n166) );
  INVX1 U139 ( .A(n12), .Y(n52) );
  NAND21X1 U140 ( .B(i_rdat[7]), .A(n24), .Y(n12) );
  INVX1 U141 ( .A(ptx_txact), .Y(n75) );
  NAND32X1 U142 ( .B(n37), .C(n124), .A(n59), .Y(n158) );
  INVX1 U143 ( .A(n258), .Y(n248) );
  NOR21XL U144 ( .B(n77), .A(n76), .Y(n78) );
  NOR32XL U145 ( .B(n75), .C(i_txreq), .A(n74), .Y(n76) );
  NOR2X1 U146 ( .A(r_txauto[3]), .B(n189), .Y(n74) );
  OAI211X1 U147 ( .C(n67), .D(n124), .A(n66), .B(n65), .Y(n259) );
  AOI221XL U148 ( .A(n248), .B(n70), .C(n246), .D(n72), .E(n61), .Y(n67) );
  OA22X1 U149 ( .A(n64), .B(n158), .C(n70), .D(n63), .Y(n65) );
  INVX1 U150 ( .A(n240), .Y(n261) );
  AOI211X1 U151 ( .C(n99), .D(n98), .A(n170), .B(n97), .Y(N272) );
  AOI211X1 U152 ( .C(n251), .D(n89), .A(n170), .B(n88), .Y(N270) );
  INVX1 U153 ( .A(n91), .Y(n88) );
  INVX1 U154 ( .A(n90), .Y(n264) );
  AO21X1 U155 ( .B(n244), .C(n224), .A(n263), .Y(n241) );
  INVX1 U156 ( .A(n35), .Y(n242) );
  NAND32X1 U157 ( .B(n225), .C(n224), .A(n244), .Y(n35) );
  NAND2X1 U158 ( .A(n265), .B(n170), .Y(N268) );
  AND2X1 U159 ( .A(srstz), .B(n240), .Y(N297) );
  NOR5XL U160 ( .A(n256), .B(n255), .C(n258), .D(n254), .E(n253), .Y(
        ptx_crcstart) );
  INVX1 U161 ( .A(n252), .Y(n255) );
  NAND21X1 U162 ( .B(n89), .A(n43), .Y(n72) );
  OAI211X1 U163 ( .C(n60), .D(n59), .A(n77), .B(n70), .Y(n257) );
  AND2X1 U164 ( .A(n47), .B(n71), .Y(n60) );
  INVX1 U165 ( .A(n69), .Y(n47) );
  INVX1 U166 ( .A(n45), .Y(n61) );
  NAND43X1 U167 ( .B(n166), .C(n248), .D(n246), .A(n44), .Y(n45) );
  AOI31X1 U168 ( .A(n197), .B(n43), .C(n89), .D(ptx_goidle), .Y(n44) );
  INVX1 U169 ( .A(n62), .Y(n46) );
  INVX1 U170 ( .A(n49), .Y(n43) );
  OAI22X1 U171 ( .A(n159), .B(n158), .C(n210), .D(n162), .Y(n160) );
  AND2X1 U172 ( .A(n146), .B(n206), .Y(n161) );
  AOI211X1 U173 ( .C(n157), .D(n3), .A(n153), .B(n198), .Y(n159) );
  NAND21X1 U174 ( .B(n188), .A(n100), .Y(n55) );
  NAND32XL U175 ( .B(n58), .C(n258), .A(n57), .Y(n70) );
  NAND21X1 U176 ( .B(n231), .A(ptx_txact), .Y(n232) );
  MUX2X1 U177 ( .D0(n230), .D1(n229), .S(n228), .Y(n231) );
  XOR2X1 U178 ( .A(n227), .B(n226), .Y(n228) );
  GEN2XL U179 ( .D(n193), .E(n192), .C(n191), .B(n188), .A(n187), .Y(n230) );
  AOI211X1 U180 ( .C(n222), .D(n221), .A(n220), .B(n219), .Y(n229) );
  MUX2X1 U181 ( .D0(n196), .D1(n195), .S(n216), .Y(n221) );
  MUX2X1 U182 ( .D0(n218), .D1(n217), .S(n216), .Y(n220) );
  MUX2BXL U183 ( .D0(n173), .D1(n172), .S(n194), .Y(n191) );
  NAND32X1 U184 ( .B(n171), .C(n169), .A(n185), .Y(n172) );
  OA21X1 U185 ( .B(n215), .C(n214), .A(n213), .Y(n218) );
  OAI31XL U186 ( .A(n212), .B(n211), .C(n210), .D(n209), .Y(n214) );
  GEN2XL U187 ( .D(n203), .E(n202), .C(n201), .B(n200), .A(n199), .Y(n204) );
  AND4X1 U188 ( .A(n186), .B(n213), .C(n185), .D(n184), .Y(n187) );
  AOI221XL U189 ( .A(n183), .B(n182), .C(i_rdat[1]), .D(n222), .E(n181), .Y(
        n184) );
  OAI22X1 U190 ( .A(n176), .B(n211), .C(n175), .D(n174), .Y(n182) );
  MUX2X1 U191 ( .D0(n180), .D1(n179), .S(n203), .Y(n181) );
  OAI22X1 U192 ( .A(n72), .B(n71), .C(n70), .D(r_txauto[4]), .Y(n73) );
  AOI221XL U193 ( .A(n175), .B(n183), .C(i_rdat[2]), .D(n222), .E(n136), .Y(
        n192) );
  MUX2X1 U194 ( .D0(n132), .D1(n131), .S(n178), .Y(n136) );
  AND2X1 U195 ( .A(n208), .B(n250), .Y(n132) );
  OAI211X1 U196 ( .C(n139), .D(n158), .A(n138), .B(n167), .Y(n142) );
  AOI221XL U197 ( .A(n3), .B(n147), .C(n135), .D(n149), .E(n122), .Y(n139) );
  INVX1 U198 ( .A(n205), .Y(n138) );
  AOI31XL U199 ( .A(n208), .B(n207), .C(n206), .D(n205), .Y(n209) );
  AO21X1 U200 ( .B(n223), .C(n225), .A(n121), .Y(n167) );
  NAND21X1 U201 ( .B(r_txauto[6]), .A(n125), .Y(n145) );
  MUX2X1 U202 ( .D0(i_rdat[5]), .D1(i_rdat[7]), .S(n194), .Y(n195) );
  OR2XL U203 ( .A(n225), .B(n2), .Y(n110) );
  AND4X1 U204 ( .A(n194), .B(n165), .C(n186), .D(n167), .Y(n193) );
  INVX1 U205 ( .A(n213), .Y(n194) );
  INVX1 U206 ( .A(n140), .Y(n203) );
  NAND31X1 U207 ( .C(n166), .A(n9), .B(n165), .Y(n217) );
  NAND3XL U208 ( .A(r_txauto[6]), .B(n164), .C(n2), .Y(n9) );
  AND4X1 U209 ( .A(n105), .B(n112), .C(n104), .D(n188), .Y(n106) );
  INVX1 U210 ( .A(r_txauto[0]), .Y(n272) );
  AO21X1 U211 ( .B(n225), .C(n224), .A(n223), .Y(n226) );
  AO21X1 U212 ( .B(n134), .C(r_txauto[0]), .A(n156), .Y(n152) );
  OA21X1 U213 ( .B(n198), .C(n3), .A(n197), .Y(n199) );
  INVX1 U214 ( .A(n202), .Y(n178) );
  INVX1 U215 ( .A(r_txauto[1]), .Y(n271) );
  NAND3X1 U216 ( .A(r_txauto[2]), .B(n271), .C(r_txauto[0]), .Y(n155) );
  INVX1 U217 ( .A(n201), .Y(n176) );
  INVX1 U218 ( .A(r_txauto[2]), .Y(n269) );
  INVX1 U219 ( .A(n162), .Y(n211) );
  INVX1 U220 ( .A(n206), .Y(n175) );
  NOR3XL U221 ( .A(r_txauto[0]), .B(r_txauto[1]), .C(n269), .Y(n156) );
  NOR2X1 U222 ( .A(n271), .B(r_txauto[2]), .Y(n134) );
  NOR3XL U223 ( .A(n271), .B(r_txauto[0]), .C(n269), .Y(n122) );
  NAND32X1 U224 ( .B(n124), .C(n59), .A(n37), .Y(n71) );
  OAI22X1 U225 ( .A(n149), .B(n272), .C(n251), .D(r_txauto[0]), .Y(n117) );
  INVX1 U226 ( .A(n157), .Y(n147) );
  INVX1 U227 ( .A(r_txauto[4]), .Y(n63) );
  INVX1 U228 ( .A(r_txauto[3]), .Y(n267) );
  OR2X1 U229 ( .A(n98), .B(n99), .Y(n95) );
  AND4X1 U230 ( .A(n261), .B(n260), .C(n259), .D(n258), .Y(ptx_pspyld) );
  NAND43X1 U231 ( .B(n14), .C(n15), .D(n13), .A(r_txnumk[3]), .Y(n22) );
  OA21X1 U232 ( .B(n19), .C(n254), .A(n48), .Y(n20) );
  XNOR2XL U233 ( .A(n2), .B(bitcnt[2]), .Y(n10) );
  NAND21X1 U234 ( .B(n58), .A(r_txendk), .Y(n48) );
  NAND6XL U235 ( .A(n54), .B(n53), .C(n144), .D(n52), .E(n51), .F(n50), .Y(
        n262) );
  NOR6XL U236 ( .A(i_rdat[5]), .B(i_rdat[4]), .C(bytcnt[1]), .D(n49), .E(n158), 
        .F(n48), .Y(n50) );
  OA21X1 U237 ( .B(bytcnt[3]), .C(n18), .A(n17), .Y(n19) );
  INVX1 U238 ( .A(r_txnumk[3]), .Y(n18) );
  OAI22X1 U239 ( .A(bytcnt[1]), .B(n15), .C(bytcnt[0]), .D(n14), .Y(n16) );
  INVX1 U240 ( .A(i_rdat[3]), .Y(n144) );
  MUX2X1 U241 ( .D0(n54), .D1(n26), .S(hinib), .Y(n123) );
  NAND32X1 U242 ( .B(ptx_fsm[0]), .C(n124), .A(n59), .Y(n258) );
  INVX1 U243 ( .A(bytcnt[2]), .Y(n39) );
  INVX1 U244 ( .A(bytcnt[4]), .Y(n86) );
  INVX1 U245 ( .A(bitcnt[0]), .Y(n225) );
  INVX1 U246 ( .A(n28), .Y(n105) );
  NAND21X1 U247 ( .B(bitcnt[3]), .A(bitcnt[2]), .Y(n28) );
  NAND42X1 U248 ( .C(n81), .D(n80), .A(n79), .B(n78), .Y(n240) );
  NAND21X1 U249 ( .B(r_txauto[5]), .A(n73), .Y(n79) );
  NOR21XL U250 ( .B(n234), .A(n85), .Y(n265) );
  NAND31X1 U251 ( .C(n84), .A(n83), .B(n82), .Y(n85) );
  NOR21XL U252 ( .B(n257), .A(ptx_fsm[2]), .Y(n84) );
  XNOR2XL U253 ( .A(ptx_fsm[1]), .B(n259), .Y(n83) );
  NAND21X1 U254 ( .B(n94), .A(n93), .Y(N271) );
  NAND21X1 U255 ( .B(n170), .A(n92), .Y(n93) );
  NOR21XL U256 ( .B(bytcnt[2]), .A(n90), .Y(n94) );
  INVX1 U257 ( .A(n33), .Y(n263) );
  NAND21X1 U258 ( .B(bitcnt[0]), .A(n244), .Y(n33) );
  GEN2XL U259 ( .D(n244), .E(n227), .C(n241), .B(bitcnt[3]), .A(n36), .Y(N255)
         );
  AND2X1 U260 ( .A(n242), .B(n105), .Y(n36) );
  MUX2X1 U261 ( .D0(n242), .D1(n241), .S(bitcnt[2]), .Y(N254) );
  AND3XL U262 ( .A(n101), .B(n100), .C(n234), .Y(n109) );
  MUX2X1 U263 ( .D0(n239), .D1(ptx_cc), .S(n236), .Y(n238) );
  NAND21X1 U264 ( .B(n11), .A(ptx_cc), .Y(n239) );
  AND3X1 U265 ( .A(srstz), .B(n235), .C(n234), .Y(n236) );
  MUX2X1 U266 ( .D0(n233), .D1(n232), .S(prx_cccnt[1]), .Y(n235) );
  MUX2X1 U267 ( .D0(n34), .D1(n263), .S(bitcnt[1]), .Y(n266) );
  AND2X1 U268 ( .A(n244), .B(bitcnt[0]), .Y(n34) );
  GEN2XL U269 ( .D(n270), .E(hinib), .C(n153), .B(n197), .A(n219), .Y(n205) );
  INVX1 U270 ( .A(n111), .Y(n121) );
  AND2X1 U271 ( .A(n4), .B(n110), .Y(n113) );
  MUX2BXL U272 ( .D0(n123), .D1(pcc_crc30[1]), .S(n246), .Y(n206) );
  MUX2BXL U273 ( .D0(n126), .D1(pcc_crc30[2]), .S(n246), .Y(n162) );
  MUX2BXL U274 ( .D0(n130), .D1(pcc_crc30[0]), .S(n246), .Y(n202) );
  NAND21X1 U275 ( .B(n151), .A(n150), .Y(n198) );
  MUX2X1 U276 ( .D0(n148), .D1(n122), .S(n147), .Y(n151) );
  AOI22X1 U277 ( .A(n152), .B(n149), .C(n154), .D(n251), .Y(n150) );
  INVX1 U278 ( .A(n137), .Y(n153) );
  OAI21X1 U279 ( .B(n120), .C(n119), .A(n197), .Y(n186) );
  GEN2XL U280 ( .D(n270), .E(bytcnt[0]), .C(n135), .B(n149), .A(n118), .Y(n119) );
  MUX2X1 U281 ( .D0(n122), .D1(n116), .S(n147), .Y(n120) );
  AND2X1 U282 ( .A(n134), .B(n117), .Y(n118) );
  INVX1 U283 ( .A(n42), .Y(ptx_goidle) );
  NAND5XL U284 ( .A(ptx_fsm[2]), .B(ptx_fsm[0]), .C(n41), .D(n124), .E(n40), 
        .Y(n42) );
  INVX1 U285 ( .A(ptx_cc), .Y(n40) );
  INVX1 U286 ( .A(n233), .Y(n41) );
  INVX1 U287 ( .A(bitcnt[1]), .Y(n224) );
  INVX1 U288 ( .A(bitcnt[2]), .Y(n227) );
  GEN2XL U289 ( .D(n212), .E(n162), .C(n250), .B(n161), .A(n160), .Y(n169) );
  OAI22XL U290 ( .A(n206), .B(n129), .C(n250), .D(n177), .Y(n131) );
  NAND21XL U291 ( .B(n2), .A(hinib), .Y(n223) );
  NAND21XL U292 ( .B(n250), .A(n175), .Y(n140) );
  NAND32XL U293 ( .B(n124), .C(n2), .A(n158), .Y(n127) );
  NAND21XL U294 ( .B(n166), .A(n2), .Y(n114) );
  OAI211XL U295 ( .C(r_txnumk[0]), .D(n251), .A(n250), .B(n249), .Y(n256) );
  XOR2XL U296 ( .A(n2), .B(bitcnt[0]), .Y(n103) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyidd_a0 ( i_trans, i_goidle, o_ccidle, o_goidle, o_gobusy, clk, srstz, 
        test_si, test_so, test_se );
  input i_trans, i_goidle, clk, srstz, test_si, test_se;
  output o_ccidle, o_goidle, o_gobusy, test_so;
  wire   n30, ttranwin_6_, ttranwin_5_, ttranwin_4_, ttranwin_3_, ttranwin_2_,
         ttranwin_1_, ttranwin_0_, N11, N12, N13, N14, N15, N16, N17, N18, N46,
         N47, N48, N49, N50, N51, N52, N53, N55, N56, N57, N58, N59, N60, N61,
         N62, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, net10685, net10691, net10696, n55, n56,
         n57, n18, n19, n20, n21, n22, n23, n24, n25, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n58, n2, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n26, n27, n28, n29;
  wire   [1:0] ntrancnt;
  wire   [7:0] trans0;
  wire   [7:0] ttranwin_minus;
  wire   [7:0] trans1;

  SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 clk_gate_trans1_reg ( .CLK(clk), .EN(N90), 
        .ENCLK(net10685), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 clk_gate_trans0_reg ( .CLK(clk), .EN(N91), 
        .ENCLK(net10691), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 clk_gate_ttranwin_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net10696), .TE(test_se) );
  phyidd_a0_DW01_sub_0 sub_47 ( .A(trans1), .B(trans0), .CI(1'b0), .DIFF({N53, 
        N52, N51, N50, N49, N48, N47, N46}), .CO() );
  phyidd_a0_DW01_sub_1 sub_24 ( .A({n25, n24, n23, n22, n21, n20, n19, n18}), 
        .B(trans0), .CI(1'b0), .DIFF(ttranwin_minus), .CO() );
  phyidd_a0_DW01_inc_0 add_23 ( .A({test_so, ttranwin_6_, ttranwin_5_, 
        ttranwin_4_, ttranwin_3_, ttranwin_2_, ttranwin_1_, ttranwin_0_}), 
        .SUM({N18, N17, N16, N15, N14, N13, N12, N11}) );
  SDFFQX1 trans1_reg_7_ ( .D(N80), .SIN(trans1[6]), .SMC(test_se), .C(net10685), .Q(trans1[7]) );
  SDFFQX1 trans0_reg_7_ ( .D(N62), .SIN(trans0[6]), .SMC(test_se), .C(net10691), .Q(trans0[7]) );
  SDFFQX1 trans1_reg_6_ ( .D(N79), .SIN(trans1[5]), .SMC(test_se), .C(net10685), .Q(trans1[6]) );
  SDFFQX1 trans1_reg_5_ ( .D(N78), .SIN(trans1[4]), .SMC(test_se), .C(net10685), .Q(trans1[5]) );
  SDFFQX1 trans0_reg_6_ ( .D(N61), .SIN(trans0[5]), .SMC(test_se), .C(net10691), .Q(trans0[6]) );
  SDFFQX1 trans1_reg_4_ ( .D(N77), .SIN(trans1[3]), .SMC(test_se), .C(net10685), .Q(trans1[4]) );
  SDFFQX1 ntrancnt_reg_1_ ( .D(n56), .SIN(ntrancnt[0]), .SMC(test_se), .C(clk), 
        .Q(ntrancnt[1]) );
  SDFFQX1 ntrancnt_reg_0_ ( .D(n57), .SIN(n30), .SMC(test_se), .C(clk), .Q(
        ntrancnt[0]) );
  SDFFQX1 trans0_reg_5_ ( .D(N60), .SIN(trans0[4]), .SMC(test_se), .C(net10691), .Q(trans0[5]) );
  SDFFQX1 trans0_reg_4_ ( .D(N59), .SIN(trans0[3]), .SMC(test_se), .C(net10691), .Q(trans0[4]) );
  SDFFQX1 trans1_reg_3_ ( .D(N76), .SIN(trans1[2]), .SMC(test_se), .C(net10685), .Q(trans1[3]) );
  SDFFQX1 trans1_reg_2_ ( .D(N75), .SIN(trans1[1]), .SMC(test_se), .C(net10685), .Q(trans1[2]) );
  SDFFQX1 trans0_reg_3_ ( .D(N58), .SIN(trans0[2]), .SMC(test_se), .C(net10691), .Q(trans0[3]) );
  SDFFQX1 trans1_reg_1_ ( .D(N74), .SIN(trans1[0]), .SMC(test_se), .C(net10685), .Q(trans1[1]) );
  SDFFQX1 trans1_reg_0_ ( .D(N73), .SIN(trans0[7]), .SMC(test_se), .C(net10685), .Q(trans1[0]) );
  SDFFQX1 trans0_reg_2_ ( .D(N57), .SIN(trans0[1]), .SMC(test_se), .C(net10691), .Q(trans0[2]) );
  SDFFQX1 trans0_reg_1_ ( .D(N56), .SIN(trans0[0]), .SMC(test_se), .C(net10691), .Q(trans0[1]) );
  SDFFQX1 ttranwin_reg_7_ ( .D(N89), .SIN(ttranwin_6_), .SMC(test_se), .C(
        net10696), .Q(test_so) );
  SDFFQX1 ttranwin_reg_6_ ( .D(N88), .SIN(ttranwin_5_), .SMC(test_se), .C(
        net10696), .Q(ttranwin_6_) );
  SDFFQX1 trans0_reg_0_ ( .D(N55), .SIN(ntrancnt[1]), .SMC(test_se), .C(
        net10691), .Q(trans0[0]) );
  SDFFQX1 ttranwin_reg_5_ ( .D(N87), .SIN(ttranwin_4_), .SMC(test_se), .C(
        net10696), .Q(ttranwin_5_) );
  SDFFQX1 ttranwin_reg_4_ ( .D(N86), .SIN(ttranwin_3_), .SMC(test_se), .C(
        net10696), .Q(ttranwin_4_) );
  SDFFQX1 ttranwin_reg_1_ ( .D(N83), .SIN(ttranwin_0_), .SMC(test_se), .C(
        net10696), .Q(ttranwin_1_) );
  SDFFQX1 ttranwin_reg_2_ ( .D(N84), .SIN(ttranwin_1_), .SMC(test_se), .C(
        net10696), .Q(ttranwin_2_) );
  SDFFQX1 ttranwin_reg_3_ ( .D(N85), .SIN(ttranwin_2_), .SMC(test_se), .C(
        net10696), .Q(ttranwin_3_) );
  SDFFQX1 ttranwin_reg_0_ ( .D(N82), .SIN(trans1[7]), .SMC(test_se), .C(
        net10696), .Q(ttranwin_0_) );
  SDFFQX1 ccidle_reg ( .D(n55), .SIN(test_si), .SMC(test_se), .C(clk), .Q(n30)
         );
  INVX1 U5 ( .A(n29), .Y(o_ccidle) );
  NAND2X1 U6 ( .A(ntrancnt[0]), .B(n14), .Y(n2) );
  NAND2X1 U7 ( .A(ntrancnt[1]), .B(n15), .Y(n5) );
  INVX1 U8 ( .A(n52), .Y(n8) );
  INVX1 U9 ( .A(srstz), .Y(n6) );
  INVX1 U10 ( .A(n47), .Y(o_goidle) );
  OAI22X1 U11 ( .A(n8), .B(n11), .C(n49), .D(n33), .Y(N87) );
  OAI22X1 U12 ( .A(n8), .B(n10), .C(n32), .D(n49), .Y(N88) );
  NOR3XL U13 ( .A(n6), .B(o_goidle), .C(o_gobusy), .Y(n46) );
  OAI22X1 U14 ( .A(n8), .B(n12), .C(n49), .D(n34), .Y(N86) );
  NOR2X1 U15 ( .A(n13), .B(n48), .Y(n52) );
  OAI22X1 U16 ( .A(n8), .B(n16), .C(n49), .D(n35), .Y(N85) );
  OAI22X1 U17 ( .A(n8), .B(n17), .C(n49), .D(n36), .Y(N84) );
  OAI22X1 U18 ( .A(n8), .B(n26), .C(n49), .D(n37), .Y(N83) );
  INVX1 U19 ( .A(n45), .Y(n13) );
  NAND2X1 U20 ( .A(N12), .B(n44), .Y(n37) );
  OAI22X1 U21 ( .A(n13), .B(n9), .C(n31), .D(n5), .Y(N80) );
  OAI22X1 U22 ( .A(n8), .B(n9), .C(n31), .D(n49), .Y(N89) );
  INVX1 U23 ( .A(n38), .Y(n18) );
  AOI21X1 U24 ( .B(n28), .C(n29), .A(i_goidle), .Y(n47) );
  NOR3XL U25 ( .A(n7), .B(n42), .C(n29), .Y(o_gobusy) );
  INVX1 U26 ( .A(ttranwin_minus[5]), .Y(n11) );
  INVX1 U27 ( .A(ttranwin_minus[6]), .Y(n10) );
  NAND2X1 U28 ( .A(N13), .B(n44), .Y(n36) );
  NAND2X1 U29 ( .A(N14), .B(n44), .Y(n35) );
  OAI22X1 U30 ( .A(n13), .B(n11), .C(n5), .D(n33), .Y(N78) );
  OAI22X1 U31 ( .A(n13), .B(n10), .C(n32), .D(n42), .Y(N79) );
  INVX1 U32 ( .A(i_trans), .Y(n7) );
  INVX1 U33 ( .A(ttranwin_minus[4]), .Y(n12) );
  NOR2X1 U34 ( .A(N17), .B(n28), .Y(n32) );
  NAND2X1 U35 ( .A(N16), .B(n44), .Y(n33) );
  NAND2X1 U36 ( .A(N15), .B(n44), .Y(n34) );
  OAI221X1 U37 ( .A(i_trans), .B(n44), .C(n45), .D(n39), .E(n46), .Y(n40) );
  OAI22X1 U38 ( .A(n13), .B(n12), .C(n42), .D(n34), .Y(N77) );
  OAI22X1 U39 ( .A(n14), .B(n40), .C(n41), .D(n39), .Y(n56) );
  AND2X1 U40 ( .A(n42), .B(n2), .Y(n41) );
  ENOX1 U41 ( .A(n32), .B(n43), .C(N52), .D(n45), .Y(N61) );
  INVX1 U42 ( .A(n44), .Y(n28) );
  NAND2X1 U43 ( .A(n46), .B(i_trans), .Y(n39) );
  AOI31X1 U44 ( .A(n50), .B(n7), .C(n44), .D(n51), .Y(n49) );
  INVX1 U45 ( .A(ttranwin_minus[2]), .Y(n17) );
  INVX1 U46 ( .A(ttranwin_minus[3]), .Y(n16) );
  AOI21X1 U47 ( .B(n5), .C(n43), .A(n48), .Y(n51) );
  OAI22X1 U48 ( .A(n8), .B(n27), .C(n49), .D(n38), .Y(N82) );
  OAI22X1 U49 ( .A(n13), .B(n17), .C(n5), .D(n36), .Y(N75) );
  OAI22X1 U50 ( .A(n13), .B(n16), .C(n42), .D(n35), .Y(N76) );
  NAND2X1 U51 ( .A(n50), .B(i_trans), .Y(n48) );
  ENOX1 U52 ( .A(n43), .B(n33), .C(N51), .D(n45), .Y(N60) );
  OAI211X1 U53 ( .C(i_trans), .D(n28), .A(n50), .B(n53), .Y(N81) );
  NOR2X1 U54 ( .A(n52), .B(n51), .Y(n53) );
  INVX1 U55 ( .A(ttranwin_minus[1]), .Y(n26) );
  OAI22X1 U56 ( .A(n13), .B(n27), .C(n5), .D(n38), .Y(N73) );
  OAI22X1 U57 ( .A(n13), .B(n26), .C(n42), .D(n37), .Y(N74) );
  OAI21X1 U58 ( .B(n43), .C(n48), .A(n8), .Y(N91) );
  OAI21X1 U59 ( .B(n5), .C(n48), .A(n8), .Y(N90) );
  ENOX1 U60 ( .A(n2), .B(n35), .C(N49), .D(n45), .Y(N58) );
  ENOX1 U61 ( .A(n43), .B(n34), .C(N50), .D(n45), .Y(N59) );
  OAI211X1 U62 ( .C(o_gobusy), .D(n29), .A(n47), .B(srstz), .Y(n55) );
  ENOX1 U63 ( .A(n2), .B(n37), .C(N47), .D(n45), .Y(N56) );
  ENOX1 U64 ( .A(n43), .B(n36), .C(N48), .D(n45), .Y(N57) );
  NOR2X1 U65 ( .A(n15), .B(n14), .Y(n45) );
  INVX1 U66 ( .A(n36), .Y(n20) );
  INVX1 U67 ( .A(n35), .Y(n21) );
  INVX1 U68 ( .A(n34), .Y(n22) );
  INVX1 U69 ( .A(n33), .Y(n23) );
  INVX1 U70 ( .A(n37), .Y(n19) );
  INVX1 U71 ( .A(n32), .Y(n24) );
  NAND4X1 U72 ( .A(test_so), .B(ttranwin_6_), .C(n54), .D(n58), .Y(n44) );
  NOR2X1 U73 ( .A(ttranwin_1_), .B(ttranwin_0_), .Y(n54) );
  NOR4XL U74 ( .A(ttranwin_5_), .B(ttranwin_4_), .C(ttranwin_3_), .D(
        ttranwin_2_), .Y(n58) );
  NAND2X1 U75 ( .A(N11), .B(n44), .Y(n38) );
  INVX1 U76 ( .A(ttranwin_minus[7]), .Y(n9) );
  INVX1 U77 ( .A(n31), .Y(n25) );
  ENOX1 U78 ( .A(n31), .B(n2), .C(N53), .D(n45), .Y(N62) );
  OAI22X1 U79 ( .A(ntrancnt[0]), .B(n39), .C(n15), .D(n40), .Y(n57) );
  NOR2X1 U80 ( .A(N18), .B(n28), .Y(n31) );
  AOI31X1 U81 ( .A(n30), .B(n15), .C(i_trans), .D(n6), .Y(n50) );
  INVX1 U82 ( .A(n30), .Y(n29) );
  NAND2X1 U83 ( .A(ntrancnt[1]), .B(n15), .Y(n42) );
  INVX1 U84 ( .A(ttranwin_minus[0]), .Y(n27) );
  INVX1 U85 ( .A(ntrancnt[0]), .Y(n15) );
  NAND2X1 U86 ( .A(ntrancnt[0]), .B(n14), .Y(n43) );
  ENOX1 U87 ( .A(n2), .B(n38), .C(N46), .D(n45), .Y(N55) );
  INVX1 U88 ( .A(ntrancnt[1]), .Y(n14) );
endmodule


module phyidd_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module phyidd_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n17), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n10), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(A[0]), .Y(n18) );
  INVX1 U2 ( .A(B[2]), .Y(n14) );
  INVX1 U3 ( .A(B[3]), .Y(n15) );
  INVX1 U4 ( .A(B[4]), .Y(n13) );
  INVX1 U5 ( .A(B[5]), .Y(n11) );
  INVX1 U6 ( .A(B[1]), .Y(n17) );
  NAND21X1 U7 ( .B(n16), .A(n18), .Y(carry[1]) );
  INVX1 U8 ( .A(B[6]), .Y(n12) );
  INVX1 U9 ( .A(B[7]), .Y(n10) );
  INVX1 U10 ( .A(B[0]), .Y(n16) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module phyidd_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n18), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n10), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(B[2]), .Y(n14) );
  INVX1 U2 ( .A(B[3]), .Y(n15) );
  INVX1 U3 ( .A(B[4]), .Y(n13) );
  INVX1 U4 ( .A(B[5]), .Y(n11) );
  INVX1 U5 ( .A(B[1]), .Y(n18) );
  NAND21X1 U6 ( .B(n17), .A(n16), .Y(carry[1]) );
  INVX1 U7 ( .A(A[0]), .Y(n16) );
  INVX1 U8 ( .A(B[6]), .Y(n12) );
  INVX1 U9 ( .A(B[7]), .Y(n10) );
  INVX1 U10 ( .A(B[0]), .Y(n17) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_a0 ( i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, 
        r_rxdb_opt, r_ords_ena, r_pshords, r_rgdcrc, prx_cccnt, prx_rst, 
        prx_setsta, prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, 
        prx_fifopsh, prx_fifowdat, pff_txreq, pid_gobusy, pid_goidle, 
        pid_ccidle, pcc_rxgood, prx_crcstart, prx_crcshfi4, prx_crcsidat, 
        prx_rxcode, prx_adpn, prx_rcvdords, prx_eoprcvd, prx_fsm, clk, srstz, 
        test_si, test_so, test_se );
  input [1:0] r_rxdb_opt;
  input [6:0] r_ords_ena;
  output [1:0] prx_cccnt;
  output [1:0] prx_rst;
  output [6:0] prx_setsta;
  output [7:0] prx_fifowdat;
  output [3:0] prx_crcsidat;
  output [4:0] prx_rxcode;
  output [5:0] prx_adpn;
  output [2:0] prx_rcvdords;
  output [3:0] prx_fsm;
  input i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_pshords,
         r_rgdcrc, pff_txreq, pid_gobusy, pid_goidle, pid_ccidle, pcc_rxgood,
         clk, srstz, test_si, test_se;
  output prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, prx_fifopsh,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd, test_so;
  wire   N32, db_gohi, db_golo, cctrans, shrtrans, N70, N71, N72, N73, N74,
         N75, N76, N96, N153, N154, N155, N156, N157, N236, N239, N246, N247,
         N248, N249, N250, N275, N276, N278, N279, net10713, net10719,
         net10724, net10729, net10734, net10739, net10744, n214, n300, n299,
         n284, n285, n286, n292, n6, n76, n127, n139, n141, n153, n154, n155,
         n164, n165, n224, n226, n2, n4, n5, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n23, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n140, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n156, n157, n158, n159, n160, n161, n162, n163, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n225, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n287, n288, n289, n290, n291, n294, n295, n296,
         n297, n298;
  wire   [5:0] cccnt;
  wire   [2:0] ps_dat5b;
  wire   [2:0] bcnt;
  wire   [7:3] ordsbuf;

  phyrx_db u0_phyrx_db ( .clk(clk), .srstz(n30), .x_cc(i_cc), .ptx_txact(n5), 
        .r_rxdb_opt(r_rxdb_opt), .gohi(db_gohi), .golo(db_golo), .gotrans(
        prx_trans), .test_si(n292), .test_so(test_so), .test_se(test_se) );
  phyrx_adp u0_phyrx_adp ( .clk(clk), .srstz(n31), .gohi(db_gohi), .golo(
        db_golo), .gobusy(pid_gobusy), .goidle(pid_goidle), .i_ccidle(
        pid_ccidle), .k0_det(n226), .r_adprx_en(r_adprx_en), .r_adp2nd(
        r_adp2nd), .adp_val(prx_adpn), .d_cc(prx_d_cc), .cctrans(cctrans), 
        .test_si(shrtrans), .test_so(n292), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 clk_gate_cccnt_reg ( .CLK(clk), .EN(N70), 
        .ENCLK(net10713), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 clk_gate_cs_dat5b_reg ( .CLK(clk), .EN(N153), 
        .ENCLK(net10719), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 clk_gate_bcnt_reg ( .CLK(clk), .EN(N236), 
        .ENCLK(net10724), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 clk_gate_cs_dat4b_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net10729), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 clk_gate_ordsbuf_reg ( .CLK(clk), .EN(n224), 
        .ENCLK(net10734), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 clk_gate_ordsbuf_reg_0 ( .CLK(clk), .EN(N250), .ENCLK(net10739), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 clk_gate_cs_bmni_reg ( .CLK(clk), .EN(N275), 
        .ENCLK(net10744), .TE(test_se) );
  SDFFQX1 ordsbuf_reg_4_ ( .D(n26), .SIN(ordsbuf[3]), .SMC(test_se), .C(
        net10734), .Q(ordsbuf[4]) );
  SDFFQX1 ordsbuf_reg_7_ ( .D(prx_fifowdat[7]), .SIN(ordsbuf[6]), .SMC(test_se), .C(net10734), .Q(ordsbuf[7]) );
  SDFFQX1 ordsbuf_reg_5_ ( .D(prx_fifowdat[5]), .SIN(ordsbuf[4]), .SMC(test_se), .C(net10734), .Q(ordsbuf[5]) );
  SDFFQX1 ordsbuf_reg_6_ ( .D(prx_fifowdat[6]), .SIN(ordsbuf[5]), .SMC(test_se), .C(net10734), .Q(ordsbuf[6]) );
  SDFFQX1 cs_dat4b_reg_1_ ( .D(prx_fifowdat[5]), .SIN(prx_rxcode[0]), .SMC(
        test_se), .C(net10729), .Q(prx_fifowdat[1]) );
  SDFFQX1 cs_dat4b_reg_2_ ( .D(prx_fifowdat[6]), .SIN(n7), .SMC(test_se), .C(
        net10729), .Q(n300) );
  SDFFQX1 ordsbuf_reg_3_ ( .D(N249), .SIN(prx_rcvdords[2]), .SMC(test_se), .C(
        net10739), .Q(ordsbuf[3]) );
  SDFFQX1 cs_dat4b_reg_0_ ( .D(prx_fifowdat[4]), .SIN(n4), .SMC(test_se), .C(
        net10729), .Q(prx_fifowdat[0]) );
  SDFFQX1 cs_dat4b_reg_3_ ( .D(prx_crcsidat[3]), .SIN(prx_fifowdat[2]), .SMC(
        test_se), .C(net10729), .Q(prx_rxcode[3]) );
  SDFFQX1 cs_dat4b_reg_4_ ( .D(N96), .SIN(prx_rxcode[3]), .SMC(test_se), .C(
        net10729), .Q(prx_rxcode[4]) );
  SDFFQX1 bcnt_reg_1_ ( .D(n294), .SIN(bcnt[0]), .SMC(test_se), .C(net10724), 
        .Q(bcnt[1]) );
  SDFFQX1 bcnt_reg_0_ ( .D(n289), .SIN(test_si), .SMC(test_se), .C(net10724), 
        .Q(bcnt[0]) );
  SDFFQX1 bcnt_reg_2_ ( .D(N239), .SIN(bcnt[1]), .SMC(test_se), .C(net10724), 
        .Q(bcnt[2]) );
  SDFFQX1 cs_bmni_reg_0_ ( .D(N276), .SIN(cccnt[5]), .SMC(test_se), .C(
        net10744), .Q(prx_fsm[0]) );
  SDFFQX1 cs_bmni_reg_2_ ( .D(N278), .SIN(prx_fsm[1]), .SMC(test_se), .C(
        net10744), .Q(prx_fsm[2]) );
  SDFFQX1 cs_dat5b_reg_0_ ( .D(N154), .SIN(prx_rxcode[4]), .SMC(test_se), .C(
        net10719), .Q(ps_dat5b[0]) );
  SDFFQX1 cs_bmni_reg_1_ ( .D(n295), .SIN(prx_fsm[0]), .SMC(test_se), .C(
        net10744), .Q(prx_fsm[1]) );
  SDFFQX1 cs_dat5b_reg_3_ ( .D(N157), .SIN(ps_dat5b[2]), .SMC(test_se), .C(
        net10719), .Q(prx_bmc) );
  SDFFQX1 cs_bmni_reg_3_ ( .D(N279), .SIN(prx_fsm[2]), .SMC(test_se), .C(
        net10744), .Q(prx_fsm[3]) );
  SDFFQX1 cs_dat5b_reg_2_ ( .D(N156), .SIN(ps_dat5b[1]), .SMC(test_se), .C(
        net10719), .Q(ps_dat5b[2]) );
  SDFFQX1 cs_dat5b_reg_1_ ( .D(N155), .SIN(ps_dat5b[0]), .SMC(test_se), .C(
        net10719), .Q(ps_dat5b[1]) );
  SDFFQX1 cccnt_reg_1_ ( .D(N72), .SIN(cccnt[0]), .SMC(test_se), .C(net10713), 
        .Q(cccnt[1]) );
  SDFFQX1 cccnt_reg_3_ ( .D(N74), .SIN(cccnt[2]), .SMC(test_se), .C(net10713), 
        .Q(cccnt[3]) );
  SDFFQX1 cccnt_reg_5_ ( .D(N76), .SIN(cccnt[4]), .SMC(test_se), .C(net10713), 
        .Q(cccnt[5]) );
  SDFFQX1 shrtrans_reg ( .D(n214), .SIN(ordsbuf[7]), .SMC(test_se), .C(clk), 
        .Q(shrtrans) );
  SDFFQX1 cccnt_reg_4_ ( .D(N75), .SIN(cccnt[3]), .SMC(test_se), .C(net10713), 
        .Q(cccnt[4]) );
  SDFFQX1 cccnt_reg_0_ ( .D(N71), .SIN(bcnt[2]), .SMC(test_se), .C(net10713), 
        .Q(cccnt[0]) );
  SDFFQX1 cccnt_reg_2_ ( .D(N73), .SIN(cccnt[1]), .SMC(test_se), .C(net10713), 
        .Q(cccnt[2]) );
  SDFFQX1 ordsbuf_reg_1_ ( .D(N247), .SIN(prx_rcvdords[0]), .SMC(test_se), .C(
        net10739), .Q(prx_rcvdords[1]) );
  SDFFQX1 ordsbuf_reg_2_ ( .D(N248), .SIN(prx_rcvdords[1]), .SMC(test_se), .C(
        net10739), .Q(prx_rcvdords[2]) );
  MUX2X1 U274 ( .D0(r_ords_ena[1]), .D1(r_ords_ena[2]), .S(n296), .Y(n285) );
  NOR21XL U273 ( .B(r_ords_ena[0]), .A(n291), .Y(n286) );
  MUX4X1 U272 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[4]), .D2(r_ords_ena[5]), 
        .D3(r_ords_ena[6]), .S0(n296), .S1(N32), .Y(n284) );
  SDFFQX1 ordsbuf_reg_0_ ( .D(N246), .SIN(prx_bmc), .SMC(test_se), .C(net10739), .Q(prx_rcvdords[0]) );
  NAND31XL U3 ( .C(n49), .A(n48), .B(n54), .Y(n50) );
  AO21X1 U4 ( .B(n282), .C(n118), .A(n117), .Y(n81) );
  AO21X1 U5 ( .B(prx_fsm[1]), .C(n257), .A(n256), .Y(n259) );
  NAND21X1 U6 ( .B(n251), .A(n234), .Y(n235) );
  AND2X1 U7 ( .A(n66), .B(n61), .Y(n53) );
  MUX2IX1 U8 ( .D0(n51), .D1(n50), .S(ps_dat5b[0]), .Y(n52) );
  NOR43XL U9 ( .B(prx_bmc), .C(n72), .D(n46), .A(ps_dat5b[1]), .Y(n51) );
  AND2X1 U10 ( .A(n31), .B(n218), .Y(n214) );
  AND2X1 U11 ( .A(prx_bmc), .B(n74), .Y(n64) );
  NAND32X1 U12 ( .B(n78), .C(n57), .A(n56), .Y(prx_fifowdat[5]) );
  AO21X1 U13 ( .B(ps_dat5b[0]), .C(n61), .A(n55), .Y(n56) );
  NOR3XL U14 ( .A(n205), .B(n35), .C(n36), .Y(prx_cccnt[0]) );
  NAND21X1 U15 ( .B(n53), .A(n52), .Y(n299) );
  INVXL U16 ( .A(n300), .Y(n2) );
  INVXL U17 ( .A(n2), .Y(prx_fifowdat[2]) );
  NAND3X4 U18 ( .A(cctrans), .B(shrtrans), .C(n217), .Y(n261) );
  AND3XL U19 ( .A(ps_dat5b[0]), .B(n72), .C(n74), .Y(n57) );
  INVX1 U20 ( .A(n16), .Y(n4) );
  BUFX3 U21 ( .A(ptx_txact), .Y(n5) );
  INVX1 U22 ( .A(n114), .Y(n7) );
  BUFX3 U23 ( .A(n7), .Y(prx_rxcode[1]) );
  BUFX3 U24 ( .A(prx_fifowdat[2]), .Y(prx_rxcode[2]) );
  BUFX3 U25 ( .A(prx_fifowdat[0]), .Y(prx_rxcode[0]) );
  INVX1 U26 ( .A(n261), .Y(n29) );
  INVX1 U27 ( .A(n54), .Y(n78) );
  INVX2 U28 ( .A(n43), .Y(n63) );
  INVX3 U29 ( .A(prx_fifowdat[5]), .Y(n80) );
  NAND32XL U30 ( .B(n71), .C(n238), .A(n189), .Y(n237) );
  NOR2X2 U31 ( .A(n251), .B(n221), .Y(n10) );
  NAND21X2 U32 ( .B(n80), .A(prx_fifowdat[6]), .Y(n67) );
  AND2XL U33 ( .A(n205), .B(n204), .Y(n207) );
  OR2XL U34 ( .A(prx_fifowdat[6]), .B(n103), .Y(n86) );
  AO21XL U35 ( .B(n15), .C(n253), .A(n9), .Y(prx_crcshfi4) );
  OR2XL U36 ( .A(n204), .B(n205), .Y(n206) );
  INVX1 U37 ( .A(prx_fsm[3]), .Y(n16) );
  AND2XL U38 ( .A(cccnt[4]), .B(cccnt[2]), .Y(n42) );
  AO21XL U39 ( .B(cccnt[4]), .C(cccnt[3]), .A(cccnt[5]), .Y(n38) );
  NAND2XL U40 ( .A(cccnt[2]), .B(n213), .Y(n205) );
  INVXL U41 ( .A(shrtrans), .Y(n216) );
  INVXL U42 ( .A(cccnt[1]), .Y(n211) );
  INVXL U43 ( .A(cccnt[5]), .Y(n35) );
  XOR2XL U44 ( .A(cccnt[2]), .B(n213), .Y(n203) );
  XOR2XL U45 ( .A(cccnt[4]), .B(n210), .Y(n208) );
  INVXL U46 ( .A(prx_rcvdords[1]), .Y(n159) );
  OR2XL U47 ( .A(prx_rcvdords[2]), .B(n100), .Y(n83) );
  INVXL U48 ( .A(prx_rcvdords[2]), .Y(n89) );
  MUX2BXL U49 ( .D0(n248), .D1(n8), .S(prx_rcvdords[2]), .Y(n270) );
  AOI21X1 U50 ( .B(r_ords_ena[5]), .C(n247), .A(n246), .Y(n8) );
  NAND21XL U51 ( .B(n100), .A(prx_rcvdords[2]), .Y(n101) );
  MUX3XL U52 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[4]), .D2(n245), .S0(
        prx_rcvdords[0]), .S1(prx_rcvdords[1]), .Y(n246) );
  AND2XL U53 ( .A(r_ords_ena[6]), .B(prx_rcvdords[0]), .Y(n245) );
  NAND43XL U54 ( .B(n125), .C(n244), .D(n124), .A(prx_rcvdords[2]), .Y(n138)
         );
  INVXL U55 ( .A(prx_rcvdords[0]), .Y(n241) );
  MUX2IXL U56 ( .D0(r_ords_ena[0]), .D1(r_ords_ena[2]), .S(prx_rcvdords[1]), 
        .Y(n242) );
  NAND21XL U57 ( .B(prx_rcvdords[0]), .A(prx_rcvdords[1]), .Y(n244) );
  NAND2XL U58 ( .A(n217), .B(n216), .Y(n17) );
  INVXL U59 ( .A(cccnt[4]), .Y(n272) );
  NOR5XL U60 ( .A(cccnt[2]), .B(cccnt[3]), .C(cccnt[5]), .D(n272), .E(n271), 
        .Y(prx_cccnt[1]) );
  INVX1 U61 ( .A(n274), .Y(n280) );
  INVX1 U62 ( .A(n32), .Y(n31) );
  INVX1 U63 ( .A(n32), .Y(n30) );
  INVX1 U64 ( .A(n92), .Y(n93) );
  INVX1 U65 ( .A(n88), .Y(n133) );
  NAND21X1 U66 ( .B(n131), .A(n136), .Y(n274) );
  INVX1 U67 ( .A(N32), .Y(n297) );
  INVX1 U68 ( .A(n156), .Y(n174) );
  NAND21X1 U69 ( .B(n297), .A(n156), .Y(n76) );
  INVX1 U70 ( .A(n238), .Y(n227) );
  INVX1 U71 ( .A(n237), .Y(n73) );
  AND2XL U72 ( .A(n73), .B(n72), .Y(N157) );
  INVX1 U73 ( .A(srstz), .Y(n32) );
  INVX1 U74 ( .A(pid_goidle), .Y(n225) );
  NAND21X1 U75 ( .B(n75), .A(n63), .Y(n54) );
  INVXL U76 ( .A(n55), .Y(n66) );
  INVX1 U77 ( .A(n152), .Y(n234) );
  NAND32X1 U78 ( .B(n240), .C(n32), .A(n239), .Y(N70) );
  INVX1 U79 ( .A(n239), .Y(n209) );
  NAND21X1 U80 ( .B(n86), .A(n137), .Y(n88) );
  OR2X1 U81 ( .A(n162), .B(n144), .Y(n288) );
  OAI32X1 U82 ( .A(n85), .B(n131), .C(n88), .D(n84), .E(n119), .Y(n96) );
  INVX1 U83 ( .A(n118), .Y(n85) );
  AND2X1 U84 ( .A(n252), .B(n10), .Y(n9) );
  AO21X1 U85 ( .B(n166), .C(n163), .A(n162), .Y(n167) );
  AO21X1 U86 ( .B(n112), .C(n288), .A(n149), .Y(N32) );
  INVX1 U87 ( .A(n151), .Y(n112) );
  NAND21X1 U88 ( .B(n119), .A(n280), .Y(n129) );
  NAND21X1 U89 ( .B(n274), .A(n278), .Y(n277) );
  OR2X1 U90 ( .A(n147), .B(n111), .Y(n149) );
  INVX1 U91 ( .A(n86), .Y(n136) );
  INVX1 U92 ( .A(n169), .Y(n147) );
  OAI21X1 U93 ( .B(n139), .C(n151), .A(n150), .Y(n156) );
  NAND21X1 U94 ( .B(n141), .A(n290), .Y(n139) );
  INVX1 U95 ( .A(n149), .Y(n150) );
  INVX1 U96 ( .A(n288), .Y(n290) );
  INVX1 U97 ( .A(n296), .Y(n291) );
  INVX1 U98 ( .A(n253), .Y(n175) );
  AO21X1 U99 ( .B(n6), .C(n265), .A(prx_setsta[6]), .Y(prx_fiforst) );
  NAND2X1 U100 ( .A(n76), .B(n233), .Y(n186) );
  INVX1 U101 ( .A(n84), .Y(n137) );
  NAND2X1 U102 ( .A(n249), .B(n30), .Y(n238) );
  AO21X1 U103 ( .B(n126), .C(n118), .A(n117), .Y(n132) );
  INVX1 U104 ( .A(n119), .Y(n117) );
  INVX1 U105 ( .A(n120), .Y(n135) );
  NAND21X1 U106 ( .B(n119), .A(n126), .Y(n120) );
  NAND32X1 U107 ( .B(pid_gobusy), .C(n238), .A(n237), .Y(N153) );
  INVX1 U108 ( .A(n229), .Y(n193) );
  INVX1 U109 ( .A(n236), .Y(n197) );
  NAND32X1 U110 ( .B(n6), .C(n32), .A(n236), .Y(N236) );
  INVXL U111 ( .A(n235), .Y(n224) );
  INVX1 U112 ( .A(n254), .Y(n255) );
  INVX1 U113 ( .A(n232), .Y(n191) );
  INVX1 U114 ( .A(pid_gobusy), .Y(n189) );
  INVX1 U115 ( .A(n206), .Y(n210) );
  AND2X1 U116 ( .A(n234), .B(prx_fifowdat[3]), .Y(N249) );
  INVX1 U117 ( .A(n264), .Y(n71) );
  INVX1 U118 ( .A(n59), .Y(n75) );
  INVX1 U119 ( .A(n271), .Y(n213) );
  INVX1 U120 ( .A(n113), .Y(n178) );
  NAND32X1 U121 ( .B(n177), .C(n258), .A(n257), .Y(n113) );
  INVX1 U122 ( .A(n221), .Y(n233) );
  NAND32X1 U123 ( .B(n257), .C(n177), .A(n79), .Y(n152) );
  INVX1 U124 ( .A(n123), .Y(prx_fifowdat[3]) );
  NAND21X1 U125 ( .B(pff_txreq), .A(n33), .Y(n240) );
  OAI31XL U126 ( .A(n206), .B(n272), .C(n35), .D(n34), .Y(n239) );
  INVX1 U127 ( .A(n240), .Y(n34) );
  AO21X1 U128 ( .B(n209), .C(n212), .A(n32), .Y(N71) );
  OAI31XL U129 ( .A(n207), .B(n210), .C(n239), .D(n31), .Y(N74) );
  OAI31XL U130 ( .A(n215), .B(n213), .C(n239), .D(n31), .Y(N72) );
  AND2X1 U131 ( .A(n212), .B(n211), .Y(n215) );
  AO21X1 U132 ( .B(n255), .C(n6), .A(n9), .Y(prx_crcstart) );
  NAND21XL U133 ( .B(n80), .A(prx_fifowdat[7]), .Y(n103) );
  NAND43X1 U134 ( .B(n111), .C(n288), .D(n110), .A(n153), .Y(n169) );
  NAND2X1 U135 ( .A(n154), .B(n155), .Y(n153) );
  INVX1 U136 ( .A(n141), .Y(n110) );
  OA21X1 U137 ( .B(n276), .C(n277), .A(n275), .Y(n154) );
  NAND43X1 U138 ( .B(n173), .C(n172), .D(n171), .A(n170), .Y(n252) );
  INVX1 U139 ( .A(n158), .Y(n172) );
  INVX1 U140 ( .A(n157), .Y(n173) );
  OAI211X1 U141 ( .C(n275), .D(n169), .A(n168), .B(n167), .Y(n171) );
  NAND21X1 U142 ( .B(n97), .A(n163), .Y(n144) );
  GEN2XL U143 ( .D(n96), .E(n114), .C(n95), .B(n94), .A(n93), .Y(n97) );
  INVX1 U144 ( .A(n140), .Y(n94) );
  INVX1 U145 ( .A(n129), .Y(n95) );
  NOR2X1 U146 ( .A(n164), .B(n165), .Y(n141) );
  OAI221X1 U147 ( .A(n91), .B(n90), .C(n114), .D(n92), .E(n157), .Y(n162) );
  OA21X1 U148 ( .B(n87), .C(n114), .A(n129), .Y(n91) );
  INVX1 U149 ( .A(n96), .Y(n87) );
  NAND32X1 U150 ( .B(n151), .C(n147), .A(n146), .Y(n296) );
  NAND21X1 U151 ( .B(n162), .A(n145), .Y(n146) );
  NAND21X1 U152 ( .B(n144), .A(n143), .Y(n145) );
  NAND21X1 U153 ( .B(n164), .A(n165), .Y(n143) );
  NOR2X1 U154 ( .A(n291), .B(n76), .Y(prx_rst[0]) );
  NOR2X1 U155 ( .A(n296), .B(n76), .Y(prx_rst[1]) );
  OAI211X1 U156 ( .C(n287), .D(n283), .A(n282), .B(n281), .Y(n155) );
  INVX1 U157 ( .A(n276), .Y(n287) );
  AO21X1 U158 ( .B(n280), .C(n279), .A(n278), .Y(n281) );
  INVX1 U159 ( .A(n277), .Y(n283) );
  NAND43XL U160 ( .B(n23), .C(n69), .D(prx_fifowdat[4]), .A(n80), .Y(n253) );
  NAND21X1 U161 ( .B(n109), .A(n158), .Y(n111) );
  OAI33XL U162 ( .A(n160), .B(n276), .C(n273), .D(n104), .E(n26), .F(n103), 
        .Y(n109) );
  GEN2XL U163 ( .D(n160), .E(n276), .C(n273), .B(n102), .A(n23), .Y(n104) );
  NAND32X1 U164 ( .B(n160), .C(n276), .A(n279), .Y(n102) );
  AND3X1 U165 ( .A(prx_eoprcvd), .B(pcc_rxgood), .C(n268), .Y(prx_setsta[3])
         );
  INVX1 U166 ( .A(n250), .Y(prx_eoprcvd) );
  NAND32X1 U167 ( .B(n249), .C(n16), .A(n270), .Y(n250) );
  INVX1 U168 ( .A(n266), .Y(n267) );
  OA21X1 U169 ( .B(n185), .C(n184), .A(n193), .Y(N279) );
  INVX1 U170 ( .A(n188), .Y(n185) );
  NAND3X1 U171 ( .A(n11), .B(n12), .C(n170), .Y(n151) );
  NAND4X1 U172 ( .A(n133), .B(n131), .C(n81), .D(n114), .Y(n11) );
  NAND3X1 U173 ( .A(n282), .B(n117), .C(n82), .Y(n12) );
  INVX1 U174 ( .A(n260), .Y(prx_setsta[6]) );
  NAND32X1 U175 ( .B(n268), .C(n269), .A(prx_eoprcvd), .Y(n260) );
  AOI31X1 U176 ( .A(n183), .B(n223), .C(n196), .D(n229), .Y(n295) );
  INVX1 U177 ( .A(n184), .Y(n183) );
  GEN2XL U178 ( .D(n194), .E(n267), .C(n220), .B(n193), .A(n192), .Y(N276) );
  AND4X1 U179 ( .A(n191), .B(n227), .C(prx_idle), .D(n225), .Y(n192) );
  INVX1 U180 ( .A(n186), .Y(n194) );
  INVX1 U181 ( .A(n231), .Y(prx_idle) );
  AOI21X1 U182 ( .B(n176), .C(n181), .A(n229), .Y(N278) );
  AO21X1 U183 ( .B(n252), .C(n266), .A(n186), .Y(n176) );
  OAI22X1 U184 ( .A(n114), .B(n152), .C(n297), .D(n221), .Y(N247) );
  OAI22X1 U185 ( .A(n148), .B(n152), .C(n291), .D(n221), .Y(N246) );
  OAI22X1 U186 ( .A(n174), .B(n221), .C(n2), .D(n152), .Y(N248) );
  NAND32X1 U187 ( .B(n123), .C(n148), .A(n2), .Y(n84) );
  NAND21X1 U188 ( .B(n83), .A(n298), .Y(n119) );
  NAND21X1 U189 ( .B(n298), .A(n83), .Y(n118) );
  NAND32X1 U190 ( .B(n124), .C(n241), .A(n159), .Y(n100) );
  NAND32X1 U191 ( .B(n140), .C(n161), .A(n159), .Y(n157) );
  NAND32X1 U192 ( .B(n140), .C(n138), .A(n148), .Y(n168) );
  NAND32X1 U193 ( .B(n161), .C(n159), .A(n282), .Y(n163) );
  NAND32X1 U194 ( .B(n148), .C(n138), .A(n126), .Y(n166) );
  INVX1 U195 ( .A(n101), .Y(n108) );
  NAND32X1 U196 ( .B(n99), .C(n98), .A(n116), .Y(n160) );
  NAND32X1 U197 ( .B(n99), .C(n116), .A(n98), .Y(n140) );
  NAND6XL U198 ( .A(n108), .B(n107), .C(n106), .D(prx_fifowdat[3]), .E(n105), 
        .F(n148), .Y(n158) );
  INVX1 U199 ( .A(n122), .Y(n106) );
  INVX1 U200 ( .A(n160), .Y(n107) );
  NAND21X1 U201 ( .B(n298), .A(n101), .Y(n279) );
  NAND32X1 U202 ( .B(n161), .C(n160), .A(n159), .Y(n275) );
  INVX1 U203 ( .A(n130), .Y(n126) );
  INVX1 U204 ( .A(n273), .Y(n278) );
  OAI221X1 U205 ( .A(n232), .B(n231), .C(n230), .D(n229), .E(n228), .Y(N275)
         );
  AND4X1 U206 ( .A(n223), .B(n222), .C(n254), .D(n221), .Y(n230) );
  AND2X1 U207 ( .A(n227), .B(n225), .Y(n228) );
  INVX1 U208 ( .A(n220), .Y(n222) );
  OAI2B11X1 U209 ( .D(n262), .C(n196), .A(n231), .B(n195), .Y(n236) );
  INVX1 U210 ( .A(n90), .Y(n282) );
  INVX1 U211 ( .A(n244), .Y(n247) );
  INVX1 U212 ( .A(n200), .Y(n289) );
  INVX1 U213 ( .A(pcc_rxgood), .Y(n269) );
  INVX1 U214 ( .A(n196), .Y(n265) );
  NAND21X1 U215 ( .B(n16), .A(n178), .Y(n254) );
  OR2X1 U216 ( .A(n189), .B(n5), .Y(n232) );
  NAND2X1 U217 ( .A(n187), .B(n188), .Y(n220) );
  INVX1 U218 ( .A(n182), .Y(n223) );
  NAND21X1 U219 ( .B(n234), .A(n181), .Y(n182) );
  NAND32X1 U220 ( .B(n16), .C(n177), .A(n258), .Y(n188) );
  AND4XL U221 ( .A(n265), .B(n264), .C(n263), .D(n262), .Y(prx_setsta[0]) );
  OAI21BBX1 U222 ( .A(ps_dat5b[0]), .B(n66), .C(n13), .Y(prx_fifowdat[6]) );
  MUX2IX1 U223 ( .D0(n65), .D1(n64), .S(n63), .Y(n13) );
  MUX2IXL U224 ( .D0(n27), .D1(n28), .S(n63), .Y(n44) );
  NAND2X1 U225 ( .A(n75), .B(ps_dat5b[0]), .Y(n28) );
  MUX2IX1 U226 ( .D0(n75), .D1(n47), .S(n72), .Y(n48) );
  AND2X1 U227 ( .A(ps_dat5b[1]), .B(n46), .Y(n47) );
  OR3XL U228 ( .A(bcnt[0]), .B(n201), .C(bcnt[1]), .Y(n70) );
  OAI21BBX1 U229 ( .A(r_pshords), .B(N250), .C(n14), .Y(prx_fifopsh) );
  NAND3X1 U230 ( .A(n259), .B(n258), .C(n15), .Y(n14) );
  NOR2XL U231 ( .A(n251), .B(n16), .Y(n15) );
  NAND21X1 U232 ( .B(cccnt[4]), .A(n204), .Y(n36) );
  AO21X1 U233 ( .B(cccnt[1]), .C(cccnt[2]), .A(cccnt[5]), .Y(n39) );
  INVX1 U234 ( .A(n41), .Y(n217) );
  GEN2XL U235 ( .D(cccnt[2]), .E(n40), .C(n39), .B(n38), .A(n37), .Y(n41) );
  NAND21X1 U236 ( .B(cccnt[0]), .A(shrtrans), .Y(n40) );
  AOI211X1 U237 ( .C(cccnt[0]), .D(cccnt[2]), .A(n36), .B(n39), .Y(n37) );
  INVX1 U238 ( .A(cccnt[3]), .Y(n204) );
  NAND21X1 U239 ( .B(n74), .A(prx_bmc), .Y(n59) );
  NAND21X1 U240 ( .B(n211), .A(cccnt[0]), .Y(n271) );
  INVX1 U241 ( .A(ps_dat5b[1]), .Y(n74) );
  INVX1 U242 ( .A(ps_dat5b[2]), .Y(n46) );
  NAND21X1 U243 ( .B(n190), .A(prx_fsm[0]), .Y(n196) );
  NAND21X1 U244 ( .B(prx_fsm[1]), .A(n79), .Y(n190) );
  INVX1 U245 ( .A(prx_fsm[2]), .Y(n258) );
  INVX1 U246 ( .A(n45), .Y(n79) );
  NAND21X1 U247 ( .B(prx_fsm[3]), .A(n258), .Y(n45) );
  INVX1 U248 ( .A(prx_bmc), .Y(n61) );
  INVX1 U249 ( .A(ps_dat5b[0]), .Y(n60) );
  NAND21X1 U250 ( .B(prx_fsm[3]), .A(n178), .Y(n221) );
  INVX1 U251 ( .A(bcnt[2]), .Y(n201) );
  INVX1 U252 ( .A(prx_fsm[1]), .Y(n177) );
  INVX1 U253 ( .A(prx_fsm[0]), .Y(n257) );
  INVX1 U254 ( .A(n179), .Y(n256) );
  NAND21X1 U255 ( .B(prx_fsm[1]), .A(prx_fsm[0]), .Y(n179) );
  MUX2IX1 U256 ( .D0(prx_rxcode[4]), .D1(prx_rxcode[3]), .S(prx_fsm[3]), .Y(
        n123) );
  GEN2XL U257 ( .D(n210), .E(cccnt[4]), .C(cccnt[5]), .B(n209), .A(n32), .Y(
        N76) );
  AO21X1 U258 ( .B(n203), .C(n209), .A(n32), .Y(N73) );
  AO21X1 U259 ( .B(n208), .C(n209), .A(n32), .Y(N75) );
  AO21XL U260 ( .B(n78), .C(prx_bmc), .A(n77), .Y(prx_crcsidat[3]) );
  NAND21X1 U261 ( .B(n142), .A(n168), .Y(n165) );
  GEN2XL U262 ( .D(prx_fifowdat[1]), .E(n137), .C(n136), .B(n135), .A(n134), 
        .Y(n142) );
  AND4X1 U263 ( .A(prx_fifowdat[1]), .B(n133), .C(n132), .D(n131), .Y(n134) );
  AND2XL U264 ( .A(n10), .B(n266), .Y(prx_setsta[1]) );
  MUX2BXL U265 ( .D0(n284), .D1(n127), .S(n174), .Y(n266) );
  AOI22X1 U266 ( .A(n286), .B(n297), .C(n285), .D(N32), .Y(n127) );
  OAI211X1 U267 ( .C(n130), .D(n129), .A(n128), .B(n166), .Y(n164) );
  NAND43X1 U268 ( .B(n123), .C(n122), .D(prx_rxcode[0]), .A(n121), .Y(n128) );
  AO21X1 U269 ( .B(n280), .C(n132), .A(n135), .Y(n121) );
  AND2XL U270 ( .A(n10), .B(n267), .Y(prx_setsta[2]) );
  OAI211X1 U271 ( .C(prx_fsm[0]), .D(n188), .A(n254), .B(n180), .Y(n184) );
  OA22X1 U275 ( .A(n265), .B(n187), .C(n267), .D(n186), .Y(n180) );
  OAI22X1 U276 ( .A(n7), .B(n84), .C(n26), .D(n86), .Y(n82) );
  AND2X1 U277 ( .A(prx_eoprcvd), .B(n269), .Y(prx_setsta[4]) );
  NAND43X1 U278 ( .B(prx_fifowdat[1]), .C(n123), .D(n148), .A(prx_fifowdat[2]), 
        .Y(n276) );
  NAND43X1 U279 ( .B(r_exist1st), .C(prx_fifowdat[2]), .D(n123), .A(n7), .Y(
        n125) );
  NAND21X1 U280 ( .B(r_ordrs4), .A(n108), .Y(n273) );
  NAND6XL U281 ( .A(prx_fifowdat[1]), .B(ordsbuf[3]), .C(prx_rcvdords[0]), .D(
        n137), .E(n105), .F(n89), .Y(n161) );
  INVX1 U282 ( .A(prx_fifowdat[0]), .Y(n148) );
  INVX1 U283 ( .A(ordsbuf[3]), .Y(n124) );
  NAND43X1 U284 ( .B(ordsbuf[4]), .C(n116), .D(n115), .A(ordsbuf[6]), .Y(n130)
         );
  OAI22X1 U285 ( .A(n244), .B(n243), .C(n242), .D(n241), .Y(n248) );
  INVX1 U286 ( .A(r_ords_ena[1]), .Y(n243) );
  NAND21X1 U287 ( .B(n115), .A(ordsbuf[4]), .Y(n99) );
  INVX1 U288 ( .A(ordsbuf[6]), .Y(n98) );
  AND2X1 U289 ( .A(n73), .B(prx_bmc), .Y(N156) );
  AND2X1 U290 ( .A(n73), .B(ps_dat5b[1]), .Y(N154) );
  AND2X1 U291 ( .A(n73), .B(ps_dat5b[2]), .Y(N155) );
  INVX1 U292 ( .A(r_ordrs4), .Y(n298) );
  INVX1 U293 ( .A(ordsbuf[5]), .Y(n116) );
  INVX1 U294 ( .A(r_exist1st), .Y(n105) );
  INVX1 U295 ( .A(ordsbuf[7]), .Y(n115) );
  NAND32X1 U296 ( .B(ordsbuf[5]), .C(n99), .A(n98), .Y(n90) );
  NAND21X1 U297 ( .B(n114), .A(prx_fifowdat[2]), .Y(n122) );
  NAND21X1 U298 ( .B(bcnt[0]), .A(n197), .Y(n200) );
  MUX2X1 U299 ( .D0(n198), .D1(n289), .S(bcnt[1]), .Y(n294) );
  AND2X1 U300 ( .A(bcnt[0]), .B(n197), .Y(n198) );
  INVX1 U301 ( .A(prx_fifowdat[1]), .Y(n114) );
  INVX1 U302 ( .A(r_rgdcrc), .Y(n268) );
  OAI22X1 U303 ( .A(n202), .B(n236), .C(n201), .D(n200), .Y(N239) );
  MUX2BXL U304 ( .D0(n201), .D1(n199), .S(bcnt[1]), .Y(n202) );
  AND2X1 U305 ( .A(bcnt[0]), .B(n201), .Y(n199) );
  OR4X1 U306 ( .A(prx_fifowdat[0]), .B(n83), .C(n90), .D(n125), .Y(n170) );
  AND3X1 U307 ( .A(pid_goidle), .B(prx_fsm[3]), .C(n270), .Y(prx_setsta[5]) );
  MUX2BXL U308 ( .D0(shrtrans), .D1(n17), .S(cctrans), .Y(n218) );
  OR2X1 U309 ( .A(prx_fsm[0]), .B(n190), .Y(n231) );
  NAND21X1 U310 ( .B(bcnt[1]), .A(n201), .Y(n262) );
  NAND21X1 U311 ( .B(prx_fsm[2]), .A(n256), .Y(n187) );
  NAND43X1 U312 ( .B(n4), .C(prx_fsm[0]), .D(prx_fsm[2]), .A(prx_fsm[1]), .Y(
        n181) );
  INVX1 U313 ( .A(cccnt[0]), .Y(n212) );
  INVX1 U314 ( .A(n23), .Y(prx_crcsidat[2]) );
  INVXL U315 ( .A(prx_fifowdat[6]), .Y(n23) );
  BUFXL U316 ( .A(prx_fifowdat[5]), .Y(prx_crcsidat[1]) );
  BUFX3 U317 ( .A(prx_fifowdat[4]), .Y(prx_crcsidat[0]) );
  INVX2 U318 ( .A(n58), .Y(n62) );
  NOR21XL U319 ( .B(prx_bmc), .A(n58), .Y(n49) );
  NAND21X2 U320 ( .B(n46), .A(n29), .Y(n43) );
  NAND2XL U321 ( .A(n58), .B(n74), .Y(n27) );
  XOR2XL U322 ( .A(n261), .B(prx_bmc), .Y(n263) );
  AOI211XL U323 ( .C(n75), .D(ps_dat5b[2]), .A(n74), .B(n261), .Y(n77) );
  NAND32X1 U324 ( .B(n46), .C(n74), .A(n261), .Y(n55) );
  NAND21X2 U325 ( .B(ps_dat5b[2]), .A(n261), .Y(n58) );
  INVXL U326 ( .A(N96), .Y(n69) );
  BUFXL U327 ( .A(n299), .Y(prx_fifowdat[4]) );
  BUFXL U328 ( .A(n299), .Y(n26) );
  INVXL U329 ( .A(n251), .Y(n6) );
  AND3XL U330 ( .A(n31), .B(n264), .C(n251), .Y(n195) );
  NAND43X1 U331 ( .B(pid_goidle), .C(n175), .D(n251), .A(n30), .Y(n229) );
  NAND21XL U332 ( .B(n251), .A(n175), .Y(n249) );
  INVXL U333 ( .A(n219), .Y(n226) );
  NAND21X2 U334 ( .B(n299), .A(n67), .Y(n68) );
  INVX1 U335 ( .A(n26), .Y(n131) );
  NAND32X1 U336 ( .B(n88), .C(n119), .A(n26), .Y(n92) );
  INVX1 U337 ( .A(n261), .Y(n72) );
  OAI31XL U338 ( .A(n62), .B(n61), .C(n60), .D(n59), .Y(n65) );
  NAND21X1 U339 ( .B(n10), .A(n235), .Y(N250) );
  MUX2IXL U340 ( .D0(cctrans), .D1(prx_cccnt[0]), .S(n5), .Y(n33) );
  NAND32X2 U341 ( .B(n69), .C(n196), .A(n68), .Y(n219) );
  GEN2XL U342 ( .D(n42), .E(cccnt[3]), .C(cccnt[5]), .B(cctrans), .A(n72), .Y(
        n264) );
  MUX2XL U343 ( .D0(N96), .D1(prx_crcsidat[3]), .S(prx_fsm[3]), .Y(
        prx_fifowdat[7]) );
  GEN2X1 U344 ( .D(n74), .E(n60), .C(n61), .B(n261), .A(n44), .Y(N96) );
  AO21X4 U345 ( .B(n70), .C(n219), .A(n71), .Y(n251) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_adp ( clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, 
        r_adprx_en, r_adp2nd, adp_val, d_cc, cctrans, test_si, test_so, 
        test_se );
  output [5:0] adp_val;
  input clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, r_adprx_en,
         r_adp2nd, test_si, test_se;
  output d_cc, cctrans, test_so;
  wire   dcnt_n_2_, dcnt_n_1_, dcnt_n_0_, N49, N51, N52, N53, N55, N97, N98,
         N99, N100, N101, N102, N103, N104, N130, N131, N132, N133, N134, N135,
         N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N169,
         N170, N171, N172, N173, net10761, net10767, net10772, net10777, n115,
         n39, n41, n63, n65, n66, n67, n68, n69, n70, n71, n76, n92, n93, n113,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n40, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n64, n72, n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n114, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7;
  wire   [7:0] dcnt_h;
  wire   [5:0] adp_v0;
  wire   [5:0] dcnt_e;

  SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 clk_gate_adp_n_reg ( .CLK(clk), .EN(N49), 
        .ENCLK(net10761), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 clk_gate_dcnt_e_reg ( .CLK(clk), .EN(N130), 
        .ENCLK(net10767), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 clk_gate_dcnt_h_reg ( .CLK(clk), .EN(N137), 
        .ENCLK(net10772), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 clk_gate_dcnt_n_reg ( .CLK(clk), .EN(N169), 
        .ENCLK(net10777), .TE(test_se) );
  phyrx_adp_DW01_inc_0 add_385 ( .A(dcnt_h), .SUM({N104, N103, N102, N101, 
        N100, N99, N98, N97}) );
  phyrx_adp_DW_div_tc_6 div_338 ( .a({n4, dcnt_h}), .b({1'b0, 1'b1, 1'b1, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, adp_v0}), .remainder({SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7}), .divide_by_0() );
  SDFFQX1 dcnt_h_reg_6_ ( .D(N144), .SIN(dcnt_h[5]), .SMC(test_se), .C(
        net10772), .Q(dcnt_h[6]) );
  SDFFQX1 dcnt_h_reg_3_ ( .D(N141), .SIN(dcnt_h[2]), .SMC(test_se), .C(
        net10772), .Q(dcnt_h[3]) );
  SDFFQX1 dcnt_h_reg_4_ ( .D(N142), .SIN(dcnt_h[3]), .SMC(test_se), .C(
        net10772), .Q(dcnt_h[4]) );
  SDFFQX1 dcnt_h_reg_5_ ( .D(N143), .SIN(dcnt_h[4]), .SMC(test_se), .C(
        net10772), .Q(dcnt_h[5]) );
  SDFFQX1 dcnt_h_reg_1_ ( .D(N139), .SIN(dcnt_h[0]), .SMC(test_se), .C(
        net10772), .Q(dcnt_h[1]) );
  SDFFQX1 dcnt_h_reg_2_ ( .D(N140), .SIN(dcnt_h[1]), .SMC(test_se), .C(
        net10772), .Q(dcnt_h[2]) );
  SDFFQX1 dcnt_h_reg_0_ ( .D(N138), .SIN(dcnt_e[5]), .SMC(test_se), .C(
        net10772), .Q(dcnt_h[0]) );
  SDFFQX1 dcnt_h_reg_7_ ( .D(N145), .SIN(dcnt_h[6]), .SMC(test_se), .C(
        net10772), .Q(dcnt_h[7]) );
  SDFFQX1 adp_n_reg_5_ ( .D(N55), .SIN(adp_val[4]), .SMC(test_se), .C(net10761), .Q(adp_val[5]) );
  SDFFQX1 adp_n_reg_3_ ( .D(N53), .SIN(adp_val[2]), .SMC(test_se), .C(net10761), .Q(adp_val[3]) );
  SDFFQX1 adp_n_reg_0_ ( .D(n139), .SIN(test_si), .SMC(test_se), .C(net10761), 
        .Q(adp_val[0]) );
  SDFFQX1 dcnt_n_reg_0_ ( .D(N170), .SIN(n4), .SMC(test_se), .C(net10777), .Q(
        dcnt_n_0_) );
  SDFFQX1 adp_n_reg_1_ ( .D(N51), .SIN(adp_val[0]), .SMC(test_se), .C(net10761), .Q(adp_val[1]) );
  SDFFQX1 dcnt_n_reg_1_ ( .D(N171), .SIN(dcnt_n_0_), .SMC(test_se), .C(
        net10777), .Q(dcnt_n_1_) );
  SDFFQX1 adp_n_reg_2_ ( .D(N52), .SIN(adp_val[1]), .SMC(test_se), .C(net10761), .Q(adp_val[2]) );
  SDFFQX1 dcnt_n_reg_3_ ( .D(N173), .SIN(dcnt_n_2_), .SMC(test_se), .C(
        net10777), .Q(test_so) );
  SDFFQX1 adp_n_reg_4_ ( .D(n113), .SIN(adp_val[3]), .SMC(test_se), .C(
        net10761), .Q(adp_val[4]) );
  SDFFQX1 dcnt_n_reg_2_ ( .D(N172), .SIN(dcnt_n_1_), .SMC(test_se), .C(
        net10777), .Q(dcnt_n_2_) );
  SDFFQX1 dcnt_e_reg_5_ ( .D(N136), .SIN(dcnt_e[4]), .SMC(test_se), .C(
        net10767), .Q(dcnt_e[5]) );
  SDFFQX1 dcnt_e_reg_1_ ( .D(N132), .SIN(dcnt_e[0]), .SMC(test_se), .C(
        net10767), .Q(dcnt_e[1]) );
  SDFFQX1 dcnt_e_reg_4_ ( .D(N135), .SIN(dcnt_e[3]), .SMC(test_se), .C(
        net10767), .Q(dcnt_e[4]) );
  SDFFQX1 dcnt_e_reg_2_ ( .D(N133), .SIN(dcnt_e[1]), .SMC(test_se), .C(
        net10767), .Q(dcnt_e[2]) );
  SDFFQX1 dcnt_e_reg_3_ ( .D(N134), .SIN(dcnt_e[2]), .SMC(test_se), .C(
        net10767), .Q(dcnt_e[3]) );
  SDFFQX1 dcnt_e_reg_0_ ( .D(N131), .SIN(d_cc), .SMC(test_se), .C(net10767), 
        .Q(dcnt_e[0]) );
  SDFFQX1 cs_d_cc_reg ( .D(n115), .SIN(adp_val[5]), .SMC(test_se), .C(clk), 
        .Q(d_cc) );
  NAND2X1 U5 ( .A(n6), .B(n26), .Y(n136) );
  INVX1 U6 ( .A(dcnt_h[7]), .Y(n3) );
  INVX1 U7 ( .A(n3), .Y(n4) );
  INVX3 U8 ( .A(gohi), .Y(n22) );
  OR3XL U9 ( .A(n27), .B(n121), .C(n125), .Y(n6) );
  OR3XL U10 ( .A(dcnt_e[3]), .B(dcnt_e[2]), .C(dcnt_e[1]), .Y(n58) );
  INVX1 U11 ( .A(dcnt_e[0]), .Y(n101) );
  NAND21XL U12 ( .B(n12), .A(n104), .Y(n120) );
  NAND32XL U13 ( .B(n128), .C(n77), .A(n130), .Y(n78) );
  NAND32XL U14 ( .B(n128), .C(n75), .A(n77), .Y(n74) );
  NAND32XL U15 ( .B(n17), .C(n101), .A(n127), .Y(n30) );
  NAND2X1 U16 ( .A(n137), .B(n21), .Y(n125) );
  XOR2XL U17 ( .A(test_so), .B(adp_val[3]), .Y(n15) );
  NAND42X1 U18 ( .C(n16), .D(n15), .A(n5), .B(n14), .Y(n121) );
  XNOR2XL U19 ( .A(dcnt_n_0_), .B(adp_val[0]), .Y(n5) );
  NAND21XL U20 ( .B(n62), .A(dcnt_e[2]), .Y(n135) );
  NAND21XL U21 ( .B(n101), .A(dcnt_e[1]), .Y(n62) );
  INVXL U22 ( .A(adp_val[4]), .Y(n23) );
  NOR32XL U23 ( .B(n10), .C(n135), .A(dcnt_e[3]), .Y(n64) );
  AND3XL U24 ( .A(dcnt_e[0]), .B(n127), .C(n126), .Y(n129) );
  MUX2XL U25 ( .D0(n112), .D1(golo), .S(d_cc), .Y(n56) );
  OAI22XL U26 ( .A(n120), .B(n124), .C(dcnt_n_0_), .D(n123), .Y(N170) );
  INVXL U27 ( .A(test_so), .Y(n114) );
  MUX2XL U28 ( .D0(n112), .D1(golo), .S(adp_val[4]), .Y(n116) );
  NAND31X1 U29 ( .C(n120), .A(n121), .B(n106), .Y(n123) );
  OR2XL U30 ( .A(dcnt_e[5]), .B(n30), .Y(n60) );
  NAND21XL U31 ( .B(dcnt_e[5]), .A(n18), .Y(n131) );
  XOR2XL U32 ( .A(test_so), .B(n107), .Y(n108) );
  INVXL U33 ( .A(dcnt_e[5]), .Y(n73) );
  NAND21XL U34 ( .B(dcnt_e[1]), .A(n101), .Y(n32) );
  NAND21XL U35 ( .B(dcnt_e[3]), .A(n34), .Y(n51) );
  OR2XL U36 ( .A(dcnt_e[2]), .B(n32), .Y(n48) );
  NAND21XL U37 ( .B(dcnt_e[4]), .A(n49), .Y(n50) );
  NAND21XL U38 ( .B(n105), .A(dcnt_n_0_), .Y(n109) );
  INVXL U39 ( .A(dcnt_n_2_), .Y(n117) );
  NAND21XL U40 ( .B(dcnt_n_0_), .A(n105), .Y(n110) );
  INVXL U41 ( .A(dcnt_n_1_), .Y(n105) );
  NAND21XL U42 ( .B(n109), .A(dcnt_n_2_), .Y(n103) );
  INVX1 U43 ( .A(srstz), .Y(n12) );
  OR2X1 U44 ( .A(n89), .B(n88), .Y(n95) );
  INVX1 U45 ( .A(n76), .Y(n128) );
  NAND21X1 U46 ( .B(n99), .A(n140), .Y(n88) );
  NAND21X1 U47 ( .B(n96), .A(n95), .Y(n39) );
  MUX2X1 U48 ( .D0(n94), .D1(n91), .S(n90), .Y(n96) );
  INVX1 U49 ( .A(n93), .Y(n90) );
  AND2X1 U50 ( .A(n89), .B(n88), .Y(n94) );
  INVX1 U51 ( .A(n41), .Y(n99) );
  INVX1 U52 ( .A(n91), .Y(n89) );
  OAI31XL U53 ( .A(n93), .B(n140), .C(n41), .D(n39), .Y(n92) );
  INVX1 U54 ( .A(n37), .Y(n38) );
  NAND21X1 U55 ( .B(n140), .A(n93), .Y(n98) );
  NOR3XL U56 ( .A(goidle), .B(gobusy), .C(n12), .Y(n76) );
  NAND21X1 U57 ( .B(n18), .A(n126), .Y(n137) );
  INVX1 U58 ( .A(n125), .Y(n104) );
  NAND21X1 U59 ( .B(adp_v0[5]), .A(adp_v0[4]), .Y(n42) );
  AO21X1 U60 ( .B(adp_v0[4]), .C(n42), .A(n38), .Y(n93) );
  AO21X1 U61 ( .B(n42), .C(n33), .A(n38), .Y(n41) );
  INVX1 U62 ( .A(adp_v0[1]), .Y(n33) );
  AO21X1 U63 ( .B(n42), .C(n40), .A(n38), .Y(n91) );
  INVX1 U64 ( .A(adp_v0[2]), .Y(n40) );
  OAI21BBX1 U65 ( .A(n7), .B(adp_v0[4]), .C(adp_v0[5]), .Y(n37) );
  OR3XL U66 ( .A(adp_v0[1]), .B(adp_v0[3]), .C(adp_v0[2]), .Y(n7) );
  INVX1 U67 ( .A(n35), .Y(n140) );
  NAND32X1 U68 ( .B(n38), .C(adp_v0[0]), .A(n42), .Y(n35) );
  XOR2X1 U69 ( .A(n44), .B(n43), .Y(n87) );
  AO21X1 U70 ( .B(adp_v0[3]), .C(n37), .A(n36), .Y(n44) );
  AND2X1 U71 ( .A(n95), .B(n93), .Y(n43) );
  INVX1 U72 ( .A(n42), .Y(n36) );
  MUX2IX1 U73 ( .D0(n8), .D1(n9), .S(n99), .Y(N51) );
  NAND2X1 U74 ( .A(n139), .B(n93), .Y(n8) );
  NAND2X1 U75 ( .A(n134), .B(n98), .Y(n9) );
  AND2X1 U76 ( .A(n134), .B(n87), .Y(N53) );
  NOR21XL U77 ( .B(n134), .A(n39), .Y(N52) );
  INVX1 U78 ( .A(n97), .Y(n139) );
  NAND21X1 U79 ( .B(n140), .A(n134), .Y(n97) );
  AND2X1 U80 ( .A(n134), .B(n93), .Y(n113) );
  NAND2X1 U81 ( .A(n132), .B(n61), .Y(n133) );
  INVX1 U82 ( .A(n100), .Y(n52) );
  INVX1 U83 ( .A(n53), .Y(n102) );
  AOI21BX1 U84 ( .C(n60), .B(n61), .A(k0_det), .Y(n10) );
  AO21X1 U85 ( .B(n102), .C(n101), .A(n100), .Y(N131) );
  OR2X1 U86 ( .A(n100), .B(n11), .Y(N132) );
  AOI21X1 U87 ( .B(n32), .C(n62), .A(n53), .Y(n11) );
  INVX1 U88 ( .A(n78), .Y(n86) );
  INVX1 U89 ( .A(n74), .Y(n85) );
  OAI31XL U90 ( .A(n54), .B(n73), .C(n53), .D(n52), .Y(N136) );
  INVX1 U91 ( .A(n75), .Y(n130) );
  OAI2B11X1 U92 ( .D(n131), .C(n133), .A(n76), .B(n132), .Y(N130) );
  INVX1 U93 ( .A(n59), .Y(n61) );
  INVX1 U94 ( .A(n146), .Y(n112) );
  NAND21X1 U95 ( .B(n134), .A(srstz), .Y(N49) );
  AND2X1 U96 ( .A(n134), .B(n73), .Y(N55) );
  OAI211X1 U97 ( .C(n125), .D(n124), .A(n123), .B(n122), .Y(N169) );
  AND2X1 U98 ( .A(n121), .B(srstz), .Y(n122) );
  AND3X1 U99 ( .A(n111), .B(n110), .C(n109), .Y(N171) );
  INVX1 U100 ( .A(n123), .Y(n111) );
  AOI211X1 U101 ( .C(n109), .D(n117), .A(n107), .B(n123), .Y(N172) );
  INVX1 U102 ( .A(n58), .Y(n127) );
  INVX1 U103 ( .A(n69), .Y(n144) );
  INVX1 U104 ( .A(n67), .Y(n143) );
  INVX1 U105 ( .A(n71), .Y(n141) );
  INVX1 U106 ( .A(n65), .Y(n142) );
  INVX1 U107 ( .A(n110), .Y(n119) );
  INVX1 U108 ( .A(n51), .Y(n49) );
  INVX1 U109 ( .A(n48), .Y(n34) );
  NOR32XL U110 ( .B(dcnt_e[4]), .C(dcnt_e[3]), .A(n135), .Y(n138) );
  OAI21BBX1 U111 ( .A(adp_val[4]), .B(n104), .C(golo), .Y(n24) );
  INVX1 U112 ( .A(n118), .Y(n27) );
  AO21X1 U113 ( .B(n104), .C(n23), .A(n22), .Y(n25) );
  NAND42X1 U114 ( .C(adp_val[3]), .D(adp_val[0]), .A(n20), .B(n19), .Y(n21) );
  INVX1 U115 ( .A(adp_val[2]), .Y(n19) );
  INVX1 U116 ( .A(n13), .Y(n18) );
  NAND32X1 U117 ( .B(dcnt_e[4]), .C(n58), .A(n101), .Y(n13) );
  XOR2X1 U118 ( .A(n17), .B(dcnt_e[5]), .Y(n126) );
  INVX1 U119 ( .A(dcnt_e[4]), .Y(n17) );
  XOR2X1 U120 ( .A(n20), .B(dcnt_n_1_), .Y(n14) );
  XOR2X1 U121 ( .A(dcnt_n_2_), .B(adp_val[2]), .Y(n16) );
  XOR2X1 U122 ( .A(n77), .B(adp_val[4]), .Y(n118) );
  INVX1 U123 ( .A(d_cc), .Y(n77) );
  INVX1 U124 ( .A(adp_val[1]), .Y(n20) );
  GEN2XL U125 ( .D(dcnt_e[3]), .E(n48), .C(n49), .B(n102), .A(n47), .Y(N134)
         );
  OAI31XL U126 ( .A(n46), .B(n133), .C(n60), .D(n52), .Y(n47) );
  AOI211X1 U127 ( .C(n45), .D(n41), .A(n92), .B(n87), .Y(n46) );
  INVX1 U128 ( .A(n98), .Y(n45) );
  AO21X1 U129 ( .B(n102), .C(n31), .A(n128), .Y(n100) );
  INVX1 U130 ( .A(r_adprx_en), .Y(n31) );
  OAI211X1 U131 ( .C(r_adp2nd), .D(n30), .A(n131), .B(n29), .Y(n53) );
  AND2X1 U132 ( .A(n28), .B(n60), .Y(n29) );
  INVX1 U133 ( .A(n133), .Y(n28) );
  NAND2X1 U134 ( .A(r_adprx_en), .B(k0_det), .Y(n132) );
  OAI211X1 U135 ( .C(dcnt_e[4]), .D(n73), .A(n72), .B(n64), .Y(n75) );
  AO21X1 U136 ( .B(dcnt_e[0]), .C(n59), .A(n58), .Y(n72) );
  GEN2XL U137 ( .D(n142), .E(dcnt_h[6]), .C(n63), .B(n85), .A(n79), .Y(N144)
         );
  AND2X1 U138 ( .A(N103), .B(n86), .Y(n79) );
  GEN2XL U139 ( .D(dcnt_h[1]), .E(dcnt_h[0]), .C(n82), .B(n85), .A(n81), .Y(
        N139) );
  INVX1 U140 ( .A(n145), .Y(n82) );
  AND2X1 U141 ( .A(N98), .B(n86), .Y(n81) );
  GEN2XL U142 ( .D(dcnt_e[4]), .E(n51), .C(n54), .B(n102), .A(n100), .Y(N135)
         );
  GEN2XL U143 ( .D(dcnt_e[2]), .E(n32), .C(n34), .B(n102), .A(n100), .Y(N133)
         );
  GEN2XL U144 ( .D(dcnt_h[2]), .E(n145), .C(n71), .B(n85), .A(n83), .Y(N140)
         );
  AND2X1 U145 ( .A(N99), .B(n86), .Y(n83) );
  AO22AXL U146 ( .A(N102), .B(n86), .C(n85), .D(n66), .Y(N143) );
  AOI21X1 U147 ( .B(dcnt_h[5]), .C(n143), .A(n65), .Y(n66) );
  AO22AXL U148 ( .A(N101), .B(n86), .C(n85), .D(n68), .Y(N142) );
  AOI21X1 U149 ( .B(dcnt_h[4]), .C(n144), .A(n67), .Y(n68) );
  AO22AXL U150 ( .A(N100), .B(n86), .C(n85), .D(n70), .Y(N141) );
  AOI21X1 U151 ( .B(dcnt_h[3]), .C(n141), .A(n69), .Y(n70) );
  AO22X1 U152 ( .A(N97), .B(n86), .C(n85), .D(n80), .Y(N138) );
  AO22X1 U153 ( .A(N104), .B(n86), .C(n85), .D(n84), .Y(N145) );
  XOR2X1 U154 ( .A(dcnt_h[7]), .B(n63), .Y(n84) );
  NAND43X1 U155 ( .B(n130), .C(n129), .D(n128), .A(n10), .Y(N137) );
  INVX1 U156 ( .A(n57), .Y(n134) );
  NAND5XL U157 ( .A(dcnt_e[0]), .B(srstz), .C(n127), .D(n126), .E(n56), .Y(n57) );
  NAND5XL U158 ( .A(n119), .B(n118), .C(n117), .D(n116), .E(n114), .Y(n124) );
  AND2X1 U159 ( .A(n55), .B(srstz), .Y(n115) );
  NAND31X1 U160 ( .C(test_so), .A(n117), .B(n119), .Y(n106) );
  AND2X1 U161 ( .A(n108), .B(n111), .Y(N173) );
  NAND21X1 U162 ( .B(dcnt_h[1]), .A(n80), .Y(n145) );
  NOR2X1 U163 ( .A(n141), .B(dcnt_h[3]), .Y(n69) );
  NOR2X1 U164 ( .A(n144), .B(dcnt_h[4]), .Y(n67) );
  NOR2X1 U165 ( .A(n143), .B(dcnt_h[5]), .Y(n65) );
  NOR2X1 U166 ( .A(n145), .B(dcnt_h[2]), .Y(n71) );
  INVX1 U167 ( .A(dcnt_h[0]), .Y(n80) );
  NOR2X1 U168 ( .A(n142), .B(dcnt_h[6]), .Y(n63) );
  INVX1 U169 ( .A(n103), .Y(n107) );
  INVX1 U170 ( .A(n50), .Y(n54) );
  NAND21XL U171 ( .B(i_ccidle), .A(n136), .Y(n59) );
  XOR2XL U172 ( .A(n136), .B(d_cc), .Y(n55) );
  MUX2X2 U173 ( .D0(n25), .D1(n24), .S(d_cc), .Y(n26) );
  INVXL U174 ( .A(gohi), .Y(n146) );
  OA21X1 U175 ( .B(n138), .C(n137), .A(n136), .Y(cctrans) );
endmodule


module phyrx_adp_DW_div_tc_6 ( a, b, quotient, remainder, divide_by_0 );
  input [8:0] a;
  input [3:0] b;
  output [8:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   u_div_SumTmp_1__0_, u_div_SumTmp_1__2_, u_div_SumTmp_2__0_,
         u_div_SumTmp_3__0_, u_div_SumTmp_4__0_, u_div_SumTmp_5__0_,
         u_div_CryTmp_0__2_, u_div_CryTmp_0__3_, u_div_CryTmp_0__4_,
         u_div_CryTmp_1__4_, u_div_CryTmp_2__4_, u_div_CryTmp_3__4_,
         u_div_CryTmp_4__4_, u_div_CryTmp_5__4_, u_div_PartRem_1__2_,
         u_div_PartRem_1__3_, u_div_PartRem_2__3_, u_div_PartRem_3__3_,
         u_div_PartRem_4__3_, u_div_PartRem_5__3_, u_div_PartRem_7__0_,
         u_div_PartRem_7__1_, n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12,
         n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32;
  wire   [5:1] u_div_QIncCry;
  wire   [5:0] u_div_QInv;
  wire   [6:1] u_div_AIncCry;
  wire   [6:0] u_div_AInv;

  HAD1X1 u_div_u_ha_AInc_6 ( .A(u_div_AInv[6]), .B(u_div_AIncCry[6]), .CO(
        u_div_PartRem_7__1_), .SO(u_div_PartRem_7__0_) );
  HAD1X1 u_div_u_ha_AInc_5 ( .A(u_div_AInv[5]), .B(u_div_AIncCry[5]), .CO(
        u_div_AIncCry[6]), .SO(u_div_SumTmp_5__0_) );
  HAD1X1 u_div_u_ha_AInc_4 ( .A(u_div_AInv[4]), .B(u_div_AIncCry[4]), .CO(
        u_div_AIncCry[5]), .SO(u_div_SumTmp_4__0_) );
  HAD1X1 u_div_u_ha_AInc_3 ( .A(u_div_AInv[3]), .B(u_div_AIncCry[3]), .CO(
        u_div_AIncCry[4]), .SO(u_div_SumTmp_3__0_) );
  HAD1X1 u_div_u_ha_AInc_2 ( .A(u_div_AInv[2]), .B(u_div_AIncCry[2]), .CO(
        u_div_AIncCry[3]), .SO(u_div_SumTmp_2__0_) );
  HAD1X1 u_div_u_ha_AInc_1 ( .A(u_div_AInv[1]), .B(u_div_AIncCry[1]), .CO(
        u_div_AIncCry[2]), .SO(u_div_SumTmp_1__0_) );
  HAD1X1 u_div_u_ha_QInc_4 ( .A(u_div_QInv[4]), .B(u_div_QIncCry[4]), .CO(
        u_div_QIncCry[5]), .SO(quotient[4]) );
  HAD1X1 u_div_u_ha_QInc_3 ( .A(u_div_QInv[3]), .B(u_div_QIncCry[3]), .CO(
        u_div_QIncCry[4]), .SO(quotient[3]) );
  HAD1X1 u_div_u_ha_QInc_2 ( .A(u_div_QInv[2]), .B(u_div_QIncCry[2]), .CO(
        u_div_QIncCry[3]), .SO(quotient[2]) );
  HAD1X1 u_div_u_ha_QInc_1 ( .A(u_div_QInv[1]), .B(u_div_QIncCry[1]), .CO(
        u_div_QIncCry[2]), .SO(quotient[1]) );
  HAD1X1 u_div_u_ha_QInc_0 ( .A(u_div_QInv[0]), .B(a[7]), .CO(u_div_QIncCry[1]), .SO(quotient[0]) );
  AND2X1 u_div_u_ha_AInc_0 ( .A(u_div_AInv[0]), .B(a[8]), .Y(u_div_AIncCry[1])
         );
  XOR2X1 u_div_u_ha_QInc_5 ( .A(u_div_QInv[5]), .B(u_div_QIncCry[5]), .Y(
        quotient[5]) );
  XOR2X1 U1 ( .A(n26), .B(n25), .Y(u_div_SumTmp_1__2_) );
  INVX1 U2 ( .A(n18), .Y(n28) );
  INVX1 U3 ( .A(n19), .Y(n27) );
  INVX1 U4 ( .A(n20), .Y(n25) );
  NAND21X1 U5 ( .B(u_div_PartRem_3__3_), .A(n2), .Y(u_div_CryTmp_2__4_) );
  MUX2IX1 U6 ( .D0(n18), .D1(n6), .S(u_div_CryTmp_3__4_), .Y(
        u_div_PartRem_3__3_) );
  NAND2X1 U7 ( .A(n27), .B(n12), .Y(n2) );
  XNOR2XL U8 ( .A(n11), .B(n28), .Y(n6) );
  MUX2AXL U9 ( .D0(n10), .D1(n10), .S(u_div_CryTmp_4__4_), .Y(n18) );
  MUX2AXL U10 ( .D0(n11), .D1(n11), .S(u_div_CryTmp_3__4_), .Y(n19) );
  NAND21X1 U11 ( .B(u_div_PartRem_4__3_), .A(n1), .Y(u_div_CryTmp_3__4_) );
  MUX2IX1 U12 ( .D0(n17), .D1(n5), .S(u_div_CryTmp_4__4_), .Y(
        u_div_PartRem_4__3_) );
  NAND2X1 U13 ( .A(n28), .B(n11), .Y(n1) );
  XNOR2XL U14 ( .A(n10), .B(n31), .Y(n5) );
  MUX2AXL U15 ( .D0(n12), .D1(n12), .S(u_div_CryTmp_2__4_), .Y(n20) );
  MUX2AXL U16 ( .D0(n21), .D1(n21), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__2_) );
  INVX1 U17 ( .A(n21), .Y(n26) );
  INVX1 U18 ( .A(u_div_CryTmp_0__3_), .Y(n23) );
  NOR21XL U19 ( .B(u_div_CryTmp_0__2_), .A(n24), .Y(u_div_CryTmp_0__3_) );
  MUX2IX1 U20 ( .D0(n32), .D1(n32), .S(u_div_CryTmp_1__4_), .Y(
        u_div_CryTmp_0__2_) );
  INVX1 U21 ( .A(u_div_PartRem_1__2_), .Y(n24) );
  INVX1 U22 ( .A(n17), .Y(n31) );
  NAND21X1 U23 ( .B(u_div_PartRem_2__3_), .A(n4), .Y(u_div_CryTmp_1__4_) );
  MUX2IX1 U24 ( .D0(n19), .D1(n7), .S(u_div_CryTmp_2__4_), .Y(
        u_div_PartRem_2__3_) );
  NAND2X1 U25 ( .A(n25), .B(n26), .Y(n4) );
  XNOR2XL U26 ( .A(n12), .B(n27), .Y(n7) );
  MUX2IX1 U27 ( .D0(u_div_SumTmp_2__0_), .D1(u_div_SumTmp_2__0_), .S(
        u_div_CryTmp_2__4_), .Y(n21) );
  MUX2AXL U28 ( .D0(u_div_PartRem_7__0_), .D1(u_div_PartRem_7__0_), .S(
        u_div_CryTmp_5__4_), .Y(n17) );
  AND2X1 U29 ( .A(u_div_PartRem_7__1_), .B(u_div_PartRem_7__0_), .Y(
        u_div_CryTmp_5__4_) );
  NAND21X1 U30 ( .B(u_div_PartRem_5__3_), .A(n3), .Y(u_div_CryTmp_4__4_) );
  MUX2IX1 U31 ( .D0(n29), .D1(n8), .S(u_div_CryTmp_5__4_), .Y(
        u_div_PartRem_5__3_) );
  NAND2X1 U32 ( .A(n31), .B(n10), .Y(n3) );
  INVX1 U33 ( .A(u_div_PartRem_7__1_), .Y(n29) );
  MUX2X1 U34 ( .D0(u_div_SumTmp_5__0_), .D1(u_div_SumTmp_5__0_), .S(
        u_div_CryTmp_5__4_), .Y(n10) );
  MUX2X1 U35 ( .D0(u_div_SumTmp_4__0_), .D1(u_div_SumTmp_4__0_), .S(
        u_div_CryTmp_4__4_), .Y(n11) );
  MUX2X1 U36 ( .D0(u_div_SumTmp_3__0_), .D1(u_div_SumTmp_3__0_), .S(
        u_div_CryTmp_3__4_), .Y(n12) );
  XNOR2XL U37 ( .A(u_div_PartRem_7__0_), .B(u_div_PartRem_7__1_), .Y(n8) );
  INVX1 U38 ( .A(u_div_SumTmp_1__0_), .Y(n32) );
  XOR2X1 U39 ( .A(a[7]), .B(u_div_CryTmp_4__4_), .Y(u_div_QInv[4]) );
  XOR2X1 U40 ( .A(a[8]), .B(a[6]), .Y(u_div_AInv[6]) );
  XNOR2XL U41 ( .A(a[7]), .B(n30), .Y(u_div_QInv[5]) );
  INVX1 U42 ( .A(u_div_CryTmp_5__4_), .Y(n30) );
  XOR2X1 U43 ( .A(a[7]), .B(u_div_CryTmp_0__4_), .Y(u_div_QInv[0]) );
  NAND21X1 U44 ( .B(u_div_PartRem_1__3_), .A(n23), .Y(u_div_CryTmp_0__4_) );
  MUX2AXL U45 ( .D0(n20), .D1(u_div_SumTmp_1__2_), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__3_) );
  XOR2X1 U46 ( .A(a[8]), .B(a[1]), .Y(u_div_AInv[1]) );
  XOR2X1 U47 ( .A(a[8]), .B(a[0]), .Y(u_div_AInv[0]) );
  XOR2X1 U48 ( .A(a[8]), .B(a[2]), .Y(u_div_AInv[2]) );
  XOR2X1 U49 ( .A(a[8]), .B(a[3]), .Y(u_div_AInv[3]) );
  XOR2X1 U50 ( .A(a[8]), .B(a[4]), .Y(u_div_AInv[4]) );
  XOR2X1 U51 ( .A(a[8]), .B(a[5]), .Y(u_div_AInv[5]) );
  XOR2X1 U52 ( .A(a[7]), .B(u_div_CryTmp_1__4_), .Y(u_div_QInv[1]) );
  XOR2X1 U53 ( .A(a[7]), .B(u_div_CryTmp_2__4_), .Y(u_div_QInv[2]) );
  XOR2X1 U54 ( .A(a[7]), .B(u_div_CryTmp_3__4_), .Y(u_div_QInv[3]) );
endmodule


module phyrx_adp_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_db ( clk, srstz, x_cc, ptx_txact, r_rxdb_opt, gohi, golo, gotrans, 
        test_si, test_so, test_se );
  input [1:0] r_rxdb_opt;
  input clk, srstz, x_cc, ptx_txact, test_si, test_se;
  output gohi, golo, gotrans, test_so;
  wire   cc_buf_6_, cc_buf_5_, cc_buf_4_, cc_buf_3_, cc_buf_2_, cc_buf_1_,
         cc_buf_0_, N11, N12, N13, N14, N15, N16, N17, N18, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48;

  SDFFQX1 cc_buf_reg_6_ ( .D(N17), .SIN(cc_buf_5_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_6_) );
  SDFFQX1 cc_buf_reg_3_ ( .D(N14), .SIN(cc_buf_2_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_3_) );
  SDFFQX1 cc_buf_reg_5_ ( .D(N16), .SIN(cc_buf_4_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_5_) );
  SDFFQX1 cc_buf_reg_7_ ( .D(N18), .SIN(cc_buf_6_), .SMC(test_se), .C(clk), 
        .Q(test_so) );
  SDFFQX1 cc_buf_reg_4_ ( .D(N15), .SIN(cc_buf_3_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_4_) );
  SDFFQX1 cc_buf_reg_2_ ( .D(N13), .SIN(cc_buf_1_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_2_) );
  SDFFQX1 cc_buf_reg_1_ ( .D(N12), .SIN(cc_buf_0_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_1_) );
  SDFFQX1 cc_buf_reg_0_ ( .D(N11), .SIN(test_si), .SMC(test_se), .C(clk), .Q(
        cc_buf_0_) );
  NAND2X1 U3 ( .A(n20), .B(n7), .Y(n8) );
  INVX1 U4 ( .A(cc_buf_6_), .Y(n22) );
  EORX1 U5 ( .A(cc_buf_2_), .B(n10), .C(n21), .D(n19), .Y(n14) );
  OA22X1 U6 ( .A(n31), .B(n34), .C(n30), .D(n33), .Y(n1) );
  NAND2X1 U7 ( .A(n12), .B(n13), .Y(n23) );
  INVX1 U8 ( .A(n23), .Y(n6) );
  INVX1 U9 ( .A(cc_buf_1_), .Y(n20) );
  AND2X2 U10 ( .A(n31), .B(n34), .Y(n30) );
  INVXL U11 ( .A(n29), .Y(n16) );
  NAND2X1 U12 ( .A(n23), .B(n2), .Y(n3) );
  NAND2X1 U13 ( .A(n3), .B(n4), .Y(n29) );
  NAND2X1 U14 ( .A(n6), .B(test_so), .Y(n4) );
  INVXL U15 ( .A(test_so), .Y(n2) );
  INVX2 U16 ( .A(n21), .Y(n11) );
  ENOX1 U17 ( .A(n29), .B(n22), .C(test_so), .D(n6), .Y(n5) );
  ENOXL U18 ( .A(n29), .B(n22), .C(test_so), .D(n6), .Y(n27) );
  NAND2X1 U19 ( .A(cc_buf_1_), .B(cc_buf_2_), .Y(n9) );
  NAND2X2 U20 ( .A(n8), .B(n9), .Y(n21) );
  INVX3 U21 ( .A(cc_buf_2_), .Y(n7) );
  INVXL U22 ( .A(n20), .Y(n10) );
  INVX1 U23 ( .A(cc_buf_4_), .Y(n26) );
  INVXL U24 ( .A(cc_buf_0_), .Y(n19) );
  INVX2 U25 ( .A(n35), .Y(n31) );
  NAND21XL U26 ( .B(n15), .A(n32), .Y(n38) );
  AND2XL U27 ( .A(n17), .B(n42), .Y(n18) );
  INVXL U28 ( .A(cc_buf_5_), .Y(n25) );
  INVXL U29 ( .A(cc_buf_3_), .Y(n24) );
  XOR2XL U30 ( .A(n28), .B(cc_buf_3_), .Y(n32) );
  INVXL U31 ( .A(n17), .Y(gotrans) );
  AND2XL U32 ( .A(srstz), .B(cc_buf_0_), .Y(N12) );
  AND2XL U33 ( .A(srstz), .B(cc_buf_4_), .Y(N16) );
  AND2XL U34 ( .A(srstz), .B(cc_buf_3_), .Y(N15) );
  AND2XL U35 ( .A(srstz), .B(cc_buf_6_), .Y(N18) );
  AND2XL U36 ( .A(srstz), .B(cc_buf_5_), .Y(N17) );
  NAND2X1 U37 ( .A(n21), .B(n19), .Y(n12) );
  NAND2X2 U38 ( .A(n11), .B(cc_buf_0_), .Y(n13) );
  NAND2X1 U39 ( .A(n46), .B(n1), .Y(n43) );
  AND2X1 U40 ( .A(x_cc), .B(srstz), .Y(N11) );
  NAND21X1 U41 ( .B(n32), .A(n15), .Y(n33) );
  XOR2X1 U42 ( .A(n5), .B(n14), .Y(n34) );
  XOR3X1 U43 ( .A(n37), .B(n36), .C(n35), .Y(n44) );
  INVXL U44 ( .A(n33), .Y(n37) );
  OAI21BBXL U45 ( .A(n19), .B(n20), .C(n42), .Y(n17) );
  MUX2IX1 U46 ( .D0(n41), .D1(n40), .S(r_rxdb_opt[1]), .Y(golo) );
  NAND21XL U47 ( .B(n43), .A(n39), .Y(n40) );
  OAI22X1 U48 ( .A(n26), .B(n25), .C(n28), .D(n24), .Y(n35) );
  XOR2X1 U49 ( .A(n26), .B(cc_buf_5_), .Y(n28) );
  XOR2X1 U50 ( .A(n16), .B(cc_buf_6_), .Y(n15) );
  AND2XL U51 ( .A(srstz), .B(cc_buf_2_), .Y(N14) );
  NAND31X1 U52 ( .C(n37), .A(n38), .B(n44), .Y(n39) );
  INVX1 U53 ( .A(n34), .Y(n36) );
  AND2X2 U54 ( .A(n44), .B(n43), .Y(n45) );
  NOR32XL U55 ( .B(srstz), .C(cc_buf_1_), .A(ptx_txact), .Y(N13) );
  NAND21XL U56 ( .B(n19), .A(cc_buf_1_), .Y(n42) );
  NAND31XL U57 ( .C(n42), .A(cc_buf_2_), .B(cc_buf_3_), .Y(n48) );
  NAND32XL U58 ( .B(cc_buf_3_), .C(cc_buf_2_), .A(n18), .Y(n41) );
  NAND21XL U59 ( .B(n14), .A(n27), .Y(n46) );
  AOI21BBX4 U60 ( .B(n1), .C(n46), .A(n45), .Y(n47) );
  MUX2IX4 U61 ( .D0(n48), .D1(n47), .S(r_rxdb_opt[0]), .Y(gohi) );
endmodule


module i2cslv_a0 ( i_sda, i_scl, o_sda, i_deva, i_inc, i_fwnak, i_fwack, o_we, 
        o_re, o_r_early, o_idle, o_dec, o_busev, o_ofs, o_lt_ofs, o_wdat, 
        o_lt_buf, o_dbgpo, i_rdat, i_rd_mem, i_clk, i_rstz, i_prefetch, 
        test_si, test_se );
  input [7:1] i_deva;
  output [3:0] o_busev;
  output [7:0] o_ofs;
  output [7:0] o_lt_ofs;
  output [7:0] o_wdat;
  output [7:0] o_lt_buf;
  output [7:0] o_dbgpo;
  input [7:0] i_rdat;
  input i_sda, i_scl, i_inc, i_fwnak, i_fwack, i_rd_mem, i_clk, i_rstz,
         i_prefetch, test_si, test_se;
  output o_sda, o_we, o_re, o_r_early, o_idle, o_dec;
  wire   i2c_scl, sdafall, cs_rwb, N74, N75, N76, N77, N78, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, ps_rwbuf_0_, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, net10794, net10800, net10805, net10810,
         net10815, n118, n119, n120, n121, n15, n16, n17, n18, n19, n64, n87,
         n88, n89, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178;
  wire   [1:0] cs_sta;

  INVX1 U5 ( .A(n19), .Y(n16) );
  INVX1 U6 ( .A(n19), .Y(n17) );
  INVX1 U7 ( .A(n19), .Y(n18) );
  INVX1 U9 ( .A(n19), .Y(n15) );
  INVX1 U10 ( .A(i_rstz), .Y(n19) );
  i2cdbnc_a0_1 db_scl ( .i_clk(i_clk), .i_rstz(n15), .i_i2c(i_scl), .r_opt({
        1'b1, 1'b0}), .o_i2c(i2c_scl), .rise(o_dbgpo[6]), .fall(o_dbgpo[7]), 
        .test_si(cs_sta[1]), .test_se(test_se) );
  i2cdbnc_a0_0 db_sda ( .i_clk(i_clk), .i_rstz(n15), .i_i2c(i_sda), .r_opt({
        1'b0, 1'b0}), .o_i2c(ps_rwbuf_0_), .rise(o_dbgpo[5]), .fall(sdafall), 
        .test_si(i2c_scl), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 clk_gate_cs_bit_reg ( .CLK(i_clk), .EN(N74), 
        .ENCLK(net10794), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 clk_gate_adcnt_reg ( .CLK(i_clk), .EN(N114), 
        .ENCLK(net10800), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 clk_gate_rwbuf_reg ( .CLK(i_clk), .EN(N144), 
        .ENCLK(net10805), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 clk_gate_lt_buf_reg ( .CLK(i_clk), .EN(N179), .ENCLK(net10810), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 clk_gate_lt_ofs_reg ( .CLK(i_clk), .EN(
        o_busev[2]), .ENCLK(net10815), .TE(test_se) );
  SDFFSQXL rwbuf_reg_3_ ( .D(N139), .SIN(o_wdat[2]), .SMC(test_se), .C(
        net10805), .XS(n16), .Q(o_wdat[3]) );
  SDFFSQXL rwbuf_reg_4_ ( .D(N140), .SIN(o_wdat[3]), .SMC(test_se), .C(
        net10805), .XS(n16), .Q(o_wdat[4]) );
  SDFFQX1 lt_ofs_reg_7_ ( .D(o_wdat[7]), .SIN(o_lt_ofs[6]), .SMC(test_se), .C(
        net10815), .Q(o_lt_ofs[7]) );
  SDFFQX1 lt_ofs_reg_6_ ( .D(o_wdat[6]), .SIN(o_lt_ofs[5]), .SMC(test_se), .C(
        net10815), .Q(o_lt_ofs[6]) );
  SDFFQX1 lt_ofs_reg_3_ ( .D(o_wdat[3]), .SIN(o_lt_ofs[2]), .SMC(test_se), .C(
        net10815), .Q(o_lt_ofs[3]) );
  SDFFQX1 lt_ofs_reg_0_ ( .D(o_wdat[0]), .SIN(o_lt_buf[7]), .SMC(test_se), .C(
        net10815), .Q(o_lt_ofs[0]) );
  SDFFQX1 lt_buf_reg_7_ ( .D(N187), .SIN(o_lt_buf[6]), .SMC(test_se), .C(
        net10810), .Q(o_lt_buf[7]) );
  SDFFQX1 lt_buf_reg_6_ ( .D(N186), .SIN(o_lt_buf[5]), .SMC(test_se), .C(
        net10810), .Q(o_lt_buf[6]) );
  SDFFQX1 lt_buf_reg_3_ ( .D(N183), .SIN(o_lt_buf[2]), .SMC(test_se), .C(
        net10810), .Q(o_lt_buf[3]) );
  SDFFQX1 lt_buf_reg_0_ ( .D(N180), .SIN(ps_rwbuf_0_), .SMC(test_se), .C(
        net10810), .Q(o_lt_buf[0]) );
  SDFFQX1 lt_ofs_reg_5_ ( .D(o_wdat[5]), .SIN(o_lt_ofs[4]), .SMC(test_se), .C(
        net10815), .Q(o_lt_ofs[5]) );
  SDFFQX1 lt_ofs_reg_4_ ( .D(o_wdat[4]), .SIN(o_lt_ofs[3]), .SMC(test_se), .C(
        net10815), .Q(o_lt_ofs[4]) );
  SDFFQX1 lt_ofs_reg_2_ ( .D(o_wdat[2]), .SIN(o_lt_ofs[1]), .SMC(test_se), .C(
        net10815), .Q(o_lt_ofs[2]) );
  SDFFQX1 lt_ofs_reg_1_ ( .D(o_wdat[1]), .SIN(o_lt_ofs[0]), .SMC(test_se), .C(
        net10815), .Q(o_lt_ofs[1]) );
  SDFFQX1 lt_buf_reg_5_ ( .D(N185), .SIN(o_lt_buf[4]), .SMC(test_se), .C(
        net10810), .Q(o_lt_buf[5]) );
  SDFFQX1 lt_buf_reg_4_ ( .D(N184), .SIN(o_lt_buf[3]), .SMC(test_se), .C(
        net10810), .Q(o_lt_buf[4]) );
  SDFFQX1 lt_buf_reg_2_ ( .D(N182), .SIN(o_lt_buf[1]), .SMC(test_se), .C(
        net10810), .Q(o_lt_buf[2]) );
  SDFFQX1 lt_buf_reg_1_ ( .D(N181), .SIN(o_lt_buf[0]), .SMC(test_se), .C(
        net10810), .Q(o_lt_buf[1]) );
  SDFFRQX1 adcnt_reg_6_ ( .D(N112), .SIN(o_ofs[5]), .SMC(test_se), .C(net10800), .XR(n18), .Q(o_ofs[6]) );
  SDFFRQX1 adcnt_reg_1_ ( .D(N107), .SIN(o_ofs[0]), .SMC(test_se), .C(net10800), .XR(n17), .Q(o_ofs[1]) );
  SDFFRQX1 adcnt_reg_5_ ( .D(N111), .SIN(o_ofs[4]), .SMC(test_se), .C(net10800), .XR(n17), .Q(o_ofs[5]) );
  SDFFRQX1 adcnt_reg_3_ ( .D(N109), .SIN(o_ofs[2]), .SMC(test_se), .C(net10800), .XR(n17), .Q(o_ofs[3]) );
  SDFFRQX1 adcnt_reg_2_ ( .D(N108), .SIN(o_ofs[1]), .SMC(test_se), .C(net10800), .XR(n17), .Q(o_ofs[2]) );
  SDFFRQX1 adcnt_reg_0_ ( .D(N106), .SIN(test_si), .SMC(test_se), .C(net10800), 
        .XR(n17), .Q(o_ofs[0]) );
  SDFFRQX1 adcnt_reg_4_ ( .D(N110), .SIN(o_ofs[3]), .SMC(test_se), .C(net10800), .XR(n17), .Q(o_ofs[4]) );
  SDFFRQX1 adcnt_reg_7_ ( .D(N113), .SIN(o_ofs[6]), .SMC(test_se), .C(net10800), .XR(n17), .Q(o_ofs[7]) );
  SDFFSQX1 sdat_reg ( .D(n118), .SIN(o_wdat[7]), .SMC(test_se), .C(i_clk), 
        .XS(n16), .Q(o_sda) );
  SDFFRQX1 cs_rwb_reg ( .D(n119), .SIN(o_dbgpo[3]), .SMC(test_se), .C(i_clk), 
        .XR(n17), .Q(cs_rwb) );
  SDFFSQX1 rwbuf_reg_6_ ( .D(N142), .SIN(o_wdat[5]), .SMC(test_se), .C(
        net10805), .XS(n16), .Q(o_wdat[6]) );
  SDFFSQX1 cs_bit_reg_0_ ( .D(N75), .SIN(o_ofs[7]), .SMC(test_se), .C(net10794), .XS(n16), .Q(o_dbgpo[0]) );
  SDFFSQX1 rwbuf_reg_7_ ( .D(N143), .SIN(o_wdat[6]), .SMC(test_se), .C(
        net10805), .XS(n15), .Q(o_wdat[7]) );
  SDFFRQX1 cs_sta_reg_1_ ( .D(n121), .SIN(cs_sta[0]), .SMC(test_se), .C(i_clk), 
        .XR(n18), .Q(cs_sta[1]) );
  SDFFSQX1 cs_bit_reg_2_ ( .D(N77), .SIN(o_dbgpo[1]), .SMC(test_se), .C(
        net10794), .XS(n16), .Q(o_dbgpo[2]) );
  SDFFSQX1 cs_bit_reg_3_ ( .D(N78), .SIN(o_dbgpo[2]), .SMC(test_se), .C(
        net10794), .XS(n16), .Q(o_dbgpo[3]) );
  SDFFSQX1 rwbuf_reg_1_ ( .D(N137), .SIN(o_wdat[0]), .SMC(test_se), .C(
        net10805), .XS(n17), .Q(o_wdat[1]) );
  SDFFSQX1 rwbuf_reg_0_ ( .D(N136), .SIN(o_lt_ofs[7]), .SMC(test_se), .C(
        net10805), .XS(n15), .Q(o_wdat[0]) );
  SDFFSQX1 rwbuf_reg_2_ ( .D(N138), .SIN(o_wdat[1]), .SMC(test_se), .C(
        net10805), .XS(n16), .Q(o_wdat[2]) );
  SDFFSQX1 rwbuf_reg_5_ ( .D(N141), .SIN(o_wdat[4]), .SMC(test_se), .C(
        net10805), .XS(n16), .Q(o_wdat[5]) );
  SDFFSQX1 cs_bit_reg_1_ ( .D(N76), .SIN(o_dbgpo[0]), .SMC(test_se), .C(
        net10794), .XS(n16), .Q(o_dbgpo[1]) );
  SDFFRQX1 cs_sta_reg_0_ ( .D(n120), .SIN(cs_rwb), .SMC(test_se), .C(i_clk), 
        .XR(n17), .Q(cs_sta[0]) );
  AO21X1 U3 ( .B(n125), .C(o_wdat[7]), .A(n74), .Y(N113) );
  INVX1 U4 ( .A(n58), .Y(n1) );
  INVX1 U8 ( .A(n137), .Y(o_busev[2]) );
  INVX1 U11 ( .A(n153), .Y(n139) );
  NAND2X1 U12 ( .A(n175), .B(n178), .Y(N74) );
  INVX1 U13 ( .A(n35), .Y(n128) );
  NAND21X1 U14 ( .B(n176), .A(n160), .Y(n126) );
  INVX1 U15 ( .A(o_dbgpo[7]), .Y(n176) );
  INVX1 U16 ( .A(n142), .Y(o_idle) );
  INVX1 U17 ( .A(n37), .Y(n131) );
  NAND21X1 U18 ( .B(n126), .A(n125), .Y(n137) );
  NAND21X1 U19 ( .B(n176), .A(n140), .Y(n153) );
  AND2X1 U20 ( .A(n160), .B(n154), .Y(n155) );
  INVX1 U21 ( .A(n115), .Y(n175) );
  NAND32X1 U22 ( .B(n176), .C(n168), .A(n142), .Y(n178) );
  INVX1 U23 ( .A(n75), .Y(n14) );
  BUFX3 U24 ( .A(o_busev[3]), .Y(o_dbgpo[4]) );
  NAND5XL U25 ( .A(o_busev[1]), .B(n86), .C(n84), .D(n90), .E(n30), .Y(n35) );
  AND4X1 U26 ( .A(n81), .B(n85), .C(n83), .D(n82), .Y(n30) );
  INVX1 U27 ( .A(o_dbgpo[6]), .Y(n105) );
  INVX1 U28 ( .A(n22), .Y(o_busev[1]) );
  NAND32X1 U29 ( .B(n163), .C(n105), .A(n140), .Y(n22) );
  INVX1 U30 ( .A(n104), .Y(n140) );
  AND3X1 U31 ( .A(n145), .B(o_dec), .C(n150), .Y(n147) );
  INVX1 U32 ( .A(n141), .Y(o_dec) );
  INVX1 U33 ( .A(n143), .Y(n145) );
  NAND21X1 U34 ( .B(n162), .A(n140), .Y(n141) );
  AND3X1 U35 ( .A(n152), .B(n151), .C(n150), .Y(o_re) );
  MUX2X1 U36 ( .D0(n147), .D1(n146), .S(i_prefetch), .Y(o_r_early) );
  MUX2X1 U37 ( .D0(n149), .D1(n160), .S(i_prefetch), .Y(n151) );
  INVX1 U38 ( .A(n36), .Y(n146) );
  NAND21X1 U39 ( .B(n161), .A(n128), .Y(n36) );
  INVX1 U40 ( .A(n163), .Y(n160) );
  INVX1 U41 ( .A(n162), .Y(n148) );
  INVX1 U42 ( .A(n144), .Y(n150) );
  NAND21X1 U43 ( .B(n164), .A(o_dbgpo[6]), .Y(n144) );
  INVX1 U44 ( .A(n21), .Y(n25) );
  AND2X1 U45 ( .A(n148), .B(n161), .Y(n149) );
  INVX1 U46 ( .A(n127), .Y(o_we) );
  INVX1 U47 ( .A(n58), .Y(n152) );
  OR3XL U48 ( .A(n133), .B(n28), .C(n77), .Y(n142) );
  INVX1 U49 ( .A(i_rdat[7]), .Y(n174) );
  INVX1 U50 ( .A(n87), .Y(n170) );
  EORX1 U51 ( .A(i_fwnak), .B(n88), .C(n89), .D(i_fwack), .Y(n87) );
  NAND2X1 U52 ( .A(i_fwack), .B(n89), .Y(n88) );
  NAND21X1 U53 ( .B(n172), .A(n171), .Y(n118) );
  NOR32XL U54 ( .B(n139), .C(n156), .A(n155), .Y(n172) );
  MUX2IX1 U55 ( .D0(n170), .D1(n169), .S(o_dbgpo[7]), .Y(n171) );
  INVX1 U56 ( .A(i_rd_mem), .Y(n177) );
  OAI22AX1 U57 ( .D(n130), .C(n174), .A(n97), .B(n37), .Y(N143) );
  NAND32X1 U58 ( .B(n105), .C(n130), .A(n162), .Y(n37) );
  OA21X1 U59 ( .B(n131), .C(n130), .A(n129), .Y(N144) );
  OR4X1 U60 ( .A(o_dbgpo[7]), .B(n105), .C(n104), .D(n154), .Y(n108) );
  NAND21X1 U61 ( .B(i_prefetch), .A(n143), .Y(n154) );
  AO21X1 U62 ( .B(n152), .C(n70), .A(n69), .Y(n72) );
  AO21X1 U63 ( .B(n152), .C(n67), .A(n140), .Y(n69) );
  INVX1 U64 ( .A(n112), .Y(n123) );
  GEN2XL U65 ( .D(o_dbgpo[7]), .E(n111), .C(n110), .B(n148), .A(n109), .Y(n112) );
  NAND21X1 U66 ( .B(n139), .A(n175), .Y(n109) );
  INVX1 U67 ( .A(n108), .Y(n110) );
  INVX1 U68 ( .A(n23), .Y(o_busev[0]) );
  INVX1 U69 ( .A(n64), .Y(o_busev[3]) );
  INVX1 U70 ( .A(n47), .Y(n54) );
  NAND21X1 U71 ( .B(o_busev[0]), .A(n64), .Y(n115) );
  AO21X1 U72 ( .B(n152), .C(n55), .A(n50), .Y(n53) );
  AND4X1 U73 ( .A(n90), .B(n86), .C(n85), .D(n84), .Y(n91) );
  AO21X1 U74 ( .B(n152), .C(n47), .A(n140), .Y(n50) );
  INVX1 U75 ( .A(n57), .Y(n125) );
  INVX1 U76 ( .A(n82), .Y(n93) );
  INVX1 U77 ( .A(n83), .Y(n92) );
  AO21X1 U78 ( .B(n152), .C(n38), .A(n140), .Y(n41) );
  INVX1 U79 ( .A(i_inc), .Y(n38) );
  NAND21X1 U80 ( .B(n178), .A(n162), .Y(n75) );
  AO21X1 U81 ( .B(n14), .C(n79), .A(n115), .Y(N75) );
  NAND21X1 U82 ( .B(n128), .A(n127), .Y(N179) );
  OR2X1 U83 ( .A(n78), .B(n2), .Y(N76) );
  AOI21X1 U84 ( .B(n77), .C(n76), .A(n75), .Y(n2) );
  OAI22X1 U85 ( .A(n164), .B(n163), .C(n162), .D(n161), .Y(n165) );
  INVX1 U86 ( .A(n129), .Y(n168) );
  OAI22X1 U87 ( .A(n127), .B(n43), .C(n35), .D(n34), .Y(N181) );
  OAI22X1 U88 ( .A(n127), .B(n33), .C(n35), .D(n43), .Y(N182) );
  OAI22X1 U89 ( .A(n127), .B(n32), .C(n35), .D(n33), .Y(N183) );
  OAI22X1 U90 ( .A(n127), .B(n56), .C(n35), .D(n32), .Y(N184) );
  OAI22X1 U91 ( .A(n127), .B(n31), .C(n35), .D(n56), .Y(N185) );
  OAI22X1 U92 ( .A(n127), .B(n97), .C(n35), .D(n31), .Y(N186) );
  OAI22X1 U93 ( .A(n96), .B(n127), .C(n35), .D(n97), .Y(N187) );
  INVX1 U94 ( .A(n68), .Y(n71) );
  NAND32X1 U95 ( .B(n67), .C(n70), .A(n152), .Y(n68) );
  INVX1 U96 ( .A(n13), .Y(n78) );
  NAND21X1 U97 ( .B(n64), .A(n23), .Y(n13) );
  NAND4X1 U98 ( .A(n3), .B(n4), .C(n5), .D(n103), .Y(n143) );
  XNOR2XL U99 ( .A(i_deva[1]), .B(o_wdat[1]), .Y(n3) );
  XNOR2XL U100 ( .A(i_deva[3]), .B(o_wdat[3]), .Y(n4) );
  XNOR2XL U101 ( .A(o_wdat[2]), .B(i_deva[2]), .Y(n5) );
  NAND43X1 U102 ( .B(o_dbgpo[2]), .C(o_dbgpo[1]), .D(o_dbgpo[3]), .A(
        o_dbgpo[0]), .Y(n163) );
  XOR2X1 U103 ( .A(n33), .B(i_deva[3]), .Y(n82) );
  XOR2X1 U104 ( .A(n31), .B(i_deva[6]), .Y(n83) );
  XOR2X1 U105 ( .A(n34), .B(i_deva[1]), .Y(n81) );
  NAND21X1 U106 ( .B(cs_sta[0]), .A(n111), .Y(n104) );
  INVX1 U107 ( .A(o_wdat[4]), .Y(n56) );
  INVX1 U108 ( .A(o_wdat[3]), .Y(n32) );
  XNOR2XL U109 ( .A(i_deva[4]), .B(o_wdat[4]), .Y(n98) );
  NOR32XL U110 ( .B(n102), .C(n101), .A(n100), .Y(n103) );
  XOR2X1 U111 ( .A(n96), .B(i_deva[7]), .Y(n102) );
  XOR2X1 U112 ( .A(n97), .B(i_deva[6]), .Y(n101) );
  NAND21X1 U113 ( .B(n99), .A(n98), .Y(n100) );
  XOR2X1 U114 ( .A(n56), .B(i_deva[5]), .Y(n84) );
  XOR2X1 U115 ( .A(n32), .B(i_deva[4]), .Y(n90) );
  XOR2X1 U116 ( .A(n43), .B(i_deva[2]), .Y(n85) );
  INVX1 U117 ( .A(o_wdat[1]), .Y(n43) );
  INVX1 U118 ( .A(o_wdat[5]), .Y(n31) );
  INVX1 U119 ( .A(o_wdat[2]), .Y(n33) );
  INVX1 U120 ( .A(o_wdat[0]), .Y(n34) );
  NAND21X1 U121 ( .B(o_dbgpo[3]), .A(n25), .Y(n162) );
  NAND21X1 U122 ( .B(o_dbgpo[1]), .A(n79), .Y(n76) );
  OR2X1 U123 ( .A(o_dbgpo[2]), .B(n76), .Y(n21) );
  XOR2X1 U124 ( .A(n97), .B(i_deva[7]), .Y(n86) );
  XOR2X1 U125 ( .A(i_deva[5]), .B(o_wdat[5]), .Y(n99) );
  INVX1 U126 ( .A(cs_sta[1]), .Y(n111) );
  INVX1 U127 ( .A(o_dbgpo[0]), .Y(n79) );
  INVX1 U128 ( .A(o_wdat[6]), .Y(n97) );
  INVX1 U129 ( .A(o_wdat[7]), .Y(n96) );
  OR3XL U130 ( .A(cs_rwb), .B(n58), .C(n126), .Y(n127) );
  NAND21X1 U131 ( .B(cs_sta[0]), .A(cs_sta[1]), .Y(n58) );
  INVX1 U132 ( .A(cs_rwb), .Y(n164) );
  INVX1 U133 ( .A(ps_rwbuf_0_), .Y(n161) );
  NAND21X1 U134 ( .B(n79), .A(o_dbgpo[1]), .Y(n77) );
  INVX1 U135 ( .A(o_dbgpo[3]), .Y(n133) );
  INVX1 U136 ( .A(o_dbgpo[2]), .Y(n28) );
  MUX2AXL U137 ( .D0(o_sda), .D1(n174), .S(n173), .Y(n89) );
  NAND42X1 U138 ( .C(cs_sta[0]), .D(n164), .A(n158), .B(n157), .Y(n159) );
  NAND21X1 U139 ( .B(i_rd_mem), .A(o_wdat[7]), .Y(n157) );
  NAND21X1 U140 ( .B(n177), .A(i_rdat[7]), .Y(n158) );
  NAND31X1 U141 ( .C(n168), .A(n167), .B(n166), .Y(n169) );
  NAND21X1 U142 ( .B(n111), .A(n165), .Y(n166) );
  NAND21X1 U143 ( .B(n160), .A(n159), .Y(n167) );
  INVX1 U144 ( .A(n26), .Y(n173) );
  NAND6XL U145 ( .A(cs_rwb), .B(o_dbgpo[3]), .C(n25), .D(n129), .E(n24), .F(
        i_rd_mem), .Y(n26) );
  NAND21X1 U146 ( .B(n173), .A(n29), .Y(n130) );
  NAND6XL U147 ( .A(i_rd_mem), .B(cs_rwb), .C(n129), .D(n28), .E(n133), .F(n27), .Y(n29) );
  INVX1 U148 ( .A(o_dbgpo[1]), .Y(n27) );
  AO22X1 U149 ( .A(n131), .B(o_wdat[4]), .C(i_rdat[5]), .D(n130), .Y(N141) );
  OAI21BBX1 U150 ( .A(i_rdat[0]), .B(n130), .C(n6), .Y(N136) );
  NAND4X1 U151 ( .A(o_dbgpo[6]), .B(ps_rwbuf_0_), .C(n162), .D(n164), .Y(n6)
         );
  AO22X1 U152 ( .A(n131), .B(o_wdat[0]), .C(i_rdat[1]), .D(n130), .Y(N137) );
  AO22X1 U153 ( .A(n131), .B(o_wdat[5]), .C(i_rdat[6]), .D(n130), .Y(N142) );
  AO22X1 U154 ( .A(n131), .B(o_wdat[1]), .C(i_rdat[2]), .D(n130), .Y(N138) );
  NAND32X1 U155 ( .B(n24), .C(o_dbgpo[7]), .A(sdafall), .Y(n23) );
  NAND21X1 U156 ( .B(n62), .A(o_ofs[4]), .Y(n67) );
  NAND31X1 U157 ( .C(n46), .A(o_ofs[0]), .B(i_inc), .Y(n47) );
  MUX2X1 U158 ( .D0(n113), .D1(cs_sta[0]), .S(n123), .Y(n120) );
  NAND21X1 U159 ( .B(n107), .A(n114), .Y(n113) );
  AND4X1 U160 ( .A(n175), .B(n148), .C(n116), .D(n164), .Y(n107) );
  MUX2X1 U161 ( .D0(n124), .D1(cs_sta[1]), .S(n123), .Y(n121) );
  NAND21X1 U162 ( .B(n122), .A(n117), .Y(n124) );
  AO21X1 U163 ( .B(n156), .C(n116), .A(n115), .Y(n117) );
  INVX1 U164 ( .A(n114), .Y(n122) );
  NAND31X1 U165 ( .C(n55), .A(o_ofs[3]), .B(n54), .Y(n62) );
  MUX2IX1 U166 ( .D0(n7), .D1(n8), .S(o_ofs[7]), .Y(n74) );
  NAND2X1 U167 ( .A(o_ofs[6]), .B(n71), .Y(n7) );
  AOI21X1 U168 ( .B(n152), .C(n73), .A(n72), .Y(n8) );
  NAND3X1 U169 ( .A(i2c_scl), .B(n176), .C(o_dbgpo[5]), .Y(n64) );
  INVX1 U170 ( .A(o_ofs[1]), .Y(n46) );
  AO21X1 U171 ( .B(n106), .C(n108), .A(n115), .Y(n114) );
  NAND5XL U172 ( .A(i_prefetch), .B(o_dbgpo[1]), .C(n133), .D(n132), .E(n95), 
        .Y(n106) );
  NAND43X1 U173 ( .B(n94), .C(n93), .D(n92), .A(n91), .Y(n95) );
  INVX1 U174 ( .A(n81), .Y(n94) );
  NAND21X1 U175 ( .B(n111), .A(cs_sta[0]), .Y(n129) );
  NAND21X1 U176 ( .B(cs_sta[1]), .A(cs_sta[0]), .Y(n57) );
  AO21X1 U177 ( .B(o_wdat[3]), .C(n125), .A(n52), .Y(N109) );
  MUX2X1 U178 ( .D0(n51), .D1(n53), .S(o_ofs[3]), .Y(n52) );
  AND3X1 U179 ( .A(n54), .B(o_ofs[2]), .C(n152), .Y(n51) );
  OAI21BBX1 U180 ( .A(o_wdat[6]), .B(n125), .C(n9), .Y(N112) );
  MUX2IX1 U181 ( .D0(n71), .D1(n72), .S(o_ofs[6]), .Y(n9) );
  AO21X1 U182 ( .B(o_wdat[5]), .C(n125), .A(n66), .Y(N111) );
  MUX2X1 U183 ( .D0(n65), .D1(n69), .S(o_ofs[5]), .Y(n66) );
  AND2X1 U184 ( .A(n63), .B(n1), .Y(n65) );
  INVX1 U185 ( .A(n67), .Y(n63) );
  OAI222XL U186 ( .A(n61), .B(n60), .C(n59), .D(n58), .E(n57), .F(n56), .Y(
        N110) );
  INVX1 U187 ( .A(o_ofs[4]), .Y(n60) );
  MUX2X1 U188 ( .D0(n62), .D1(o_ofs[3]), .S(o_ofs[4]), .Y(n59) );
  INVX1 U189 ( .A(n53), .Y(n61) );
  INVX1 U190 ( .A(i2c_scl), .Y(n24) );
  INVX1 U191 ( .A(o_ofs[2]), .Y(n55) );
  GEN2XL U192 ( .D(o_dbgpo[3]), .E(n21), .C(n148), .B(n20), .A(n115), .Y(N78)
         );
  INVX1 U193 ( .A(n178), .Y(n20) );
  GEN2XL U194 ( .D(o_dbgpo[2]), .E(n76), .C(n25), .B(n14), .A(n78), .Y(N77) );
  MUX2BXL U195 ( .D0(ps_rwbuf_0_), .D1(n10), .S(n11), .Y(n119) );
  NAND2X1 U196 ( .A(cs_rwb), .B(n23), .Y(n10) );
  NAND2X1 U197 ( .A(o_busev[1]), .B(n23), .Y(n11) );
  NAND21X1 U198 ( .B(n162), .A(cs_rwb), .Y(n156) );
  AO21X1 U199 ( .B(o_wdat[0]), .C(o_we), .A(n146), .Y(N180) );
  AO21X1 U200 ( .B(o_wdat[0]), .C(n125), .A(n40), .Y(N106) );
  MUX2X1 U201 ( .D0(n39), .D1(n41), .S(o_ofs[0]), .Y(n40) );
  AND2X1 U202 ( .A(i_inc), .B(n152), .Y(n39) );
  AO21X1 U203 ( .B(o_wdat[2]), .C(n125), .A(n49), .Y(N108) );
  MUX2X1 U204 ( .D0(n48), .D1(n50), .S(o_ofs[2]), .Y(n49) );
  AND2X1 U205 ( .A(n54), .B(n1), .Y(n48) );
  NAND32X1 U206 ( .B(n139), .C(n138), .A(n137), .Y(N114) );
  AND3X1 U207 ( .A(n1), .B(o_dbgpo[7]), .C(n136), .Y(n138) );
  MUX2X1 U208 ( .D0(n148), .D1(n135), .S(cs_rwb), .Y(n136) );
  MUX2X1 U209 ( .D0(n160), .D1(n134), .S(i_prefetch), .Y(n135) );
  AND3X1 U210 ( .A(o_dbgpo[1]), .B(n133), .C(n132), .Y(n134) );
  OAI222XL U211 ( .A(n45), .B(n46), .C(n44), .D(n58), .E(n57), .F(n43), .Y(
        N107) );
  MUX2BXL U212 ( .D0(n46), .D1(n42), .S(o_ofs[0]), .Y(n44) );
  INVX1 U213 ( .A(n41), .Y(n45) );
  AND2X1 U214 ( .A(i_inc), .B(n46), .Y(n42) );
  INVX1 U215 ( .A(n80), .Y(n132) );
  NAND21X1 U216 ( .B(o_dbgpo[2]), .A(n79), .Y(n80) );
  INVX1 U217 ( .A(o_ofs[6]), .Y(n73) );
  INVX1 U218 ( .A(o_ofs[5]), .Y(n70) );
  INVX1 U219 ( .A(cs_sta[0]), .Y(n116) );
  AO22XL U220 ( .A(n131), .B(o_wdat[3]), .C(i_rdat[4]), .D(n130), .Y(N140) );
  AO22XL U221 ( .A(n131), .B(o_wdat[2]), .C(i_rdat[3]), .D(n130), .Y(N139) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2cdbnc_a0_0 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall, test_si, 
        test_se );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c, test_si, test_se;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n9, n1, n2, n3, n4, n5, n6, n7;

  SDFFSQX1 d_i2c_reg_2_ ( .D(N19), .SIN(N19), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(d_i2c_2_) );
  SDFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .SIN(test_si), .SMC(test_se), .C(i_clk), 
        .XS(i_rstz), .Q(N18) );
  SDFFSQX1 d_i2c_reg_1_ ( .D(N18), .SIN(N18), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(N19) );
  SDFFSQXX1 r_i2c_reg ( .D(n9), .SIN(d_i2c_2_), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(o_i2c), .XQ(n1) );
  AND2X1 U3 ( .A(o_i2c), .B(n7), .Y(fall) );
  INVX1 U4 ( .A(n6), .Y(n7) );
  NOR43XL U5 ( .B(N19), .C(N18), .D(n1), .A(n5), .Y(rise) );
  NOR2X1 U6 ( .A(r_opt[0]), .B(d_i2c_2_), .Y(n5) );
  OAI211X1 U7 ( .C(r_opt[1]), .D(n4), .A(n3), .B(n2), .Y(n6) );
  INVX1 U8 ( .A(N18), .Y(n3) );
  INVX1 U9 ( .A(N19), .Y(n2) );
  INVX1 U10 ( .A(d_i2c_2_), .Y(n4) );
  AO21X1 U11 ( .B(o_i2c), .C(n6), .A(rise), .Y(n9) );
endmodule


module i2cdbnc_a0_1 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall, test_si, 
        test_se );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c, test_si, test_se;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n6, n1, n2, n3, n4;

  SDFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .SIN(test_si), .SMC(test_se), .C(i_clk), 
        .XS(i_rstz), .Q(N18) );
  SDFFSQX1 d_i2c_reg_1_ ( .D(N18), .SIN(N18), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(N19) );
  SDFFSQX1 d_i2c_reg_2_ ( .D(N19), .SIN(N19), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(d_i2c_2_) );
  SDFFSQXX1 r_i2c_reg ( .D(n6), .SIN(d_i2c_2_), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(o_i2c), .XQ(n3) );
  INVX1 U3 ( .A(n4), .Y(fall) );
  NOR43XL U4 ( .B(N19), .C(N18), .D(n3), .A(n2), .Y(rise) );
  NOR2X1 U5 ( .A(d_i2c_2_), .B(r_opt[0]), .Y(n2) );
  NAND42X1 U6 ( .C(N18), .D(N19), .A(n1), .B(o_i2c), .Y(n4) );
  NAND21X1 U7 ( .B(r_opt[1]), .A(d_i2c_2_), .Y(n1) );
  AO21X1 U8 ( .B(o_i2c), .C(n4), .A(rise), .Y(n6) );
endmodule


module regbank_a0 ( srci, lg_pulse_len, dm_fault, cc1_di, cc2_di, di_rd_det, 
        i_tmrf, i_vcbyval, dnchk_en, r_pwrv_upd, aswkup, lg_dischg, frc_hg_off, 
        ps_pwrdn, r_sleep, r_pwrdn, r_ocdrv_enz, r_osc_stop, r_osc_lo, 
        r_osc_gate, r_fw_pwrv, r_cvcwr, r_cvofs, r_otpi_gate, r_pwrctl, 
        r_pwr_i, r_cvctl, r_srcctl, r_dpdmctl, r_ccrx, r_cctrx, r_ccctl, 
        r_fcpwr, r_fcpre, fcp_r_dat, fcp_r_sta, fcp_r_msk, fcp_r_ctl, 
        fcp_r_crc, fcp_r_acc, fcp_r_tui, r_accctl, r_bclk_sel, r_dacwr, 
        r_dac_en, r_sar_en, r_adofs, r_isofs, x_daclsb, r_comp_opt, dac_r_ctl, 
        dac_r_comp, dac_r_cmpsta, dac_r_vs, REVID, atpg_en, sfr_r, sfr_w, 
        set_hold, bkpt_hold, cpurst, sfr_addr, sfr_wdat, sfr_rdat, ff_p0, 
        di_p0, ictlr_idle, ictlr_inc, r_inst_ofs, r_psrd, r_pswr, r_fortxdat, 
        r_fortxrdy, r_fortxen, r_ana_tm, r_gpio_tm, r_gpio_ie, r_gpio_oe, 
        r_gpio_pu, r_gpio_pd, r_gpio_s0, r_gpio_s1, r_gpio_s2, r_gpio_s3, 
        r_regtrm, i_pc, i_goidle, i_gobusy, i_i2c_idle, bus_idle, i2c_stretch, 
        i_i2c_rwbuf, i_i2c_ltbuf, i_i2c_ofs, o_intr, r_auto_gdcrc, r_exist1st, 
        r_ordrs4, r_fifopsh, r_fifopop, r_unlock, r_first, r_last, r_fiforst, 
        r_set_cpmsgid, r_txendk, r_txnumk, r_txshrt, r_auto_discard, 
        r_hold_mcu, r_txauto, r_rxords_ena, r_spec, r_dat_spec, r_dat_portrole, 
        r_dat_datarole, r_discard, r_pshords, r_pg0_sel, r_strtch, r_i2c_attr, 
        r_i2c_ninc, r_hwi2c_en, r_i2c_fwnak, r_i2c_fwack, r_i2c_deva, i2c_ev, 
        prl_c0set, prl_cany0, prl_discard, prl_GCTxDone, prl_cpmsgid, pff_ack, 
        prx_rst, pff_obsd, pff_full, pff_empty, ptx_ack, pff_ptr, prx_adpn, 
        pff_rdat, pff_rxpart, prx_rcvinf, ptx_fsm, prx_fsm, prl_fsm, 
        prx_setsta, clk_1p0m, clk_500, clk, xrstz, xclk, dbgpo, srstz, prstz, 
        test_si2, test_si1, test_so2, test_so1, test_se );
  input [5:0] srci;
  input [1:0] lg_pulse_len;
  output [11:0] r_fw_pwrv;
  output [1:0] r_cvcwr;
  input [15:0] r_cvofs;
  output [7:4] r_pwrctl;
  output [7:0] r_pwr_i;
  output [7:0] r_cvctl;
  output [7:0] r_srcctl;
  output [7:0] r_dpdmctl;
  output [7:0] r_ccrx;
  output [7:0] r_cctrx;
  output [7:0] r_ccctl;
  output [6:0] r_fcpwr;
  input [7:0] fcp_r_dat;
  input [7:0] fcp_r_sta;
  input [7:0] fcp_r_msk;
  input [7:0] fcp_r_ctl;
  input [7:0] fcp_r_crc;
  input [7:0] fcp_r_acc;
  input [7:0] fcp_r_tui;
  input [7:0] r_accctl;
  output [14:0] r_dacwr;
  input [7:0] r_dac_en;
  input [7:0] r_sar_en;
  input [7:0] r_adofs;
  input [7:0] r_isofs;
  input [5:0] x_daclsb;
  output [7:0] r_comp_opt;
  input [7:0] dac_r_ctl;
  input [7:0] dac_r_comp;
  input [7:0] dac_r_cmpsta;
  input [63:0] dac_r_vs;
  input [6:0] REVID;
  input [7:0] sfr_addr;
  input [7:0] sfr_wdat;
  output [7:0] sfr_rdat;
  input [7:0] ff_p0;
  input [7:0] di_p0;
  output [14:0] r_inst_ofs;
  output [3:0] r_ana_tm;
  output [1:0] r_gpio_ie;
  output [6:0] r_gpio_oe;
  output [6:0] r_gpio_pu;
  output [6:0] r_gpio_pd;
  output [2:0] r_gpio_s0;
  output [2:0] r_gpio_s1;
  output [2:0] r_gpio_s2;
  output [2:0] r_gpio_s3;
  output [55:0] r_regtrm;
  input [15:0] i_pc;
  input [7:0] i_i2c_rwbuf;
  input [7:0] i_i2c_ltbuf;
  input [7:0] i_i2c_ofs;
  output [4:0] o_intr;
  output [1:0] r_auto_gdcrc;
  output [4:0] r_txnumk;
  output [6:0] r_txauto;
  output [6:0] r_rxords_ena;
  output [1:0] r_spec;
  output [1:0] r_dat_spec;
  output [3:0] r_pg0_sel;
  output [7:1] r_i2c_deva;
  input [7:0] i2c_ev;
  input [2:0] prl_cpmsgid;
  input [1:0] pff_ack;
  input [1:0] prx_rst;
  input [5:0] pff_ptr;
  input [5:0] prx_adpn;
  input [7:0] pff_rdat;
  input [15:0] pff_rxpart;
  input [4:0] prx_rcvinf;
  input [2:0] ptx_fsm;
  input [3:0] prx_fsm;
  input [3:0] prl_fsm;
  input [6:0] prx_setsta;
  output [31:0] dbgpo;
  input dm_fault, cc1_di, cc2_di, di_rd_det, i_tmrf, i_vcbyval, dnchk_en,
         atpg_en, sfr_r, sfr_w, set_hold, bkpt_hold, cpurst, ictlr_idle,
         ictlr_inc, i_goidle, i_gobusy, i_i2c_idle, prl_c0set, prl_cany0,
         prl_discard, prl_GCTxDone, pff_obsd, pff_full, pff_empty, ptx_ack,
         clk_1p0m, clk_500, clk, xrstz, xclk, test_si2, test_si1, test_se;
  output r_pwrv_upd, aswkup, lg_dischg, frc_hg_off, ps_pwrdn, r_sleep, r_pwrdn,
         r_ocdrv_enz, r_osc_stop, r_osc_lo, r_osc_gate, r_otpi_gate, r_fcpre,
         r_bclk_sel, r_psrd, r_pswr, r_fortxdat, r_fortxrdy, r_fortxen,
         r_gpio_tm, bus_idle, i2c_stretch, r_exist1st, r_ordrs4, r_fifopsh,
         r_fifopop, r_unlock, r_first, r_last, r_fiforst, r_set_cpmsgid,
         r_txendk, r_txshrt, r_auto_discard, r_hold_mcu, r_dat_portrole,
         r_dat_datarole, r_discard, r_pshords, r_strtch, r_i2c_attr,
         r_i2c_ninc, r_hwi2c_en, r_i2c_fwnak, r_i2c_fwack, srstz, prstz,
         test_so2, test_so1;
  wire   we_246, we_245, we_232, we_231, we_230, we_228, we_227, we_222,
         we_217, we_215, we_214, we_213, we_211, we_209, we_203, we_191,
         we_187, we_182, we_181, we_176, we_175, we_172, we_171, we_148,
         we_143, regF4_7_, regF4_3, regE3_0, regD4_6_, regD4_5_, regD4_4_,
         regD4_3_, regD4_2_, regD4_1_, regD4_0_, regD3_7_, regD3_3, reg25_0_,
         reg19_7_, reg12_1, reg11_7_, reg11_4, regAD_7, N26, N27, N28, N29,
         N30, N32, N33, N34, N35, N36, N37, N38, N39, upd01, phyrst, upd12,
         upd18, upd19, upd20, upd21, lt_reg26_0, i2c_mode_upd, i2c_mode_wdat,
         upd31, N84, as_p0_chg, dmf_wkup, p0_chg_clr, di_rd_det_clr,
         dm_fault_clr, pwrdn_rstz, osc_low_clr, osc_low_rstz, r_pos_gate,
         osc_gate_n_2_, osc_gate_n_1_, osc_gate_n_0_, m_ovp, m_ovp_sta,
         setAE_7, m_scp, m_scp_sta, s_ovp, s_ovp_sta, s_scp, s_scp_sta,
         lg_pulse_12m, N108, N109, N110, N111, N112, N113, net10832, net10838,
         n1219, n1220, n1221, n1222, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n77, n109, n111, n112,
         n113, n115, n117, n118, n119, n120, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n134, n135, n140, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n170,
         n171, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n1, n2, n3, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n110, n114, n116, n121, n133, n136,
         n137, n138, n139, n141, n142, n143, n144, n168, n169, n172, n183,
         n184, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462,
         SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464,
         SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466,
         SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468,
         SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470,
         SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472,
         SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474,
         SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476,
         SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478,
         SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480,
         SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482,
         SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484,
         SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486,
         SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488,
         SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490,
         SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492,
         SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494,
         SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496,
         SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498,
         SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500,
         SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502,
         SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504,
         SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506,
         SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508,
         SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510,
         SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512,
         SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514,
         SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516,
         SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518,
         SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520,
         SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522,
         SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524,
         SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526,
         SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528,
         SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530,
         SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532,
         SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534,
         SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536,
         SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538,
         SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540,
         SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542,
         SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544,
         SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546,
         SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548,
         SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550,
         SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552,
         SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554,
         SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556,
         SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558,
         SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560,
         SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562,
         SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564,
         SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566,
         SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568,
         SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570,
         SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572,
         SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574,
         SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576,
         SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578,
         SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580,
         SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582,
         SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584,
         SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586,
         SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588,
         SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590,
         SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592,
         SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594,
         SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596,
         SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598,
         SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600,
         SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602,
         SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604,
         SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606,
         SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608,
         SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610,
         SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612,
         SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614,
         SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616,
         SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618,
         SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620,
         SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622,
         SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624,
         SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626,
         SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628,
         SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630,
         SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632,
         SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634,
         SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636,
         SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638,
         SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640,
         SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642,
         SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644,
         SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646,
         SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648,
         SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650,
         SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652,
         SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654,
         SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656,
         SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658,
         SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660,
         SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662,
         SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664,
         SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666,
         SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668,
         SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670,
         SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672,
         SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674,
         SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676,
         SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678,
         SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680,
         SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682,
         SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684,
         SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686,
         SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688,
         SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690,
         SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692,
         SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694,
         SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696,
         SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698,
         SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700,
         SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702,
         SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704,
         SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706,
         SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708,
         SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710,
         SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712,
         SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714,
         SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716,
         SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718,
         SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720,
         SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722,
         SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724,
         SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726,
         SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728,
         SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730,
         SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732,
         SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734,
         SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736,
         SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738,
         SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740,
         SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742,
         SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744,
         SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746,
         SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748,
         SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750,
         SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752,
         SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754,
         SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756,
         SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758,
         SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760,
         SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762,
         SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764,
         SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766,
         SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768,
         SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770,
         SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772,
         SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774,
         SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776,
         SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778,
         SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780,
         SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782,
         SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784,
         SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786,
         SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788,
         SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790,
         SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792,
         SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794,
         SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796,
         SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798,
         SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800,
         SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802,
         SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804,
         SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806,
         SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808,
         SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810,
         SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812,
         SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814,
         SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816,
         SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818,
         SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820,
         SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822,
         SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824,
         SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826,
         SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828,
         SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830,
         SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832,
         SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834,
         SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836,
         SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838,
         SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840,
         SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842,
         SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844,
         SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846,
         SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848,
         SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850,
         SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852,
         SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854,
         SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856,
         SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858,
         SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860,
         SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862,
         SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864,
         SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866,
         SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868,
         SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870,
         SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872,
         SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874,
         SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876,
         SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878,
         SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880,
         SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882,
         SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884,
         SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886,
         SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888,
         SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890,
         SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892,
         SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894,
         SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896,
         SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898,
         SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900,
         SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902,
         SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904,
         SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906,
         SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908,
         SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910,
         SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912,
         SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914,
         SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916,
         SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918,
         SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920,
         SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922,
         SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924,
         SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926,
         SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928,
         SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930,
         SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932,
         SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934,
         SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936,
         SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938,
         SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940,
         SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942,
         SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944,
         SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946,
         SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948,
         SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950,
         SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952,
         SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954,
         SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956,
         SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958,
         SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960,
         SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962,
         SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964,
         SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966,
         SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968,
         SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970,
         SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972,
         SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974,
         SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976,
         SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978,
         SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980,
         SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982,
         SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984,
         SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986,
         SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988,
         SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990,
         SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992,
         SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994,
         SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996,
         SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998,
         SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000,
         SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002,
         SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004,
         SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006,
         SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008,
         SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010,
         SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012,
         SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014,
         SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016,
         SYNOPSYS_UNCONNECTED_1017;
  wire   [167:161] we;
  wire   [3:2] regE3;
  wire   [7:0] regDF;
  wire   [7:0] regDE;
  wire   [7:0] reg31;
  wire   [7:0] reg30;
  wire   [7:0] reg28;
  wire   [7:0] reg27;
  wire   [7:1] reg21;
  wire   [4:0] reg20;
  wire   [7:3] reg12;
  wire   [7:0] reg06;
  wire   [7:0] reg05;
  wire   [7:0] regAF;
  wire   [7:0] regAE;
  wire   [5:0] regAD;
  wire   [7:0] regAC;
  wire   [7:0] regAB;
  wire   [7:0] reg94;
  wire   [7:0] irqAE;
  wire   [7:0] irqDF;
  wire   [7:0] irq28;
  wire   [7:0] irq04;
  wire   [7:0] irq03;
  wire   [1:0] drstz;
  wire   [4:0] rstcnt;
  wire   [1:0] r_phyrst;
  wire   [7:0] wd01;
  wire   [7:0] clr03;
  wire   [7:0] set03;
  wire   [7:0] clr04;
  wire   [7:0] set04;
  wire   [7:0] wd12;
  wire   [14:0] inst_ofs_plus;
  wire   [7:0] wd18;
  wire   [7:0] wd19;
  wire   [7:0] wd20;
  wire   [7:0] wd21;
  wire   [7:0] clr28;
  wire   [2:0] oscdwn_shft;
  wire   [7:0] d_p0;
  wire   [7:0] setDF;
  wire   [7:0] clrDF;
  wire   [7:0] clrAE;
  wire   [5:0] setAE;
  wire   [4:0] lg_pulse_cnt;
  wire   [3:0] lt_regE4_3_0;
  wire   [4:2] add_180_carry;

  AND2X1 U0_MASK_0 ( .A(oscdwn_shft[2]), .B(as_p0_chg), .Y(p0_chg_clr) );
  AND2X1 U0_MASK_2 ( .A(regD4_6_), .B(di_rd_det), .Y(di_rd_det_clr) );
  AND2X1 U0_MASK_3 ( .A(r_srcctl[6]), .B(dmf_wkup), .Y(dm_fault_clr) );
  AND2X1 U0_MASK_4 ( .A(regD4_5_), .B(aswkup), .Y(osc_low_clr) );
  HAD1X1 add_180_U1_1_1 ( .A(N29), .B(N30), .CO(add_180_carry[2]), .SO(N32) );
  HAD1X1 add_180_U1_1_2 ( .A(N28), .B(add_180_carry[2]), .CO(add_180_carry[3]), 
        .SO(N33) );
  HAD1X1 add_180_U1_1_3 ( .A(N27), .B(add_180_carry[3]), .CO(add_180_carry[4]), 
        .SO(N34) );
  glreg_a0_79 u0_reg00 ( .clk(clk), .arstz(n65), .we(we_176), .wdat({n249, 
        n241, n229, n222, n216, n168, n138, n116}), .rdat({r_txendk, r_txauto}), .test_si(n316), .test_se(test_se) );
  glreg_a0_78 u0_reg01 ( .clk(clk), .arstz(n64), .we(upd01), .wdat(wd01), 
        .rdat({r_last, r_first, r_unlock, r_txnumk}), .test_si(r_txendk), 
        .test_se(test_se) );
  glsta_a0_6 u0_reg03 ( .clk(clk), .arstz(n36), .rst0(n16), .set2({set03[7:4], 
        n77, set03[2:0]}), .clr1(clr03), .rdat(dbgpo[7:0]), .irq(irq03), 
        .test_si(r_last), .test_se(test_se) );
  glsta_a0_5 u0_reg04 ( .clk(clk), .arstz(n37), .rst0(n17), .set2(set04), 
        .clr1(clr04), .rdat(dbgpo[15:8]), .irq(irq04), .test_si(dbgpo[7]), 
        .test_se(test_se) );
  glreg_a0_77 u0_reg05 ( .clk(clk), .arstz(n45), .we(we_181), .wdat({n250, 
        n241, n229, n222, n217, n169, n138, n114}), .rdat(reg05), .test_si(
        dbgpo[15]), .test_se(test_se) );
  glreg_a0_76 u0_reg06 ( .clk(clk), .arstz(n38), .we(we_182), .wdat({n250, 
        n238, n228, n222, n216, n168, n138, n116}), .rdat(reg06), .test_si(
        reg05[7]), .test_se(test_se) );
  glreg_a0_75 u0_reg11 ( .clk(clk), .arstz(n39), .we(we_187), .wdat({n250, 
        sfr_wdat[6], n228, n222, n217, n169, n139, n116}), .rdat({reg11_7_, 
        r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0]}), .test_si(r_dpdmctl[7]), .test_se(test_se) );
  glreg_a0_74 u0_reg12 ( .clk(clk), .arstz(n63), .we(upd12), .wdat(wd12), 
        .rdat({reg12, r_txshrt, reg12_1, r_pshords}), .test_si(reg11_7_), 
        .test_se(test_se) );
  glreg_WIDTH5_2 u0_reg14 ( .clk(clk), .arstz(n79), .we(r_set_cpmsgid), .wdat(
        {n250, n239, n229, n222, n217}), .rdat({r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1]}), .test_si(reg12[7]), 
        .test_se(test_se) );
  glreg_a0_73 u0_reg15 ( .clk(clk), .arstz(n40), .we(we_191), .wdat({n250, 
        n238, n229, n223, n217, n169, n139, n121}), .rdat(dbgpo[31:24]), 
        .test_si(r_auto_gdcrc[0]), .test_se(test_se) );
  glreg_a0_72 u0_reg18 ( .clk(clk), .arstz(n46), .we(upd18), .wdat(wd18), 
        .rdat(r_inst_ofs[7:0]), .test_si(dbgpo[31]), .test_se(test_se) );
  glreg_a0_71 u0_reg19 ( .clk(clk), .arstz(n41), .we(upd19), .wdat(wd19), 
        .rdat({reg19_7_, r_inst_ofs[14:8]}), .test_si(r_inst_ofs[7]), 
        .test_se(test_se) );
  glreg_a0_70 u0_reg20 ( .clk(clk), .arstz(n61), .we(upd20), .wdat(wd20), 
        .rdat({r_dat_spec, r_dat_datarole, reg20}), .test_si(reg19_7_), 
        .test_se(test_se) );
  glreg_a0_69 u0_reg21 ( .clk(clk), .arstz(n51), .we(upd21), .wdat(wd21), 
        .rdat({reg21, r_dat_portrole}), .test_si(r_dat_spec[1]), .test_se(
        test_se) );
  glreg_6_00000018 u0_reg25 ( .clk(clk), .arstz(n74), .we(n212), .wdat({
        sfr_wdat[5:4], n216, n172, n139, n116}), .rdat({r_i2c_attr, r_pg0_sel, 
        reg25_0_}), .test_si(reg21[7]), .test_se(test_se) );
  glreg_1_1_1 u0_reg26 ( .clk(clk), .arstz(n86), .we(n213), .wdat(n114), 
        .rdat(lt_reg26_0), .test_si(r_i2c_attr), .test_se(test_se) );
  glreg_1_1_0 u1_reg26 ( .clk(clk), .arstz(n86), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat(r_hwi2c_en), .test_si(n311), .test_se(test_se)
         );
  glreg_7_70 u2_reg26 ( .clk(clk), .arstz(n71), .we(n213), .wdat({n249, 
        sfr_wdat[6], n228, n222, n217, n169, n139}), .rdat(r_i2c_deva), 
        .test_si(n308), .test_se(test_se) );
  glreg_a0_68 u0_reg27 ( .clk(clk), .arstz(n50), .we(we_203), .wdat({n250, 
        n238, n229, n222, n217, n169, n139, n116}), .rdat(reg27), .test_si(
        lt_reg26_0), .test_se(test_se) );
  glsta_a0_4 u0_reg28 ( .clk(clk), .arstz(n43), .rst0(1'b0), .set2(i2c_ev), 
        .clr1(clr28), .rdat(reg28), .irq(irq28), .test_si(reg27[7]), .test_se(
        test_se) );
  glreg_a0_67 u0_reg31 ( .clk(clk), .arstz(n44), .we(upd31), .wdat(i_pc[15:8]), 
        .rdat(reg31), .test_si(reg28[7]), .test_se(test_se) );
  glreg_8_00000001 u0_regD1 ( .clk(clk), .arstz(n35), .we(we_209), .wdat({n250, 
        n238, n229, n222, n217, n169, n139, n114}), .rdat({r_exist1st, 
        r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, r_gpio_oe[6], r_gpio_pu[6], 
        r_gpio_pd[6]}), .test_si(regAF[7]), .test_se(test_se) );
  glreg_8_00000011 u0_regD3 ( .clk(clk), .arstz(n32), .we(we_211), .wdat({n250, 
        n238, n229, n225, n217, n169, n139, n114}), .rdat({regD3_7_, 
        r_gpio_oe[5], r_gpio_pu[5], r_gpio_pd[5], regD3_3, r_gpio_oe[4], 
        r_gpio_pu[4], r_gpio_pd[4]}), .test_si(r_exist1st), .test_se(test_se)
         );
  glreg_WIDTH3 u4_regD4 ( .clk(clk), .arstz(n86), .we(n10), .wdat({n250, n238, 
        n229}), .rdat({test_so2, regD4_6_, regD4_5_}), .test_si(regD4_4_), 
        .test_se(test_se) );
  glreg_WIDTH2_2 u3_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n10), .wdat({
        n225, n216}), .rdat({regD4_4_, regD4_3_}), .test_si(regD4_2_), 
        .test_se(test_se) );
  glreg_WIDTH1_5 u2_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n10), .wdat(
        n168), .rdat(regD4_2_), .test_si(r_i2c_deva[7]), .test_se(test_se) );
  glreg_WIDTH1_4 u1_regD4 ( .clk(clk), .arstz(osc_low_rstz), .we(n10), .wdat(
        n138), .rdat(regD4_1_), .test_si(r_hwi2c_en), .test_se(test_se) );
  glreg_WIDTH1_3 u0_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n10), .wdat(
        n114), .rdat(regD4_0_), .test_si(regD3_7_), .test_se(test_se) );
  glreg_8_000000f0 u0_regD5 ( .clk(clk), .arstz(n29), .we(we_213), .wdat({n249, 
        n241, n228, n225, n217, n169, n139, n116}), .rdat({r_gpio_pu[3:0], 
        r_gpio_pd[3:0]}), .test_si(regD4_0_), .test_se(test_se) );
  glreg_8_00000098 u0_regD6 ( .clk(clk), .arstz(n31), .we(we_214), .wdat({n249, 
        n238, n229, n225, n216, n169, n139, n116}), .rdat({r_gpio_oe[1], 
        r_gpio_s1, r_gpio_oe[0], r_gpio_s0}), .test_si(r_gpio_pu[3]), 
        .test_se(test_se) );
  glreg_8_00000032 u0_regD7 ( .clk(clk), .arstz(n30), .we(we_215), .wdat({n250, 
        n238, n228, n225, n218, n169, n138, n116}), .rdat({r_gpio_oe[3], 
        r_gpio_s3, r_gpio_oe[2], r_gpio_s2}), .test_si(r_gpio_oe[1]), 
        .test_se(test_se) );
  glreg_a0_66 u0_regD9 ( .clk(clk), .arstz(n47), .we(we_217), .wdat({n251, 
        n238, n229, n222, n218, n172, n139, n116}), .rdat({r_ana_tm, 
        r_fortxdat, r_fortxrdy, r_fortxen, r_sleep}), .test_si(r_gpio_oe[3]), 
        .test_se(test_se) );
  glreg_a0_65 u0_regDE ( .clk(clk), .arstz(n48), .we(we_222), .wdat({n251, 
        n238, n231, n223, n218, n172, n141, n116}), .rdat(regDE), .test_si(
        r_ana_tm[3]), .test_se(test_se) );
  glsta_a0_3 u0_regDF ( .clk(clk), .arstz(n49), .rst0(1'b0), .set2(setDF), 
        .clr1(clrDF), .rdat(regDF), .irq(irqDF), .test_si(regDE[7]), .test_se(
        test_se) );
  glreg_a0_64 u0_reg8F ( .clk(clk), .arstz(n54), .we(we_143), .wdat({n251, 
        n239, n231, n223, n218, n172, n141, n121}), .rdat(r_dpdmctl), 
        .test_si(reg06[7]), .test_se(test_se) );
  glreg_WIDTH4 u0_reg94 ( .clk(clk), .arstz(n83), .we(we_148), .wdat({n239, 
        n231, n223, n218}), .rdat(reg94[6:3]), .test_si(reg31[7]), .test_se(
        test_se) );
  glreg_a0_63 u0_regA1 ( .clk(clk), .arstz(n52), .we(we[161]), .wdat({n251, 
        n239, n231, n223, n218, n172, n141, n121}), .rdat(r_regtrm[7:0]), 
        .test_si(reg94[6]), .test_se(test_se) );
  glreg_a0_62 u0_regA2 ( .clk(clk), .arstz(n53), .we(we[162]), .wdat({n251, 
        n239, n231, n223, n218, n172, n141, n121}), .rdat(r_regtrm[15:8]), 
        .test_si(r_regtrm[7]), .test_se(test_se) );
  glreg_a0_61 u0_regA3 ( .clk(clk), .arstz(n58), .we(we[163]), .wdat({n251, 
        n239, n231, n223, n218, n172, n141, n121}), .rdat(r_regtrm[23:16]), 
        .test_si(r_regtrm[15]), .test_se(test_se) );
  glreg_a0_60 u0_regA4 ( .clk(clk), .arstz(n55), .we(we[164]), .wdat({n251, 
        n239, n231, n223, n218, n172, n141, n121}), .rdat(r_regtrm[31:24]), 
        .test_si(r_regtrm[23]), .test_se(test_se) );
  glreg_a0_59 u0_regA5 ( .clk(clk), .arstz(n56), .we(we[165]), .wdat({n251, 
        n239, n231, n223, n219, n172, n141, n121}), .rdat(r_regtrm[39:32]), 
        .test_si(r_regtrm[31]), .test_se(test_se) );
  glreg_a0_58 u0_regA6 ( .clk(clk), .arstz(n57), .we(we[166]), .wdat({n251, 
        n239, n231, n223, n218, n172, n141, n121}), .rdat(r_regtrm[47:40]), 
        .test_si(r_regtrm[39]), .test_se(test_se) );
  glreg_a0_57 u0_regA7 ( .clk(clk), .arstz(n60), .we(we[167]), .wdat({n252, 
        n239, n230, n224, n219, n183, n141, n121}), .rdat(r_regtrm[55:48]), 
        .test_si(r_regtrm[47]), .test_se(test_se) );
  glreg_a0_56 u0_regAB ( .clk(clk), .arstz(n59), .we(we_171), .wdat({n252, 
        n240, n230, n224, n219, n183, n141, n121}), .rdat(regAB), .test_si(
        r_regtrm[55]), .test_se(test_se) );
  glreg_8_00000028 u0_regAC ( .clk(clk), .arstz(n33), .we(we_172), .wdat({n252, 
        n240, n228, n224, n216, n183, n142, n133}), .rdat(regAC), .test_si(
        regAB[7]), .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_2 u2_ovp_db ( .o_dbc(reg94[2]), .o_chg(), .i_org(
        srci[2]), .clk(clk_500), .rstz(n75), .test_si(n309), .test_so(n308), 
        .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_1 u1_ocp_db ( .o_dbc(reg94[1]), .o_chg(), .i_org(
        srci[1]), .clk(clk_500), .rstz(n78), .test_si(n313), .test_so(n312), 
        .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_0 u1_uvp_db ( .o_dbc(reg94[0]), .o_chg(), .i_org(
        srci[0]), .clk(clk_500), .rstz(n76), .test_si(n310), .test_so(n309), 
        .test_se(test_se) );
  dbnc_WIDTH5_TIMEOUT30 u1_ovp_db ( .o_dbc(m_ovp), .o_chg(m_ovp_sta), .i_org(
        srci[2]), .clk(clk_1p0m), .rstz(n72), .test_si(n312), .test_so(n311), 
        .test_se(test_se) );
  dbnc_WIDTH2_4 u0_otpi_db ( .o_dbc(regAD[3]), .o_chg(setAE[3]), .i_org(
        srci[5]), .clk(clk_1p0m), .rstz(n85), .test_si(n319), .test_so(n318), 
        .test_se(test_se) );
  dbnc_WIDTH2_3 u0_ocp_db ( .o_dbc(regAD[1]), .o_chg(setAE[1]), .i_org(srci[1]), .clk(clk_1p0m), .rstz(n85), .test_si(n320), .test_so(n319), .test_se(test_se) );
  dbnc_WIDTH2_2 u0_uvp_db ( .o_dbc(regAD[0]), .o_chg(setAE[0]), .i_org(srci[0]), .clk(clk_1p0m), .rstz(n84), .test_si(n315), .test_so(n314), .test_se(test_se) );
  dbnc_WIDTH2_1 u1_scp_db ( .o_dbc(m_scp), .o_chg(m_scp_sta), .i_org(srci[3]), 
        .clk(clk_1p0m), .rstz(n84), .test_si(r_fw_pwrv[3]), .test_so(n310), 
        .test_se(test_se) );
  dbnc_WIDTH2_0 u0_dmf_db ( .o_dbc(regAD_7), .o_chg(setAE_7), .i_org(dm_fault), 
        .clk(clk_1p0m), .rstz(n83), .test_si(n321), .test_so(n320), .test_se(
        test_se) );
  dbnc_WIDTH2_TIMEOUT2_13 u0_otps_db ( .o_dbc(reg94[7]), .o_chg(), .i_org(
        srci[5]), .clk(clk), .rstz(n80), .test_si(n318), .test_so(n317), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_12 u0_cc1_db ( .o_dbc(regF4_3), .o_chg(), .i_org(cc1_di), .clk(clk), .rstz(n82), .test_si(rstcnt[4]), .test_so(n322), .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_11 u0_cc2_db ( .o_dbc(regF4_7_), .o_chg(), .i_org(
        cc2_di), .clk(clk), .rstz(n82), .test_si(n322), .test_so(n321), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_10 u0_ovp_db ( .o_dbc(s_ovp), .o_chg(s_ovp_sta), 
        .i_org(srci[2]), .clk(clk), .rstz(n81), .test_si(n317), .test_so(n316), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_9 u0_scp_db ( .o_dbc(s_scp), .o_chg(s_scp_sta), .i_org(
        srci[3]), .clk(clk), .rstz(n81), .test_si(r_cctrx[7]), .test_so(n315), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_8 u0_v5oc_db ( .o_dbc(regAD[5]), .o_chg(setAE[5]), 
        .i_org(srci[4]), .clk(clk), .rstz(n80), .test_si(n314), .test_so(n313), 
        .test_se(test_se) );
  glsta_a0_2 u0_regAE ( .clk(clk), .arstz(n69), .rst0(1'b0), .set2({setAE_7, 
        1'b0, setAE}), .clr1(clrAE), .rdat(regAE), .irq(irqAE), .test_si(
        regAC[7]), .test_se(test_se) );
  glreg_a0_55 u0_regAF ( .clk(clk), .arstz(n70), .we(we_175), .wdat({n252, 
        n240, n230, n224, n219, n183, n142, n133}), .rdat(regAF), .test_si(
        regAE[7]), .test_se(test_se) );
  glreg_WIDTH7_2 u0_regE3 ( .clk(clk), .arstz(n73), .we(we_227), .wdat({n252, 
        n240, n230, n224, n219, n183, n133}), .rdat({r_srcctl[7:4], regE3, 
        regE3_0}), .test_si(regDF[7]), .test_se(test_se) );
  glreg_4_00000004 u1_regE4 ( .clk(clk), .arstz(n79), .we(r_pwrv_upd), .wdat(
        lt_regE4_3_0), .rdat(r_fw_pwrv[3:0]), .test_si(regD4_1_), .test_se(
        test_se) );
  glreg_8_00000004 u0_regE4 ( .clk(clk), .arstz(n34), .we(we_228), .wdat({n252, 
        n240, n230, n224, n219, n168, n142, n133}), .rdat({r_pwrctl, 
        lt_regE4_3_0}), .test_si(r_srcctl[7]), .test_se(test_se) );
  glreg_8_0000001f u0_regE5 ( .clk(clk), .arstz(n28), .we(r_pwrv_upd), .wdat({
        n252, n240, n230, n225, n216, n168, n138, n114}), .rdat(
        r_fw_pwrv[11:4]), .test_si(r_pwrctl[7]), .test_se(test_se) );
  glreg_a0_54 u0_regE6 ( .clk(clk), .arstz(n42), .we(we_230), .wdat({n252, 
        n240, n230, n224, n219, n183, n142, n133}), .rdat(r_ccrx), .test_si(
        r_fw_pwrv[11]), .test_se(test_se) );
  glreg_a0_53 u0_regE7 ( .clk(clk), .arstz(n68), .we(we_231), .wdat({n252, 
        n240, n230, n224, n219, n183, n142, n133}), .rdat(r_ccctl), .test_si(
        r_ccrx[7]), .test_se(test_se) );
  glreg_a0_52 u0_regE8 ( .clk(clk), .arstz(n67), .we(we_232), .wdat({n252, 
        n240, n230, n224, n219, n183, n142, n133}), .rdat(r_comp_opt), 
        .test_si(r_ccctl[7]), .test_se(test_se) );
  glreg_a0_51 u0_regF5 ( .clk(clk), .arstz(n66), .we(we_245), .wdat({n249, 
        n240, n230, n224, n216, n183, n142, n133}), .rdat(r_cvctl), .test_si(
        r_comp_opt[7]), .test_se(test_se) );
  glreg_a0_50 u0_regF6 ( .clk(clk), .arstz(n62), .we(we_246), .wdat({n251, 
        n241, n228, n222, n217, n168, n138, n114}), .rdat(r_cctrx), .test_si(
        r_cvctl[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_regbank_a0_1 clk_gate_rstcnt_reg ( .CLK(clk), .EN(N26), 
        .ENCLK(net10832), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_regbank_a0_0 clk_gate_lg_pulse_cnt_reg ( .CLK(clk_1p0m), 
        .EN(N108), .ENCLK(net10838), .TE(test_se) );
  regbank_a0_DW01_add_0 add_525 ( .A(regAC), .B(regAB), .CI(1'b0), .SUM(
        r_pwr_i), .CO() );
  regbank_a0_DW01_inc_0 add_304 ( .A({1'b0, r_inst_ofs}), .SUM({
        SYNOPSYS_UNCONNECTED_1, inst_ofs_plus}) );
  regbank_a0_DW_rightsh_1 srl_133 ( .A({dac_r_vs, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, r_cctrx, r_cvctl, regF4_7_, x_daclsb[5:3], regF4_3, 
        x_daclsb[2:0], r_sar_en, r_dac_en, dac_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_comp_opt, r_ccctl, r_ccrx, r_fw_pwrv[11:4], r_pwrctl, r_fw_pwrv[3:0], 
        r_srcctl[7:4], regE3, r_srcctl[1], regE3_0, dac_r_cmpsta, dac_r_comp, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, regDF, regDE, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_ana_tm, r_fortxdat, 
        r_fortxrdy, r_fortxen, r_sleep, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, r_gpio_oe[3], r_gpio_s3, r_gpio_oe[2], r_gpio_s2, 
        r_gpio_oe[1], r_gpio_s1, r_gpio_oe[0], r_gpio_s0, r_gpio_pu[3:0], 
        r_gpio_pd[3:0], test_so2, regD4_6_, regD4_5_, regD4_4_, regD4_3_, 
        regD4_2_, regD4_1_, regD4_0_, regD3_7_, r_gpio_oe[5], r_gpio_pu[5], 
        r_gpio_pd[5], regD3_3, r_gpio_oe[4], r_gpio_pu[4], r_gpio_pd[4], 
        i_i2c_rwbuf, r_exist1st, r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, 
        r_gpio_oe[6], r_gpio_pu[6], r_gpio_pd[6], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, reg31, reg30, i_i2c_ltbuf, reg28, reg27, r_i2c_deva, 
        r_hwi2c_en, 1'b0, 1'b0, r_i2c_attr, r_pg0_sel, reg25_0_, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, prx_rcvinf[4], REVID, 
        prx_rcvinf[3], ptx_fsm, prx_fsm, reg21, r_dat_portrole, r_dat_spec, 
        r_dat_datarole, reg20, reg19_7_, r_inst_ofs, i_i2c_ofs, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, dbgpo[31:24], r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1], prl_cpmsgid, n12, 
        prx_rcvinf[2:0], prl_fsm, reg12, r_txshrt, reg12_1, r_pshords, 
        reg11_7_, r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0], 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, pff_empty, 
        pff_full, pff_ptr, reg06, reg05, dbgpo[15:0], pff_rdat, r_last, 
        r_first, r_unlock, r_txnumk, r_txendk, r_txauto, regAF, regAE, regAD_7, 
        1'b0, regAD, regAC, regAB, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_regtrm, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, fcp_r_crc, fcp_r_dat, fcp_r_msk, fcp_r_sta, 
        fcp_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, fcp_r_acc, r_accctl, fcp_r_tui, reg94, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, r_isofs, r_adofs, r_dpdmctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_cvofs, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .DATA_TC(1'b0), .SH({n107, sfr_addr[5:0], 
        1'b0, 1'b0, 1'b0}), .B({SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, 
        SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, 
        SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, 
        SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, 
        SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, 
        SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, 
        SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, 
        SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, 
        SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, 
        SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, 
        SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, 
        SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, 
        SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, 
        SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, 
        SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, 
        SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, 
        SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, 
        SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, 
        SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, 
        SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, 
        SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, 
        SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, 
        SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, 
        SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, 
        SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, 
        SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, 
        SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, 
        SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, 
        SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, 
        SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, 
        SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, 
        SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, 
        SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, 
        SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, 
        SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, 
        SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, 
        SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, 
        SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, 
        SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, 
        SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, 
        SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, 
        SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, 
        SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, 
        SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, 
        SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, 
        SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, 
        SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, 
        SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, 
        SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, 
        SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, 
        SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, 
        SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, 
        SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, 
        SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, 
        SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, 
        SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, 
        SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, 
        SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, 
        SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, 
        SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, 
        SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, 
        SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, 
        SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, 
        SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, 
        SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, 
        SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, 
        SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, 
        SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, 
        SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, 
        SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, 
        SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, 
        SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, 
        SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, 
        SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, 
        SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, 
        SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, 
        SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, 
        SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, 
        SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, 
        SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, 
        SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, 
        SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, 
        SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, 
        SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, 
        SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, 
        SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, 
        SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, 
        SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, 
        SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, 
        SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, 
        SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, 
        SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, 
        SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, 
        SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, 
        SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, 
        SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, 
        SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, 
        SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, 
        SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, 
        SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, 
        SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, 
        SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, 
        SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, 
        SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, 
        SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, 
        SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, 
        SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, 
        SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, 
        SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, 
        SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, 
        SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, 
        SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, 
        SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, 
        SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, 
        SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, 
        SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, 
        SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, 
        SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, 
        SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, 
        SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, 
        SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, 
        SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, 
        SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, 
        SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, 
        SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, 
        SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, 
        SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, 
        SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, 
        SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, 
        SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, 
        SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, 
        SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, 
        SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, 
        SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, 
        SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, 
        SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, 
        SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, 
        SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, 
        SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, 
        SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, 
        SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, 
        SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, 
        SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, 
        SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, 
        SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, 
        SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, 
        SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, 
        SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, 
        SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, 
        SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, 
        SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, 
        SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, 
        SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, 
        SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, 
        SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, 
        SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, 
        SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, 
        SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, 
        SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, 
        SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, 
        SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, 
        SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, 
        SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, 
        SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, 
        SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, 
        SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, 
        SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, 
        SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, 
        SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, 
        SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, 
        SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, 
        SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, 
        SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, 
        SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, 
        SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, 
        SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, 
        SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, 
        SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, 
        SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, 
        SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, 
        SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, 
        SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, 
        SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, 
        SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, 
        SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, 
        SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, 
        SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, 
        SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, 
        SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, 
        SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, 
        SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, 
        SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, 
        SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, 
        SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, 
        SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, 
        SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, 
        SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, 
        SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, 
        SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, 
        SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, 
        SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, 
        SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, 
        SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, 
        SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, 
        SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, 
        SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, 
        SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, 
        SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, 
        SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, 
        SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, 
        SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, 
        SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, 
        SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, 
        SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, 
        SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, 
        SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, 
        SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, 
        SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, 
        SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, 
        SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, 
        SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, 
        SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, 
        SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, 
        SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, 
        SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, 
        SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, 
        SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, 
        SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, 
        SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, 
        SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, 
        SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, 
        SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, 
        SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, 
        SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, 
        SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, 
        SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, 
        SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, 
        SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, 
        SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, 
        SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, 
        SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, 
        SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, 
        SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, 
        SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, 
        SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, 
        SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, 
        SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, 
        SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, 
        SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, 
        SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, 
        SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, 
        SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, 
        SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, 
        SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, 
        SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, 
        SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, 
        SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, 
        SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, 
        SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, 
        SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, 
        SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, 
        SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, 
        SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, 
        SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, 
        SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, 
        SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, 
        SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, 
        SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, 
        SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, 
        SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, 
        SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, 
        SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, 
        SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, 
        SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, 
        SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, 
        SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, 
        SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, 
        SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, 
        SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, 
        SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017, sfr_rdat}) );
  SDFFRQX1 r_phyrst_reg_0_ ( .D(n1222), .SIN(oscdwn_shft[2]), .SMC(test_se), 
        .C(clk), .XR(n2), .Q(r_phyrst[0]) );
  SDFFRQX1 lg_pulse_cnt_reg_3_ ( .D(N112), .SIN(lg_pulse_cnt[2]), .SMC(test_se), .C(net10838), .XR(n86), .Q(lg_pulse_cnt[3]) );
  SDFFRQX1 lg_pulse_cnt_reg_4_ ( .D(N113), .SIN(lg_pulse_cnt[3]), .SMC(test_se), .C(net10838), .XR(n86), .Q(lg_pulse_cnt[4]) );
  SDFFRQX1 lg_pulse_cnt_reg_1_ ( .D(N110), .SIN(lg_pulse_cnt[0]), .SMC(test_se), .C(net10838), .XR(n87), .Q(lg_pulse_cnt[1]) );
  SDFFRQX1 lg_pulse_cnt_reg_2_ ( .D(N111), .SIN(lg_pulse_cnt[1]), .SMC(test_se), .C(net10838), .XR(n101), .Q(lg_pulse_cnt[2]) );
  SDFFRQX1 rstcnt_reg_0_ ( .D(N39), .SIN(r_phyrst[1]), .SMC(test_se), .C(
        net10832), .XR(n3), .Q(rstcnt[0]) );
  SDFFRQX1 lg_pulse_cnt_reg_0_ ( .D(N109), .SIN(lg_pulse_12m), .SMC(test_se), 
        .C(net10838), .XR(n86), .Q(lg_pulse_cnt[0]) );
  SDFFRQX1 d_p0_reg_7_ ( .D(ff_p0[7]), .SIN(d_p0[6]), .SMC(test_se), .C(clk), 
        .XR(n87), .Q(d_p0[7]) );
  SDFFRQX1 d_p0_reg_6_ ( .D(ff_p0[6]), .SIN(d_p0[5]), .SMC(test_se), .C(clk), 
        .XR(n87), .Q(d_p0[6]) );
  SDFFRQX1 d_p0_reg_5_ ( .D(ff_p0[5]), .SIN(d_p0[4]), .SMC(test_se), .C(clk), 
        .XR(n87), .Q(d_p0[5]) );
  SDFFRQX1 d_p0_reg_4_ ( .D(ff_p0[4]), .SIN(d_p0[3]), .SMC(test_se), .C(clk), 
        .XR(n87), .Q(d_p0[4]) );
  SDFFRQX1 d_p0_reg_3_ ( .D(ff_p0[3]), .SIN(d_p0[2]), .SMC(test_se), .C(clk), 
        .XR(n87), .Q(d_p0[3]) );
  SDFFRQX1 d_p0_reg_2_ ( .D(ff_p0[2]), .SIN(d_p0[1]), .SMC(test_se), .C(clk), 
        .XR(n87), .Q(d_p0[2]) );
  SDFFRQX1 d_p0_reg_1_ ( .D(ff_p0[1]), .SIN(d_p0[0]), .SMC(test_se), .C(clk), 
        .XR(n87), .Q(d_p0[1]) );
  SDFFRQX1 d_p0_reg_0_ ( .D(ff_p0[0]), .SIN(test_si2), .SMC(test_se), .C(clk), 
        .XR(n87), .Q(d_p0[0]) );
  SDFFRQX1 r_phyrst_reg_1_ ( .D(n1221), .SIN(r_phyrst[0]), .SMC(test_se), .C(
        clk), .XR(n2), .Q(r_phyrst[1]) );
  SDFFNRQX1 osc_gate_n_reg_3_ ( .D(osc_gate_n_2_), .SIN(osc_gate_n_2_), .SMC(
        test_se), .XC(xclk), .XR(n3), .Q(test_so1) );
  SDFFNRQX1 osc_gate_n_reg_0_ ( .D(r_pos_gate), .SIN(test_si1), .SMC(test_se), 
        .XC(xclk), .XR(n2), .Q(osc_gate_n_0_) );
  SDFFNRQX1 osc_gate_n_reg_1_ ( .D(osc_gate_n_0_), .SIN(osc_gate_n_0_), .SMC(
        test_se), .XC(xclk), .XR(n3), .Q(osc_gate_n_1_) );
  SDFFNRQX1 osc_gate_n_reg_2_ ( .D(osc_gate_n_1_), .SIN(osc_gate_n_1_), .SMC(
        test_se), .XC(xclk), .XR(n2), .Q(osc_gate_n_2_) );
  SDFFQX1 oscdwn_shft_reg_1_ ( .D(oscdwn_shft[0]), .SIN(oscdwn_shft[0]), .SMC(
        test_se), .C(clk), .Q(oscdwn_shft[1]) );
  SDFFRQX1 rstcnt_reg_3_ ( .D(N36), .SIN(rstcnt[2]), .SMC(test_se), .C(
        net10832), .XR(n3), .Q(rstcnt[3]) );
  SDFFRQX1 lg_pulse_reg ( .D(n1220), .SIN(lg_pulse_cnt[4]), .SMC(test_se), .C(
        clk_1p0m), .XR(n86), .Q(lg_dischg) );
  SDFFRQX1 drstz_reg_1_ ( .D(drstz[0]), .SIN(drstz[0]), .SMC(test_se), .C(clk), 
        .XR(n2), .Q(drstz[1]) );
  SDFFRQX1 lg_pulse_12m_reg ( .D(n1219), .SIN(drstz[1]), .SMC(test_se), .C(clk), .XR(n87), .Q(lg_pulse_12m) );
  SDFFRQX1 rstcnt_reg_1_ ( .D(N38), .SIN(rstcnt[0]), .SMC(test_se), .C(
        net10832), .XR(n3), .Q(rstcnt[1]) );
  SDFFRQX1 rstcnt_reg_2_ ( .D(N37), .SIN(rstcnt[1]), .SMC(test_se), .C(
        net10832), .XR(n2), .Q(rstcnt[2]) );
  SDFFRQX1 rstcnt_reg_4_ ( .D(N35), .SIN(rstcnt[3]), .SMC(test_se), .C(
        net10832), .XR(n3), .Q(rstcnt[4]) );
  SDFFQX1 oscdwn_shft_reg_2_ ( .D(n377), .SIN(oscdwn_shft[1]), .SMC(test_se), 
        .C(clk), .Q(oscdwn_shft[2]) );
  OAI21X1 U434 ( .B(n211), .C(n413), .A(n259), .Y(srstz) );
  SDFFQX1 oscdwn_shft_reg_0_ ( .D(N84), .SIN(lg_dischg), .SMC(test_se), .C(clk), .Q(oscdwn_shft[0]) );
  SDFFRQX1 drstz_reg_0_ ( .D(1'b1), .SIN(d_p0[7]), .SMC(test_se), .C(clk), 
        .XR(n2), .Q(drstz[0]) );
  NOR3X1 U8 ( .A(n334), .B(n304), .C(n299), .Y(n18) );
  INVX1 U9 ( .A(sfr_addr[6]), .Y(n110) );
  INVX2 U10 ( .A(n110), .Y(n107) );
  MUX2X1 U11 ( .D0(pff_rxpart[6]), .D1(n241), .S(n270), .Y(wd20[6]) );
  INVXL U12 ( .A(xrstz), .Y(n1) );
  INVXL U13 ( .A(n1), .Y(n2) );
  INVXL U14 ( .A(n1), .Y(n3) );
  INVXL U15 ( .A(n18), .Y(n9) );
  INVXL U16 ( .A(n9), .Y(n10) );
  NAND43X1 U17 ( .B(sfr_addr[5]), .C(sfr_addr[6]), .D(n372), .A(n371), .Y(n373) );
  INVX1 U18 ( .A(prl_cany0), .Y(n11) );
  INVX1 U19 ( .A(n11), .Y(n12) );
  INVX1 U20 ( .A(n380), .Y(n13) );
  INVX1 U21 ( .A(n388), .Y(n14) );
  BUFX3 U22 ( .A(n109), .Y(n15) );
  NOR2X1 U23 ( .A(n146), .B(prl_c0set), .Y(phyrst) );
  INVX1 U24 ( .A(phyrst), .Y(n16) );
  INVX1 U25 ( .A(phyrst), .Y(n17) );
  BUFX3 U26 ( .A(pff_ptr[0]), .Y(dbgpo[16]) );
  BUFX3 U27 ( .A(pff_ptr[4]), .Y(dbgpo[20]) );
  BUFX3 U28 ( .A(pff_ptr[2]), .Y(dbgpo[18]) );
  BUFX3 U29 ( .A(pff_ptr[5]), .Y(dbgpo[21]) );
  BUFX3 U30 ( .A(pff_ptr[3]), .Y(dbgpo[19]) );
  BUFX3 U31 ( .A(pff_ptr[1]), .Y(dbgpo[17]) );
  NAND21XL U32 ( .B(n305), .A(n341), .Y(n306) );
  NAND21XL U33 ( .B(n341), .A(n302), .Y(n303) );
  NAND21XL U34 ( .B(n300), .A(n341), .Y(n263) );
  NAND21XL U35 ( .B(n268), .A(n341), .Y(n260) );
  INVXL U36 ( .A(sfr_addr[5]), .Y(n106) );
  INVXL U37 ( .A(sfr_addr[6]), .Y(n108) );
  NAND21XL U38 ( .B(n262), .A(sfr_addr[2]), .Y(n268) );
  NAND21XL U39 ( .B(n262), .A(sfr_addr[1]), .Y(n346) );
  NAND21XL U40 ( .B(n262), .A(sfr_addr[4]), .Y(n294) );
  NAND21XL U41 ( .B(n262), .A(sfr_addr[0]), .Y(n279) );
  NAND21XL U42 ( .B(n262), .A(sfr_addr[3]), .Y(n371) );
  NAND43XL U43 ( .B(n391), .C(n343), .D(n342), .A(n341), .Y(n344) );
  MUX2XL U44 ( .D0(i_pc[4]), .D1(prx_adpn[4]), .S(reg19_7_), .Y(reg30[4]) );
  MUX2XL U45 ( .D0(i_pc[3]), .D1(prx_adpn[3]), .S(reg19_7_), .Y(reg30[3]) );
  MUX2XL U46 ( .D0(i_pc[1]), .D1(prx_adpn[1]), .S(reg19_7_), .Y(reg30[1]) );
  MUX2XL U47 ( .D0(i_pc[0]), .D1(prx_adpn[0]), .S(reg19_7_), .Y(reg30[0]) );
  MUX2XL U48 ( .D0(i_pc[2]), .D1(prx_adpn[2]), .S(reg19_7_), .Y(reg30[2]) );
  NAND41X1 U49 ( .D(n12), .A(prx_rcvinf[4]), .B(i_i2c_idle), .C(n204), .Y(n180) );
  ENOXL U50 ( .A(n214), .B(n117), .C(r_txnumk[2]), .D(n117), .Y(wd01[2]) );
  ENOXL U51 ( .A(n144), .B(n14), .C(r_txnumk[1]), .D(n117), .Y(wd01[1]) );
  ENOXL U52 ( .A(n226), .B(n14), .C(r_txnumk[4]), .D(n117), .Y(wd01[4]) );
  MUX2XL U53 ( .D0(r_txnumk[3]), .D1(n220), .S(n388), .Y(wd01[3]) );
  INVX1 U54 ( .A(n253), .Y(n249) );
  INVX1 U55 ( .A(n246), .Y(n240) );
  INVX1 U56 ( .A(n256), .Y(n252) );
  INVX1 U57 ( .A(n255), .Y(n251) );
  INVX1 U58 ( .A(n245), .Y(n239) );
  INVX1 U59 ( .A(n244), .Y(n238) );
  INVX1 U60 ( .A(n254), .Y(n250) );
  INVX1 U61 ( .A(n221), .Y(n215) );
  INVX1 U62 ( .A(n221), .Y(n216) );
  BUFX3 U63 ( .A(n248), .Y(n243) );
  BUFX3 U64 ( .A(n258), .Y(n253) );
  NAND2X1 U65 ( .A(n136), .B(n184), .Y(n135) );
  NOR3XL U66 ( .A(n140), .B(n227), .C(n184), .Y(r_discard) );
  INVX1 U67 ( .A(n351), .Y(we_227) );
  INVX1 U68 ( .A(n381), .Y(n379) );
  AND2X1 U69 ( .A(n359), .B(n358), .Y(r_dacwr[12]) );
  INVX1 U70 ( .A(n214), .Y(n168) );
  INVX1 U71 ( .A(n389), .Y(n213) );
  INVX1 U72 ( .A(n137), .Y(n114) );
  INVX1 U73 ( .A(n144), .Y(n138) );
  AND2X1 U74 ( .A(n367), .B(n366), .Y(r_fcpwr[0]) );
  AND2X1 U75 ( .A(n286), .B(n366), .Y(we_171) );
  AND2X1 U76 ( .A(n366), .B(n329), .Y(we_187) );
  INVX1 U77 ( .A(n214), .Y(n183) );
  INVX1 U78 ( .A(n221), .Y(n219) );
  INVX1 U79 ( .A(n137), .Y(n133) );
  INVX1 U80 ( .A(n144), .Y(n142) );
  BUFX3 U81 ( .A(n254), .Y(n256) );
  BUFX3 U82 ( .A(n242), .Y(n245) );
  BUFX3 U83 ( .A(n258), .Y(n254) );
  BUFX3 U84 ( .A(n242), .Y(n244) );
  BUFX3 U85 ( .A(n242), .Y(n246) );
  BUFX3 U86 ( .A(n254), .Y(n255) );
  BUFX3 U87 ( .A(n244), .Y(n247) );
  BUFX3 U88 ( .A(n254), .Y(n257) );
  INVX1 U89 ( .A(n226), .Y(n225) );
  INVX1 U90 ( .A(n221), .Y(n220) );
  INVX1 U91 ( .A(n242), .Y(n241) );
  INVX1 U92 ( .A(n227), .Y(n224) );
  INVX1 U93 ( .A(n144), .Y(n141) );
  INVX1 U94 ( .A(n221), .Y(n218) );
  INVX1 U95 ( .A(n214), .Y(n172) );
  INVX1 U96 ( .A(n227), .Y(n223) );
  INVX1 U97 ( .A(n137), .Y(n121) );
  INVX1 U98 ( .A(n144), .Y(n139) );
  INVX1 U99 ( .A(n214), .Y(n169) );
  INVX1 U100 ( .A(n221), .Y(n217) );
  INVX1 U101 ( .A(n227), .Y(n222) );
  INVX1 U102 ( .A(n137), .Y(n116) );
  INVX1 U103 ( .A(n98), .Y(n86) );
  INVX1 U104 ( .A(n89), .Y(n87) );
  INVX1 U105 ( .A(n90), .Y(n79) );
  INVX1 U106 ( .A(n88), .Y(n84) );
  INVX1 U107 ( .A(n93), .Y(n69) );
  INVX1 U108 ( .A(n93), .Y(n49) );
  INVX1 U109 ( .A(n102), .Y(n43) );
  INVX1 U110 ( .A(n98), .Y(n37) );
  INVX1 U111 ( .A(n102), .Y(n62) );
  INVX1 U112 ( .A(n91), .Y(n66) );
  INVX1 U113 ( .A(n93), .Y(n67) );
  INVX1 U114 ( .A(n93), .Y(n68) );
  INVX1 U115 ( .A(n97), .Y(n42) );
  INVX1 U116 ( .A(n92), .Y(n70) );
  INVX1 U117 ( .A(n89), .Y(n81) );
  INVX1 U118 ( .A(n89), .Y(n82) );
  INVX1 U119 ( .A(n89), .Y(n80) );
  INVX1 U120 ( .A(n88), .Y(n85) );
  INVX1 U121 ( .A(n94), .Y(n59) );
  INVX1 U122 ( .A(n94), .Y(n60) );
  INVX1 U123 ( .A(n95), .Y(n57) );
  INVX1 U124 ( .A(n95), .Y(n56) );
  INVX1 U125 ( .A(n95), .Y(n55) );
  INVX1 U126 ( .A(n94), .Y(n58) );
  INVX1 U127 ( .A(n96), .Y(n53) );
  INVX1 U128 ( .A(n96), .Y(n52) );
  INVX1 U129 ( .A(n88), .Y(n83) );
  INVX1 U130 ( .A(n96), .Y(n54) );
  INVX1 U131 ( .A(n102), .Y(n48) );
  INVX1 U132 ( .A(n97), .Y(n47) );
  INVX1 U133 ( .A(n89), .Y(n44) );
  INVX1 U134 ( .A(n92), .Y(n50) );
  INVX1 U135 ( .A(n88), .Y(n51) );
  INVX1 U136 ( .A(n98), .Y(n61) );
  INVX1 U137 ( .A(n97), .Y(n41) );
  INVX1 U138 ( .A(n95), .Y(n46) );
  INVX1 U139 ( .A(n97), .Y(n40) );
  INVX1 U140 ( .A(n90), .Y(n63) );
  INVX1 U141 ( .A(n98), .Y(n39) );
  INVX1 U142 ( .A(n98), .Y(n38) );
  INVX1 U143 ( .A(n91), .Y(n45) );
  INVX1 U144 ( .A(n90), .Y(n64) );
  INVX1 U145 ( .A(n94), .Y(n65) );
  INVX1 U146 ( .A(n92), .Y(n71) );
  INVX1 U147 ( .A(n91), .Y(n73) );
  INVX1 U148 ( .A(n92), .Y(n72) );
  INVX1 U149 ( .A(n91), .Y(n74) );
  INVX1 U150 ( .A(n90), .Y(n76) );
  INVX1 U151 ( .A(n90), .Y(n78) );
  INVX1 U152 ( .A(n91), .Y(n75) );
  INVX1 U153 ( .A(atpg_en), .Y(n259) );
  INVX1 U154 ( .A(sfr_wdat[3]), .Y(n221) );
  AND2X1 U155 ( .A(n356), .B(n374), .Y(r_dacwr[4]) );
  AND2X1 U156 ( .A(n356), .B(n366), .Y(r_dacwr[3]) );
  AND2X1 U157 ( .A(n356), .B(n375), .Y(r_dacwr[5]) );
  AND2X1 U158 ( .A(n357), .B(n361), .Y(r_dacwr[8]) );
  INVX1 U159 ( .A(n326), .Y(n366) );
  AND2X1 U160 ( .A(n356), .B(n359), .Y(r_dacwr[2]) );
  AND2X1 U161 ( .A(n356), .B(n361), .Y(r_dacwr[1]) );
  AND2X1 U162 ( .A(n356), .B(n368), .Y(r_dacwr[7]) );
  AND2X1 U163 ( .A(n356), .B(n370), .Y(r_dacwr[6]) );
  INVX1 U164 ( .A(n289), .Y(n359) );
  INVX1 U165 ( .A(n304), .Y(n272) );
  INVX1 U166 ( .A(n342), .Y(n333) );
  INVX1 U167 ( .A(n232), .Y(n228) );
  INVX1 U168 ( .A(sfr_wdat[7]), .Y(n258) );
  INVX1 U169 ( .A(sfr_wdat[1]), .Y(n143) );
  INVX1 U170 ( .A(sfr_wdat[4]), .Y(n227) );
  INVX1 U171 ( .A(sfr_wdat[2]), .Y(n184) );
  INVX1 U172 ( .A(sfr_wdat[0]), .Y(n136) );
  AND2X1 U173 ( .A(n367), .B(n370), .Y(r_fcpwr[3]) );
  NAND5XL U174 ( .A(n241), .B(n249), .C(n215), .D(n137), .E(n378), .Y(n140) );
  INVX1 U175 ( .A(n134), .Y(n378) );
  INVX1 U176 ( .A(n365), .Y(n367) );
  NAND21X1 U177 ( .B(n364), .A(n363), .Y(n365) );
  NAND21X1 U178 ( .B(n326), .A(n358), .Y(n351) );
  NAND21X1 U179 ( .B(n328), .A(n374), .Y(n381) );
  NAND21X1 U180 ( .B(n289), .A(n348), .Y(n389) );
  AND2X1 U181 ( .A(n369), .B(n375), .Y(r_fcpwr[4]) );
  AND2X1 U182 ( .A(n367), .B(n374), .Y(r_fcpwr[1]) );
  NAND21X1 U183 ( .B(n326), .A(n327), .Y(n123) );
  AND2X1 U184 ( .A(n325), .B(n228), .Y(clr28[5]) );
  AND2X1 U185 ( .A(n325), .B(n138), .Y(clr28[1]) );
  AND2X1 U186 ( .A(n336), .B(n228), .Y(clr04[5]) );
  AND2X1 U187 ( .A(n336), .B(n138), .Y(clr04[1]) );
  AND2X1 U188 ( .A(n325), .B(n225), .Y(clr28[4]) );
  AND2X1 U189 ( .A(n325), .B(n114), .Y(clr28[0]) );
  AND2X1 U190 ( .A(n336), .B(n225), .Y(clr04[4]) );
  AND2X1 U191 ( .A(n336), .B(n114), .Y(clr04[0]) );
  NOR2X1 U192 ( .A(n233), .B(n182), .Y(clrAE[5]) );
  NOR2X1 U193 ( .A(n143), .B(n182), .Y(clrAE[1]) );
  NOR2X1 U194 ( .A(n232), .B(n181), .Y(clrDF[5]) );
  NOR2X1 U195 ( .A(n143), .B(n181), .Y(clrDF[1]) );
  NOR2X1 U196 ( .A(n234), .B(n185), .Y(clr03[5]) );
  NOR2X1 U197 ( .A(n144), .B(n185), .Y(clr03[1]) );
  NOR2X1 U198 ( .A(n254), .B(n390), .Y(r_i2c_fwack) );
  NOR2X1 U199 ( .A(n226), .B(n182), .Y(clrAE[4]) );
  NOR2X1 U200 ( .A(n137), .B(n182), .Y(clrAE[0]) );
  NOR2X1 U201 ( .A(n226), .B(n181), .Y(clrDF[4]) );
  NOR2X1 U202 ( .A(n136), .B(n181), .Y(clrDF[0]) );
  NOR2X1 U203 ( .A(n226), .B(n185), .Y(clr03[4]) );
  NOR2X1 U204 ( .A(n137), .B(n185), .Y(clr03[0]) );
  NOR2X1 U205 ( .A(n245), .B(n182), .Y(clrAE[6]) );
  NOR2X1 U206 ( .A(n214), .B(n182), .Y(clrAE[2]) );
  NOR2X1 U207 ( .A(n244), .B(n181), .Y(clrDF[6]) );
  NOR2X1 U208 ( .A(n184), .B(n181), .Y(clrDF[2]) );
  NOR2X1 U209 ( .A(n246), .B(n185), .Y(clr03[6]) );
  NOR2X1 U210 ( .A(n214), .B(n185), .Y(clr03[2]) );
  AND2X1 U211 ( .A(n357), .B(n374), .Y(r_dacwr[11]) );
  INVX1 U212 ( .A(n280), .Y(n358) );
  AND2X1 U213 ( .A(n325), .B(n241), .Y(clr28[6]) );
  AND2X1 U214 ( .A(n325), .B(n168), .Y(clr28[2]) );
  AND2X1 U215 ( .A(n336), .B(n241), .Y(clr04[6]) );
  AND2X1 U216 ( .A(n336), .B(n168), .Y(clr04[2]) );
  AND2X1 U217 ( .A(n325), .B(n249), .Y(clr28[7]) );
  AND2X1 U218 ( .A(n325), .B(n215), .Y(clr28[3]) );
  AND2X1 U219 ( .A(n336), .B(n249), .Y(clr04[7]) );
  AND2X1 U220 ( .A(n336), .B(n215), .Y(clr04[3]) );
  NOR21XL U221 ( .B(n215), .A(n182), .Y(clrAE[3]) );
  NOR21XL U222 ( .B(n215), .A(n181), .Y(clrDF[3]) );
  NOR21XL U223 ( .B(n215), .A(n185), .Y(clr03[3]) );
  AND2X1 U224 ( .A(n368), .B(n367), .Y(r_fcpwr[5]) );
  INVX1 U225 ( .A(n271), .Y(r_set_cpmsgid) );
  NAND21X1 U226 ( .B(n328), .A(n370), .Y(n271) );
  INVX1 U227 ( .A(n281), .Y(r_pwrv_upd) );
  NAND21X1 U228 ( .B(n280), .A(n375), .Y(n281) );
  INVX1 U229 ( .A(sfr_wdat[0]), .Y(n137) );
  INVX1 U230 ( .A(sfr_wdat[2]), .Y(n214) );
  NOR2X1 U231 ( .A(n254), .B(n182), .Y(clrAE[7]) );
  NOR2X1 U232 ( .A(n253), .B(n181), .Y(clrDF[7]) );
  NOR2X1 U233 ( .A(n255), .B(n185), .Y(clr03[7]) );
  AO21X1 U234 ( .B(n327), .C(n359), .A(n103), .Y(upd18) );
  AND2X1 U235 ( .A(n358), .B(n374), .Y(we_228) );
  AND2X1 U236 ( .A(n286), .B(n374), .Y(we_172) );
  AND2X1 U237 ( .A(n291), .B(n374), .Y(we[164]) );
  AND2X1 U238 ( .A(n369), .B(n374), .Y(we_148) );
  INVX1 U239 ( .A(n284), .Y(n286) );
  NAND21X1 U240 ( .B(n364), .A(n283), .Y(n284) );
  AND2X1 U241 ( .A(n367), .B(n375), .Y(r_fcpwr[2]) );
  AND2X1 U242 ( .A(n357), .B(n375), .Y(we_245) );
  AND2X1 U243 ( .A(n291), .B(n375), .Y(we[165]) );
  AND2X1 U244 ( .A(n361), .B(n369), .Y(r_dacwr[14]) );
  AND2X1 U245 ( .A(n291), .B(n361), .Y(we[161]) );
  AND2X1 U246 ( .A(n298), .B(n361), .Y(we_217) );
  INVX1 U247 ( .A(sfr_wdat[4]), .Y(n226) );
  AND2X1 U248 ( .A(n332), .B(n331), .Y(we_181) );
  AND2X1 U249 ( .A(n298), .B(n370), .Y(we_222) );
  AND2X1 U250 ( .A(n330), .B(n331), .Y(we_182) );
  AND2X1 U251 ( .A(n357), .B(n366), .Y(r_dacwr[10]) );
  AND2X1 U252 ( .A(n357), .B(n359), .Y(r_dacwr[9]) );
  AND2X1 U253 ( .A(n357), .B(n370), .Y(we_246) );
  AND2X1 U254 ( .A(n286), .B(n368), .Y(we_175) );
  AND2X1 U255 ( .A(n368), .B(n358), .Y(we_231) );
  AND2X1 U256 ( .A(n368), .B(n329), .Y(we_191) );
  AND2X1 U257 ( .A(n291), .B(n368), .Y(we[167]) );
  AND2X1 U258 ( .A(n291), .B(n370), .Y(we[166]) );
  AND2X1 U259 ( .A(n291), .B(n366), .Y(we[163]) );
  AND2X1 U260 ( .A(n291), .B(n359), .Y(we[162]) );
  AND2X1 U261 ( .A(n370), .B(n369), .Y(r_fcpwr[6]) );
  AND2X1 U262 ( .A(n370), .B(n358), .Y(we_230) );
  AND2X1 U263 ( .A(n348), .B(n366), .Y(we_203) );
  INVX1 U264 ( .A(n390), .Y(n212) );
  BUFX3 U265 ( .A(n248), .Y(n242) );
  INVX1 U266 ( .A(sfr_wdat[6]), .Y(n248) );
  INVX1 U267 ( .A(sfr_wdat[1]), .Y(n144) );
  INVX1 U268 ( .A(n235), .Y(n230) );
  INVX1 U269 ( .A(n234), .Y(n229) );
  INVX1 U270 ( .A(n328), .Y(n329) );
  INVX1 U271 ( .A(n99), .Y(n28) );
  INVX1 U272 ( .A(n99), .Y(n29) );
  INVX1 U273 ( .A(n99), .Y(n30) );
  INVX1 U274 ( .A(n102), .Y(n31) );
  INVX1 U275 ( .A(n99), .Y(n33) );
  INVX1 U276 ( .A(n147), .Y(n32) );
  INVX1 U277 ( .A(n96), .Y(n34) );
  INVX1 U278 ( .A(n96), .Y(n35) );
  INVX1 U279 ( .A(n94), .Y(n36) );
  INVX1 U280 ( .A(n100), .Y(n93) );
  INVX1 U281 ( .A(n101), .Y(n89) );
  INVX1 U282 ( .A(n100), .Y(n95) );
  INVX1 U283 ( .A(n382), .Y(n94) );
  INVX1 U284 ( .A(n382), .Y(n88) );
  INVX1 U285 ( .A(n101), .Y(n96) );
  INVX1 U286 ( .A(n100), .Y(n92) );
  INVX1 U287 ( .A(n101), .Y(n91) );
  INVX1 U288 ( .A(n382), .Y(n97) );
  INVX1 U289 ( .A(n101), .Y(n90) );
  INVX1 U290 ( .A(n101), .Y(n98) );
  INVX1 U291 ( .A(n299), .Y(n363) );
  INVX1 U292 ( .A(n274), .Y(n375) );
  NAND21X1 U293 ( .B(n305), .A(n282), .Y(n326) );
  INVX1 U294 ( .A(n290), .Y(n361) );
  NAND21X1 U295 ( .B(n343), .A(n282), .Y(n289) );
  AND2X1 U296 ( .A(n356), .B(n360), .Y(r_dacwr[0]) );
  INVX1 U297 ( .A(n285), .Y(n370) );
  INVX1 U298 ( .A(n297), .Y(n368) );
  INVX1 U299 ( .A(n273), .Y(n357) );
  NAND21X1 U300 ( .B(n354), .A(n272), .Y(n273) );
  INVX1 U301 ( .A(n305), .Y(n307) );
  NAND21X1 U302 ( .B(n340), .A(n392), .Y(r_fiforst) );
  INVX1 U303 ( .A(prl_c0set), .Y(n392) );
  NOR6XL U304 ( .A(n135), .B(n216), .C(n134), .D(n249), .E(sfr_wdat[4]), .F(
        n241), .Y(n340) );
  NAND43X1 U305 ( .B(n347), .C(n339), .D(n228), .A(n143), .Y(n134) );
  INVX1 U306 ( .A(n355), .Y(n356) );
  NAND21X1 U307 ( .B(n354), .A(n353), .Y(n355) );
  INVX1 U308 ( .A(n339), .Y(n362) );
  INVX1 U309 ( .A(n261), .Y(n330) );
  NAND21X1 U310 ( .B(n265), .A(n278), .Y(n261) );
  INVX1 U311 ( .A(n275), .Y(n353) );
  INVX1 U312 ( .A(n127), .Y(r_fifopsh) );
  INVX1 U313 ( .A(n343), .Y(n345) );
  BUFX3 U314 ( .A(n237), .Y(n232) );
  INVX1 U315 ( .A(n264), .Y(n348) );
  NAND32X1 U316 ( .B(n372), .C(n275), .A(n106), .Y(n264) );
  INVX1 U317 ( .A(n324), .Y(n325) );
  INVX1 U318 ( .A(n335), .Y(n336) );
  NAND21X1 U319 ( .B(n347), .A(n337), .Y(n185) );
  NAND21X1 U320 ( .B(n285), .A(n286), .Y(n182) );
  NAND21X1 U321 ( .B(n297), .A(n298), .Y(n181) );
  NAND21X1 U322 ( .B(n123), .A(n105), .Y(n111) );
  NAND21X1 U323 ( .B(n290), .A(n348), .Y(n390) );
  INVX1 U324 ( .A(n293), .Y(n369) );
  NAND32X1 U325 ( .B(n292), .C(n299), .A(n108), .Y(n293) );
  INVX1 U326 ( .A(n269), .Y(n270) );
  NAND21X1 U327 ( .B(n274), .A(n327), .Y(n109) );
  NAND21X1 U328 ( .B(n287), .A(n272), .Y(n280) );
  INVX1 U329 ( .A(n117), .Y(n388) );
  INVX1 U330 ( .A(n267), .Y(n327) );
  NAND32X1 U331 ( .B(n372), .C(n304), .A(n106), .Y(n267) );
  INVX1 U332 ( .A(n287), .Y(n283) );
  OR2X1 U333 ( .A(n364), .B(n354), .Y(n328) );
  AND2X1 U334 ( .A(n376), .B(n374), .Y(r_cvcwr[0]) );
  AND3X1 U335 ( .A(n353), .B(n283), .C(n360), .Y(we_232) );
  INVX1 U336 ( .A(n296), .Y(n298) );
  NAND21X1 U337 ( .B(n299), .A(n353), .Y(n296) );
  INVX1 U338 ( .A(n347), .Y(n331) );
  INVX1 U339 ( .A(n306), .Y(n337) );
  AND2X1 U340 ( .A(n376), .B(n375), .Y(r_cvcwr[1]) );
  AND2X1 U341 ( .A(n360), .B(n369), .Y(r_dacwr[13]) );
  AND2X1 U342 ( .A(n323), .B(n362), .Y(we_215) );
  AND2X1 U343 ( .A(n323), .B(n330), .Y(we_214) );
  AND2X1 U344 ( .A(n323), .B(n332), .Y(we_213) );
  AND2X1 U345 ( .A(n323), .B(n337), .Y(we_211) );
  INVX1 U346 ( .A(n288), .Y(n291) );
  NAND32X1 U347 ( .B(n292), .C(n287), .A(n108), .Y(n288) );
  BUFX3 U348 ( .A(n237), .Y(n234) );
  BUFX3 U349 ( .A(n237), .Y(n233) );
  INVX1 U350 ( .A(n303), .Y(n332) );
  BUFX3 U351 ( .A(n233), .Y(n235) );
  BUFX3 U352 ( .A(n234), .Y(n236) );
  INVX1 U353 ( .A(N33), .Y(n409) );
  INVX1 U354 ( .A(n105), .Y(n103) );
  INVX1 U355 ( .A(n105), .Y(n104) );
  INVX1 U356 ( .A(n147), .Y(n101) );
  INVX1 U357 ( .A(n88), .Y(n100) );
  INVX1 U358 ( .A(n100), .Y(n99) );
  NAND32X1 U359 ( .B(n276), .C(n268), .A(n279), .Y(n334) );
  INVX1 U360 ( .A(n371), .Y(n292) );
  INVX1 U361 ( .A(n294), .Y(n372) );
  INVX1 U362 ( .A(n346), .Y(n341) );
  INVX1 U363 ( .A(n263), .Y(n282) );
  NAND2X1 U364 ( .A(n268), .B(n265), .Y(n305) );
  NAND21X1 U365 ( .B(n300), .A(n330), .Y(n285) );
  NAND21X1 U366 ( .B(n300), .A(n362), .Y(n297) );
  INVX1 U367 ( .A(n277), .Y(n360) );
  NAND21X1 U368 ( .B(n300), .A(n333), .Y(n347) );
  NAND21X1 U369 ( .B(n279), .A(n278), .Y(n339) );
  INVX1 U370 ( .A(n279), .Y(n265) );
  INVX1 U371 ( .A(n260), .Y(n278) );
  INVX1 U372 ( .A(n266), .Y(n302) );
  NAND21X1 U373 ( .B(n268), .A(n265), .Y(n266) );
  NAND21X1 U374 ( .B(n265), .A(n268), .Y(n343) );
  NAND32X1 U375 ( .B(n347), .C(n346), .A(n345), .Y(n127) );
  AND3X1 U376 ( .A(n362), .B(sfr_r), .C(n350), .Y(r_psrd) );
  INVX1 U377 ( .A(sfr_wdat[5]), .Y(n237) );
  AND2X1 U378 ( .A(n350), .B(n368), .Y(r_pswr) );
  AND3X1 U379 ( .A(n369), .B(n362), .C(sfr_r), .Y(r_fcpre) );
  INVX1 U380 ( .A(n205), .Y(n387) );
  NAND32X1 U381 ( .B(n347), .C(n305), .A(n346), .Y(n117) );
  MUX2X1 U382 ( .D0(pff_rxpart[1]), .D1(n142), .S(n270), .Y(wd20[1]) );
  ENOX1 U383 ( .A(n109), .B(n257), .C(pff_rxpart[15]), .D(n109), .Y(wd21[7])
         );
  NAND4X1 U384 ( .A(n123), .B(n124), .C(n125), .D(n105), .Y(upd19) );
  AND4X1 U385 ( .A(n368), .B(n295), .C(n294), .D(n106), .Y(we_143) );
  INVX1 U386 ( .A(n364), .Y(n295) );
  AND3X1 U387 ( .A(n323), .B(n307), .C(n346), .Y(we_209) );
  AND3X1 U388 ( .A(n345), .B(n331), .C(n346), .Y(we_176) );
  INVX1 U389 ( .A(n301), .Y(n323) );
  NAND32X1 U390 ( .B(n300), .C(n304), .A(n363), .Y(n301) );
  INVX1 U391 ( .A(n373), .Y(n376) );
  INVX1 U392 ( .A(n122), .Y(n77) );
  XOR2X1 U393 ( .A(N34), .B(N35), .Y(N36) );
  XNOR2XL U394 ( .A(n409), .B(N32), .Y(N38) );
  XNOR2XL U395 ( .A(N34), .B(n409), .Y(N37) );
  INVX1 U396 ( .A(ictlr_inc), .Y(n105) );
  INVX1 U397 ( .A(n382), .Y(n102) );
  BUFX3 U398 ( .A(pff_empty), .Y(dbgpo[23]) );
  BUFX3 U399 ( .A(pff_full), .Y(dbgpo[22]) );
  NAND21X1 U400 ( .B(n341), .A(sfr_w), .Y(n276) );
  INVX1 U401 ( .A(n344), .Y(r_fifopop) );
  INVX1 U402 ( .A(n180), .Y(bus_idle) );
  NOR2X1 U403 ( .A(n243), .B(n390), .Y(r_i2c_fwnak) );
  INVX1 U404 ( .A(n349), .Y(n350) );
  NAND21X1 U405 ( .B(n383), .A(n348), .Y(n349) );
  NAND42X1 U406 ( .C(n140), .D(n168), .A(n171), .B(n226), .Y(n125) );
  OA21X1 U407 ( .B(prx_rst[0]), .C(prx_rst[1]), .A(set03[1]), .Y(set03[7]) );
  INVX1 U408 ( .A(n175), .Y(n386) );
  NAND2X1 U409 ( .A(n410), .B(n125), .Y(n146) );
  NAND2X1 U410 ( .A(n113), .B(n379), .Y(n112) );
  NAND2X1 U411 ( .A(n175), .B(n174), .Y(n205) );
  OAI22X1 U412 ( .A(n105), .B(n383), .C(n257), .D(n111), .Y(wd19[7]) );
  NAND4X1 U413 ( .A(n114), .B(n168), .C(n200), .D(n201), .Y(n124) );
  NOR4XL U414 ( .A(n249), .B(n215), .C(n242), .D(n226), .Y(n201) );
  NOR21XL U415 ( .B(n171), .A(n134), .Y(n200) );
  NAND43X1 U416 ( .B(set_hold), .C(cpurst), .D(n379), .A(n113), .Y(upd12) );
  MUX2X1 U417 ( .D0(n219), .D1(pff_rxpart[11]), .S(n109), .Y(wd21[3]) );
  MUX2X1 U418 ( .D0(pff_rxpart[5]), .D1(n231), .S(n270), .Y(wd20[5]) );
  INVX1 U419 ( .A(n233), .Y(n231) );
  MUX2X1 U420 ( .D0(pff_rxpart[3]), .D1(n220), .S(n270), .Y(wd20[3]) );
  MUX2X1 U421 ( .D0(pff_rxpart[4]), .D1(n225), .S(n270), .Y(wd20[4]) );
  MUX2X1 U422 ( .D0(pff_rxpart[0]), .D1(n133), .S(n270), .Y(wd20[0]) );
  MUX2X1 U423 ( .D0(pff_rxpart[2]), .D1(n183), .S(n270), .Y(wd20[2]) );
  MUX2X1 U424 ( .D0(pff_rxpart[7]), .D1(sfr_wdat[7]), .S(n270), .Y(wd20[7]) );
  AO22AXL U425 ( .A(inst_ofs_plus[11]), .B(n103), .C(n215), .D(n111), .Y(
        wd19[3]) );
  OAI32X1 U426 ( .A(n396), .B(r_fifopsh), .C(n388), .D(n256), .E(n117), .Y(
        wd01[7]) );
  ENOX1 U427 ( .A(n15), .B(n226), .C(pff_rxpart[12]), .D(n109), .Y(wd21[4]) );
  ENOX1 U428 ( .A(n15), .B(n214), .C(pff_rxpart[10]), .D(n109), .Y(wd21[2]) );
  ENOX1 U429 ( .A(n15), .B(n235), .C(pff_rxpart[13]), .D(n109), .Y(wd21[5]) );
  ENOX1 U430 ( .A(n15), .B(n143), .C(pff_rxpart[9]), .D(n109), .Y(wd21[1]) );
  ENOX1 U431 ( .A(n15), .B(n247), .C(pff_rxpart[14]), .D(n109), .Y(wd21[6]) );
  ENOX1 U432 ( .A(n236), .B(n111), .C(inst_ofs_plus[13]), .D(n104), .Y(wd19[5]) );
  ENOX1 U433 ( .A(n226), .B(n111), .C(inst_ofs_plus[12]), .D(n104), .Y(wd19[4]) );
  ENOX1 U435 ( .A(n144), .B(n111), .C(inst_ofs_plus[9]), .D(n104), .Y(wd19[1])
         );
  ENOX1 U436 ( .A(n136), .B(n111), .C(inst_ofs_plus[8]), .D(n104), .Y(wd19[0])
         );
  ENOX1 U437 ( .A(n184), .B(n111), .C(inst_ofs_plus[10]), .D(n104), .Y(wd19[2]) );
  OAI211X1 U438 ( .C(n396), .D(n127), .A(n14), .B(n118), .Y(upd01) );
  NAND2X1 U439 ( .A(n120), .B(n15), .Y(upd21) );
  NAND2X1 U440 ( .A(n175), .B(n205), .Y(N108) );
  NAND21X1 U441 ( .B(n270), .A(n120), .Y(upd20) );
  MUX2X1 U442 ( .D0(n216), .D1(inst_ofs_plus[3]), .S(n103), .Y(wd18[3]) );
  AND4X1 U443 ( .A(n348), .B(n383), .C(n330), .D(sfr_r), .Y(upd31) );
  ENOX1 U444 ( .A(n103), .B(n256), .C(inst_ofs_plus[7]), .D(n104), .Y(wd18[7])
         );
  ENOX1 U445 ( .A(n103), .B(n247), .C(inst_ofs_plus[6]), .D(n104), .Y(wd18[6])
         );
  ENOX1 U446 ( .A(n103), .B(n226), .C(inst_ofs_plus[4]), .D(ictlr_inc), .Y(
        wd18[4]) );
  ENOX1 U447 ( .A(n103), .B(n214), .C(inst_ofs_plus[2]), .D(ictlr_inc), .Y(
        wd18[2]) );
  ENOX1 U448 ( .A(n103), .B(n144), .C(inst_ofs_plus[1]), .D(ictlr_inc), .Y(
        wd18[1]) );
  ENOX1 U449 ( .A(n103), .B(n236), .C(inst_ofs_plus[5]), .D(n104), .Y(wd18[5])
         );
  AND2X1 U450 ( .A(prx_setsta[6]), .B(n11), .Y(set03[6]) );
  NAND2X1 U451 ( .A(prx_setsta[3]), .B(n11), .Y(n122) );
  XNOR2XL U452 ( .A(N27), .B(n412), .Y(N28) );
  XNOR2XL U453 ( .A(N28), .B(n411), .Y(N29) );
  AND2X1 U454 ( .A(i_goidle), .B(n11), .Y(set04[1]) );
  XNOR2XL U455 ( .A(n414), .B(add_180_carry[4]), .Y(N35) );
  XNOR2XL U456 ( .A(N30), .B(N32), .Y(N39) );
  NOR2X1 U457 ( .A(n11), .B(i_goidle), .Y(n173) );
  NAND2X1 U458 ( .A(n206), .B(n406), .Y(n174) );
  INVX1 U459 ( .A(n209), .Y(n407) );
  INVX1 U460 ( .A(n210), .Y(n408) );
  NAND2X1 U461 ( .A(n132), .B(n384), .Y(N84) );
  XNOR2XL U462 ( .A(di_p0[3]), .B(n403), .Y(n193) );
  XNOR2XL U463 ( .A(di_p0[5]), .B(n402), .Y(n195) );
  XNOR2XL U464 ( .A(di_p0[7]), .B(n397), .Y(n197) );
  XNOR2XL U465 ( .A(di_p0[4]), .B(n398), .Y(n196) );
  XNOR2XL U466 ( .A(di_p0[6]), .B(n401), .Y(n198) );
  XNOR2XL U467 ( .A(di_p0[2]), .B(n404), .Y(n194) );
  NAND2X1 U468 ( .A(n259), .B(aswkup), .Y(pwrdn_rstz) );
  AND2X1 U469 ( .A(dnchk_en), .B(dm_fault), .Y(dmf_wkup) );
  INVX1 U470 ( .A(n147), .Y(n382) );
  MUX2X1 U471 ( .D0(s_scp), .D1(m_scp), .S(reg94[5]), .Y(regAD[4]) );
  AND2X1 U472 ( .A(i_pc[6]), .B(n383), .Y(reg30[6]) );
  AND2X1 U473 ( .A(i_pc[7]), .B(n383), .Y(reg30[7]) );
  MUX2X1 U474 ( .D0(s_ovp), .D1(m_ovp), .S(reg94[4]), .Y(regAD[2]) );
  AND3X1 U475 ( .A(n18), .B(n215), .C(n377), .Y(ps_pwrdn) );
  INVX1 U476 ( .A(n145), .Y(n377) );
  AOI222XL U477 ( .A(reg28[7]), .B(reg27[7]), .C(reg28[4]), .D(reg27[4]), .E(
        reg28[6]), .F(reg27[6]), .Y(n178) );
  NAND3X1 U478 ( .A(n176), .B(n177), .C(n178), .Y(i2c_stretch) );
  AOI22X1 U479 ( .A(reg28[2]), .B(reg27[2]), .C(reg28[3]), .D(reg27[3]), .Y(
        n176) );
  AOI22X1 U480 ( .A(reg28[0]), .B(reg27[0]), .C(reg28[1]), .D(reg27[1]), .Y(
        n177) );
  NAND32X1 U481 ( .B(bkpt_hold), .C(reg12[3]), .A(n132), .Y(r_hold_mcu) );
  OAI211X1 U482 ( .C(ictlr_idle), .D(n338), .A(oscdwn_shft[1]), .B(bus_idle), 
        .Y(n145) );
  AND2X1 U483 ( .A(n132), .B(regD4_1_), .Y(n338) );
  AND2X1 U484 ( .A(regD4_0_), .B(oscdwn_shft[2]), .Y(r_osc_stop) );
  NOR21XL U485 ( .B(oscdwn_shft[2]), .A(n384), .Y(r_osc_lo) );
  NOR2X1 U486 ( .A(regD4_2_), .B(regD4_0_), .Y(n132) );
  INVX1 U487 ( .A(regD4_1_), .Y(n384) );
  AND2X1 U488 ( .A(regE3_0), .B(n129), .Y(r_srcctl[0]) );
  AND2X1 U489 ( .A(regE3[3]), .B(n128), .Y(r_srcctl[3]) );
  AND2X1 U490 ( .A(regE3[2]), .B(n128), .Y(r_srcctl[2]) );
  NOR2X1 U491 ( .A(r_srcctl[7]), .B(n129), .Y(frc_hg_off) );
  AOI22X1 U492 ( .A(regAF[4]), .B(regAE[4]), .C(regAF[2]), .D(regAE[2]), .Y(
        n129) );
  MUX2X1 U493 ( .D0(i_pc[5]), .D1(prx_adpn[5]), .S(reg19_7_), .Y(reg30[5]) );
  AOI22X1 U494 ( .A(regAF[5]), .B(regAE[5]), .C(regAD[5]), .D(i_vcbyval), .Y(
        n128) );
  INVX1 U495 ( .A(regD3_7_), .Y(r_gpio_ie[1]) );
  NOR21XL U496 ( .B(pff_ack[1]), .A(prl_cany0), .Y(set04[5]) );
  NOR4XL U497 ( .A(prl_fsm[3]), .B(prl_fsm[2]), .C(prl_fsm[1]), .D(prl_fsm[0]), 
        .Y(n204) );
  AND2X1 U498 ( .A(reg94[7]), .B(reg94[6]), .Y(r_otpi_gate) );
  NAND21X1 U499 ( .B(lg_dischg), .A(n352), .Y(r_srcctl[1]) );
  NOR21XL U500 ( .B(pff_ack[0]), .A(prl_cany0), .Y(set04[4]) );
  AND2X1 U501 ( .A(regD4_4_), .B(oscdwn_shft[2]), .Y(r_ocdrv_enz) );
  INVX1 U502 ( .A(reg19_7_), .Y(n383) );
  NAND4X1 U503 ( .A(n160), .B(n161), .C(n162), .D(n163), .Y(o_intr[1]) );
  AOI22X1 U504 ( .A(reg06[6]), .B(irq04[6]), .C(reg06[7]), .D(irq04[7]), .Y(
        n160) );
  AOI22X1 U505 ( .A(reg06[0]), .B(irq04[0]), .C(reg06[1]), .D(irq04[1]), .Y(
        n163) );
  AOI211X1 U506 ( .C(n412), .D(n411), .A(rstcnt[3]), .B(n414), .Y(n211) );
  AOI22X1 U507 ( .A(reg06[4]), .B(irq04[4]), .C(reg06[5]), .D(irq04[5]), .Y(
        n161) );
  INVX1 U508 ( .A(rstcnt[4]), .Y(n414) );
  INVX1 U509 ( .A(lg_pulse_12m), .Y(n352) );
  INVX1 U510 ( .A(rstcnt[2]), .Y(n412) );
  INVX1 U511 ( .A(rstcnt[1]), .Y(n411) );
  AND2X1 U512 ( .A(regD4_3_), .B(oscdwn_shft[2]), .Y(r_pwrdn) );
  INVX1 U513 ( .A(drstz[1]), .Y(n413) );
  INVX1 U514 ( .A(sfr_r), .Y(n391) );
  NOR21XL U515 ( .B(prx_setsta[1]), .A(n12), .Y(set03[1]) );
  AOI21X1 U516 ( .B(n138), .C(we_227), .A(lg_pulse_12m), .Y(n175) );
  OR4X1 U517 ( .A(osc_gate_n_1_), .B(osc_gate_n_0_), .C(test_so1), .D(
        osc_gate_n_2_), .Y(r_osc_gate) );
  OAI21X1 U518 ( .B(lg_pulse_len[1]), .C(lg_pulse_len[0]), .A(n386), .Y(n207)
         );
  NAND4X1 U519 ( .A(n164), .B(n165), .C(n166), .D(n167), .Y(o_intr[0]) );
  AOI22X1 U520 ( .A(reg05[4]), .B(irq03[4]), .C(reg05[5]), .D(irq03[5]), .Y(
        n165) );
  AOI22X1 U521 ( .A(reg05[2]), .B(irq03[2]), .C(reg05[3]), .D(irq03[3]), .Y(
        n166) );
  OAI33XL U522 ( .A(n205), .B(n206), .C(n406), .D(n394), .E(n393), .F(n207), 
        .Y(N113) );
  INVX1 U523 ( .A(lg_pulse_len[0]), .Y(n394) );
  OAI32X1 U524 ( .A(n405), .B(r_phyrst[1]), .C(n395), .D(r_phyrst[0]), .E(n170), .Y(n1222) );
  INVX1 U525 ( .A(n173), .Y(n395) );
  AOI21X1 U526 ( .B(reg11_7_), .C(set03[7]), .A(n146), .Y(n170) );
  AOI22X1 U527 ( .A(reg05[6]), .B(irq03[6]), .C(reg05[7]), .D(irq03[7]), .Y(
        n164) );
  AND2X1 U528 ( .A(regD4_2_), .B(oscdwn_shft[2]), .Y(r_pos_gate) );
  NOR21XL U529 ( .B(prx_setsta[2]), .A(prl_cany0), .Y(set03[2]) );
  GEN2XL U530 ( .D(lg_pulse_cnt[1]), .E(lg_pulse_cnt[0]), .C(n210), .B(n387), 
        .A(n386), .Y(N110) );
  ENOX1 U531 ( .A(n137), .B(n389), .C(n389), .D(lt_reg26_0), .Y(i2c_mode_wdat)
         );
  AOI21X1 U532 ( .B(n179), .C(n389), .A(n180), .Y(i2c_mode_upd) );
  XNOR2XL U533 ( .A(r_hwi2c_en), .B(lt_reg26_0), .Y(n179) );
  AOI22X1 U534 ( .A(reg05[0]), .B(irq03[0]), .C(reg05[1]), .D(irq03[1]), .Y(
        n167) );
  OAI22X1 U535 ( .A(n208), .B(n205), .C(n393), .D(n207), .Y(N112) );
  AOI21X1 U536 ( .B(lg_pulse_cnt[3]), .C(n407), .A(n206), .Y(n208) );
  OAI21BBX1 U537 ( .A(n174), .B(lg_dischg), .C(n175), .Y(n1220) );
  OAI21X1 U538 ( .B(lg_pulse_cnt[0]), .C(n205), .A(n175), .Y(N109) );
  OAI21BX1 U539 ( .C(reg12[3]), .B(n113), .A(n115), .Y(wd12[3]) );
  AOI32X1 U540 ( .A(set_hold), .B(n113), .C(n381), .D(n215), .E(n380), .Y(n115) );
  INVX1 U541 ( .A(n112), .Y(n380) );
  GEN2XL U542 ( .D(lg_pulse_cnt[2]), .E(n408), .C(n209), .B(n387), .A(n385), 
        .Y(N111) );
  INVX1 U543 ( .A(n207), .Y(n385) );
  NAND2X1 U544 ( .A(n19), .B(n113), .Y(wd12[4]) );
  MUX2IX1 U545 ( .D0(reg12[4]), .D1(n225), .S(n379), .Y(n19) );
  NOR21XL U546 ( .B(n118), .A(n119), .Y(wd01[6]) );
  AOI22X1 U547 ( .A(n388), .B(n241), .C(r_first), .D(n117), .Y(n119) );
  OAI21X1 U548 ( .B(r_fifopsh), .C(r_fifopop), .A(r_first), .Y(n118) );
  OAI22X1 U549 ( .A(n351), .B(n144), .C(lg_dischg), .D(n352), .Y(n1219) );
  OAI21X1 U550 ( .B(n199), .C(n180), .A(n124), .Y(N26) );
  NOR21XL U551 ( .B(n126), .A(rstcnt[4]), .Y(n199) );
  ENOX1 U552 ( .A(n15), .B(n137), .C(pff_rxpart[8]), .D(n109), .Y(wd21[0]) );
  ENOX1 U553 ( .A(n247), .B(n111), .C(inst_ofs_plus[14]), .D(n104), .Y(wd19[6]) );
  ENOX1 U554 ( .A(n214), .B(n112), .C(r_txshrt), .D(n112), .Y(wd12[2]) );
  ENOX1 U555 ( .A(n136), .B(n112), .C(r_pshords), .D(n112), .Y(wd12[0]) );
  ENOX1 U556 ( .A(n144), .B(n112), .C(reg12_1), .D(n112), .Y(wd12[1]) );
  ENOX1 U557 ( .A(n236), .B(n13), .C(reg12[5]), .D(n112), .Y(wd12[5]) );
  ENOX1 U558 ( .A(n247), .B(n13), .C(reg12[6]), .D(n112), .Y(wd12[6]) );
  ENOX1 U559 ( .A(n257), .B(n13), .C(reg12[7]), .D(n112), .Y(wd12[7]) );
  AO22AXL U560 ( .A(r_txnumk[0]), .B(n117), .C(sfr_wdat[0]), .D(n117), .Y(
        wd01[0]) );
  ENOX1 U561 ( .A(n236), .B(n14), .C(r_unlock), .D(n117), .Y(wd01[5]) );
  NOR21XL U562 ( .B(pff_obsd), .A(n12), .Y(set04[3]) );
  AOI22X1 U563 ( .A(reg06[2]), .B(irq04[2]), .C(reg06[3]), .D(irq04[3]), .Y(
        n162) );
  ENOX1 U564 ( .A(n103), .B(n137), .C(inst_ofs_plus[0]), .D(n104), .Y(wd18[0])
         );
  NOR21XL U565 ( .B(prx_setsta[4]), .A(prl_cany0), .Y(set03[4]) );
  AOI21BBXL U566 ( .B(r_auto_gdcrc[1]), .C(n122), .A(set03[6]), .Y(n120) );
  AO21X1 U567 ( .B(n130), .C(n131), .A(reg11_4), .Y(r_rxords_ena[4]) );
  NOR3XL U568 ( .A(r_rxords_ena[3]), .B(r_rxords_ena[6]), .C(r_rxords_ena[5]), 
        .Y(n131) );
  NOR3XL U569 ( .A(r_rxords_ena[0]), .B(r_rxords_ena[2]), .C(r_rxords_ena[1]), 
        .Y(n130) );
  INVX1 U570 ( .A(regD3_3), .Y(r_gpio_ie[0]) );
  OAI31XL U571 ( .A(n211), .B(r_phyrst[1]), .C(n413), .D(n259), .Y(prstz) );
  NOR21XL U572 ( .B(i_gobusy), .A(prl_cany0), .Y(set04[2]) );
  NOR21XL U573 ( .B(prx_setsta[5]), .A(prl_cany0), .Y(set03[5]) );
  AOI22X1 U574 ( .A(reg27[6]), .B(irq28[6]), .C(reg27[7]), .D(irq28[7]), .Y(
        n156) );
  NAND4X1 U575 ( .A(n156), .B(n157), .C(n158), .D(n159), .Y(o_intr[2]) );
  AOI22X1 U576 ( .A(reg27[4]), .B(irq28[4]), .C(reg27[5]), .D(irq28[5]), .Y(
        n157) );
  AOI22X1 U577 ( .A(reg27[0]), .B(irq28[0]), .C(reg27[1]), .D(irq28[1]), .Y(
        n159) );
  NOR21XL U578 ( .B(ptx_ack), .A(prl_cany0), .Y(set04[0]) );
  XNOR2XL U579 ( .A(n414), .B(rstcnt[3]), .Y(N27) );
  XOR2X1 U580 ( .A(N29), .B(rstcnt[0]), .Y(N30) );
  NOR21XL U581 ( .B(prl_GCTxDone), .A(n12), .Y(set04[6]) );
  AO22AXL U582 ( .A(reg94[4]), .B(m_ovp_sta), .C(s_ovp_sta), .D(reg94[4]), .Y(
        setAE[2]) );
  AO22AXL U583 ( .A(reg94[5]), .B(m_scp_sta), .C(s_scp_sta), .D(reg94[5]), .Y(
        setAE[4]) );
  NOR21XL U584 ( .B(prl_discard), .A(prl_cany0), .Y(set04[7]) );
  INVX1 U585 ( .A(reg25_0_), .Y(r_i2c_ninc) );
  NAND4X1 U586 ( .A(n148), .B(n149), .C(n150), .D(n151), .Y(o_intr[4]) );
  AOI22X1 U587 ( .A(regAF[6]), .B(irqAE[6]), .C(regAF[7]), .D(irqAE[7]), .Y(
        n148) );
  AOI22X1 U588 ( .A(regAF[0]), .B(irqAE[0]), .C(regAF[1]), .D(irqAE[1]), .Y(
        n151) );
  AOI22X1 U589 ( .A(irqAE[2]), .B(regAF[2]), .C(regAF[3]), .D(irqAE[3]), .Y(
        n150) );
  AOI22X1 U590 ( .A(irqAE[4]), .B(regAF[4]), .C(irqAE[5]), .D(regAF[5]), .Y(
        n149) );
  AOI22X1 U591 ( .A(reg27[2]), .B(irq28[2]), .C(reg27[3]), .D(irq28[3]), .Y(
        n158) );
  NOR21XL U592 ( .B(prx_setsta[0]), .A(prl_cany0), .Y(set03[0]) );
  XNOR2XL U593 ( .A(d_p0[0]), .B(n400), .Y(setDF[0]) );
  XNOR2XL U594 ( .A(d_p0[1]), .B(n399), .Y(setDF[1]) );
  XNOR2XL U595 ( .A(d_p0[2]), .B(n404), .Y(setDF[2]) );
  XNOR2XL U596 ( .A(d_p0[3]), .B(n403), .Y(setDF[3]) );
  XNOR2XL U597 ( .A(d_p0[4]), .B(n398), .Y(setDF[4]) );
  NAND2X1 U598 ( .A(rstcnt[4]), .B(n126), .Y(n113) );
  NOR42XL U599 ( .C(n202), .D(r_inst_ofs[10]), .A(r_inst_ofs[8]), .B(n203), 
        .Y(n171) );
  NAND4X1 U600 ( .A(r_inst_ofs[14]), .B(r_inst_ofs[13]), .C(r_inst_ofs[12]), 
        .D(r_inst_ofs[11]), .Y(n203) );
  NOR2X1 U601 ( .A(reg19_7_), .B(r_inst_ofs[9]), .Y(n202) );
  AOI22X1 U602 ( .A(regDE[0]), .B(irqDF[0]), .C(regDE[1]), .D(irqDF[1]), .Y(
        n155) );
  NOR4XL U603 ( .A(rstcnt[0]), .B(rstcnt[1]), .C(rstcnt[2]), .D(rstcnt[3]), 
        .Y(n126) );
  AOI22X1 U604 ( .A(regDE[2]), .B(irqDF[2]), .C(regDE[3]), .D(irqDF[3]), .Y(
        n154) );
  OAI32X1 U605 ( .A(n405), .B(r_phyrst[1]), .C(n173), .D(r_phyrst[0]), .E(n410), .Y(n1221) );
  XNOR2XL U606 ( .A(d_p0[6]), .B(n401), .Y(setDF[6]) );
  XNOR2XL U607 ( .A(d_p0[7]), .B(n397), .Y(setDF[7]) );
  XNOR2XL U608 ( .A(d_p0[5]), .B(n402), .Y(setDF[5]) );
  INVX1 U609 ( .A(ff_p0[6]), .Y(n401) );
  INVX1 U610 ( .A(ff_p0[7]), .Y(n397) );
  INVX1 U611 ( .A(ff_p0[1]), .Y(n399) );
  INVX1 U612 ( .A(ff_p0[0]), .Y(n400) );
  INVX1 U613 ( .A(ff_p0[3]), .Y(n403) );
  INVX1 U614 ( .A(ff_p0[2]), .Y(n404) );
  INVX1 U615 ( .A(ff_p0[5]), .Y(n402) );
  INVX1 U616 ( .A(ff_p0[4]), .Y(n398) );
  NAND4X1 U617 ( .A(n152), .B(n153), .C(n154), .D(n155), .Y(o_intr[3]) );
  AOI22X1 U618 ( .A(regDE[6]), .B(irqDF[6]), .C(regDE[7]), .D(irqDF[7]), .Y(
        n152) );
  AOI22X1 U619 ( .A(regDE[4]), .B(irqDF[4]), .C(regDE[5]), .D(irqDF[5]), .Y(
        n153) );
  NOR2X1 U620 ( .A(n408), .B(lg_pulse_cnt[2]), .Y(n209) );
  NOR2X1 U621 ( .A(lg_pulse_cnt[1]), .B(lg_pulse_cnt[0]), .Y(n210) );
  NOR2X1 U622 ( .A(n407), .B(lg_pulse_cnt[3]), .Y(n206) );
  INVX1 U623 ( .A(r_phyrst[1]), .Y(n410) );
  INVX1 U624 ( .A(lg_pulse_cnt[4]), .Y(n406) );
  INVX1 U625 ( .A(r_last), .Y(n396) );
  INVX1 U626 ( .A(r_phyrst[0]), .Y(n405) );
  INVX1 U627 ( .A(lg_pulse_len[1]), .Y(n393) );
  NAND42X1 U628 ( .C(di_rd_det_clr), .D(dm_fault_clr), .A(n86), .B(n186), .Y(
        aswkup) );
  NOR2X1 U629 ( .A(p0_chg_clr), .B(i_tmrf), .Y(n186) );
  OAI21X1 U630 ( .B(osc_low_clr), .C(n147), .A(n259), .Y(osc_low_rstz) );
  NAND2X1 U631 ( .A(n3), .B(srstz), .Y(n147) );
  AOI22X1 U632 ( .A(regDE[1]), .B(n191), .C(regDE[0]), .D(n192), .Y(n190) );
  XNOR2XL U633 ( .A(di_p0[0]), .B(n400), .Y(n192) );
  XNOR2XL U634 ( .A(di_p0[1]), .B(n399), .Y(n191) );
  NAND4X1 U635 ( .A(n187), .B(n188), .C(n189), .D(n190), .Y(as_p0_chg) );
  AOI22X1 U636 ( .A(regDE[7]), .B(n197), .C(regDE[6]), .D(n198), .Y(n187) );
  AOI22X1 U637 ( .A(regDE[5]), .B(n195), .C(regDE[4]), .D(n196), .Y(n188) );
  AOI22X1 U638 ( .A(regDE[3]), .B(n193), .C(regDE[2]), .D(n194), .Y(n189) );
  INVX1 U639 ( .A(sfr_addr[7]), .Y(n262) );
  INVXL U640 ( .A(n334), .Y(n374) );
  INVXL U641 ( .A(sfr_w), .Y(n300) );
  NAND21XL U642 ( .B(n334), .A(n327), .Y(n269) );
  NAND21XL U643 ( .B(n334), .A(n348), .Y(n324) );
  NAND21XL U644 ( .B(n334), .A(n333), .Y(n335) );
  NAND21XL U645 ( .B(n276), .A(n345), .Y(n277) );
  NAND21XL U646 ( .B(n276), .A(n302), .Y(n274) );
  NAND21XL U647 ( .B(n276), .A(n307), .Y(n290) );
  NAND32XL U648 ( .B(n292), .C(n354), .A(n110), .Y(n342) );
  NAND21XL U649 ( .B(n372), .A(sfr_addr[5]), .Y(n287) );
  NAND21XL U650 ( .B(n294), .A(sfr_addr[5]), .Y(n354) );
  NAND21XL U651 ( .B(sfr_addr[5]), .A(n372), .Y(n299) );
  NAND21XL U652 ( .B(n107), .A(n292), .Y(n364) );
  NAND21XL U653 ( .B(n371), .A(n107), .Y(n275) );
  NAND21XL U654 ( .B(n292), .A(n107), .Y(n304) );
endmodule


module regbank_a0_DW_rightsh_1 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n114, n115, n116, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n183, n184, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n305, n309, n310, n312, n313, n314, n315, n316, n317,
         n319, n320, n328, n478, n497, n498, n503, n509, n510, n515, n516,
         n522, n527, n528, n533, n534, n539, n540, n545, n546, n557, n558,
         n563, n564, n569, n570, n575, n585, n586, n589, n590, n593, n594,
         n597, n598, n609, n610, n613, n614, n617, n618, n625, n626, n629,
         n630, n633, n634, n637, n638, n645, n646, n653, n654, n669, n670,
         n673, n674, n677, n678, n681, n684, n687, n690, n693, n696, n699,
         n702, n705, n706, n709, n710, n713, n714, n717, n718, n721, n722,
         n725, n726, n729, n730, n733, n734, n737, n740, n743, n746, n749,
         n752, n755, n758, n761, n762, n765, n766, n769, n770, n773, n774,
         n781, n782, n789, n790, n795, n796, n801, n802, n807, n808, n813,
         n814, n819, n820, n831, n837, n838, n843, n855, n856, n861, n862,
         n867, n868, n874, n879, n880, n885, n886, n891, n892, n897, n898,
         n903, n909, n910, n915, n916, n921, n922, n937, n938, n941, n942,
         n945, n946, n949, n950, n953, n954, n957, n958, n961, n962, n965,
         n966, n969, n970, n973, n974, n977, n978, n981, n982, n985, n986,
         n989, n990, n993, n994, n997, n998, n1015, n1021, n1022, n1027, n1028,
         n1034, n1039, n1040, n1045, n1046, n1049, n1050, n1053, n1054, n1057,
         n1058, n1061, n1062, n1065, n1066, n1069, n1070, n1073, n1074, n1077,
         n1078, n1081, n1082, n1085, n1086, n1089, n1090, n1093, n1094, n1097,
         n1098, n1101, n1102, n1105, n1106, n1109, n1110, n1113, n1114, n1117,
         n1118, n1121, n1122, n1125, n1126, n1129, n1130, n1134, n1137, n1138,
         n1141, n1142, n1145, n1146, n1149, n1153, n1154, n1157, n1158, n1161,
         n1162, n1165, n1166, n1169, n1170, n1173, n1174, n1177, n1178, n1181,
         n1182, n1185, n1186, n1189, n1190, n1193, n1194, n1197, n1198, n1201,
         n1205, n1206, n1209, n1213, n1217, n1218, n1221, n1222, n1225, n1226,
         n1229, n1230, n1233, n1234, n1237, n1238, n1241, n1244, n1247, n1250,
         n1253, n1256, n1259, n1262, n1269, n1272, n1275, n1278, n1281, n1284,
         n1287, n1290, n1293, n1296, n1299, n1302, n1305, n1308, n1311, n1312,
         n1315, n1316, n1319, n1320, n1323, n1324, n1327, n1328, n1331, n1332,
         n1335, n1336, n1339, n1340, n1343, n1344, n1347, n1348, n1351, n1352,
         n1355, n1356, n1359, n1360, n1363, n1364, n1367, n1368, n1371, n1372,
         n1377, n1378, n1389, n1390, n1395, n1396, n1401, n1402, n1407, n1408,
         n1413, n1414, n1419, n1425, n1426, n1431, n1432, n1437, n1438, n1443,
         n1444, n1450, n1456, n1467, n1468, n1471, n1472, n1475, n1476, n1479,
         n1480, n1483, n1484, n1487, n1488, n1491, n1492, n1495, n1496, n1499,
         n1500, n1503, n1504, n1507, n1511, n1512, n1515, n1516, n1519, n1520,
         n1523, n1524, n1527, n1528, n1531, n1532, n1535, n1536, n1539, n1540,
         n1543, n1544, n1547, n1548, n1551, n1552, n1555, n1556, n1559, n1560,
         n1563, n1564, n1583, n1584, n1592, n1597, n1598, n1599, n1600, n1602,
         n1603, n1605, n1607, n1613, n1615, n1616, n1618, n1624, n1628, n1629,
         n1630, n1631, n1632, n1634, n1637, n1639, n1642, n1643, n1646, n1647,
         n1648, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1669, n1670, n1671, n1672, n1679, n1685,
         n1686, n1687, n1688, n1693, n1694, n1695, n1696, n1709, n1711, n1712,
         n1720, n1725, n1726, n1727, n1728, n1730, n1731, n1733, n1735, n1741,
         n1743, n1744, n1746, n1751, n1752, n1756, n1757, n1758, n1759, n1760,
         n1762, n1766, n1767, n1770, n1771, n1774, n1776, n1778, n1797, n1807,
         n1814, n1815, n1816, n1820, n1821, n1822, n1823, n1824, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037;

  MUX2IX4 U13 ( .D0(n28), .D1(n44), .S(n3895), .Y(n12) );
  MUX2IX4 U21 ( .D0(n20), .D1(n36), .S(n3896), .Y(n4) );
  MUX2IX4 U39 ( .D0(n66), .D1(n98), .S(SH[5]), .Y(n34) );
  MUX2IX4 U70 ( .D0(n163), .D1(n227), .S(n3903), .Y(n99) );
  MUX2IX4 U71 ( .D0(n162), .D1(n226), .S(n3903), .Y(n98) );
  MUX2IX4 U102 ( .D0(n131), .D1(n195), .S(n3906), .Y(n67) );
  MUX2IX4 U110 ( .D0(n123), .D1(n187), .S(n3907), .Y(n59) );
  MUX2IX4 U166 ( .D0(n315), .D1(n3734), .S(n3913), .Y(n195) );
  MUX2IX4 U174 ( .D0(n3880), .D1(n3882), .S(n3914), .Y(n187) );
  MUX2IX4 U238 ( .D0(n3891), .D1(n3889), .S(n3920), .Y(n123) );
  AO22X1 U514 ( .A(n4015), .B(A[510]), .C(n3971), .D(A[1022]), .Y(n498) );
  AO22X1 U525 ( .A(n4022), .B(A[253]), .C(n3700), .D(A[765]), .Y(n503) );
  AO22X1 U534 ( .A(n4015), .B(A[508]), .C(n3997), .D(A[1020]), .Y(n510) );
  AO22X1 U535 ( .A(n4016), .B(A[252]), .C(n3999), .D(A[764]), .Y(n509) );
  AO22X1 U544 ( .A(n4022), .B(A[507]), .C(n3701), .D(A[1019]), .Y(n516) );
  AO22X1 U554 ( .A(n4016), .B(A[506]), .C(n3997), .D(A[1018]), .Y(n522) );
  AO22X1 U560 ( .A(n528), .B(n3945), .C(n527), .D(n3954), .Y(n1824) );
  AO22X1 U570 ( .A(n534), .B(n3945), .C(n533), .D(n3961), .Y(n1823) );
  AO22X1 U575 ( .A(n4016), .B(A[248]), .C(n3999), .D(A[760]), .Y(n533) );
  AO22X1 U580 ( .A(n540), .B(n3944), .C(n539), .D(n3954), .Y(n1822) );
  AO22X1 U584 ( .A(n4022), .B(A[503]), .C(n3997), .D(A[1015]), .Y(n540) );
  AO22X1 U590 ( .A(n546), .B(n3944), .C(n545), .D(n3961), .Y(n1821) );
  AO22X1 U594 ( .A(n4023), .B(A[502]), .C(n3984), .D(A[1014]), .Y(n546) );
  AO22X1 U614 ( .A(n4018), .B(A[500]), .C(n3700), .D(A[1012]), .Y(n558) );
  AO22X1 U615 ( .A(n3853), .B(A[244]), .C(n3999), .D(A[756]), .Y(n557) );
  AO22X1 U624 ( .A(n4019), .B(A[499]), .C(n3997), .D(A[1011]), .Y(n564) );
  AO22X1 U635 ( .A(n4013), .B(A[242]), .C(n4029), .D(A[754]), .Y(n569) );
  AO22X1 U645 ( .A(n4023), .B(A[241]), .C(n3999), .D(A[753]), .Y(n575) );
  NOR2X1 U664 ( .A(n3992), .B(A[239]), .Y(n585) );
  NOR2X1 U672 ( .A(n3992), .B(A[238]), .Y(n589) );
  NOR2X1 U680 ( .A(n3991), .B(A[237]), .Y(n593) );
  NOR2X1 U688 ( .A(n3991), .B(A[236]), .Y(n597) );
  NOR2X1 U712 ( .A(n3991), .B(A[233]), .Y(n609) );
  NOR2X1 U720 ( .A(n3990), .B(A[232]), .Y(n613) );
  NOR2X1 U728 ( .A(n3991), .B(A[231]), .Y(n617) );
  NOR2X1 U744 ( .A(n3989), .B(A[229]), .Y(n625) );
  NOR2X1 U752 ( .A(n3989), .B(A[228]), .Y(n629) );
  NOR2X1 U760 ( .A(n3991), .B(A[227]), .Y(n633) );
  NOR2X1 U784 ( .A(n3989), .B(A[224]), .Y(n645) );
  NOR2X1 U800 ( .A(n3989), .B(A[222]), .Y(n653) );
  NOR2X1 U840 ( .A(n3989), .B(A[217]), .Y(n673) );
  NOR2X1 U848 ( .A(n3989), .B(A[216]), .Y(n677) );
  NOR2X1 U1031 ( .A(n3990), .B(A[447]), .Y(n762) );
  NOR2X1 U1039 ( .A(n3990), .B(A[446]), .Y(n766) );
  NOR2X1 U1047 ( .A(n3990), .B(A[445]), .Y(n770) );
  NOR2X1 U1055 ( .A(n3990), .B(A[444]), .Y(n774) );
  NOR2X1 U1071 ( .A(n3990), .B(A[442]), .Y(n782) );
  NOR2X1 U1087 ( .A(n3991), .B(A[440]), .Y(n790) );
  AO22X1 U1092 ( .A(n796), .B(n3943), .C(n795), .D(n3953), .Y(n1758) );
  AO22X1 U1096 ( .A(n4023), .B(A[439]), .C(n3996), .D(A[951]), .Y(n796) );
  AO22X1 U1097 ( .A(n4016), .B(A[183]), .C(n4005), .D(A[695]), .Y(n795) );
  AO22X1 U1102 ( .A(n802), .B(n3942), .C(n801), .D(n3962), .Y(n1757) );
  AO22X1 U1106 ( .A(n4017), .B(A[438]), .C(n3987), .D(A[950]), .Y(n802) );
  AO22X1 U1107 ( .A(n4017), .B(A[182]), .C(n4033), .D(A[694]), .Y(n801) );
  AO22X1 U1116 ( .A(n4016), .B(A[437]), .C(n3979), .D(A[949]), .Y(n808) );
  AO22X1 U1117 ( .A(n4016), .B(A[181]), .C(n4002), .D(A[693]), .Y(n807) );
  AO22X1 U1126 ( .A(n4017), .B(A[436]), .C(n3984), .D(A[948]), .Y(n814) );
  AO22X1 U1127 ( .A(n4017), .B(A[180]), .C(n3974), .D(A[692]), .Y(n813) );
  AO22X1 U1136 ( .A(n4023), .B(A[435]), .C(n3999), .D(A[947]), .Y(n820) );
  AO22X1 U1137 ( .A(n4024), .B(A[179]), .C(n4001), .D(A[691]), .Y(n819) );
  AO22X1 U1157 ( .A(n4024), .B(A[177]), .C(n4001), .D(A[689]), .Y(n831) );
  AO22X1 U1162 ( .A(n838), .B(n3942), .C(n837), .D(n3711), .Y(n1751) );
  AO22X1 U1166 ( .A(n4018), .B(A[432]), .C(n4001), .D(A[944]), .Y(n838) );
  AO22X1 U1167 ( .A(n4018), .B(A[176]), .C(n4001), .D(A[688]), .Y(n837) );
  AO22X1 U1177 ( .A(n4024), .B(A[175]), .C(n4001), .D(A[687]), .Y(n843) );
  AO22X1 U1196 ( .A(n4024), .B(A[429]), .C(n4000), .D(A[941]), .Y(n856) );
  AO22X1 U1197 ( .A(n4025), .B(A[173]), .C(n4000), .D(A[685]), .Y(n855) );
  AO22X1 U1206 ( .A(n4019), .B(A[428]), .C(n4000), .D(A[940]), .Y(n862) );
  AO22X1 U1207 ( .A(n4016), .B(A[172]), .C(n4000), .D(A[684]), .Y(n861) );
  AO22X1 U1212 ( .A(n868), .B(n3942), .C(n867), .D(n3951), .Y(n1746) );
  AO22X1 U1216 ( .A(n4025), .B(A[427]), .C(n4000), .D(A[939]), .Y(n868) );
  AO22X1 U1217 ( .A(n4025), .B(A[171]), .C(n4000), .D(A[683]), .Y(n867) );
  AO22X1 U1226 ( .A(n4019), .B(A[426]), .C(n4000), .D(A[938]), .Y(n874) );
  AO22X1 U1232 ( .A(n880), .B(n3941), .C(n879), .D(n3951), .Y(n1744) );
  AO22X1 U1236 ( .A(n4025), .B(A[425]), .C(n3701), .D(A[937]), .Y(n880) );
  AO22X1 U1237 ( .A(n4025), .B(A[169]), .C(n4002), .D(A[681]), .Y(n879) );
  AO22X1 U1242 ( .A(n886), .B(n3942), .C(n885), .D(n3963), .Y(n1743) );
  AO22X1 U1246 ( .A(n4022), .B(A[424]), .C(n3700), .D(A[936]), .Y(n886) );
  AO22X1 U1247 ( .A(n4019), .B(A[168]), .C(n3999), .D(A[680]), .Y(n885) );
  AO22X1 U1256 ( .A(n4025), .B(A[423]), .C(n3999), .D(A[935]), .Y(n892) );
  AO22X1 U1257 ( .A(n4026), .B(A[167]), .C(n4002), .D(A[679]), .Y(n891) );
  AO22X1 U1262 ( .A(n898), .B(n3942), .C(n897), .D(n3963), .Y(n1741) );
  AO22X1 U1266 ( .A(n4019), .B(A[422]), .C(n3973), .D(A[934]), .Y(n898) );
  AO22X1 U1267 ( .A(n4019), .B(A[166]), .C(n3701), .D(A[678]), .Y(n897) );
  AO22X1 U1277 ( .A(n4026), .B(A[165]), .C(n3701), .D(A[677]), .Y(n903) );
  AO22X1 U1286 ( .A(n4019), .B(A[420]), .C(n3997), .D(A[932]), .Y(n910) );
  AO22X1 U1287 ( .A(n4019), .B(A[164]), .C(n3701), .D(A[676]), .Y(n909) );
  AO22X1 U1296 ( .A(n4026), .B(A[419]), .C(n3998), .D(A[931]), .Y(n916) );
  AO22X1 U1297 ( .A(n4026), .B(A[163]), .C(n4002), .D(A[675]), .Y(n915) );
  AO22X1 U1306 ( .A(n4019), .B(A[418]), .C(n3998), .D(A[930]), .Y(n922) );
  AO22X1 U1307 ( .A(n4015), .B(A[162]), .C(n3700), .D(A[674]), .Y(n921) );
  AO22X1 U1494 ( .A(n4017), .B(A[396]), .C(n3987), .D(A[908]), .Y(n1022) );
  AO22X1 U1504 ( .A(n4013), .B(A[395]), .C(n3979), .D(A[907]), .Y(n1028) );
  AO22X1 U1505 ( .A(n4013), .B(A[139]), .C(n3981), .D(A[651]), .Y(n1027) );
  AO22X1 U1514 ( .A(n4020), .B(A[394]), .C(n3988), .D(A[906]), .Y(n1034) );
  AO22X1 U1520 ( .A(n1040), .B(n3940), .C(n1039), .D(n3957), .Y(n1712) );
  AO22X1 U1524 ( .A(n4013), .B(A[393]), .C(n3988), .D(A[905]), .Y(n1040) );
  AO22X1 U1525 ( .A(n4013), .B(A[137]), .C(n4032), .D(A[649]), .Y(n1039) );
  AO22X1 U1530 ( .A(n1046), .B(n3942), .C(n1045), .D(n3959), .Y(n1711) );
  AO22X1 U1534 ( .A(n4020), .B(A[392]), .C(n4027), .D(A[904]), .Y(n1046) );
  AO22X1 U1535 ( .A(n4020), .B(A[136]), .C(n4005), .D(A[648]), .Y(n1045) );
  NOR2X1 U1544 ( .A(n3996), .B(A[135]), .Y(n1049) );
  NOR2X1 U1551 ( .A(n3996), .B(A[390]), .Y(n1054) );
  NOR2X1 U1552 ( .A(n3995), .B(A[134]), .Y(n1053) );
  NOR2X1 U1559 ( .A(n3995), .B(A[389]), .Y(n1058) );
  NOR2X1 U1560 ( .A(n3995), .B(A[133]), .Y(n1057) );
  NOR2X1 U1567 ( .A(n3995), .B(A[388]), .Y(n1062) );
  NOR2X1 U1575 ( .A(n3995), .B(A[387]), .Y(n1066) );
  NOR2X1 U1583 ( .A(n3995), .B(A[386]), .Y(n1070) );
  NOR2X1 U1584 ( .A(n3995), .B(A[130]), .Y(n1069) );
  NOR2X1 U1591 ( .A(n3996), .B(A[385]), .Y(n1074) );
  NOR2X1 U1599 ( .A(n3994), .B(A[384]), .Y(n1078) );
  NOR2X1 U1623 ( .A(n3994), .B(A[381]), .Y(n1090) );
  NOR2X1 U1631 ( .A(n3994), .B(A[380]), .Y(n1094) );
  NOR2X1 U1639 ( .A(n3994), .B(A[379]), .Y(n1098) );
  NOR2X1 U1647 ( .A(n3865), .B(A[378]), .Y(n1102) );
  NOR2X1 U1655 ( .A(n3992), .B(A[377]), .Y(n1106) );
  NOR2X1 U1663 ( .A(n4027), .B(A[376]), .Y(n1110) );
  NOR2X1 U1671 ( .A(n3979), .B(A[375]), .Y(n1114) );
  NOR2X1 U1679 ( .A(n4027), .B(A[374]), .Y(n1118) );
  NOR2X1 U1687 ( .A(n3866), .B(A[373]), .Y(n1122) );
  NOR2X1 U1695 ( .A(n4005), .B(A[372]), .Y(n1126) );
  NOR2X1 U1703 ( .A(n3993), .B(A[371]), .Y(n1130) );
  NOR2X1 U1719 ( .A(n3993), .B(A[369]), .Y(n1138) );
  NOR2X1 U1727 ( .A(n3993), .B(A[368]), .Y(n1142) );
  NOR2X1 U1735 ( .A(n3993), .B(A[367]), .Y(n1146) );
  NOR2X1 U1751 ( .A(n3993), .B(A[365]), .Y(n1154) );
  NOR2X1 U1759 ( .A(n3993), .B(A[364]), .Y(n1158) );
  NOR2X1 U1767 ( .A(n3992), .B(A[363]), .Y(n1162) );
  NOR2X1 U1783 ( .A(n3992), .B(A[361]), .Y(n1170) );
  NOR2X1 U1791 ( .A(n3992), .B(A[360]), .Y(n1174) );
  NOR2X1 U1799 ( .A(n3992), .B(A[359]), .Y(n1178) );
  NOR2X1 U1807 ( .A(n3995), .B(A[358]), .Y(n1182) );
  NOR2X1 U1815 ( .A(n3992), .B(A[357]), .Y(n1186) );
  NOR2X1 U1823 ( .A(n3992), .B(A[356]), .Y(n1190) );
  NOR2X1 U1831 ( .A(n3993), .B(A[355]), .Y(n1194) );
  NOR2X1 U1855 ( .A(n3987), .B(A[352]), .Y(n1206) );
  NOR2X1 U1887 ( .A(n3994), .B(A[348]), .Y(n1222) );
  NOR2X1 U1895 ( .A(n3994), .B(A[347]), .Y(n1226) );
  NOR2X1 U1903 ( .A(n3996), .B(A[346]), .Y(n1230) );
  NOR2X1 U1911 ( .A(n3996), .B(A[345]), .Y(n1234) );
  NOR2X1 U1919 ( .A(n3996), .B(A[344]), .Y(n1238) );
  NAND21X1 U1924 ( .B(n3937), .A(n1241), .Y(n1662) );
  NAND21X1 U1931 ( .B(n3925), .A(n1244), .Y(n1661) );
  NAND21X1 U1938 ( .B(n3966), .A(n1247), .Y(n1660) );
  NAND21X1 U1945 ( .B(n3966), .A(n1250), .Y(n1659) );
  NAND21X1 U1952 ( .B(n3945), .A(n1253), .Y(n1658) );
  NAND21X1 U1966 ( .B(n3966), .A(n1259), .Y(n1656) );
  NAND21X1 U1973 ( .B(n3945), .A(n1262), .Y(n1655) );
  NAND21X1 U1980 ( .B(n3942), .A(n3977), .Y(n1654) );
  NAND21X1 U1986 ( .B(n3931), .A(n3977), .Y(n1653) );
  NAND21X1 U1992 ( .B(n3967), .A(n1269), .Y(n1652) );
  NAND21X1 U1999 ( .B(n3940), .A(n1272), .Y(n1651) );
  NAND21X1 U2006 ( .B(n3940), .A(n1275), .Y(n1650) );
  NAND21X1 U2020 ( .B(n3940), .A(n1281), .Y(n1648) );
  NAND21X1 U2027 ( .B(n3940), .A(n1284), .Y(n1647) );
  AO22X1 U2222 ( .A(n4020), .B(A[303]), .C(n4005), .D(A[815]), .Y(n1378) );
  AO22X1 U2223 ( .A(n3853), .B(A[47]), .C(n4028), .D(A[559]), .Y(n1377) );
  AO22X1 U2242 ( .A(n4025), .B(A[301]), .C(n4005), .D(A[813]), .Y(n1390) );
  AO22X1 U2252 ( .A(n3853), .B(A[300]), .C(n4004), .D(A[812]), .Y(n1396) );
  AO22X1 U2253 ( .A(n4017), .B(A[44]), .C(n4004), .D(A[556]), .Y(n1395) );
  AO22X1 U2258 ( .A(n1402), .B(n3943), .C(n1401), .D(n3956), .Y(n1618) );
  AO22X1 U2262 ( .A(n4026), .B(A[299]), .C(n4004), .D(A[811]), .Y(n1402) );
  AO22X1 U2263 ( .A(n4025), .B(A[43]), .C(n4004), .D(A[555]), .Y(n1401) );
  AO22X1 U2272 ( .A(n4013), .B(A[298]), .C(n4004), .D(A[810]), .Y(n1408) );
  AO22X1 U2273 ( .A(n4023), .B(A[42]), .C(n4004), .D(A[554]), .Y(n1407) );
  AO22X1 U2278 ( .A(n1414), .B(n3965), .C(n1413), .D(n3956), .Y(n1616) );
  AO22X1 U2282 ( .A(n4025), .B(A[297]), .C(n4004), .D(A[809]), .Y(n1414) );
  AO22X1 U2283 ( .A(n4021), .B(A[41]), .C(n4004), .D(A[553]), .Y(n1413) );
  AO22X1 U2293 ( .A(n4014), .B(A[40]), .C(n4003), .D(A[552]), .Y(n1419) );
  AO22X1 U2302 ( .A(n4021), .B(A[295]), .C(n4003), .D(A[807]), .Y(n1426) );
  AO22X1 U2303 ( .A(n4021), .B(A[39]), .C(n4003), .D(A[551]), .Y(n1425) );
  AO22X1 U2308 ( .A(n1432), .B(n3966), .C(n1431), .D(n3960), .Y(n1613) );
  AO22X1 U2312 ( .A(n4014), .B(A[294]), .C(n4003), .D(A[806]), .Y(n1432) );
  AO22X1 U2313 ( .A(n4014), .B(A[38]), .C(n4003), .D(A[550]), .Y(n1431) );
  AO22X1 U2322 ( .A(n4021), .B(A[293]), .C(n4003), .D(A[805]), .Y(n1438) );
  AO22X1 U2323 ( .A(n4021), .B(A[37]), .C(n4003), .D(A[549]), .Y(n1437) );
  AO22X1 U2332 ( .A(n4014), .B(A[292]), .C(n4003), .D(A[804]), .Y(n1444) );
  AO22X1 U2333 ( .A(n4014), .B(A[36]), .C(n4003), .D(A[548]), .Y(n1443) );
  AO22X1 U2352 ( .A(n4014), .B(A[290]), .C(n4002), .D(A[802]), .Y(n1456) );
  AO22X1 U2368 ( .A(n1468), .B(n3944), .C(n1467), .D(n3960), .Y(n1607) );
  AO22X1 U2372 ( .A(n4015), .B(A[288]), .C(n3999), .D(A[800]), .Y(n1468) );
  AO22X1 U2373 ( .A(n4015), .B(A[32]), .C(n4001), .D(A[544]), .Y(n1467) );
  NOR21X1 U2470 ( .B(n3986), .A(A[532]), .Y(n1515) );
  NOR21XL U2611 ( .B(n3980), .A(A[717]), .Y(n713) );
  NOR21XL U2612 ( .B(n3980), .A(A[973]), .Y(n714) );
  NOR21XL U2613 ( .B(n3981), .A(A[621]), .Y(n1153) );
  NOR21XL U2614 ( .B(n3980), .A(A[661]), .Y(n977) );
  NOR21XL U2615 ( .B(n3987), .A(A[610]), .Y(n1197) );
  NOR21XL U2616 ( .B(n3982), .A(A[834]), .Y(n1302) );
  NOR21XL U2617 ( .B(n3987), .A(A[660]), .Y(n981) );
  NOR21XL U2618 ( .B(n3865), .A(A[628]), .Y(n1125) );
  MUX2IX1 U2619 ( .D0(n1483), .D1(n1484), .S(n3933), .Y(n1603) );
  MUX2IX1 U2620 ( .D0(n3722), .D1(n3670), .S(n3915), .Y(n173) );
  MUX2IX1 U2621 ( .D0(n309), .D1(n3794), .S(n3914), .Y(n189) );
  MUX2IX1 U2622 ( .D0(n3709), .D1(n3682), .S(n3911), .Y(n213) );
  MUX2IX1 U2623 ( .D0(n3673), .D1(n3714), .S(n3918), .Y(n142) );
  MUX2XL U2624 ( .D0(n945), .D1(n946), .S(n3929), .Y(n3714) );
  MUX2IX1 U2625 ( .D0(n3801), .D1(n3835), .S(n3912), .Y(n206) );
  MUX2X1 U2626 ( .D0(n1217), .D1(n1218), .S(n3929), .Y(n3801) );
  MUX2IX1 U2627 ( .D0(n3715), .D1(n3671), .S(n3915), .Y(n174) );
  MUX2XL U2628 ( .D0(n1319), .D1(n1320), .S(n3930), .Y(n3715) );
  NOR21XL U2629 ( .B(n3865), .A(A[606]), .Y(n1213) );
  MUX2IX1 U2630 ( .D0(n3731), .D1(n3679), .S(n3911), .Y(n212) );
  MUX2IX1 U2631 ( .D0(n3733), .D1(n3663), .S(n3920), .Y(n124) );
  MUX2XL U2632 ( .D0(n1551), .D1(n1552), .S(n3938), .Y(n3733) );
  MUX2X1 U2633 ( .D0(n1648), .D1(n1776), .S(n3914), .Y(n186) );
  MUX2X1 U2634 ( .D0(n1584), .D1(n1712), .S(n3920), .Y(n122) );
  MUX2IXL U2635 ( .D0(n115), .D1(n179), .S(n3907), .Y(n51) );
  MUX2IX1 U2636 ( .D0(n147), .D1(n211), .S(n3904), .Y(n83) );
  MUX2IX1 U2637 ( .D0(n139), .D1(n203), .S(n3905), .Y(n75) );
  MUX2IXL U2638 ( .D0(n3893), .D1(n3660), .S(n3912), .Y(n203) );
  MUX2IX1 U2639 ( .D0(n22), .D1(n38), .S(n3896), .Y(n6) );
  MUX2IX1 U2640 ( .D0(n3651), .D1(n86), .S(n3870), .Y(n22) );
  MUX2IX1 U2641 ( .D0(n17), .D1(n33), .S(n3896), .Y(n1) );
  NOR21XL U2642 ( .B(n3985), .A(A[540]), .Y(n1483) );
  NOR21XL U2643 ( .B(n3865), .A(A[524]), .Y(n1547) );
  NOR21XL U2644 ( .B(n3980), .A(A[972]), .Y(n718) );
  NOR21XL U2645 ( .B(n3978), .A(A[965]), .Y(n743) );
  MUX2IX1 U2646 ( .D0(A[285]), .D1(A[797]), .S(n3976), .Y(n1480) );
  NOR21XL U2647 ( .B(n3985), .A(A[541]), .Y(n1479) );
  MUX2IX1 U2648 ( .D0(A[413]), .D1(A[925]), .S(n3984), .Y(n946) );
  OR2X1 U2649 ( .A(n3990), .B(A[221]), .Y(n3836) );
  MUX2IX1 U2650 ( .D0(A[317]), .D1(A[829]), .S(n3866), .Y(n1320) );
  AOI22AXL U2651 ( .A(n3700), .B(A[546]), .D(n3850), .C(n4015), .Y(n3861) );
  MUX2X1 U2652 ( .D0(n714), .D1(n713), .S(n3856), .Y(n3855) );
  MUX2X1 U2653 ( .D0(n1153), .D1(n1154), .S(n3924), .Y(n3725) );
  MUX2IX1 U2654 ( .D0(n3831), .D1(n478), .S(n3910), .Y(n230) );
  MUX2X1 U2655 ( .D0(n1121), .D1(n1122), .S(n3925), .Y(n3831) );
  MUX2X1 U2656 ( .D0(n1628), .D1(n1756), .S(n3916), .Y(n166) );
  MUX2IX1 U2657 ( .D0(n3672), .D1(n3649), .S(n3919), .Y(n134) );
  MUX2AXL U2658 ( .D0(n1209), .D1(n3789), .S(n3929), .Y(n1670) );
  NOR21XL U2659 ( .B(n3983), .A(A[575]), .Y(n1311) );
  AOI22BXL U2660 ( .B(n3843), .A(n3945), .D(n3844), .C(n3955), .Y(n3842) );
  NOR21XL U2661 ( .B(n3988), .A(A[534]), .Y(n1507) );
  NOR21XL U2662 ( .B(n3981), .A(A[622]), .Y(n1149) );
  MUX2AXL U2663 ( .D0(n1201), .D1(n3783), .S(n3927), .Y(n1672) );
  AOI22BXL U2664 ( .B(n3809), .A(n3942), .D(n3810), .C(n3950), .Y(n3808) );
  AND2X1 U2665 ( .A(n699), .B(n3925), .Y(n3740) );
  MUX2X1 U2666 ( .D0(n3792), .D1(n3793), .S(n3931), .Y(n1760) );
  NOR21XL U2667 ( .B(n3982), .A(A[618]), .Y(n1165) );
  MUX2X1 U2668 ( .D0(n3873), .D1(n3874), .S(n3958), .Y(n3886) );
  NOR21XL U2669 ( .B(n4021), .A(A[234]), .Y(n3874) );
  NOR21XL U2670 ( .B(n3981), .A(A[586]), .Y(n1278) );
  MUX2X1 U2671 ( .D0(n1556), .D1(n1555), .S(n3952), .Y(n3891) );
  NOR21XL U2672 ( .B(n3987), .A(A[522]), .Y(n1555) );
  MUX2X1 U2673 ( .D0(n726), .D1(n725), .S(n3960), .Y(n3882) );
  MUX2X1 U2674 ( .D0(n1070), .D1(n1069), .S(n3955), .Y(n3852) );
  MUX2IX1 U2675 ( .D0(n3868), .D1(n3656), .S(n3911), .Y(n211) );
  MUX2X1 U2676 ( .D0(n1198), .D1(n1197), .S(n3951), .Y(n3868) );
  MUX2IX1 U2677 ( .D0(n3658), .D1(n3648), .S(n3915), .Y(n179) );
  INVX1 U2678 ( .A(n1657), .Y(n315) );
  NAND21X1 U2679 ( .B(n3967), .A(n1256), .Y(n1657) );
  NOR21XL U2680 ( .B(n3983), .A(A[594]), .Y(n1256) );
  MUX2IX1 U2681 ( .D0(n3665), .D1(n3887), .S(n3916), .Y(n163) );
  MUX2IX1 U2682 ( .D0(n3652), .D1(n3869), .S(n3910), .Y(n227) );
  MUX2IX1 U2683 ( .D0(n3878), .D1(n3875), .S(n3919), .Y(n131) );
  MUX2X1 U2684 ( .D0(n1524), .D1(n1523), .S(n3960), .Y(n3878) );
  MUX2X1 U2685 ( .D0(n990), .D1(n989), .S(n3958), .Y(n3875) );
  MUX2X1 U2686 ( .D0(n1230), .D1(n1229), .S(n3952), .Y(n3893) );
  NOR21XL U2687 ( .B(n3984), .A(A[602]), .Y(n1229) );
  MUX2IX1 U2688 ( .D0(n3881), .D1(n3777), .S(n3923), .Y(n235) );
  MUX2IX1 U2689 ( .D0(n3657), .D1(n3883), .S(n3919), .Y(n139) );
  MUX2X1 U2690 ( .D0(n958), .D1(n957), .S(n3952), .Y(n3883) );
  NOR21XL U2691 ( .B(n3986), .A(A[539]), .Y(n1487) );
  MUX2X1 U2692 ( .D0(n3786), .D1(n3787), .S(n3931), .Y(n1762) );
  MUX2IX1 U2693 ( .D0(n3730), .D1(n3687), .S(n3909), .Y(n236) );
  MUX2X1 U2694 ( .D0(n1225), .D1(n1226), .S(n3930), .Y(n3752) );
  MUX2IX1 U2695 ( .D0(n133), .D1(n197), .S(n3906), .Y(n69) );
  AND2X1 U2696 ( .A(n690), .B(n3939), .Y(n3737) );
  MUX2IX1 U2697 ( .D0(n165), .D1(n229), .S(n3903), .Y(n101) );
  MUX2IX1 U2698 ( .D0(n3712), .D1(n3686), .S(n3910), .Y(n229) );
  MUX2IX1 U2699 ( .D0(n77), .D1(n109), .S(n3898), .Y(n45) );
  MUX2IX1 U2700 ( .D0(n173), .D1(n237), .S(n3902), .Y(n109) );
  MUX2IX1 U2701 ( .D0(n3713), .D1(n3662), .S(n3909), .Y(n237) );
  MUX2IX1 U2702 ( .D0(n61), .D1(n93), .S(n3900), .Y(n29) );
  MUX2IX1 U2703 ( .D0(n125), .D1(n189), .S(SH[6]), .Y(n61) );
  MUX2IX1 U2704 ( .D0(n3706), .D1(n181), .S(SH[6]), .Y(n53) );
  MUX2IX1 U2705 ( .D0(n149), .D1(n213), .S(n3904), .Y(n85) );
  MUX2IX1 U2706 ( .D0(n3708), .D1(n3681), .S(n3911), .Y(n214) );
  MUX2IX1 U2707 ( .D0(n3779), .D1(n3780), .S(n3907), .Y(n3778) );
  MUX2X1 U2708 ( .D0(n1185), .D1(n1186), .S(n3927), .Y(n3708) );
  AOI22AXL U2709 ( .A(n1437), .B(n3956), .D(n3711), .C(n1438), .Y(n3710) );
  MUX2IX1 U2710 ( .D0(n174), .D1(n238), .S(n3902), .Y(n110) );
  MUX2IX1 U2711 ( .D0(n142), .D1(n206), .S(n3905), .Y(n78) );
  MUX2IX1 U2712 ( .D0(n3719), .D1(n3664), .S(n3909), .Y(n238) );
  MUX2IX1 U2713 ( .D0(n70), .D1(n102), .S(n3900), .Y(n38) );
  MUX2IX1 U2714 ( .D0(n134), .D1(n198), .S(n3906), .Y(n70) );
  MUX2IX1 U2715 ( .D0(n166), .D1(n230), .S(n3903), .Y(n102) );
  MUX2IX1 U2716 ( .D0(n3716), .D1(n3717), .S(n3913), .Y(n198) );
  INVX1 U2717 ( .A(n3950), .Y(n3924) );
  MUX2X1 U2718 ( .D0(n1669), .D1(n1797), .S(n3912), .Y(n207) );
  MUX2BXL U2719 ( .D0(n1653), .D1(n3761), .S(n3913), .Y(n191) );
  AOI22BXL U2720 ( .B(n3812), .A(n3940), .D(n3813), .C(n3958), .Y(n3811) );
  MUX2BXL U2721 ( .D0(n1637), .D1(n3762), .S(n3915), .Y(n175) );
  MUX2IX1 U2722 ( .D0(n148), .D1(n212), .S(n3904), .Y(n84) );
  MUX2IX1 U2723 ( .D0(n68), .D1(n100), .S(n3900), .Y(n36) );
  MUX2IX1 U2724 ( .D0(n132), .D1(n196), .S(n3906), .Y(n68) );
  MUX2IX1 U2725 ( .D0(n164), .D1(n228), .S(n3903), .Y(n100) );
  MUX2IX1 U2726 ( .D0(n124), .D1(n188), .S(n3907), .Y(n60) );
  MUX2IX1 U2727 ( .D0(n76), .D1(n108), .S(n3898), .Y(n44) );
  MUX2IX1 U2728 ( .D0(n140), .D1(n204), .S(n3905), .Y(n76) );
  MUX2IX1 U2729 ( .D0(n172), .D1(n236), .S(n3902), .Y(n108) );
  MUX2X1 U2730 ( .D0(n1602), .D1(n1730), .S(n3919), .Y(n140) );
  MUX2IX1 U2731 ( .D0(n5), .D1(n13), .S(SH[3]), .Y(B[4]) );
  MUX2IX1 U2732 ( .D0(n21), .D1(n37), .S(n3896), .Y(n5) );
  MUX2IX1 U2733 ( .D0(n29), .D1(n45), .S(n3895), .Y(n13) );
  MUX2IX1 U2734 ( .D0(n69), .D1(n101), .S(n3900), .Y(n37) );
  MUX2X1 U2735 ( .D0(n1607), .D1(n1735), .S(n3918), .Y(n145) );
  MUX2BXL U2736 ( .D0(n1671), .D1(n3728), .S(n3912), .Y(n209) );
  MUX2X1 U2737 ( .D0(n1237), .D1(n1238), .S(n3930), .Y(n3756) );
  MUX2IX1 U2738 ( .D0(n18), .D1(n34), .S(n3896), .Y(n2) );
  MUX2IX1 U2739 ( .D0(n3), .D1(n11), .S(SH[3]), .Y(B[2]) );
  MUX2IX1 U2740 ( .D0(n19), .D1(n35), .S(n3896), .Y(n3) );
  MUX2IX1 U2741 ( .D0(n49), .D1(n81), .S(n3900), .Y(n17) );
  MUX2BXL U2742 ( .D0(n3775), .D1(n177), .S(n3907), .Y(n49) );
  MUX2IX1 U2743 ( .D0(n145), .D1(n209), .S(n3905), .Y(n81) );
  MUX2X1 U2744 ( .D0(n1639), .D1(n1767), .S(n3915), .Y(n177) );
  MUX2IX1 U2745 ( .D0(n65), .D1(n97), .S(n3900), .Y(n33) );
  MUX2IX1 U2746 ( .D0(n129), .D1(n193), .S(n3906), .Y(n65) );
  MUX2IX1 U2747 ( .D0(n161), .D1(n225), .S(n3903), .Y(n97) );
  MUX2AXL U2748 ( .D0(n121), .D1(n3729), .S(n3907), .Y(n57) );
  MUX2X1 U2749 ( .D0(n305), .D1(n3757), .S(n3914), .Y(n3729) );
  INVX1 U2750 ( .A(SH[9]), .Y(n4035) );
  BUFX1 U2751 ( .A(SH[9]), .Y(n3845) );
  BUFX1 U2752 ( .A(SH[9]), .Y(n3854) );
  INVXL U2753 ( .A(n4006), .Y(n4004) );
  INVX1 U2754 ( .A(n4027), .Y(n4024) );
  INVX1 U2755 ( .A(n3908), .Y(n3907) );
  INVX1 U2756 ( .A(SH[8]), .Y(n3969) );
  INVX1 U2757 ( .A(n4033), .Y(n4014) );
  AND2X1 U2758 ( .A(n752), .B(n3939), .Y(n3648) );
  MUX2X1 U2759 ( .D0(n977), .D1(n978), .S(n3928), .Y(n3649) );
  MUX2X1 U2760 ( .D0(n985), .D1(n986), .S(n3928), .Y(n3650) );
  INVXL U2761 ( .A(n3854), .Y(n3853) );
  INVXL U2762 ( .A(n4027), .Y(n4026) );
  INVXL U2763 ( .A(n4027), .Y(n4025) );
  MUX2X1 U2764 ( .D0(n3710), .D1(n3680), .S(n3918), .Y(n3651) );
  MUX2X1 U2765 ( .D0(n3683), .D1(n1134), .S(n3924), .Y(n3652) );
  AND2X1 U2766 ( .A(n1293), .B(n3938), .Y(n3653) );
  AOI22X1 U2767 ( .A(n1390), .B(n3943), .C(n1389), .D(n3957), .Y(n3654) );
  AOI22X1 U2768 ( .A(n1408), .B(n3943), .C(n1407), .D(n3953), .Y(n3655) );
  INVXL U2769 ( .A(n3969), .Y(n3965) );
  INVX1 U2770 ( .A(n3966), .Y(n3952) );
  MUX2X1 U2771 ( .D0(n637), .D1(n638), .S(n3935), .Y(n3656) );
  MUX2X1 U2772 ( .D0(n1491), .D1(n1492), .S(n3934), .Y(n3657) );
  AND2X1 U2773 ( .A(n1302), .B(n3938), .Y(n3658) );
  MUX2X1 U2774 ( .D0(n1073), .D1(n1074), .S(n3926), .Y(n3659) );
  MUX2X1 U2775 ( .D0(n669), .D1(n670), .S(n3934), .Y(n3660) );
  MUX2X1 U2776 ( .D0(n593), .D1(n594), .S(n3930), .Y(n3661) );
  AOI22X1 U2777 ( .A(n510), .B(n3945), .C(n509), .D(n3960), .Y(n3662) );
  AOI22X1 U2778 ( .A(n1028), .B(n3940), .C(n1027), .D(n3957), .Y(n3663) );
  AOI22X1 U2779 ( .A(n503), .B(n3955), .C(n3945), .D(n3745), .Y(n3664) );
  MUX2X1 U2780 ( .D0(n1363), .D1(n1364), .S(n3932), .Y(n3665) );
  MUX2X1 U2781 ( .D0(n1531), .D1(n1532), .S(n3937), .Y(n3666) );
  MUX2X1 U2782 ( .D0(n673), .D1(n674), .S(n3935), .Y(n3667) );
  MUX2X1 U2783 ( .D0(n1535), .D1(n1536), .S(n3938), .Y(n3668) );
  MUX2X1 U2784 ( .D0(n937), .D1(n938), .S(n3929), .Y(n3669) );
  MUX2X1 U2785 ( .D0(n773), .D1(n774), .S(n3931), .Y(n3670) );
  MUX2X1 U2786 ( .D0(n769), .D1(n770), .S(n3931), .Y(n3671) );
  MUX2X1 U2787 ( .D0(n1511), .D1(n1512), .S(n3937), .Y(n3672) );
  MUX2X1 U2788 ( .D0(n1479), .D1(n1480), .S(n3934), .Y(n3673) );
  MUX2X1 U2789 ( .D0(n1177), .D1(n1178), .S(n3927), .Y(n3674) );
  MUX2X1 U2790 ( .D0(n1515), .D1(n1516), .S(n3937), .Y(n3675) );
  MUX2X1 U2791 ( .D0(n1355), .D1(n1356), .S(n3932), .Y(n3676) );
  MUX2X1 U2792 ( .D0(n1157), .D1(n1158), .S(n3924), .Y(n3677) );
  MUX2X1 U2793 ( .D0(n1165), .D1(n1166), .S(n3924), .Y(n3678) );
  MUX2X1 U2794 ( .D0(n633), .D1(n634), .S(n3936), .Y(n3679) );
  AOI22X1 U2795 ( .A(n903), .B(n3951), .C(n3941), .D(n3766), .Y(n3680) );
  MUX2X1 U2796 ( .D0(n625), .D1(n626), .S(n3936), .Y(n3681) );
  MUX2X1 U2797 ( .D0(n629), .D1(n630), .S(n3935), .Y(n3682) );
  NOR2X1 U2798 ( .A(n4014), .B(A[626]), .Y(n3683) );
  MUX2X1 U2799 ( .D0(n1519), .D1(n1520), .S(n3937), .Y(n3684) );
  MUX2IX1 U2800 ( .D0(n3790), .D1(n3791), .S(n3935), .Y(n3685) );
  AOI22X1 U2801 ( .A(n558), .B(n3944), .C(n557), .D(n3961), .Y(n3686) );
  AOI22X1 U2802 ( .A(n516), .B(n3945), .C(n515), .D(n3954), .Y(n3687) );
  AOI22X1 U2803 ( .A(n1444), .B(n3872), .C(n1443), .D(n3953), .Y(n3688) );
  AOI22X1 U2804 ( .A(n3817), .B(n3941), .C(n1015), .D(n3958), .Y(n3689) );
  AOI22X1 U2805 ( .A(n564), .B(n3944), .C(n563), .D(n3953), .Y(n3690) );
  AOI22X1 U2806 ( .A(n498), .B(n3945), .C(n497), .D(n3960), .Y(n3691) );
  AOI22X1 U2807 ( .A(n1022), .B(n3940), .C(n1021), .D(n3958), .Y(n3692) );
  AOI22X1 U2808 ( .A(n862), .B(n3941), .C(n861), .D(n3952), .Y(n3693) );
  AOI22X1 U2809 ( .A(n916), .B(n3941), .C(n915), .D(n3950), .Y(n3694) );
  AOI22X1 U2810 ( .A(n856), .B(n3941), .C(n855), .D(n3952), .Y(n3695) );
  AOI22X1 U2811 ( .A(n820), .B(n3942), .C(n819), .D(n3952), .Y(n3696) );
  AOI22X1 U2812 ( .A(n892), .B(n3943), .C(n891), .D(n3951), .Y(n3697) );
  AOI22X1 U2813 ( .A(n843), .B(n3952), .C(n3943), .D(n3767), .Y(n3698) );
  AND2X1 U2814 ( .A(n743), .B(n3939), .Y(n3699) );
  INVXL U2815 ( .A(n3969), .Y(n3967) );
  INVXL U2816 ( .A(n3969), .Y(n3966) );
  INVX1 U2817 ( .A(n4032), .Y(n4015) );
  INVX1 U2818 ( .A(n4030), .Y(n4019) );
  AO22XL U2819 ( .A(n4020), .B(A[509]), .C(SH[9]), .D(A[1021]), .Y(n3745) );
  INVXL U2820 ( .A(SH[9]), .Y(n4037) );
  INVX1 U2821 ( .A(n3845), .Y(n4006) );
  INVX1 U2822 ( .A(n4007), .Y(n3700) );
  NOR21XL U2823 ( .B(n4031), .A(A[607]), .Y(n1209) );
  INVXL U2824 ( .A(n4035), .Y(n4033) );
  MUX2IX1 U2825 ( .D0(n60), .D1(n92), .S(n3899), .Y(n28) );
  MUX2IX1 U2826 ( .D0(n52), .D1(n84), .S(n3899), .Y(n20) );
  MUX2IX1 U2827 ( .D0(n53), .D1(n85), .S(n3899), .Y(n21) );
  MUX2IX1 U2828 ( .D0(n51), .D1(n83), .S(n3899), .Y(n19) );
  MUX2IX1 U2829 ( .D0(n3778), .D1(n214), .S(n3899), .Y(n86) );
  AOI22BXL U2830 ( .B(n3822), .A(n3966), .D(n3823), .C(n3959), .Y(n3821) );
  EORX1 U2831 ( .A(n1450), .B(n3872), .C(n3860), .D(n3872), .Y(n3859) );
  AOI22BXL U2832 ( .B(n3819), .A(n3965), .D(n3820), .C(n3955), .Y(n3818) );
  NOR21XL U2833 ( .B(n4030), .A(A[620]), .Y(n1157) );
  NOR21XL U2834 ( .B(n4029), .A(A[609]), .Y(n1201) );
  INVXL U2835 ( .A(n4007), .Y(n3701) );
  INVX1 U2836 ( .A(n4034), .Y(n4007) );
  MUX2IX1 U2837 ( .D0(n1), .D1(n9), .S(SH[3]), .Y(B[0]) );
  INVXL U2838 ( .A(n3703), .Y(n4021) );
  INVXL U2839 ( .A(n4034), .Y(n4011) );
  INVX1 U2840 ( .A(n3935), .Y(n3702) );
  MUX2IX1 U2841 ( .D0(n141), .D1(n205), .S(n3905), .Y(n77) );
  MUX2X1 U2842 ( .D0(n1311), .D1(n1312), .S(n3930), .Y(n3747) );
  MUX2IX1 U2843 ( .D0(n3837), .D1(n3836), .S(n3702), .Y(n3835) );
  AND2XL U2844 ( .A(n687), .B(n3939), .Y(n3717) );
  INVX1 U2845 ( .A(n1660), .Y(n3716) );
  MUX2X1 U2846 ( .D0(n1193), .D1(n1194), .S(n3927), .Y(n3731) );
  AND2XL U2847 ( .A(n696), .B(n3939), .Y(n3734) );
  INVX1 U2848 ( .A(n3854), .Y(n4018) );
  INVX1 U2849 ( .A(n3922), .Y(n3919) );
  INVX1 U2850 ( .A(n3923), .Y(n3915) );
  INVX1 U2851 ( .A(n3923), .Y(n3911) );
  MUX2IX1 U2852 ( .D0(n3772), .D1(n3739), .S(n3915), .Y(n178) );
  MUX2X2 U2853 ( .D0(n1189), .D1(n1190), .S(n3927), .Y(n3709) );
  NOR2XL U2854 ( .A(n3993), .B(A[354]), .Y(n1198) );
  INVXL U2855 ( .A(n4012), .Y(n3703) );
  INVXL U2856 ( .A(SH[9]), .Y(n4012) );
  INVXL U2857 ( .A(n3853), .Y(n3994) );
  INVXL U2858 ( .A(n3950), .Y(n3944) );
  INVX1 U2859 ( .A(n3968), .Y(n3948) );
  INVXL U2860 ( .A(n3922), .Y(n3912) );
  MUX2IXL U2861 ( .D0(n941), .D1(n942), .S(n3929), .Y(n1733) );
  MUX2IXL U2862 ( .D0(A[404]), .D1(A[916]), .S(n3970), .Y(n982) );
  MUX2XL U2863 ( .D0(n717), .D1(n718), .S(n3933), .Y(n3794) );
  MUX2XL U2864 ( .D0(A[476]), .D1(A[988]), .S(n3976), .Y(n3829) );
  OR2XL U2865 ( .A(n3989), .B(A[220]), .Y(n3828) );
  INVX1 U2866 ( .A(n3933), .Y(n3856) );
  INVX1 U2867 ( .A(n4031), .Y(n4017) );
  INVX1 U2868 ( .A(n3967), .Y(n3955) );
  INVXL U2869 ( .A(n3969), .Y(n3929) );
  INVX1 U2870 ( .A(n3967), .Y(n3958) );
  MUX2XL U2871 ( .D0(n997), .D1(n998), .S(n3927), .Y(n3732) );
  MUX2IX1 U2872 ( .D0(n3754), .D1(n3749), .S(n3911), .Y(n218) );
  NAND2X1 U2873 ( .A(n3852), .B(n3921), .Y(n115) );
  MUX2IX1 U2874 ( .D0(n116), .D1(n180), .S(n3907), .Y(n52) );
  MUX2XL U2875 ( .D0(n1181), .D1(n1182), .S(n3927), .Y(n3721) );
  AND2X1 U2876 ( .A(n684), .B(n3966), .Y(n3741) );
  MUX2IXL U2877 ( .D0(n961), .D1(n962), .S(n3928), .Y(n1728) );
  MUX2XL U2878 ( .D0(A[477]), .D1(A[989]), .S(n3976), .Y(n3837) );
  NOR21XL U2879 ( .B(n3980), .A(A[716]), .Y(n717) );
  MUX2XL U2880 ( .D0(n1081), .D1(n1082), .S(n3926), .Y(n3841) );
  AO22XL U2881 ( .A(n4015), .B(A[254]), .C(n3996), .D(A[766]), .Y(n497) );
  AO22XL U2882 ( .A(n4026), .B(A[421]), .C(n3997), .D(A[933]), .Y(n3766) );
  AO22X1 U2883 ( .A(n4008), .B(A[504]), .C(n3701), .D(A[1016]), .Y(n534) );
  INVXL U2884 ( .A(n3969), .Y(n3930) );
  INVXL U2885 ( .A(n3968), .Y(n3954) );
  INVXL U2886 ( .A(n3949), .Y(n3928) );
  INVX2 U2887 ( .A(n3923), .Y(n3909) );
  MUX2IXL U2888 ( .D0(n3771), .D1(n3742), .S(n3914), .Y(n183) );
  MUX2BXL U2889 ( .D0(n1685), .D1(n3764), .S(n3910), .Y(n223) );
  MUX2X1 U2890 ( .D0(n617), .D1(n618), .S(n3936), .Y(n3735) );
  AOI22X1 U2891 ( .A(n1426), .B(n3872), .C(n1425), .D(n3956), .Y(n3723) );
  MUX2IXL U2892 ( .D0(n613), .D1(n614), .S(n3936), .Y(n1807) );
  MUX2IXL U2893 ( .D0(n789), .D1(n790), .S(n3931), .Y(n1759) );
  INVXL U2894 ( .A(n3944), .Y(n3802) );
  MUX2IXL U2895 ( .D0(A[493]), .D1(A[1005]), .S(n3973), .Y(n594) );
  MUX2XL U2896 ( .D0(n733), .D1(n734), .S(n3932), .Y(n3757) );
  OAI22XL U2897 ( .A(n3998), .B(n3863), .C(n4025), .D(n3864), .Y(n3817) );
  AO22X1 U2898 ( .A(n575), .B(n3953), .C(n3944), .D(n3770), .Y(n1816) );
  NOR21XL U2899 ( .B(n3982), .A(A[837]), .Y(n1293) );
  NOR21XL U2900 ( .B(n3866), .A(A[629]), .Y(n1121) );
  MUX2AXL U2901 ( .D0(n1213), .D1(n3788), .S(n3929), .Y(n1669) );
  AO22XL U2902 ( .A(n3853), .B(A[296]), .C(n4004), .D(A[808]), .Y(n3769) );
  INVX1 U2903 ( .A(n3968), .Y(n3949) );
  INVX1 U2904 ( .A(n3966), .Y(n3960) );
  INVX1 U2905 ( .A(n3967), .Y(n3957) );
  INVX1 U2906 ( .A(n3908), .Y(n3906) );
  INVX1 U2907 ( .A(n3908), .Y(n3902) );
  INVX1 U2908 ( .A(n3922), .Y(n3914) );
  MUX2X1 U2909 ( .D0(n1129), .D1(n1130), .S(n3925), .Y(n3736) );
  MUX2XL U2910 ( .D0(n597), .D1(n598), .S(n3935), .Y(n3707) );
  MUX2IX1 U2911 ( .D0(n1563), .D1(n1564), .S(n3930), .Y(n1583) );
  MUX2IXL U2912 ( .D0(n3821), .D1(n3824), .S(n3917), .Y(n159) );
  MUX2IX1 U2913 ( .D0(n152), .D1(n216), .S(n3904), .Y(n88) );
  MUX2IX1 U2914 ( .D0(n3688), .D1(n3718), .S(n3918), .Y(n149) );
  MUX2BX1 U2915 ( .D0(n1672), .D1(n3795), .S(n3912), .Y(n210) );
  MUX2IX1 U2916 ( .D0(n156), .D1(n220), .S(n3904), .Y(n92) );
  NAND2X1 U2917 ( .A(n3830), .B(n3921), .Y(n3706) );
  INVXL U2918 ( .A(n3965), .Y(n3711) );
  MUX2IX1 U2919 ( .D0(n157), .D1(n221), .S(n3903), .Y(n93) );
  MUX2XL U2920 ( .D0(n1097), .D1(n1098), .S(n3925), .Y(n3730) );
  MUX2XL U2921 ( .D0(n1101), .D1(n1102), .S(n3965), .Y(n3777) );
  MUX2IX1 U2922 ( .D0(n949), .D1(n950), .S(n3929), .Y(n1731) );
  MUX2X2 U2923 ( .D0(n1603), .D1(n1731), .S(n3918), .Y(n141) );
  MUX2X1 U2924 ( .D0(n1634), .D1(n1762), .S(n3915), .Y(n172) );
  MUX2X1 U2925 ( .D0(n1686), .D1(n1814), .S(n3910), .Y(n224) );
  MUX2IX1 U2926 ( .D0(n1499), .D1(n1500), .S(n3936), .Y(n1599) );
  MUX2X1 U2927 ( .D0(n1599), .D1(n1727), .S(n3919), .Y(n137) );
  INVXL U2928 ( .A(n3926), .Y(n3720) );
  AOI22XL U2929 ( .A(n1378), .B(n3943), .C(n1377), .D(n3957), .Y(n3724) );
  NAND2X1 U2930 ( .A(n3659), .B(n3921), .Y(n114) );
  AND2XL U2931 ( .A(n693), .B(n3925), .Y(n3743) );
  AND2XL U2932 ( .A(n702), .B(n3941), .Y(n3744) );
  AND2XL U2933 ( .A(n740), .B(n3925), .Y(n3742) );
  MUX2XL U2934 ( .D0(n1471), .D1(n1472), .S(n3934), .Y(n3765) );
  AOI22XL U2935 ( .A(n4018), .B(A[178]), .C(n4001), .D(A[690]), .Y(n3857) );
  MUX2IXL U2936 ( .D0(n761), .D1(n762), .S(n3932), .Y(n1766) );
  MUX2IX1 U2937 ( .D0(n25), .D1(n41), .S(n3895), .Y(n9) );
  NOR21XL U2938 ( .B(n3984), .A(A[565]), .Y(n1351) );
  MUX2IXL U2939 ( .D0(A[472]), .D1(A[984]), .S(n3972), .Y(n678) );
  MUX2XL U2940 ( .D0(n1332), .D1(n1331), .S(n3961), .Y(n3879) );
  MUX2IXL U2941 ( .D0(A[283]), .D1(A[795]), .S(n3977), .Y(n1488) );
  MUX2IXL U2942 ( .D0(A[190]), .D1(A[702]), .S(n3972), .Y(n765) );
  NAND21XL U2943 ( .B(n1709), .A(n3921), .Y(n119) );
  OR2XL U2944 ( .A(n3979), .B(A[350]), .Y(n3788) );
  NOR2XL U2945 ( .A(n3996), .B(A[391]), .Y(n1050) );
  NOR2XL U2946 ( .A(n3995), .B(A[131]), .Y(n1065) );
  NOR2XL U2947 ( .A(n3994), .B(A[128]), .Y(n1077) );
  MUX2XL U2948 ( .D0(n1085), .D1(n1086), .S(n3926), .Y(n3751) );
  NOR2XL U2949 ( .A(n3994), .B(A[382]), .Y(n1086) );
  AO22XL U2950 ( .A(n4024), .B(A[433]), .C(n4001), .D(A[945]), .Y(n3768) );
  AO22XL U2951 ( .A(n831), .B(n3952), .C(n3943), .D(n3768), .Y(n1752) );
  INVXL U2952 ( .A(n4037), .Y(n3972) );
  INVXL U2953 ( .A(n4037), .Y(n3970) );
  INVXL U2954 ( .A(n4010), .Y(n4005) );
  INVXL U2955 ( .A(n3854), .Y(n4020) );
  INVXL U2956 ( .A(n3845), .Y(n4009) );
  INVXL U2957 ( .A(n3854), .Y(n4008) );
  INVXL U2958 ( .A(n4034), .Y(n4010) );
  INVXL U2959 ( .A(n3954), .Y(n3945) );
  INVXL U2960 ( .A(n3967), .Y(n3953) );
  INVXL U2961 ( .A(n3968), .Y(n3946) );
  INVXL U2962 ( .A(SH[8]), .Y(n3947) );
  INVXL U2963 ( .A(n3967), .Y(n3959) );
  INVXL U2964 ( .A(n3968), .Y(n3951) );
  INVXL U2965 ( .A(n3967), .Y(n3956) );
  INVXL U2966 ( .A(n3966), .Y(n3962) );
  INVXL U2967 ( .A(n3965), .Y(n3963) );
  INVXL U2968 ( .A(n3965), .Y(n3964) );
  INVXL U2969 ( .A(n3923), .Y(n3917) );
  INVXL U2970 ( .A(n3922), .Y(n3921) );
  INVXL U2971 ( .A(n3908), .Y(n3904) );
  INVXL U2972 ( .A(n3901), .Y(n3900) );
  MUX2IXL U2973 ( .D0(n160), .D1(n224), .S(n3903), .Y(n96) );
  MUX2X1 U2974 ( .D0(n981), .D1(n982), .S(n3928), .Y(n3704) );
  MUX2X2 U2975 ( .D0(n1547), .D1(n1548), .S(n3937), .Y(n3705) );
  NAND2XL U2976 ( .A(n3773), .B(n3921), .Y(n120) );
  MUX2X2 U2977 ( .D0(n1125), .D1(n1126), .S(n3925), .Y(n3712) );
  MUX2X2 U2978 ( .D0(n1093), .D1(n1094), .S(n3925), .Y(n3713) );
  AOI22X1 U2979 ( .A(n910), .B(n3940), .C(n909), .D(n3963), .Y(n3718) );
  MUX2X2 U2980 ( .D0(n1090), .D1(n1089), .S(n3720), .Y(n3719) );
  MUX2IX1 U2981 ( .D0(n3721), .D1(n3685), .S(n3911), .Y(n215) );
  MUX2X2 U2982 ( .D0(n1323), .D1(n1324), .S(n3930), .Y(n3722) );
  MUX2IXL U2983 ( .D0(n653), .D1(n654), .S(n3935), .Y(n1797) );
  MUX2IX1 U2984 ( .D0(n3723), .D1(n3697), .S(n3917), .Y(n152) );
  MUX2IX1 U2985 ( .D0(n3724), .D1(n3698), .S(n3917), .Y(n160) );
  MUX2IX1 U2986 ( .D0(n3725), .D1(n3661), .S(n3910), .Y(n222) );
  AOI22X1 U2987 ( .A(n1396), .B(n3965), .C(n1395), .D(n3959), .Y(n3726) );
  MUX2IX1 U2988 ( .D0(n1559), .D1(n1560), .S(n3924), .Y(n1584) );
  MUX2AX2 U2989 ( .D0(n3727), .D1(n1751), .S(n3916), .Y(n161) );
  MUX2XL U2990 ( .D0(n1371), .D1(n1372), .S(n3933), .Y(n3727) );
  MUX2XL U2991 ( .D0(n645), .D1(n646), .S(n3934), .Y(n3728) );
  MUX2IX2 U2992 ( .D0(n130), .D1(n194), .S(n3906), .Y(n66) );
  NAND2XL U2993 ( .A(n3763), .B(n3921), .Y(n116) );
  AND2XL U2994 ( .A(n3755), .B(n3921), .Y(n3775) );
  MUX2IXL U2995 ( .D0(n73), .D1(n105), .S(n3898), .Y(n41) );
  MUX2IXL U2996 ( .D0(n137), .D1(n201), .S(n3905), .Y(n73) );
  MUX2IXL U2997 ( .D0(n169), .D1(n233), .S(n3902), .Y(n105) );
  MUX2IXL U2998 ( .D0(n3756), .D1(n3760), .S(n3912), .Y(n201) );
  MUX2IX1 U2999 ( .D0(n3666), .D1(n3732), .S(n3920), .Y(n129) );
  NAND2XL U3000 ( .A(n746), .B(n3939), .Y(n1771) );
  NAND2XL U3001 ( .A(n737), .B(n3939), .Y(n1774) );
  NAND2XL U3002 ( .A(n749), .B(n3872), .Y(n1770) );
  NOR21XL U3003 ( .B(n3978), .A(A[962]), .Y(n752) );
  MUX2IX1 U3004 ( .D0(n3674), .D1(n3735), .S(n3911), .Y(n216) );
  MUX2IX1 U3005 ( .D0(n1145), .D1(n1146), .S(n3924), .Y(n1686) );
  MUX2IXL U3006 ( .D0(n1527), .D1(n1528), .S(n3938), .Y(n1592) );
  NAND2XL U3007 ( .A(n1299), .B(n3938), .Y(n1642) );
  MUX2IXL U3008 ( .D0(n1335), .D1(n1336), .S(n3931), .Y(n1632) );
  MUX2IXL U3009 ( .D0(n1343), .D1(n1344), .S(n3932), .Y(n1630) );
  MUX2IXL U3010 ( .D0(n1347), .D1(n1348), .S(n3932), .Y(n1629) );
  NAND2XL U3011 ( .A(n1308), .B(n3938), .Y(n1639) );
  NAND2XL U3012 ( .A(n1296), .B(n3938), .Y(n1643) );
  MUX2X2 U3013 ( .D0(n1616), .D1(n1744), .S(n3917), .Y(n154) );
  AND2XL U3014 ( .A(n681), .B(n3939), .Y(n3738) );
  AND2X1 U3015 ( .A(n755), .B(n3927), .Y(n3739) );
  MUX2IX1 U3016 ( .D0(A[277]), .D1(A[789]), .S(n3975), .Y(n1512) );
  MUX2IXL U3017 ( .D0(A[268]), .D1(A[780]), .S(n3973), .Y(n1548) );
  MUX2IXL U3018 ( .D0(A[269]), .D1(A[781]), .S(n3973), .Y(n1544) );
  MUX2X2 U3019 ( .D0(n1221), .D1(n1222), .S(n3929), .Y(n3746) );
  AO22XL U3020 ( .A(n4014), .B(A[141]), .C(n4028), .D(A[653]), .Y(n1015) );
  AO22XL U3021 ( .A(n3853), .B(A[505]), .C(n3999), .D(A[1017]), .Y(n528) );
  MUX2IXL U3022 ( .D0(n1507), .D1(n3748), .S(n3936), .Y(n1597) );
  MUX2IXL U3023 ( .D0(A[278]), .D1(A[790]), .S(n3975), .Y(n3748) );
  INVXL U3024 ( .A(n3944), .Y(n3814) );
  MUX2XL U3025 ( .D0(n609), .D1(n610), .S(n3936), .Y(n3749) );
  MUX2XL U3026 ( .D0(n1539), .D1(n1540), .S(n3937), .Y(n3750) );
  NOR2XL U3027 ( .A(n3994), .B(A[383]), .Y(n1082) );
  MUX2IXL U3028 ( .D0(A[272]), .D1(A[784]), .S(n3974), .Y(n1532) );
  MUX2IXL U3029 ( .D0(n585), .D1(n586), .S(n3937), .Y(n1814) );
  MUX2IXL U3030 ( .D0(n3796), .D1(n3797), .S(n3935), .Y(n3795) );
  OR2XL U3031 ( .A(n3989), .B(A[225]), .Y(n3796) );
  MUX2IXL U3032 ( .D0(n3799), .D1(n3800), .S(n3935), .Y(n3798) );
  OR2XL U3033 ( .A(n3989), .B(A[223]), .Y(n3799) );
  MUX2IXL U3034 ( .D0(A[184]), .D1(A[696]), .S(n4032), .Y(n789) );
  OAI22AXL U3035 ( .D(n3964), .C(n3781), .A(n3782), .B(n3961), .Y(n1735) );
  MUX2XL U3036 ( .D0(n1233), .D1(n1234), .S(n3930), .Y(n3753) );
  MUX2IXL U3037 ( .D0(A[415]), .D1(A[927]), .S(n3988), .Y(n938) );
  MUX2IXL U3038 ( .D0(A[315]), .D1(A[827]), .S(n3854), .Y(n1328) );
  MUX2IXL U3039 ( .D0(A[414]), .D1(A[926]), .S(n4032), .Y(n942) );
  MUX2IXL U3040 ( .D0(A[318]), .D1(A[830]), .S(n3703), .Y(n1316) );
  MUX2IXL U3041 ( .D0(n1475), .D1(n1476), .S(n3933), .Y(n1605) );
  MUX2IXL U3042 ( .D0(n1173), .D1(n1174), .S(n3927), .Y(n1679) );
  MUX2IXL U3043 ( .D0(A[407]), .D1(A[919]), .S(n3972), .Y(n970) );
  MUX2IXL U3044 ( .D0(n965), .D1(n966), .S(n3928), .Y(n1727) );
  MUX2IXL U3045 ( .D0(A[408]), .D1(A[920]), .S(n3970), .Y(n966) );
  MUX2IXL U3046 ( .D0(A[405]), .D1(A[917]), .S(n3970), .Y(n978) );
  MUX2IXL U3047 ( .D0(A[411]), .D1(A[923]), .S(n3970), .Y(n954) );
  MUX2IXL U3048 ( .D0(A[403]), .D1(A[915]), .S(n3970), .Y(n986) );
  MUX2IXL U3049 ( .D0(A[406]), .D1(A[918]), .S(n3970), .Y(n974) );
  MUX2IXL U3050 ( .D0(A[305]), .D1(A[817]), .S(n3972), .Y(n1368) );
  MUX2IXL U3051 ( .D0(A[304]), .D1(A[816]), .S(n3972), .Y(n1372) );
  MUX2IXL U3052 ( .D0(A[307]), .D1(A[819]), .S(n3972), .Y(n1360) );
  NOR21XL U3053 ( .B(n4022), .A(A[370]), .Y(n1134) );
  MUX2IXL U3054 ( .D0(n1205), .D1(n1206), .S(n3929), .Y(n1671) );
  MUX2IXL U3055 ( .D0(n1339), .D1(n1340), .S(n3932), .Y(n1631) );
  MUX2IXL U3056 ( .D0(n1487), .D1(n1488), .S(n3934), .Y(n1602) );
  MUX2IXL U3057 ( .D0(n729), .D1(n730), .S(n3933), .Y(n1776) );
  MUX2IXL U3058 ( .D0(A[191]), .D1(A[703]), .S(n3972), .Y(n761) );
  MUX2IXL U3059 ( .D0(A[480]), .D1(A[992]), .S(n3977), .Y(n646) );
  MUX2IXL U3060 ( .D0(A[281]), .D1(A[793]), .S(n3977), .Y(n1496) );
  MUX2IXL U3061 ( .D0(A[409]), .D1(A[921]), .S(n3970), .Y(n962) );
  AO22XL U3062 ( .A(n4021), .B(A[291]), .C(n4003), .D(A[803]), .Y(n1450) );
  NOR21XL U3063 ( .B(n3986), .A(A[605]), .Y(n1217) );
  MUX2XL U3064 ( .D0(n1169), .D1(n1170), .S(n3931), .Y(n3754) );
  MUX2XL U3065 ( .D0(n1077), .D1(n1078), .S(n3926), .Y(n3755) );
  NOR2XL U3066 ( .A(n3994), .B(A[129]), .Y(n1073) );
  MUX2XL U3067 ( .D0(n1061), .D1(n1062), .S(n3926), .Y(n3830) );
  NOR2XL U3068 ( .A(n3995), .B(A[132]), .Y(n1061) );
  NOR2X1 U3069 ( .A(n3992), .B(A[362]), .Y(n1166) );
  NAND2XL U3070 ( .A(n758), .B(n3937), .Y(n1767) );
  MUX2XL U3071 ( .D0(n1161), .D1(n1162), .S(n3924), .Y(n3758) );
  MUX2XL U3072 ( .D0(n705), .D1(n706), .S(n3934), .Y(n3759) );
  MUX2XL U3073 ( .D0(n677), .D1(n678), .S(n3934), .Y(n3760) );
  MUX2XL U3074 ( .D0(n709), .D1(n710), .S(n3932), .Y(n3761) );
  MUX2XL U3075 ( .D0(n765), .D1(n766), .S(n3932), .Y(n3762) );
  NOR21XL U3076 ( .B(n3984), .A(A[570]), .Y(n1331) );
  MUX2XL U3077 ( .D0(n1065), .D1(n1066), .S(n3926), .Y(n3763) );
  MUX2XL U3078 ( .D0(n589), .D1(n590), .S(n3936), .Y(n3764) );
  MUX2IXL U3079 ( .D0(A[473]), .D1(A[985]), .S(n3972), .Y(n674) );
  AO22XL U3080 ( .A(n4020), .B(A[243]), .C(n4002), .D(A[755]), .Y(n563) );
  AO22X1 U3081 ( .A(n4024), .B(A[431]), .C(n4001), .D(A[943]), .Y(n3767) );
  AO22XL U3082 ( .A(n4022), .B(A[251]), .C(n3854), .D(A[763]), .Y(n515) );
  AO22XL U3083 ( .A(n4009), .B(A[247]), .C(n3703), .D(A[759]), .Y(n539) );
  AO22XL U3084 ( .A(n4023), .B(A[246]), .C(n4002), .D(A[758]), .Y(n545) );
  AO22X1 U3085 ( .A(n1419), .B(n3953), .C(n3944), .D(n3769), .Y(n1615) );
  AO22XL U3086 ( .A(n4022), .B(A[497]), .C(n3997), .D(A[1009]), .Y(n3770) );
  MUX2X1 U3087 ( .D0(n781), .D1(n782), .S(n3931), .Y(n3785) );
  MUX2XL U3088 ( .D0(A[187]), .D1(A[699]), .S(n3971), .Y(n3786) );
  OR2XL U3089 ( .A(n3991), .B(A[443]), .Y(n3787) );
  OR2XL U3090 ( .A(n3993), .B(A[353]), .Y(n3783) );
  AND2XL U3091 ( .A(n1290), .B(n3939), .Y(n3771) );
  AND2XL U3092 ( .A(n1305), .B(n3939), .Y(n3772) );
  MUX2IXL U3093 ( .D0(n1053), .D1(n1054), .S(n3926), .Y(n1709) );
  MUX2XL U3094 ( .D0(n1049), .D1(n1050), .S(n3927), .Y(n3773) );
  INVXL U3095 ( .A(A[498]), .Y(n3849) );
  INVX1 U3096 ( .A(n4012), .Y(n3971) );
  INVX1 U3097 ( .A(n4011), .Y(n3976) );
  INVX1 U3098 ( .A(n4012), .Y(n3973) );
  INVX1 U3099 ( .A(n4012), .Y(n3978) );
  INVX1 U3100 ( .A(n4009), .Y(n3983) );
  INVX1 U3101 ( .A(n4007), .Y(n3999) );
  INVX1 U3102 ( .A(n4012), .Y(n3974) );
  INVX1 U3103 ( .A(n4007), .Y(n3997) );
  INVX1 U3104 ( .A(n4007), .Y(n3998) );
  INVX1 U3105 ( .A(n4012), .Y(n3975) );
  INVX1 U3106 ( .A(n4010), .Y(n3987) );
  INVX1 U3107 ( .A(n4011), .Y(n3977) );
  INVX1 U3108 ( .A(n4009), .Y(n3985) );
  INVX1 U3109 ( .A(n4024), .Y(n3865) );
  INVX1 U3110 ( .A(n4010), .Y(n3981) );
  INVX1 U3111 ( .A(n4009), .Y(n3984) );
  INVX1 U3112 ( .A(n4018), .Y(n3866) );
  INVX1 U3113 ( .A(n4008), .Y(n3989) );
  INVX1 U3114 ( .A(n4007), .Y(n4002) );
  INVX1 U3115 ( .A(n4008), .Y(n3990) );
  INVX1 U3116 ( .A(n4009), .Y(n3993) );
  INVX1 U3117 ( .A(n4008), .Y(n3991) );
  INVX1 U3118 ( .A(n4008), .Y(n3992) );
  INVX1 U3119 ( .A(n4011), .Y(n3980) );
  INVX1 U3120 ( .A(n4009), .Y(n3986) );
  INVX1 U3121 ( .A(n4011), .Y(n3982) );
  INVX1 U3122 ( .A(n4018), .Y(n3995) );
  INVXL U3123 ( .A(n4033), .Y(n4013) );
  INVX1 U3124 ( .A(n3949), .Y(n3927) );
  INVX1 U3125 ( .A(n3949), .Y(n3926) );
  INVX1 U3126 ( .A(n3948), .Y(n3931) );
  INVX1 U3127 ( .A(n3949), .Y(n3925) );
  INVX1 U3128 ( .A(n3948), .Y(n3933) );
  INVX1 U3129 ( .A(n3948), .Y(n3934) );
  INVX1 U3130 ( .A(n3948), .Y(n3935) );
  INVX1 U3131 ( .A(n3948), .Y(n3936) );
  INVX1 U3132 ( .A(n3947), .Y(n3937) );
  INVX1 U3133 ( .A(n3949), .Y(n3938) );
  INVX1 U3134 ( .A(n3948), .Y(n3932) );
  INVX1 U3135 ( .A(n3946), .Y(n3939) );
  INVX1 U3136 ( .A(n4035), .Y(n4034) );
  INVX1 U3137 ( .A(n3947), .Y(n3940) );
  INVX1 U3138 ( .A(n3946), .Y(n3943) );
  INVX1 U3139 ( .A(n4006), .Y(n4001) );
  INVX1 U3140 ( .A(n4006), .Y(n3996) );
  INVX1 U3141 ( .A(n4006), .Y(n4000) );
  INVX1 U3142 ( .A(n4006), .Y(n4003) );
  INVX1 U3143 ( .A(n3946), .Y(n3941) );
  INVX1 U3144 ( .A(n3946), .Y(n3942) );
  INVX1 U3145 ( .A(n3968), .Y(n3950) );
  INVX1 U3146 ( .A(n3966), .Y(n3961) );
  INVX1 U3147 ( .A(n3923), .Y(n3913) );
  INVX1 U3148 ( .A(n3922), .Y(n3910) );
  INVX1 U3149 ( .A(n3908), .Y(n3905) );
  INVX1 U3150 ( .A(n3923), .Y(n3916) );
  INVX1 U3151 ( .A(n3922), .Y(n3920) );
  INVX1 U3152 ( .A(n3901), .Y(n3899) );
  INVX1 U3153 ( .A(n3923), .Y(n3918) );
  INVX1 U3154 ( .A(n3908), .Y(n3903) );
  INVX1 U3155 ( .A(n3969), .Y(n3968) );
  INVX1 U3156 ( .A(n3897), .Y(n3895) );
  INVX1 U3157 ( .A(n3897), .Y(n3896) );
  MUX2IX1 U3158 ( .D0(n31), .D1(n47), .S(n3895), .Y(n15) );
  MUX2IX1 U3159 ( .D0(n79), .D1(n111), .S(n3898), .Y(n47) );
  MUX2IX1 U3160 ( .D0(n63), .D1(n95), .S(n3900), .Y(n31) );
  MUX2IX1 U3161 ( .D0(n143), .D1(n207), .S(n3905), .Y(n79) );
  MUX2IX1 U3162 ( .D0(n48), .D1(n32), .S(n3897), .Y(n16) );
  MUX2IX1 U3163 ( .D0(n64), .D1(n96), .S(n3900), .Y(n32) );
  MUX2IX1 U3164 ( .D0(n50), .D1(n82), .S(n3900), .Y(n18) );
  NAND2X1 U3165 ( .A(SH[5]), .B(n3908), .Y(n3870) );
  INVX1 U3166 ( .A(n3901), .Y(n3898) );
  INVX1 U3167 ( .A(SH[7]), .Y(n3923) );
  INVX1 U3168 ( .A(SH[6]), .Y(n3908) );
  INVX1 U3169 ( .A(SH[7]), .Y(n3922) );
  INVX1 U3170 ( .A(SH[5]), .Y(n3901) );
  INVX1 U3171 ( .A(SH[3]), .Y(n3894) );
  INVX1 U3172 ( .A(SH[4]), .Y(n3897) );
  MUX2AXL U3173 ( .D0(n3747), .D1(n1766), .S(n3915), .Y(n176) );
  MUX2IX1 U3174 ( .D0(n312), .D1(n3759), .S(n3913), .Y(n192) );
  MUX2IX1 U3175 ( .D0(n3668), .D1(n3805), .S(n3920), .Y(n128) );
  INVX1 U3176 ( .A(n1654), .Y(n312) );
  MUX2XL U3177 ( .D0(n1359), .D1(n1360), .S(n3933), .Y(n3774) );
  NOR21XL U3178 ( .B(n3978), .A(A[964]), .Y(n746) );
  NOR21XL U3179 ( .B(n3978), .A(A[963]), .Y(n749) );
  NOR21XL U3180 ( .B(n3978), .A(A[967]), .Y(n737) );
  NOR21XL U3181 ( .B(n3866), .A(A[981]), .Y(n687) );
  MUX2IX1 U3182 ( .D0(n122), .D1(n186), .S(n3907), .Y(n58) );
  MUX2X1 U3183 ( .D0(n1696), .D1(n1824), .S(n3909), .Y(n234) );
  MUX2IX1 U3184 ( .D0(n1105), .D1(n1106), .S(n3872), .Y(n1696) );
  MUX2X1 U3185 ( .D0(n1694), .D1(n1822), .S(n3909), .Y(n232) );
  MUX2IX1 U3186 ( .D0(n1113), .D1(n1114), .S(n3925), .Y(n1694) );
  MUX2X1 U3187 ( .D0(n1693), .D1(n1821), .S(n3909), .Y(n231) );
  MUX2IX1 U3188 ( .D0(n1117), .D1(n1118), .S(n3872), .Y(n1693) );
  MUX2X1 U3189 ( .D0(n1695), .D1(n1823), .S(n3909), .Y(n233) );
  MUX2IX1 U3190 ( .D0(n1109), .D1(n1110), .S(n3872), .Y(n1695) );
  MUX2X1 U3191 ( .D0(n1600), .D1(n1728), .S(n3919), .Y(n138) );
  MUX2IXL U3192 ( .D0(n1495), .D1(n1496), .S(n3934), .Y(n1600) );
  MUX2X1 U3193 ( .D0(n1597), .D1(n1725), .S(n3919), .Y(n135) );
  MUX2IX1 U3194 ( .D0(n973), .D1(n974), .S(n3928), .Y(n1725) );
  MUX2X1 U3195 ( .D0(n1598), .D1(n1726), .S(n3919), .Y(n136) );
  MUX2IX1 U3196 ( .D0(n1503), .D1(n1504), .S(n3937), .Y(n1598) );
  MUX2IX1 U3197 ( .D0(n953), .D1(n954), .S(n3929), .Y(n1730) );
  MUX2IX1 U3198 ( .D0(n3675), .D1(n3704), .S(n3919), .Y(n133) );
  MUX2IX1 U3199 ( .D0(n3684), .D1(n3650), .S(n3919), .Y(n132) );
  MUX2IX1 U3200 ( .D0(n1327), .D1(n1328), .S(n3930), .Y(n1634) );
  NOR21XL U3201 ( .B(n3998), .A(A[971]), .Y(n722) );
  MUX2X1 U3202 ( .D0(n1687), .D1(n1815), .S(n3910), .Y(n225) );
  MUX2IXL U3203 ( .D0(n1141), .D1(n1142), .S(n3924), .Y(n1687) );
  MUX2X1 U3204 ( .D0(n1688), .D1(n1816), .S(n3910), .Y(n226) );
  MUX2IXL U3205 ( .D0(n1137), .D1(n1138), .S(n3924), .Y(n1688) );
  MUX2X1 U3206 ( .D0(n1642), .D1(n1770), .S(n3915), .Y(n180) );
  MUX2X1 U3207 ( .D0(n1583), .D1(n1711), .S(n3920), .Y(n121) );
  MUX2IX1 U3208 ( .D0(n1351), .D1(n1352), .S(n3932), .Y(n1628) );
  MUX2X1 U3209 ( .D0(n1631), .D1(n1759), .S(n3916), .Y(n169) );
  MUX2X1 U3210 ( .D0(n1632), .D1(n1760), .S(n3916), .Y(n170) );
  MUX2IX1 U3211 ( .D0(n3705), .D1(n3692), .S(n3920), .Y(n125) );
  MUX2IX1 U3212 ( .D0(n3676), .D1(n3858), .S(n3916), .Y(n165) );
  MUX2X1 U3213 ( .D0(n1624), .D1(n1752), .S(n3916), .Y(n162) );
  MUX2IXL U3214 ( .D0(n1367), .D1(n1368), .S(n3933), .Y(n1624) );
  MUX2X1 U3215 ( .D0(n1630), .D1(n1758), .S(n3916), .Y(n168) );
  MUX2X1 U3216 ( .D0(n1629), .D1(n1757), .S(n3916), .Y(n167) );
  MUX2IX1 U3217 ( .D0(n127), .D1(n191), .S(n3906), .Y(n63) );
  MUX2IX1 U3218 ( .D0(n3750), .D1(n3811), .S(n3920), .Y(n127) );
  MUX2X1 U3219 ( .D0(n1592), .D1(n1720), .S(n3920), .Y(n130) );
  MUX2X1 U3220 ( .D0(n1650), .D1(n1778), .S(n3914), .Y(n188) );
  MUX2IXL U3221 ( .D0(n721), .D1(n722), .S(n3933), .Y(n1778) );
  MUX2IX1 U3222 ( .D0(n146), .D1(n210), .S(n3905), .Y(n82) );
  MUX2IX1 U3223 ( .D0(n3818), .D1(n3808), .S(n3918), .Y(n146) );
  MUX2X1 U3224 ( .D0(n1643), .D1(n1771), .S(n3914), .Y(n181) );
  MUX2X1 U3225 ( .D0(n1646), .D1(n1774), .S(n3914), .Y(n184) );
  NAND2X1 U3226 ( .A(n1287), .B(n3938), .Y(n1646) );
  MUX2X1 U3227 ( .D0(n1679), .D1(n1807), .S(n3911), .Y(n217) );
  MUX2IX1 U3228 ( .D0(n57), .D1(n89), .S(n3899), .Y(n25) );
  MUX2IX1 U3229 ( .D0(n153), .D1(n217), .S(n3904), .Y(n89) );
  MUX2IX1 U3230 ( .D0(n3758), .D1(n3838), .S(n3911), .Y(n220) );
  MUX2IX1 U3231 ( .D0(n56), .D1(n88), .S(n3899), .Y(n24) );
  MUX2IX1 U3232 ( .D0(n120), .D1(n184), .S(SH[6]), .Y(n56) );
  MUX2IX1 U3233 ( .D0(n55), .D1(n87), .S(n3899), .Y(n23) );
  MUX2IX1 U3234 ( .D0(n119), .D1(n183), .S(n3907), .Y(n55) );
  MUX2IX1 U3235 ( .D0(n151), .D1(n215), .S(n3904), .Y(n87) );
  MUX2X1 U3236 ( .D0(n1615), .D1(n1743), .S(n3917), .Y(n153) );
  MUX2X2 U3237 ( .D0(n1618), .D1(n1746), .S(n3917), .Y(n156) );
  MUX2X1 U3238 ( .D0(n1613), .D1(n1741), .S(n3917), .Y(n151) );
  MUX2X1 U3239 ( .D0(n1605), .D1(n1733), .S(n3918), .Y(n143) );
  MUX2IX1 U3240 ( .D0(n175), .D1(n239), .S(n3902), .Y(n111) );
  MUX2IX1 U3241 ( .D0(n3751), .D1(n3691), .S(n3909), .Y(n239) );
  MUX2IX1 U3242 ( .D0(n313), .D1(n3744), .S(n3913), .Y(n193) );
  MUX2IX1 U3243 ( .D0(n316), .D1(n3743), .S(n3913), .Y(n196) );
  MUX2IX1 U3244 ( .D0(n317), .D1(n3737), .S(n3913), .Y(n197) );
  MUX2IX1 U3245 ( .D0(n314), .D1(n3740), .S(n3913), .Y(n194) );
  MUX2IX1 U3246 ( .D0(n3752), .D1(n3832), .S(n3912), .Y(n204) );
  MUX2IX1 U3247 ( .D0(n3746), .D1(n3827), .S(n3912), .Y(n205) );
  MUX2IX1 U3248 ( .D0(n72), .D1(n104), .S(n3898), .Y(n40) );
  MUX2IX1 U3249 ( .D0(n136), .D1(n200), .S(n3906), .Y(n72) );
  MUX2IX1 U3250 ( .D0(n168), .D1(n232), .S(n3902), .Y(n104) );
  MUX2IX1 U3251 ( .D0(n320), .D1(n3738), .S(n3913), .Y(n200) );
  MUX2IX1 U3252 ( .D0(n71), .D1(n103), .S(n3898), .Y(n39) );
  MUX2IX1 U3253 ( .D0(n135), .D1(n199), .S(n3906), .Y(n71) );
  MUX2IX1 U3254 ( .D0(n167), .D1(n231), .S(n3902), .Y(n103) );
  MUX2IX1 U3255 ( .D0(n319), .D1(n3741), .S(n3913), .Y(n199) );
  MUX2IX1 U3256 ( .D0(n159), .D1(n223), .S(n3903), .Y(n95) );
  MUX2IX1 U3257 ( .D0(n114), .D1(n178), .S(n3907), .Y(n50) );
  MUX2X1 U3258 ( .D0(n1543), .D1(n1544), .S(n3938), .Y(n3776) );
  MUX2IX1 U3259 ( .D0(n3726), .D1(n3693), .S(n3917), .Y(n157) );
  MUX2IX1 U3260 ( .D0(n3736), .D1(n3690), .S(n3910), .Y(n228) );
  MUX2IX1 U3261 ( .D0(n3677), .D1(n3707), .S(n3910), .Y(n221) );
  MUX2IX1 U3262 ( .D0(n144), .D1(n208), .S(n3905), .Y(n80) );
  MUX2IX1 U3263 ( .D0(n328), .D1(n3798), .S(n3912), .Y(n208) );
  MUX2IX1 U3264 ( .D0(n3765), .D1(n3669), .S(n3918), .Y(n144) );
  INVX1 U3265 ( .A(n1670), .Y(n328) );
  MUX2IX1 U3266 ( .D0(n310), .D1(n3855), .S(n3914), .Y(n190) );
  INVX1 U3267 ( .A(n1652), .Y(n310) );
  MUX2IX1 U3268 ( .D0(n75), .D1(n107), .S(n3898), .Y(n43) );
  MUX2IX1 U3269 ( .D0(n171), .D1(n235), .S(n3902), .Y(n107) );
  MUX2IX1 U3270 ( .D0(n3879), .D1(n3785), .S(n3915), .Y(n171) );
  MUX2IX1 U3271 ( .D0(n74), .D1(n106), .S(n3898), .Y(n42) );
  MUX2IX1 U3272 ( .D0(n138), .D1(n202), .S(n3905), .Y(n74) );
  MUX2IX1 U3273 ( .D0(n170), .D1(n234), .S(n3902), .Y(n106) );
  MUX2IX1 U3274 ( .D0(n3753), .D1(n3667), .S(n3912), .Y(n202) );
  NOR21XL U3275 ( .B(n3987), .A(A[978]), .Y(n696) );
  AND2X1 U3276 ( .A(n3784), .B(n3921), .Y(n3779) );
  MUX2X2 U3277 ( .D0(n3653), .D1(n3699), .S(n3914), .Y(n3780) );
  NOR21XL U3278 ( .B(n3978), .A(A[966]), .Y(n740) );
  NOR21XL U3279 ( .B(n3977), .A(A[961]), .Y(n755) );
  NOR21XL U3280 ( .B(n4031), .A(A[980]), .Y(n690) );
  NOR21XL U3281 ( .B(n3866), .A(A[977]), .Y(n699) );
  NOR21XL U3282 ( .B(n3981), .A(A[979]), .Y(n693) );
  NOR21XL U3283 ( .B(n3981), .A(A[976]), .Y(n702) );
  NOR21XL U3284 ( .B(n4031), .A(A[982]), .Y(n684) );
  NOR21XL U3285 ( .B(n3982), .A(A[983]), .Y(n681) );
  MUX2IX1 U3286 ( .D0(n8), .D1(n16), .S(SH[3]), .Y(B[7]) );
  MUX2IX1 U3287 ( .D0(n24), .D1(n40), .S(n3895), .Y(n8) );
  AOI22XL U3288 ( .A(n4026), .B(A[160]), .C(n3701), .D(A[672]), .Y(n3781) );
  AOI22XL U3289 ( .A(n4013), .B(A[416]), .C(n3701), .D(A[928]), .Y(n3782) );
  NOR21XL U3290 ( .B(n3980), .A(A[615]), .Y(n1177) );
  NOR21XL U3291 ( .B(n3982), .A(A[616]), .Y(n1173) );
  NOR21XL U3292 ( .B(n3981), .A(A[659]), .Y(n985) );
  MUX2X2 U3293 ( .D0(n1057), .D1(n1058), .S(n3926), .Y(n3784) );
  MUX2IX1 U3294 ( .D0(A[188]), .D1(A[700]), .S(n3971), .Y(n773) );
  NOR21XL U3295 ( .B(n3986), .A(A[608]), .Y(n1205) );
  OR2X1 U3296 ( .A(n3987), .B(A[351]), .Y(n3789) );
  NOR21XL U3297 ( .B(n3974), .A(A[713]), .Y(n729) );
  NOR21XL U3298 ( .B(n3979), .A(A[969]), .Y(n730) );
  MUX2IX1 U3299 ( .D0(A[284]), .D1(A[796]), .S(n3976), .Y(n1484) );
  NOR21XL U3300 ( .B(n3985), .A(A[542]), .Y(n1475) );
  MUX2IXL U3301 ( .D0(A[286]), .D1(A[798]), .S(n3976), .Y(n1476) );
  MUX2IX1 U3302 ( .D0(n1315), .D1(n1316), .S(n3930), .Y(n1637) );
  NOR21XL U3303 ( .B(n3983), .A(A[574]), .Y(n1315) );
  MUX2IXL U3304 ( .D0(n1149), .D1(n4024), .S(n3924), .Y(n1685) );
  MUX2IX1 U3305 ( .D0(A[485]), .D1(A[997]), .S(n3975), .Y(n626) );
  OR2XL U3306 ( .A(n3991), .B(A[230]), .Y(n3790) );
  MUX2XL U3307 ( .D0(A[486]), .D1(A[998]), .S(n3975), .Y(n3791) );
  MUX2IX1 U3308 ( .D0(A[484]), .D1(A[996]), .S(n3975), .Y(n630) );
  MUX2IXL U3309 ( .D0(A[483]), .D1(A[995]), .S(n3975), .Y(n634) );
  NOR21XL U3310 ( .B(n3980), .A(A[665]), .Y(n961) );
  NOR21XL U3311 ( .B(n3980), .A(A[664]), .Y(n965) );
  MUX2IX1 U3312 ( .D0(n969), .D1(n970), .S(n3928), .Y(n1726) );
  NOR21XL U3313 ( .B(n3980), .A(A[663]), .Y(n969) );
  NOR21XL U3314 ( .B(n4028), .A(A[533]), .Y(n1511) );
  NOR21XL U3315 ( .B(n4033), .A(A[531]), .Y(n1519) );
  MUX2IXL U3316 ( .D0(A[275]), .D1(A[787]), .S(n3975), .Y(n1520) );
  NOR21XL U3317 ( .B(n3984), .A(A[528]), .Y(n1531) );
  NOR21XL U3318 ( .B(n3979), .A(A[568]), .Y(n1339) );
  MUX2IXL U3319 ( .D0(A[312]), .D1(A[824]), .S(n3971), .Y(n1340) );
  NOR21XL U3320 ( .B(n3985), .A(A[562]), .Y(n1363) );
  NOR21XL U3321 ( .B(n3865), .A(A[587]), .Y(n1275) );
  NOR21XL U3322 ( .B(n3983), .A(A[597]), .Y(n1247) );
  NOR21XL U3323 ( .B(n3982), .A(A[836]), .Y(n1296) );
  NOR21XL U3324 ( .B(n3982), .A(A[835]), .Y(n1299) );
  NOR21XL U3325 ( .B(n3985), .A(A[832]), .Y(n1308) );
  NOR21XL U3326 ( .B(n3866), .A(A[839]), .Y(n1287) );
  MUX2IX1 U3327 ( .D0(A[189]), .D1(A[701]), .S(n3971), .Y(n769) );
  AND2XL U3328 ( .A(n4026), .B(n3862), .Y(n637) );
  INVX1 U3329 ( .A(A[226]), .Y(n3862) );
  MUX2IX1 U3330 ( .D0(A[412]), .D1(A[924]), .S(n3970), .Y(n950) );
  MUX2IX1 U3331 ( .D0(A[316]), .D1(A[828]), .S(n3988), .Y(n1324) );
  MUX2XL U3332 ( .D0(A[185]), .D1(A[697]), .S(n3971), .Y(n3792) );
  OR2XL U3333 ( .A(n3990), .B(A[441]), .Y(n3793) );
  MUX2IX1 U3334 ( .D0(A[309]), .D1(A[821]), .S(n3971), .Y(n1352) );
  MUX2IXL U3335 ( .D0(A[313]), .D1(A[825]), .S(n3971), .Y(n1336) );
  MUX2IXL U3336 ( .D0(A[311]), .D1(A[823]), .S(n3971), .Y(n1344) );
  MUX2IXL U3337 ( .D0(A[280]), .D1(A[792]), .S(n3700), .Y(n1500) );
  MUX2IXL U3338 ( .D0(A[478]), .D1(A[990]), .S(n3976), .Y(n654) );
  NOR21XL U3339 ( .B(n3985), .A(A[563]), .Y(n1359) );
  NOR21XL U3340 ( .B(n3985), .A(A[560]), .Y(n1371) );
  MUX2IXL U3341 ( .D0(A[267]), .D1(A[779]), .S(n3973), .Y(n1552) );
  MUX2IXL U3342 ( .D0(A[265]), .D1(A[777]), .S(n3973), .Y(n1560) );
  MUX2IXL U3343 ( .D0(A[264]), .D1(A[776]), .S(n3973), .Y(n1564) );
  MUX2IXL U3344 ( .D0(A[310]), .D1(A[822]), .S(n4031), .Y(n1348) );
  MUX2IX1 U3345 ( .D0(A[492]), .D1(A[1004]), .S(n3974), .Y(n598) );
  MUX2IXL U3346 ( .D0(A[273]), .D1(A[785]), .S(n3974), .Y(n1528) );
  MUX2IXL U3347 ( .D0(A[488]), .D1(A[1000]), .S(n3974), .Y(n614) );
  NOR21XL U3348 ( .B(n3985), .A(A[561]), .Y(n1367) );
  NOR21XL U3349 ( .B(n3979), .A(A[566]), .Y(n1347) );
  NOR21XL U3350 ( .B(n3866), .A(A[624]), .Y(n1141) );
  NOR21XL U3351 ( .B(n3865), .A(A[627]), .Y(n1129) );
  NOR21XL U3352 ( .B(n4029), .A(A[625]), .Y(n1137) );
  NOR21XL U3353 ( .B(n3700), .A(A[669]), .Y(n945) );
  NOR21XL U3354 ( .B(n4029), .A(A[668]), .Y(n949) );
  NOR21XL U3355 ( .B(n3986), .A(A[715]), .Y(n721) );
  NOR21XL U3356 ( .B(n3984), .A(A[667]), .Y(n953) );
  NOR21XL U3357 ( .B(n3978), .A(A[670]), .Y(n941) );
  NOR21XL U3358 ( .B(n3988), .A(A[569]), .Y(n1335) );
  NOR21XL U3359 ( .B(n4033), .A(A[613]), .Y(n1185) );
  NOR21XL U3360 ( .B(n3998), .A(A[612]), .Y(n1189) );
  NOR21XL U3361 ( .B(n4028), .A(A[523]), .Y(n1551) );
  NOR21XL U3362 ( .B(n3981), .A(A[656]), .Y(n997) );
  NOR21XL U3363 ( .B(n4032), .A(A[614]), .Y(n1181) );
  NOR21XL U3364 ( .B(n4029), .A(A[525]), .Y(n1543) );
  NOR21XL U3365 ( .B(n3986), .A(A[537]), .Y(n1495) );
  NOR21XL U3366 ( .B(n4030), .A(A[611]), .Y(n1193) );
  NOR21XL U3367 ( .B(n3866), .A(A[536]), .Y(n1499) );
  NOR21XL U3368 ( .B(n3986), .A(A[535]), .Y(n1503) );
  NOR21XL U3369 ( .B(n4030), .A(A[975]), .Y(n706) );
  NOR21XL U3370 ( .B(n4030), .A(A[719]), .Y(n705) );
  NOR21XL U3371 ( .B(n3865), .A(A[521]), .Y(n1559) );
  NOR21XL U3372 ( .B(n4031), .A(A[529]), .Y(n1527) );
  MUX2IX1 U3373 ( .D0(n993), .D1(n994), .S(n3928), .Y(n1720) );
  NOR21XL U3374 ( .B(n3865), .A(A[657]), .Y(n993) );
  NOR21XL U3375 ( .B(n3984), .A(A[571]), .Y(n1327) );
  NOR21XL U3376 ( .B(n3982), .A(A[520]), .Y(n1563) );
  NOR21XL U3377 ( .B(n3865), .A(A[630]), .Y(n1117) );
  NOR21XL U3378 ( .B(n3980), .A(A[662]), .Y(n973) );
  NOR21XL U3379 ( .B(n4030), .A(A[623]), .Y(n1145) );
  NOR21XL U3380 ( .B(n3981), .A(A[631]), .Y(n1113) );
  NOR21XL U3381 ( .B(n3989), .A(A[567]), .Y(n1343) );
  MUX2IXL U3382 ( .D0(A[279]), .D1(A[791]), .S(n3975), .Y(n1504) );
  MUX2IXL U3383 ( .D0(A[487]), .D1(A[999]), .S(n3975), .Y(n618) );
  MUX2X1 U3384 ( .D0(A[481]), .D1(A[993]), .S(n3977), .Y(n3797) );
  MUX2X1 U3385 ( .D0(A[479]), .D1(A[991]), .S(n3977), .Y(n3800) );
  MUX2IXL U3386 ( .D0(A[489]), .D1(A[1001]), .S(n3974), .Y(n610) );
  MUX2IXL U3387 ( .D0(A[495]), .D1(A[1007]), .S(n3973), .Y(n586) );
  MUX2IX1 U3388 ( .D0(n3859), .D1(n3694), .S(n3918), .Y(n148) );
  NOR21XL U3389 ( .B(n4029), .A(A[585]), .Y(n1281) );
  NOR21XL U3390 ( .B(n4029), .A(A[589]), .Y(n1269) );
  NOR21XL U3391 ( .B(n3977), .A(A[960]), .Y(n758) );
  NOR21XL U3392 ( .B(n4031), .A(A[530]), .Y(n1523) );
  NOR21XL U3393 ( .B(n3701), .A(A[714]), .Y(n725) );
  NOR21XL U3394 ( .B(n3700), .A(A[970]), .Y(n726) );
  NOR21XL U3395 ( .B(n3987), .A(A[658]), .Y(n989) );
  OAI22AX1 U3396 ( .D(n3954), .C(n3803), .A(n3804), .B(n3802), .Y(n1820) );
  AOI22XL U3397 ( .A(n3853), .B(A[245]), .C(n4002), .D(A[757]), .Y(n3803) );
  AOI22XL U3398 ( .A(n4022), .B(A[501]), .C(n3999), .D(A[1013]), .Y(n3804) );
  AOI22BX1 U3399 ( .B(n3806), .A(n3941), .D(n3807), .C(n3958), .Y(n3805) );
  AOI22XL U3400 ( .A(n4017), .B(A[399]), .C(n4005), .D(A[911]), .Y(n3806) );
  AOI22X1 U3401 ( .A(n4010), .B(A[143]), .C(n4005), .D(A[655]), .Y(n3807) );
  NOR21XL U3402 ( .B(n3985), .A(A[564]), .Y(n1355) );
  MUX2IXL U3403 ( .D0(A[474]), .D1(A[986]), .S(n4028), .Y(n670) );
  MUX2IXL U3404 ( .D0(A[786]), .D1(A[274]), .S(n3853), .Y(n1524) );
  AOI22XL U3405 ( .A(n4026), .B(A[417]), .C(n3998), .D(A[929]), .Y(n3809) );
  AOI22XL U3406 ( .A(n4024), .B(A[161]), .C(n3998), .D(A[673]), .Y(n3810) );
  AOI22XL U3407 ( .A(n4013), .B(A[398]), .C(n4005), .D(A[910]), .Y(n3812) );
  AOI22XL U3408 ( .A(n4026), .B(A[142]), .C(n4005), .D(A[654]), .Y(n3813) );
  AO22X1 U3409 ( .A(n808), .B(n3942), .C(n807), .D(n3953), .Y(n1756) );
  OAI22AXL U3410 ( .D(n3962), .C(n3815), .A(n3816), .B(n3814), .Y(n1815) );
  AOI22XL U3411 ( .A(n4017), .B(A[240]), .C(n3700), .D(A[752]), .Y(n3815) );
  AOI22XL U3412 ( .A(n4017), .B(A[496]), .C(n4000), .D(A[1008]), .Y(n3816) );
  MUX2IXL U3413 ( .D0(A[266]), .D1(A[778]), .S(n4030), .Y(n1556) );
  AOI22XL U3414 ( .A(n4013), .B(A[289]), .C(n3998), .D(A[801]), .Y(n3819) );
  AOI22XL U3415 ( .A(n4008), .B(A[33]), .C(n4002), .D(A[545]), .Y(n3820) );
  AOI22XL U3416 ( .A(n4013), .B(A[302]), .C(n4033), .D(A[814]), .Y(n3822) );
  AOI22XL U3417 ( .A(n3853), .B(A[46]), .C(n3991), .D(A[558]), .Y(n3823) );
  AOI22BXL U3418 ( .B(n3825), .A(n3943), .D(n3826), .C(n3711), .Y(n3824) );
  AOI22XL U3419 ( .A(n4018), .B(A[430]), .C(n4000), .D(A[942]), .Y(n3825) );
  AOI22XL U3420 ( .A(n4018), .B(A[174]), .C(n4000), .D(A[686]), .Y(n3826) );
  AO22X1 U3421 ( .A(n4014), .B(A[45]), .C(n3700), .D(A[557]), .Y(n1389) );
  NOR21X1 U3422 ( .B(n3986), .A(A[604]), .Y(n1221) );
  MUX2IX1 U3423 ( .D0(n3828), .D1(n3829), .S(n3934), .Y(n3827) );
  INVX1 U3424 ( .A(n1647), .Y(n305) );
  NOR21XL U3425 ( .B(n4031), .A(A[584]), .Y(n1284) );
  INVX1 U3426 ( .A(n1658), .Y(n316) );
  NOR21XL U3427 ( .B(n3983), .A(A[595]), .Y(n1253) );
  INVX1 U3428 ( .A(n1659), .Y(n317) );
  NOR21XL U3429 ( .B(n3983), .A(A[596]), .Y(n1250) );
  INVX1 U3430 ( .A(n1661), .Y(n319) );
  NOR21XL U3431 ( .B(n3983), .A(A[598]), .Y(n1244) );
  INVX1 U3432 ( .A(n1662), .Y(n320) );
  NOR21XL U3433 ( .B(n3983), .A(A[599]), .Y(n1241) );
  INVX1 U3434 ( .A(n1656), .Y(n314) );
  NOR21XL U3435 ( .B(n3866), .A(A[593]), .Y(n1259) );
  INVX1 U3436 ( .A(n1655), .Y(n313) );
  NOR21XL U3437 ( .B(n3865), .A(A[592]), .Y(n1262) );
  NOR21XL U3438 ( .B(n3985), .A(A[603]), .Y(n1225) );
  NOR21XL U3439 ( .B(n3983), .A(A[600]), .Y(n1237) );
  NOR21XL U3440 ( .B(n3983), .A(A[601]), .Y(n1233) );
  MUX2IX1 U3441 ( .D0(A[319]), .D1(A[831]), .S(n4029), .Y(n1312) );
  NOR21XL U3442 ( .B(n3978), .A(A[671]), .Y(n937) );
  NOR21XL U3443 ( .B(n3982), .A(A[617]), .Y(n1169) );
  MUX2IX1 U3444 ( .D0(n3833), .D1(n3834), .S(n3931), .Y(n3832) );
  OR2XL U3445 ( .A(n3990), .B(A[219]), .Y(n3833) );
  MUX2XL U3446 ( .D0(A[475]), .D1(A[987]), .S(n3976), .Y(n3834) );
  MUX2IXL U3447 ( .D0(A[287]), .D1(A[799]), .S(n3976), .Y(n1472) );
  NOR21XL U3448 ( .B(n3986), .A(A[543]), .Y(n1471) );
  NOR21XL U3449 ( .B(n4031), .A(A[619]), .Y(n1161) );
  MUX2IXL U3450 ( .D0(A[271]), .D1(A[783]), .S(n3974), .Y(n1536) );
  NOR21XL U3451 ( .B(n3986), .A(A[527]), .Y(n1535) );
  MUX2IX1 U3452 ( .D0(n3839), .D1(n3840), .S(n3936), .Y(n3838) );
  OR2XL U3453 ( .A(n3991), .B(A[235]), .Y(n3839) );
  MUX2XL U3454 ( .D0(A[491]), .D1(A[1003]), .S(n3974), .Y(n3840) );
  MUX2IXL U3455 ( .D0(A[494]), .D1(A[1006]), .S(n3973), .Y(n590) );
  NOR21XL U3456 ( .B(n4030), .A(A[526]), .Y(n1539) );
  MUX2IXL U3457 ( .D0(A[270]), .D1(A[782]), .S(n3974), .Y(n1540) );
  NOR21XL U3458 ( .B(n3978), .A(A[968]), .Y(n734) );
  NOR21XL U3459 ( .B(n3978), .A(A[712]), .Y(n733) );
  NOR21XL U3460 ( .B(n4031), .A(A[718]), .Y(n709) );
  NOR21XL U3461 ( .B(n3981), .A(A[974]), .Y(n710) );
  INVX1 U3462 ( .A(n1651), .Y(n309) );
  NOR21XL U3463 ( .B(n3866), .A(A[588]), .Y(n1272) );
  AOI22XL U3464 ( .A(n4008), .B(A[511]), .C(n3701), .D(A[1023]), .Y(n3843) );
  AOI22XL U3465 ( .A(n4012), .B(A[255]), .C(n3996), .D(A[767]), .Y(n3844) );
  NOR21XL U3466 ( .B(n3982), .A(A[833]), .Y(n1305) );
  NOR21XL U3467 ( .B(n4030), .A(A[838]), .Y(n1290) );
  MUX2IX1 U3468 ( .D0(n7), .D1(n15), .S(SH[3]), .Y(B[6]) );
  MUX2IX1 U3469 ( .D0(n23), .D1(n39), .S(n3895), .Y(n7) );
  INVX1 U3470 ( .A(A[34]), .Y(n3850) );
  INVX1 U3471 ( .A(A[397]), .Y(n3863) );
  INVX1 U3472 ( .A(A[909]), .Y(n3864) );
  INVX1 U3473 ( .A(A[186]), .Y(n3888) );
  INVX1 U3474 ( .A(A[282]), .Y(n3892) );
  INVX1 U3475 ( .A(A[826]), .Y(n3848) );
  INVX1 U3476 ( .A(A[314]), .Y(n3847) );
  INVX1 U3477 ( .A(A[538]), .Y(n3885) );
  NOR21XL U3478 ( .B(n3979), .A(A[572]), .Y(n1323) );
  NOR21XL U3479 ( .B(n3979), .A(A[573]), .Y(n1319) );
  INVX1 U3480 ( .A(n4037), .Y(n4029) );
  INVXL U3481 ( .A(SH[9]), .Y(n4036) );
  EORX1 U3482 ( .A(n1034), .B(n3941), .C(n3846), .D(n3967), .Y(n3889) );
  AOI22X1 U3483 ( .A(n4020), .B(A[138]), .C(n3987), .D(A[650]), .Y(n3846) );
  MUX2IXL U3484 ( .D0(n176), .D1(n240), .S(n3902), .Y(n112) );
  MUX2IX1 U3485 ( .D0(n3841), .D1(n3842), .S(n3909), .Y(n240) );
  MUX2IX1 U3486 ( .D0(n80), .D1(n112), .S(n3898), .Y(n48) );
  NOR2XL U3487 ( .A(n3979), .B(A[349]), .Y(n1218) );
  MUX2X1 U3488 ( .D0(n3848), .D1(n3847), .S(n4015), .Y(n1332) );
  MUX2IX1 U3489 ( .D0(A[120]), .D1(A[632]), .S(n4029), .Y(n1109) );
  MUX2IX1 U3490 ( .D0(A[121]), .D1(A[633]), .S(n4029), .Y(n1105) );
  MUX2IX1 U3491 ( .D0(A[122]), .D1(A[634]), .S(n3703), .Y(n1101) );
  MUX2IX1 U3492 ( .D0(A[123]), .D1(A[635]), .S(n4028), .Y(n1097) );
  MUX2IX1 U3493 ( .D0(A[124]), .D1(A[636]), .S(n4027), .Y(n1093) );
  MUX2IX1 U3494 ( .D0(A[125]), .D1(A[637]), .S(n4032), .Y(n1089) );
  MUX2IX1 U3495 ( .D0(A[126]), .D1(A[638]), .S(n4033), .Y(n1085) );
  MUX2IX1 U3496 ( .D0(A[127]), .D1(A[639]), .S(n4033), .Y(n1081) );
  MUX2IX1 U3497 ( .D0(A[400]), .D1(A[912]), .S(n3990), .Y(n998) );
  MUX2IX1 U3498 ( .D0(A[401]), .D1(A[913]), .S(n4032), .Y(n994) );
  OAI22AXL U3499 ( .D(A[1010]), .C(n4018), .A(n4002), .B(n3849), .Y(n570) );
  INVX1 U3500 ( .A(n3884), .Y(n1491) );
  EORX1 U3501 ( .A(n3872), .B(n522), .C(n3851), .D(n3967), .Y(n3881) );
  AOI22X1 U3502 ( .A(n4016), .B(A[250]), .C(n3998), .D(A[762]), .Y(n3851) );
  INVXL U3503 ( .A(n4028), .Y(n4023) );
  INVX2 U3504 ( .A(n4032), .Y(n4016) );
  INVXL U3505 ( .A(n4008), .Y(n3988) );
  INVX1 U3506 ( .A(n4037), .Y(n4030) );
  NOR21XL U3507 ( .B(n4024), .A(A[218]), .Y(n669) );
  OA22X1 U3508 ( .A(n3857), .B(n3965), .C(n3876), .D(n3952), .Y(n3887) );
  MUX2IX1 U3509 ( .D0(A[788]), .D1(A[276]), .S(n4017), .Y(n1516) );
  AOI22X1 U3510 ( .A(n814), .B(n3943), .C(n813), .D(n3962), .Y(n3858) );
  AO22XL U3511 ( .A(n4022), .B(A[249]), .C(n3998), .D(A[761]), .Y(n527) );
  AOI22XL U3512 ( .A(n4012), .B(A[35]), .C(n3997), .D(A[547]), .Y(n3860) );
  EORX1 U3513 ( .A(n1456), .B(n3965), .C(n3861), .D(n3872), .Y(n3867) );
  MUX2IX1 U3514 ( .D0(n3867), .D1(n3871), .S(n3918), .Y(n147) );
  MUX2IXL U3515 ( .D0(A[922]), .D1(A[410]), .S(n4016), .Y(n958) );
  MUX2IX1 U3516 ( .D0(A[818]), .D1(A[306]), .S(n4019), .Y(n1364) );
  MUX2IXL U3517 ( .D0(A[914]), .D1(A[402]), .S(n4016), .Y(n990) );
  INVX1 U3518 ( .A(n1820), .Y(n478) );
  INVXL U3519 ( .A(n4011), .Y(n3979) );
  MUX2IX4 U3520 ( .D0(n12), .D1(n4), .S(n3894), .Y(B[3]) );
  MUX2IX1 U3521 ( .D0(n128), .D1(n192), .S(n3906), .Y(n64) );
  AOI22X1 U3522 ( .A(n570), .B(n3944), .C(n569), .D(n3962), .Y(n3869) );
  MUX2IX1 U3523 ( .D0(n3890), .D1(n3655), .S(n3922), .Y(n155) );
  INVX1 U3524 ( .A(n4028), .Y(n4022) );
  MUX2IXL U3525 ( .D0(A[482]), .D1(A[994]), .S(n4028), .Y(n638) );
  MUX2IX1 U3526 ( .D0(n3678), .D1(n3886), .S(n3911), .Y(n219) );
  MUX2IX1 U3527 ( .D0(n155), .D1(n219), .S(n3904), .Y(n91) );
  MUX2IX1 U3528 ( .D0(n78), .D1(n110), .S(n3898), .Y(n46) );
  AOI22X1 U3529 ( .A(n922), .B(n3940), .C(n921), .D(n3964), .Y(n3871) );
  INVX1 U3530 ( .A(n4037), .Y(n4031) );
  INVX1 U3531 ( .A(n4036), .Y(n4027) );
  INVXL U3532 ( .A(n3969), .Y(n3872) );
  MUX2IX1 U3533 ( .D0(A[490]), .D1(A[1002]), .S(n4030), .Y(n3873) );
  MUX2IX1 U3534 ( .D0(n2), .D1(n10), .S(SH[3]), .Y(B[1]) );
  MUX2IX1 U3535 ( .D0(n26), .D1(n42), .S(n3895), .Y(n10) );
  AOI22X1 U3536 ( .A(n4018), .B(A[434]), .C(n4001), .D(A[946]), .Y(n3876) );
  INVX1 U3537 ( .A(n4037), .Y(n4028) );
  MUX2IX1 U3538 ( .D0(n58), .D1(n90), .S(n3899), .Y(n26) );
  MUX2IX1 U3539 ( .D0(n154), .D1(n218), .S(n3904), .Y(n90) );
  EORX1 U3540 ( .A(n874), .B(n3941), .C(n3877), .D(n3965), .Y(n3890) );
  AOI22X1 U3541 ( .A(n4022), .B(A[170]), .C(n3997), .D(A[682]), .Y(n3877) );
  MUX2IX1 U3542 ( .D0(n94), .D1(n62), .S(n3901), .Y(n30) );
  MUX2IX1 U3543 ( .D0(n30), .D1(n46), .S(n3895), .Y(n14) );
  AND2X2 U3544 ( .A(n3711), .B(n1278), .Y(n3880) );
  MUX2IX1 U3545 ( .D0(n126), .D1(n190), .S(n3904), .Y(n62) );
  MUX2IX1 U3546 ( .D0(n3776), .D1(n3689), .S(n3920), .Y(n126) );
  MUX2IX4 U3547 ( .D0(n67), .D1(n99), .S(n3900), .Y(n35) );
  NAND21XL U3548 ( .B(n4014), .A(n3885), .Y(n3884) );
  MUX2AXL U3549 ( .D0(A[698]), .D1(n3888), .S(n4007), .Y(n781) );
  MUX2IX1 U3550 ( .D0(n6), .D1(n14), .S(SH[3]), .Y(B[5]) );
  MUX2AXL U3551 ( .D0(A[794]), .D1(n3892), .S(n4020), .Y(n1492) );
  INVX1 U3552 ( .A(n4036), .Y(n4032) );
  MUX2IX1 U3553 ( .D0(n3774), .D1(n3696), .S(n3916), .Y(n164) );
  MUX2IX1 U3554 ( .D0(n158), .D1(n222), .S(n3903), .Y(n94) );
  NOR21XL U3555 ( .B(n3997), .A(A[666]), .Y(n957) );
  MUX2IX1 U3556 ( .D0(n59), .D1(n91), .S(n3899), .Y(n27) );
  MUX2IX1 U3557 ( .D0(n3654), .D1(n3695), .S(n3917), .Y(n158) );
  MUX2IX1 U3558 ( .D0(A[308]), .D1(A[820]), .S(n3972), .Y(n1356) );
  AO22XL U3559 ( .A(n4020), .B(A[140]), .C(n4027), .D(A[652]), .Y(n1021) );
  MUX2IX1 U3560 ( .D0(n27), .D1(n43), .S(n3895), .Y(n11) );
endmodule


module regbank_a0_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module regbank_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regbank_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regbank_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_50 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10855;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_50 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10855), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10855), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10855), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10855), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10855), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10855), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10855), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10855), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10855), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_51 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10873;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_51 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10873), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10873), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10873), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10873), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10873), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10873), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10873), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10873), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10873), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_52 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10891;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_52 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10891), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10891), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10891), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10891), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10891), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10891), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10891), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10891), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10891), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_53 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10909;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_53 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10909), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10909), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10909), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10909), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10909), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10909), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10909), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10909), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10909), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_54 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10927;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_54 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10927), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10927), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10927), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10927), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10927), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10927), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10927), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10927), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10927), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_0000001f ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10945;

  SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10945), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10945), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10945), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10945), .XR(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10945), .XS(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10945), .XS(arstz), .Q(rdat[2]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10945), .XS(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10945), .XS(arstz), .Q(rdat[1]) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10945), .XS(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000004 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10963;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10963), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10963), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10963), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10963), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10963), .XR(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10963), .XS(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10963), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10963), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10963), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_4_00000004 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10981;

  SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10981), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10981), .XR(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10981), .XS(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10981), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10981), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH7_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10999;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10999), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10999), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10999), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10999), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10999), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10999), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10999), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10999), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_55 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11017;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_55 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11017), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11017), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11017), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11017), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11017), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11017), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11017), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11017), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11017), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_55 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_2 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_2 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[7]), .Y(n4) );
  INVX1 U4 ( .A(set2[0]), .Y(n3) );
  INVX1 U5 ( .A(set2[1]), .Y(n14) );
  INVX1 U6 ( .A(set2[3]), .Y(n15) );
  INVX1 U7 ( .A(set2[2]), .Y(n13) );
  INVX1 U8 ( .A(set2[4]), .Y(n1) );
  INVX1 U9 ( .A(set2[5]), .Y(n2) );
  NAND3X1 U10 ( .A(n16), .B(n4), .C(n2), .Y(n21) );
  NAND4X1 U11 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U12 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U13 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U14 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U15 ( .C(n1), .D(n12), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U16 ( .A(rdat[4]), .Y(n12) );
  AOI211X1 U17 ( .C(n2), .D(n11), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U18 ( .A(rdat[5]), .Y(n11) );
  AOI211X1 U19 ( .C(n13), .D(n10), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U20 ( .A(rdat[2]), .Y(n10) );
  AOI211X1 U21 ( .C(n14), .D(n9), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U22 ( .A(rdat[1]), .Y(n9) );
  AOI211X1 U23 ( .C(n3), .D(n8), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U24 ( .A(rdat[0]), .Y(n8) );
  AOI211X1 U25 ( .C(n16), .D(n6), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U26 ( .A(rdat[6]), .Y(n6) );
  AOI211X1 U27 ( .C(n4), .D(n5), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U28 ( .A(rdat[7]), .Y(n5) );
  AOI211X1 U29 ( .C(n15), .D(n7), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U30 ( .A(rdat[3]), .Y(n7) );
  NOR2X1 U31 ( .A(rdat[3]), .B(n15), .Y(irq[3]) );
  NOR2X1 U32 ( .A(rdat[2]), .B(n13), .Y(irq[2]) );
  NOR2X1 U33 ( .A(rdat[5]), .B(n2), .Y(irq[5]) );
  NOR2X1 U34 ( .A(rdat[4]), .B(n1), .Y(irq[4]) );
  NOR2X1 U35 ( .A(rdat[0]), .B(n3), .Y(irq[0]) );
  NOR2X1 U36 ( .A(rdat[7]), .B(n4), .Y(irq[7]) );
  NOR2X1 U37 ( .A(rdat[1]), .B(n14), .Y(irq[1]) );
  NOR2X1 U38 ( .A(rdat[6]), .B(n16), .Y(irq[6]) );
  INVX1 U39 ( .A(set2[6]), .Y(n16) );
endmodule


module glreg_WIDTH8_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11035;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11035), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11035), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11035), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11035), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11035), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11035), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11035), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11035), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11035), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_8 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR3XL U7 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_9 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR3XL U7 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_10 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR3XL U7 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n2), .Y(n8) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_11 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_12 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_13 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n4, n5, n6, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n5), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n6), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n4), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n4) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n6) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n5) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n10, n1, n2, n3, n5;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n9), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n8), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n10), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n3), .B(n5), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n3) );
  INVX1 U6 ( .A(test_so), .Y(n1) );
  AO22AXL U7 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n10) );
  NOR2X1 U8 ( .A(n5), .B(db_cnt_0_), .Y(n8) );
  OAI32X1 U9 ( .A(n3), .B(test_so), .C(n5), .D(n1), .E(n2), .Y(n9) );
  INVX1 U10 ( .A(n8), .Y(n2) );
endmodule


module dbnc_WIDTH2_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n10, n1, n2, n3, n5;

  SDFFRQX1 db_cnt_reg_1_ ( .D(n9), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n8), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n10), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n3), .B(n5), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n3) );
  INVX1 U6 ( .A(test_so), .Y(n1) );
  AO22AXL U7 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n10) );
  NOR2X1 U8 ( .A(n5), .B(db_cnt_0_), .Y(n8) );
  OAI32X1 U9 ( .A(n3), .B(test_so), .C(n5), .D(n1), .E(n2), .Y(n9) );
  INVX1 U10 ( .A(n8), .Y(n2) );
endmodule


module dbnc_WIDTH2_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n10, n1, n2, n3, n5;

  SDFFRQX1 db_cnt_reg_1_ ( .D(n9), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n8), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n10), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n3), .B(n5), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n3) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n10) );
  INVX1 U7 ( .A(test_so), .Y(n1) );
  NOR2X1 U8 ( .A(n5), .B(db_cnt_0_), .Y(n8) );
  OAI32X1 U9 ( .A(n3), .B(test_so), .C(n5), .D(n1), .E(n2), .Y(n9) );
  INVX1 U10 ( .A(n8), .Y(n2) );
endmodule


module dbnc_WIDTH2_3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n10, n4, n1, n2, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n9), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n8), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n10), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n3), .B(n4), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n3) );
  INVX1 U6 ( .A(test_so), .Y(n1) );
  AO22AXL U7 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n10) );
  NOR2X1 U8 ( .A(n4), .B(db_cnt_0_), .Y(n8) );
  OAI32X1 U9 ( .A(n3), .B(test_so), .C(n4), .D(n1), .E(n2), .Y(n9) );
  INVX1 U10 ( .A(n8), .Y(n2) );
endmodule


module dbnc_WIDTH2_4 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n5, n6, n7, n4, n1, n2, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n6), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n5), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n3), .B(n4), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n3) );
  INVX1 U6 ( .A(test_so), .Y(n1) );
  AO22AXL U7 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n5) );
  NOR2X1 U8 ( .A(n4), .B(db_cnt_0_), .Y(n7) );
  OAI32X1 U9 ( .A(n3), .B(test_so), .C(n4), .D(n1), .E(n2), .Y(n6) );
  INVX1 U10 ( .A(n7), .Y(n2) );
endmodule


module dbnc_WIDTH5_TIMEOUT30 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_3_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N8, N9, N10,
         N17, N18, N19, N20, N21, N22, net11053, n6, n1, n2, n3, n4, n5, n7;
  wire   [4:2] add_165_carry;

  HAD1X1 add_165_U1_1_1 ( .A(db_cnt_1_), .B(db_cnt_0_), .CO(add_165_carry[2]), 
        .SO(N8) );
  HAD1X1 add_165_U1_1_2 ( .A(db_cnt_2_), .B(add_165_carry[2]), .CO(
        add_165_carry[3]), .SO(N9) );
  HAD1X1 add_165_U1_1_3 ( .A(db_cnt_3_), .B(add_165_carry[3]), .CO(
        add_165_carry[4]), .SO(N10) );
  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH5_TIMEOUT30 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N17), .ENCLK(net11053), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_4_ ( .D(N22), .SIN(db_cnt_3_), .SMC(test_se), .C(
        net11053), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N21), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11053), .XR(rstz), .Q(db_cnt_3_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N20), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11053), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N19), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11053), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N18), .SIN(o_dbc), .SMC(test_se), .C(net11053), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n6), .SIN(d_org_0_), .SMC(test_se), .C(net11053), 
        .XR(rstz), .Q(o_dbc) );
  NOR2X1 U3 ( .A(n1), .B(n2), .Y(o_chg) );
  NAND21X1 U4 ( .B(n2), .A(n1), .Y(n4) );
  NOR21XL U5 ( .B(N8), .A(n4), .Y(N19) );
  NOR21XL U6 ( .B(N9), .A(n4), .Y(N20) );
  NOR21XL U7 ( .B(N10), .A(n4), .Y(N21) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  NAND4X1 U9 ( .A(test_so), .B(db_cnt_3_), .C(n5), .D(db_cnt_2_), .Y(n1) );
  NOR21XL U10 ( .B(db_cnt_1_), .A(db_cnt_0_), .Y(n5) );
  AO22AXL U11 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n6) );
  NOR2X1 U12 ( .A(n3), .B(n4), .Y(N22) );
  XNOR2XL U13 ( .A(test_so), .B(add_165_carry[4]), .Y(n3) );
  NOR2X1 U14 ( .A(db_cnt_0_), .B(n4), .Y(N18) );
  NAND42X1 U15 ( .C(db_cnt_0_), .D(db_cnt_1_), .A(n2), .B(n7), .Y(N17) );
  NOR3XL U16 ( .A(db_cnt_2_), .B(test_so), .C(db_cnt_3_), .Y(n7) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH5_TIMEOUT30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N19,
         net11071, n13, n6, n7, n8, n9, n10, n11, n12, n14, n1, n2, n3, n4, n5
;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11071), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11071), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11071), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11071), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(n1), .SIN(db_cnt_1_), .SMC(test_se), .C(net11071), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11071), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n2) );
  NOR2X1 U4 ( .A(n2), .B(n11), .Y(n9) );
  NOR21XL U5 ( .B(n6), .A(n7), .Y(n8) );
  NOR2X1 U6 ( .A(n3), .B(n4), .Y(n11) );
  AOI211X1 U7 ( .C(n3), .D(n4), .A(n2), .B(n11), .Y(N17) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  GEN2XL U9 ( .D(n8), .E(n5), .C(n9), .B(test_so), .A(n10), .Y(N19) );
  NOR42XL U10 ( .C(n11), .D(db_cnt_2_), .A(n2), .B(test_so), .Y(n10) );
  INVX1 U11 ( .A(n12), .Y(n1) );
  AOI32X1 U12 ( .A(n11), .B(n5), .C(n8), .D(db_cnt_2_), .E(n9), .Y(n12) );
  AO22AXL U13 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U14 ( .A(n6), .B(n7), .Y(o_chg) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  NAND4X1 U16 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(n3), .Y(n6) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n5) );
  INVX1 U18 ( .A(db_cnt_1_), .Y(n4) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n2), .Y(N16) );
  NAND3X1 U20 ( .A(n7), .B(n3), .C(n14), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N19,
         net11089, n13, n6, n7, n8, n9, n10, n11, n12, n14, n1, n2, n3, n4, n5
;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11089), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11089), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11089), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11089), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(n1), .SIN(db_cnt_1_), .SMC(test_se), .C(net11089), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11089), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n2) );
  NOR2X1 U4 ( .A(n2), .B(n11), .Y(n9) );
  NOR21XL U5 ( .B(n6), .A(n7), .Y(n8) );
  NOR2X1 U6 ( .A(n3), .B(n4), .Y(n11) );
  AOI211X1 U7 ( .C(n3), .D(n4), .A(n2), .B(n11), .Y(N17) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  GEN2XL U9 ( .D(n8), .E(n5), .C(n9), .B(test_so), .A(n10), .Y(N19) );
  NOR42XL U10 ( .C(n11), .D(db_cnt_2_), .A(n2), .B(test_so), .Y(n10) );
  INVX1 U11 ( .A(n12), .Y(n1) );
  AOI32X1 U12 ( .A(n11), .B(n5), .C(n8), .D(db_cnt_2_), .E(n9), .Y(n12) );
  AO22AXL U13 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U14 ( .A(n6), .B(n7), .Y(o_chg) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  NAND4X1 U16 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(n3), .Y(n6) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n5) );
  INVX1 U18 ( .A(db_cnt_1_), .Y(n4) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n2), .Y(N16) );
  NAND3X1 U20 ( .A(n7), .B(n3), .C(n14), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N19,
         net11107, n13, n6, n7, n8, n9, n10, n11, n12, n14, n1, n2, n3, n4, n5
;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11107), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11107), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11107), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11107), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(n1), .SIN(db_cnt_1_), .SMC(test_se), .C(net11107), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11107), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n2) );
  NOR2X1 U4 ( .A(n2), .B(n11), .Y(n9) );
  NOR21XL U5 ( .B(n6), .A(n7), .Y(n8) );
  NOR2X1 U6 ( .A(n3), .B(n4), .Y(n11) );
  AOI211X1 U7 ( .C(n3), .D(n4), .A(n2), .B(n11), .Y(N17) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  GEN2XL U9 ( .D(n8), .E(n5), .C(n9), .B(test_so), .A(n10), .Y(N19) );
  NOR42XL U10 ( .C(n11), .D(db_cnt_2_), .A(n2), .B(test_so), .Y(n10) );
  INVX1 U11 ( .A(n12), .Y(n1) );
  AOI32X1 U12 ( .A(n11), .B(n5), .C(n8), .D(db_cnt_2_), .E(n9), .Y(n12) );
  AO22AXL U13 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U14 ( .A(n6), .B(n7), .Y(o_chg) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  NAND4X1 U16 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(n3), .Y(n6) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n5) );
  INVX1 U18 ( .A(db_cnt_1_), .Y(n4) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n2), .Y(N16) );
  NAND3X1 U20 ( .A(n7), .B(n3), .C(n14), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000028 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11125;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11125), .TE(test_se) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11125), .XS(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11125), .XS(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11125), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11125), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11125), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11125), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11125), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11125), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_56 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11143;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_56 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11143), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11143), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11143), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11143), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11143), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11143), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11143), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11143), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11143), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_56 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_57 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11161;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_57 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11161), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11161), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11161), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11161), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11161), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11161), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11161), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11161), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11161), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_57 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_58 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11179;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_58 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11179), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11179), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11179), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11179), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11179), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11179), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11179), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11179), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11179), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_58 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_59 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11197;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_59 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11197), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11197), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11197), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11197), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11197), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11197), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11197), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11197), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11197), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_59 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_60 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11215;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_60 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11215), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11215), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11215), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11215), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11215), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11215), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11215), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11215), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11215), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_60 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_61 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11233;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_61 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11233), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11233), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11233), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11233), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11233), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11233), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11233), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11233), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11233), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_61 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_62 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11251;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_62 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11251), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11251), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11251), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11251), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11251), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11251), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11251), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11251), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11251), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_62 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_63 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11269;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_63 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11269), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11269), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11269), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11269), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11269), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11269), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11269), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11269), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11269), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_63 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11287;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11287), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11287), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11287), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11287), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11287), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_64 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11305;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_64 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11305), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11305), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11305), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11305), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11305), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11305), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11305), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11305), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11305), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_64 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_3 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_3 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[0]), .Y(n12) );
  INVX1 U4 ( .A(set2[1]), .Y(n11) );
  INVX1 U5 ( .A(set2[2]), .Y(n16) );
  INVX1 U6 ( .A(set2[3]), .Y(n15) );
  INVX1 U7 ( .A(set2[4]), .Y(n10) );
  NAND3X1 U8 ( .A(n13), .B(n9), .C(n14), .Y(n21) );
  NAND4X1 U9 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U10 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U11 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U12 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U13 ( .C(n12), .D(n8), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U14 ( .A(rdat[0]), .Y(n8) );
  AOI211X1 U15 ( .C(n16), .D(n7), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U16 ( .A(rdat[2]), .Y(n7) );
  AOI211X1 U17 ( .C(n10), .D(n5), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U18 ( .A(rdat[4]), .Y(n5) );
  AOI211X1 U19 ( .C(n14), .D(n4), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U20 ( .A(rdat[5]), .Y(n4) );
  AOI211X1 U21 ( .C(n9), .D(n3), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U22 ( .A(rdat[7]), .Y(n3) );
  AOI211X1 U23 ( .C(n11), .D(n2), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U24 ( .A(rdat[1]), .Y(n2) );
  AOI211X1 U25 ( .C(n13), .D(n1), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U26 ( .A(rdat[6]), .Y(n1) );
  AOI211X1 U27 ( .C(n15), .D(n6), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U28 ( .A(rdat[3]), .Y(n6) );
  NOR2X1 U29 ( .A(rdat[0]), .B(n12), .Y(irq[0]) );
  NOR2X1 U30 ( .A(rdat[1]), .B(n11), .Y(irq[1]) );
  NOR2X1 U31 ( .A(rdat[2]), .B(n16), .Y(irq[2]) );
  NOR2X1 U32 ( .A(rdat[3]), .B(n15), .Y(irq[3]) );
  INVX1 U33 ( .A(set2[6]), .Y(n13) );
  INVX1 U34 ( .A(set2[7]), .Y(n9) );
  INVX1 U35 ( .A(set2[5]), .Y(n14) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n10), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n13), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[5]), .B(n14), .Y(irq[5]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n9), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11323;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11323), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11323), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11323), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11323), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11323), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11323), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11323), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11323), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11323), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_65 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11341;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_65 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11341), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11341), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11341), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11341), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11341), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11341), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11341), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11341), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11341), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_65 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_66 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11359;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_66 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11359), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11359), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11359), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11359), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11359), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11359), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11359), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11359), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11359), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_66 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000032 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11377;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11377), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11377), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11377), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11377), .XR(arstz), .Q(rdat[2]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11377), .XS(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11377), .XS(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11377), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11377), .XR(arstz), .Q(rdat[0]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11377), .XS(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000098 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11395;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11395), .TE(test_se) );
  SDFFSQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11395), .XS(arstz), .Q(rdat[7]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11395), .XS(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11395), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11395), .XR(arstz), .Q(rdat[2]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11395), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11395), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11395), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11395), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_000000f0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11413;

  SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11413), .TE(test_se) );
  SDFFSQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11413), .XS(arstz), .Q(rdat[7]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11413), .XS(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11413), .XS(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11413), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11413), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11413), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11413), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11413), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH1_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH1_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH2_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2, n3, n1;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(n3), .SIN(rdat[0]), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[1]) );
  AO22XL U2 ( .A(we), .B(wdat[1]), .C(rdat[1]), .D(n1), .Y(n3) );
  INVXL U3 ( .A(we), .Y(n1) );
  AO22XL U4 ( .A(wdat[0]), .B(we), .C(rdat[0]), .D(n1), .Y(n2) );
endmodule


module glreg_WIDTH3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [2:0] wdat;
  output [2:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11431;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11431), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11431), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11431), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11431), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000011 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11449;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11449), .TE(test_se) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11449), .XS(arstz), .Q(rdat[0]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11449), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11449), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11449), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11449), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11449), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11449), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11449), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000001 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11467;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11467), .TE(test_se) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11467), .XS(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11467), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11467), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11467), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11467), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11467), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11467), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11467), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_67 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11485;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_67 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11485), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11485), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11485), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11485), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11485), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11485), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11485), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11485), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11485), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_67 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_4 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_4 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[4]), .Y(n13) );
  INVX1 U4 ( .A(set2[7]), .Y(n12) );
  NAND3X1 U5 ( .A(n11), .B(n12), .C(n10), .Y(n21) );
  INVX1 U6 ( .A(set2[3]), .Y(n14) );
  INVX1 U7 ( .A(set2[0]), .Y(n9) );
  INVX1 U8 ( .A(set2[1]), .Y(n16) );
  INVX1 U9 ( .A(set2[5]), .Y(n10) );
  INVX1 U10 ( .A(set2[6]), .Y(n11) );
  INVX1 U11 ( .A(set2[2]), .Y(n15) );
  NAND4X1 U12 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U13 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U14 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U15 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U16 ( .C(n10), .D(n1), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U17 ( .A(rdat[5]), .Y(n1) );
  AOI211X1 U18 ( .C(n12), .D(n8), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U19 ( .A(rdat[7]), .Y(n8) );
  AOI211X1 U20 ( .C(n13), .D(n7), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U21 ( .A(rdat[4]), .Y(n7) );
  AOI211X1 U22 ( .C(n11), .D(n6), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U23 ( .A(rdat[6]), .Y(n6) );
  AOI211X1 U24 ( .C(n9), .D(n5), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U25 ( .A(rdat[0]), .Y(n5) );
  AOI211X1 U26 ( .C(n16), .D(n4), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U27 ( .A(rdat[1]), .Y(n4) );
  AOI211X1 U28 ( .C(n14), .D(n3), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U29 ( .A(rdat[3]), .Y(n3) );
  AOI211X1 U30 ( .C(n15), .D(n2), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U31 ( .A(rdat[2]), .Y(n2) );
  NOR2X1 U32 ( .A(rdat[7]), .B(n12), .Y(irq[7]) );
  NOR2X1 U33 ( .A(rdat[6]), .B(n11), .Y(irq[6]) );
  NOR2X1 U34 ( .A(rdat[0]), .B(n9), .Y(irq[0]) );
  NOR2X1 U35 ( .A(rdat[4]), .B(n13), .Y(irq[4]) );
  NOR2X1 U36 ( .A(rdat[3]), .B(n14), .Y(irq[3]) );
  NOR2X1 U37 ( .A(rdat[2]), .B(n15), .Y(irq[2]) );
  NOR2X1 U38 ( .A(rdat[1]), .B(n16), .Y(irq[1]) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n10), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11503;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11503), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11503), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11503), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11503), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11503), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11503), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11503), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11503), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11503), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_68 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11521;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_68 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11521), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11521), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11521), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11521), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11521), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11521), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11521), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11521), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11521), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_68 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_7_70 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11539;

  SNPS_CLOCK_GATE_HIGH_glreg_7_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11539), .TE(test_se) );
  SDFFSQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11539), .XS(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11539), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11539), .XR(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11539), .XS(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11539), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11539), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11539), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_7_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_1_1_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFSQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XS(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_1_1_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFSQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XS(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_6_00000018 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11557;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11557), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11557), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11557), .XR(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11557), .XS(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11557), .XR(arstz), .Q(rdat[1]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11557), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11557), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_69 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11575;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_69 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11575), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11575), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11575), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11575), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11575), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11575), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11575), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11575), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11575), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_69 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_70 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11593;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11593), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11593), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11593), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11593), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11593), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11593), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11593), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11593), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11593), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_71 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11611;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_71 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11611), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11611), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11611), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11611), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11611), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11611), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11611), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11611), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11611), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_71 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_72 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11629;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_72 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11629), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11629), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11629), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11629), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11629), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11629), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11629), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11629), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11629), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_72 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_73 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11647;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_73 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11647), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11647), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11647), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11647), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11647), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11647), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11647), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11647), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11647), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_73 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11665;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11665), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11665), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11665), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11665), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11665), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11665), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_74 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11683;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_74 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11683), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11683), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11683), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11683), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11683), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11683), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11683), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11683), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11683), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_74 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_75 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11701;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_75 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11701), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11701), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11701), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11701), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11701), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11701), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11701), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11701), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11701), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_75 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_76 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11719;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_76 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11719), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11719), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11719), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11719), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11719), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11719), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11719), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11719), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11719), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_76 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_77 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11737;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_77 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11737), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11737), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11737), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11737), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11737), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11737), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11737), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11737), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11737), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_77 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_5 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_5 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[1]), .Y(n14) );
  INVX1 U3 ( .A(set2[4]), .Y(n2) );
  NAND4X1 U4 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U5 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U6 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  NOR4XL U7 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U8 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NAND3X1 U9 ( .A(n16), .B(n1), .C(n3), .Y(n21) );
  INVX1 U10 ( .A(set2[3]), .Y(n4) );
  INVX1 U11 ( .A(set2[2]), .Y(n5) );
  INVX1 U12 ( .A(set2[0]), .Y(n15) );
  INVX1 U13 ( .A(set2[5]), .Y(n3) );
  NOR2X1 U14 ( .A(rdat[4]), .B(n2), .Y(irq[4]) );
  NOR2X1 U15 ( .A(rdat[5]), .B(n3), .Y(irq[5]) );
  AOI211X1 U16 ( .C(n2), .D(n9), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U17 ( .A(rdat[4]), .Y(n9) );
  AOI211X1 U18 ( .C(n3), .D(n8), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U19 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U20 ( .C(n15), .D(n13), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U21 ( .A(rdat[0]), .Y(n13) );
  AOI211X1 U22 ( .C(n14), .D(n12), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U23 ( .A(rdat[1]), .Y(n12) );
  AOI211X1 U24 ( .C(n5), .D(n11), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U25 ( .A(rdat[2]), .Y(n11) );
  AOI211X1 U26 ( .C(n4), .D(n10), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U27 ( .A(rdat[3]), .Y(n10) );
  AOI211X1 U28 ( .C(n16), .D(n7), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U29 ( .A(rdat[6]), .Y(n7) );
  AOI211X1 U30 ( .C(n1), .D(n6), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U31 ( .A(rdat[7]), .Y(n6) );
  NOR2X1 U32 ( .A(rdat[2]), .B(n5), .Y(irq[2]) );
  NOR2X1 U33 ( .A(rdat[3]), .B(n4), .Y(irq[3]) );
  INVX1 U34 ( .A(set2[6]), .Y(n16) );
  NOR2X1 U35 ( .A(rdat[6]), .B(n16), .Y(irq[6]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n15), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[1]), .B(n14), .Y(irq[1]) );
  INVX1 U38 ( .A(set2[7]), .Y(n1) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n1), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11755;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11755), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11755), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11755), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11755), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11755), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11755), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11755), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11755), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11755), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_6 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_6 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[3]), .Y(n1) );
  INVX1 U3 ( .A(set2[7]), .Y(n5) );
  INVX1 U4 ( .A(set2[6]), .Y(n2) );
  NOR4XL U5 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NAND4X1 U6 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR3XL U7 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U8 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U9 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U10 ( .A(set2[1]), .Y(n4) );
  INVX1 U11 ( .A(set2[2]), .Y(n6) );
  NAND3X1 U12 ( .A(n2), .B(n5), .C(n16), .Y(n21) );
  INVX1 U13 ( .A(set2[4]), .Y(n3) );
  INVX1 U14 ( .A(set2[0]), .Y(n15) );
  NOR2X1 U15 ( .A(rdat[6]), .B(n2), .Y(irq[6]) );
  NOR2X1 U16 ( .A(rdat[7]), .B(n5), .Y(irq[7]) );
  AOI211X1 U17 ( .C(n4), .D(n14), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U18 ( .A(rdat[1]), .Y(n14) );
  AOI211X1 U19 ( .C(n3), .D(n13), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U20 ( .A(rdat[4]), .Y(n13) );
  AOI211X1 U21 ( .C(n16), .D(n12), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U22 ( .A(rdat[5]), .Y(n12) );
  AOI211X1 U23 ( .C(n15), .D(n11), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U24 ( .A(rdat[0]), .Y(n11) );
  AOI211X1 U25 ( .C(n6), .D(n10), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U26 ( .A(rdat[2]), .Y(n10) );
  AOI211X1 U27 ( .C(n2), .D(n8), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U28 ( .A(rdat[6]), .Y(n8) );
  AOI211X1 U29 ( .C(n5), .D(n7), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U30 ( .A(rdat[7]), .Y(n7) );
  AOI211X1 U31 ( .C(n1), .D(n9), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U32 ( .A(rdat[3]), .Y(n9) );
  NOR2X1 U33 ( .A(rdat[0]), .B(n15), .Y(irq[0]) );
  NOR2X1 U34 ( .A(rdat[1]), .B(n4), .Y(irq[1]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n6), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n3), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[3]), .B(n1), .Y(irq[3]) );
  INVX1 U38 ( .A(set2[5]), .Y(n16) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_6 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11773;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11773), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11773), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11773), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11773), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11773), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11773), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11773), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11773), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11773), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_78 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11791;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_78 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11791), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11791), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11791), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11791), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11791), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11791), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11791), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11791), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11791), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_78 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_79 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11809;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_79 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11809), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11809), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11809), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11809), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11809), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11809), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11809), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11809), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11809), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_79 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ictlr_a0 ( bkpt_ena, bkpt_pc, memaddr_c, memaddr, mcu_psr_c, mcu_psw, 
        hit_ps_c, hit_ps, mempsack, memdatao, o_set_hold, o_bkp_hold, 
        o_ofs_inc, o_inst, d_inst, sfr_psrack, sfr_psofs, sfr_psr, sfr_psw, 
        dw_rst, dw_ena, sfr_wdat, pmem_pgm, pmem_re, pmem_csb, pmem_clk, 
        pmem_a, pmem_q0, pmem_q1, pmem_twlb, wd_twlb, we_twlb, pwrdn_rst, 
        r_pwdn_en, r_multi, r_hold_mcu, clk, srst, test_si3, test_si2, 
        test_si1, test_so2, test_so1, test_se );
  input [14:0] bkpt_pc;
  input [14:0] memaddr_c;
  input [14:0] memaddr;
  input [7:0] memdatao;
  output [7:0] o_inst;
  output [7:0] d_inst;
  input [14:0] sfr_psofs;
  input [7:0] sfr_wdat;
  output [1:0] pmem_clk;
  output [15:0] pmem_a;
  input [7:0] pmem_q0;
  input [7:0] pmem_q1;
  output [1:0] pmem_twlb;
  input [1:0] wd_twlb;
  input bkpt_ena, mcu_psr_c, mcu_psw, hit_ps_c, hit_ps, sfr_psr, sfr_psw,
         dw_rst, dw_ena, we_twlb, pwrdn_rst, r_pwdn_en, r_multi, r_hold_mcu,
         clk, srst, test_si3, test_si2, test_si1, test_se;
  output mempsack, o_set_hold, o_bkp_hold, o_ofs_inc, sfr_psrack, pmem_pgm,
         pmem_re, pmem_csb, test_so2, test_so1;
  wire   N152, N153, N154, c_buf_22__7_, c_buf_22__6_, c_buf_22__5_,
         c_buf_22__4_, c_buf_22__3_, c_buf_22__2_, c_buf_22__1_, c_buf_22__0_,
         c_buf_21__7_, c_buf_21__6_, c_buf_21__5_, c_buf_21__4_, c_buf_21__3_,
         c_buf_21__2_, c_buf_21__1_, c_buf_21__0_, c_buf_20__7_, c_buf_20__6_,
         c_buf_20__5_, c_buf_20__4_, c_buf_20__3_, c_buf_20__2_, c_buf_20__1_,
         c_buf_20__0_, c_buf_19__7_, c_buf_19__6_, c_buf_19__5_, c_buf_19__4_,
         c_buf_19__3_, c_buf_19__2_, c_buf_19__1_, c_buf_19__0_, c_buf_18__7_,
         c_buf_18__6_, c_buf_18__5_, c_buf_18__4_, c_buf_18__3_, c_buf_18__2_,
         c_buf_18__1_, c_buf_18__0_, c_buf_17__7_, c_buf_17__6_, c_buf_17__5_,
         c_buf_17__4_, c_buf_17__3_, c_buf_17__2_, c_buf_17__1_, c_buf_17__0_,
         c_buf_16__7_, c_buf_16__6_, c_buf_16__5_, c_buf_16__4_, c_buf_16__3_,
         c_buf_16__2_, c_buf_16__1_, c_buf_16__0_, wspp_cnt_5_, wspp_cnt_4_,
         wspp_cnt_3_, wspp_cnt_2_, wspp_cnt_1_, wspp_cnt_0_, d_psrd, r_rdy,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617,
         N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628,
         N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639,
         N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650,
         N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661,
         N662, N757, N759, N786, N787, N788, N789, N790, N791, N792, N793,
         N795, N796, N797, N798, N799, N800, N801, N820, N821, N822, N823,
         N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834,
         N835, N836, N837, N838, N839, N840, N842, N843, N844, N845, N846,
         N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863,
         N864, N865, N866, N867, N868, N874, N875, N876, N877, N878, N879,
         N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890,
         N891, N892, N893, N894, N895, N896, N897, N898, N899, un_hold,
         net11835, net11841, net11846, net11851, net11856, net11861, net11866,
         net11871, net11876, net11881, net11886, net11891, net11896, net11901,
         net11906, net11911, net11916, net11921, net11926, net11931, net11936,
         net11941, net11946, net11951, net11956, net11961, net11966, net11971,
         net11976, net11981, n93, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n874, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n285, n286, n287, n288, n289, n291, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n306, n307, n308, n309,
         n310, n311, n312, n313, n316, n317, n318, n319, n320, n321, n322,
         n323, n326, n327, n328, n329, n330, n331, n332, n333, n336, n337,
         n338, n339, n340, n341, n342, n343, n349, n350, n351, n352, n353,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n376, n377, n378, n379, n380, n383, n384,
         n385, n387, n388, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n417, n418, n465, n467, n541, n552, n553, n554, n555,
         n556, n574, n575, n576, n762, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n283, n284, n290, n292, n293, n294, n304, n305, n314, n315,
         n324, n325, n334, n335, n344, n345, n346, n347, n348, n354, n355,
         n356, n357, n358, n374, n375, n381, n382, n386, n389, n390, n391,
         n392, n414, n415, n416, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n466, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940;
  wire   [3:0] d_hold;
  wire   [1:0] dummy;
  wire   [3:0] cs_ft;
  wire   [4:0] c_ptr;
  wire   [14:0] c_adr;
  wire   [14:13] adr_p;
  wire   [7:0] rd_buf;
  wire   [7:0] dbg_01;
  wire   [7:0] dbg_02;
  wire   [7:0] dbg_03;
  wire   [7:0] dbg_04;
  wire   [7:0] dbg_05;
  wire   [7:0] dbg_06;
  wire   [7:0] dbg_07;
  wire   [7:0] dbg_08;
  wire   [7:0] dbg_09;
  wire   [7:0] dbg_0a;
  wire   [7:0] dbg_0b;
  wire   [7:0] dbg_0c;
  wire   [7:0] dbg_0d;
  wire   [7:0] dbg_0e;
  wire   [7:0] dbg_0f;
  wire   [7:0] wr_buf;
  wire   [14:0] pre_1_adr;

  SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 clk_gate_wspp_cnt_reg ( .CLK(clk), .EN(N899), 
        .ENCLK(net11835), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 clk_gate_a_bit_reg ( .CLK(clk), .EN(N898), 
        .ENCLK(net11841), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 clk_gate_adr_p_reg ( .CLK(clk), .EN(N853), 
        .ENCLK(net11846), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 clk_gate_c_buf_reg_23_ ( .CLK(clk), .EN(
        N897), .ENCLK(net11851), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 clk_gate_c_buf_reg_22_ ( .CLK(clk), .EN(
        N896), .ENCLK(net11856), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 clk_gate_c_buf_reg_21_ ( .CLK(clk), .EN(
        N895), .ENCLK(net11861), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 clk_gate_c_buf_reg_20_ ( .CLK(clk), .EN(
        N894), .ENCLK(net11866), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 clk_gate_c_buf_reg_19_ ( .CLK(clk), .EN(
        N893), .ENCLK(net11871), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 clk_gate_c_buf_reg_18_ ( .CLK(clk), .EN(
        N892), .ENCLK(net11876), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 clk_gate_c_buf_reg_17_ ( .CLK(clk), .EN(
        N891), .ENCLK(net11881), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 clk_gate_c_buf_reg_16_ ( .CLK(clk), .EN(
        N890), .ENCLK(net11886), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 clk_gate_c_buf_reg_15_ ( .CLK(clk), .EN(
        N889), .ENCLK(net11891), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 clk_gate_c_buf_reg_14_ ( .CLK(clk), .EN(
        N888), .ENCLK(net11896), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 clk_gate_c_buf_reg_13_ ( .CLK(clk), .EN(
        N887), .ENCLK(net11901), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 clk_gate_c_buf_reg_12_ ( .CLK(clk), .EN(
        N886), .ENCLK(net11906), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 clk_gate_c_buf_reg_11_ ( .CLK(clk), .EN(
        N885), .ENCLK(net11911), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 clk_gate_c_buf_reg_10_ ( .CLK(clk), .EN(
        N884), .ENCLK(net11916), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 clk_gate_c_buf_reg_9_ ( .CLK(clk), .EN(N883), .ENCLK(net11921), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 clk_gate_c_buf_reg_8_ ( .CLK(clk), .EN(N882), .ENCLK(net11926), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 clk_gate_c_buf_reg_7_ ( .CLK(clk), .EN(N881), .ENCLK(net11931), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 clk_gate_c_buf_reg_6_ ( .CLK(clk), .EN(N880), .ENCLK(net11936), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 clk_gate_c_buf_reg_5_ ( .CLK(clk), .EN(N879), 
        .ENCLK(net11941), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 clk_gate_c_buf_reg_4_ ( .CLK(clk), .EN(N878), 
        .ENCLK(net11946), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 clk_gate_c_buf_reg_3_ ( .CLK(clk), .EN(N877), 
        .ENCLK(net11951), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 clk_gate_c_buf_reg_2_ ( .CLK(clk), .EN(N876), 
        .ENCLK(net11956), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 clk_gate_c_buf_reg_1_ ( .CLK(clk), .EN(N875), 
        .ENCLK(net11961), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 clk_gate_c_buf_reg_0_ ( .CLK(clk), .EN(N874), 
        .ENCLK(net11966), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 clk_gate_c_ptr_reg ( .CLK(clk), .EN(n93), 
        .ENCLK(net11971), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 clk_gate_c_adr_reg ( .CLK(clk), .EN(N825), 
        .ENCLK(net11976), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 clk_gate_cs_ft_reg ( .CLK(clk), .EN(N820), 
        .ENCLK(net11981), .TE(test_se) );
  ictlr_a0_DW01_inc_1 add_242 ( .A(c_adr), .SUM({N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431}) );
  ictlr_a0_DW01_inc_2 r492 ( .A({adr_p, pmem_a[15:9], pmem_a[5:0]}), .SUM(
        pre_1_adr) );
  SDFFNQX1 ck_n_reg_1_ ( .D(n642), .SIN(pmem_clk[0]), .SMC(test_se), .XC(clk), 
        .Q(pmem_clk[1]) );
  SDFFNQXL ck_n_reg_0_ ( .D(n641), .SIN(test_si1), .SMC(test_se), .XC(clk), 
        .Q(pmem_clk[0]) );
  SDFFQX2 a_bit_reg_2_ ( .D(N759), .SIN(pmem_a[7]), .SMC(test_se), .C(net11841), .Q(pmem_a[8]) );
  SDFFQX2 a_bit_reg_0_ ( .D(N757), .SIN(test_si2), .SMC(test_se), .C(net11841), 
        .Q(pmem_a[6]) );
  SDFFQX1 wspp_cnt_reg_2_ ( .D(N797), .SIN(wspp_cnt_1_), .SMC(test_se), .C(
        net11835), .Q(wspp_cnt_2_) );
  SDFFQX1 wspp_cnt_reg_0_ ( .D(N795), .SIN(un_hold), .SMC(test_se), .C(
        net11835), .Q(wspp_cnt_0_) );
  SDFFQX1 wspp_cnt_reg_1_ ( .D(N796), .SIN(wspp_cnt_0_), .SMC(test_se), .C(
        net11835), .Q(wspp_cnt_1_) );
  SDFFQX1 d_hold_reg_3_ ( .D(N154), .SIN(d_hold[2]), .SMC(test_se), .C(clk), 
        .Q(d_hold[3]) );
  SDFFQX1 d_hold_reg_0_ ( .D(n874), .SIN(cs_ft[3]), .SMC(test_se), .C(clk), 
        .Q(d_hold[0]) );
  SDFFQX1 d_hold_reg_1_ ( .D(N152), .SIN(d_hold[0]), .SMC(test_se), .C(clk), 
        .Q(d_hold[1]) );
  SDFFQX1 d_hold_reg_2_ ( .D(N153), .SIN(d_hold[1]), .SMC(test_se), .C(clk), 
        .Q(d_hold[2]) );
  SDFFQX1 dummy_reg_1_ ( .D(n650), .SIN(dummy[0]), .SMC(test_se), .C(clk), .Q(
        dummy[1]) );
  SDFFQX1 dummy_reg_0_ ( .D(n651), .SIN(n24), .SMC(test_se), .C(clk), .Q(
        dummy[0]) );
  SDFFQX1 d_psrd_reg ( .D(n649), .SIN(d_hold[3]), .SMC(test_se), .C(net11981), 
        .Q(d_psrd) );
  SDFFQX2 adr_p_reg_3_ ( .D(N857), .SIN(pmem_a[2]), .SMC(test_se), .C(net11846), .Q(pmem_a[3]) );
  SDFFQX2 adr_p_reg_4_ ( .D(N858), .SIN(pmem_a[3]), .SMC(test_se), .C(net11846), .Q(pmem_a[4]) );
  SDFFQX2 adr_p_reg_5_ ( .D(N859), .SIN(pmem_a[4]), .SMC(test_se), .C(net11846), .Q(pmem_a[5]) );
  SDFFQX2 adr_p_reg_1_ ( .D(N855), .SIN(pmem_a[0]), .SMC(test_se), .C(net11846), .Q(pmem_a[1]) );
  SDFFQX2 adr_p_reg_2_ ( .D(N856), .SIN(pmem_a[1]), .SMC(test_se), .C(net11846), .Q(pmem_a[2]) );
  SDFFQX1 c_adr_reg_14_ ( .D(N840), .SIN(c_adr[13]), .SMC(test_se), .C(
        net11976), .Q(c_adr[14]) );
  SDFFQX1 c_adr_reg_13_ ( .D(N839), .SIN(c_adr[12]), .SMC(test_se), .C(
        net11976), .Q(c_adr[13]) );
  SDFFQX1 c_adr_reg_12_ ( .D(N838), .SIN(c_adr[11]), .SMC(test_se), .C(
        net11976), .Q(c_adr[12]) );
  SDFFQX1 c_adr_reg_8_ ( .D(N834), .SIN(c_adr[7]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[8]) );
  SDFFQX1 c_adr_reg_11_ ( .D(N837), .SIN(c_adr[10]), .SMC(test_se), .C(
        net11976), .Q(c_adr[11]) );
  SDFFQX1 c_adr_reg_10_ ( .D(N836), .SIN(c_adr[9]), .SMC(test_se), .C(net11976), .Q(c_adr[10]) );
  SDFFQX1 c_adr_reg_9_ ( .D(N835), .SIN(c_adr[8]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[9]) );
  SDFFQX1 c_adr_reg_7_ ( .D(N833), .SIN(c_adr[6]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[7]) );
  SDFFQX1 c_adr_reg_6_ ( .D(N832), .SIN(c_adr[5]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[6]) );
  SDFFQX1 c_adr_reg_5_ ( .D(N831), .SIN(c_adr[4]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[5]) );
  SDFFQX1 c_ptr_reg_4_ ( .D(N846), .SIN(c_ptr[3]), .SMC(test_se), .C(net11971), 
        .Q(c_ptr[4]) );
  SDFFQX1 c_ptr_reg_3_ ( .D(N845), .SIN(c_ptr[2]), .SMC(test_se), .C(net11971), 
        .Q(c_ptr[3]) );
  SDFFQX1 c_ptr_reg_2_ ( .D(N844), .SIN(c_ptr[1]), .SMC(test_se), .C(net11971), 
        .Q(c_ptr[2]) );
  SDFFQX1 c_ptr_reg_1_ ( .D(N843), .SIN(c_ptr[0]), .SMC(test_se), .C(net11971), 
        .Q(c_ptr[1]) );
  SDFFQX1 c_ptr_reg_0_ ( .D(N842), .SIN(wr_buf[7]), .SMC(test_se), .C(net11971), .Q(c_ptr[0]) );
  SDFFQX1 c_buf_reg_7__0_ ( .D(N535), .SIN(dbg_06[7]), .SMC(test_se), .C(
        net11931), .Q(dbg_07[0]) );
  SDFFQX1 c_buf_reg_6__6_ ( .D(N533), .SIN(dbg_06[5]), .SMC(test_se), .C(
        net11936), .Q(dbg_06[6]) );
  SDFFQX1 c_buf_reg_6__5_ ( .D(N532), .SIN(dbg_06[4]), .SMC(test_se), .C(
        net11936), .Q(dbg_06[5]) );
  SDFFQX1 c_buf_reg_6__4_ ( .D(N531), .SIN(dbg_06[3]), .SMC(test_se), .C(
        net11936), .Q(dbg_06[4]) );
  SDFFQX1 c_buf_reg_6__3_ ( .D(N530), .SIN(dbg_06[2]), .SMC(test_se), .C(
        net11936), .Q(dbg_06[3]) );
  SDFFQX1 c_buf_reg_5__0_ ( .D(N519), .SIN(dbg_04[7]), .SMC(test_se), .C(
        net11941), .Q(dbg_05[0]) );
  SDFFQX1 c_buf_reg_1__0_ ( .D(N487), .SIN(rd_buf[7]), .SMC(test_se), .C(
        net11961), .Q(dbg_01[0]) );
  SDFFQX1 c_buf_reg_6__0_ ( .D(N527), .SIN(dbg_05[7]), .SMC(test_se), .C(
        net11936), .Q(dbg_06[0]) );
  SDFFQX1 c_buf_reg_2__0_ ( .D(N495), .SIN(dbg_01[7]), .SMC(test_se), .C(
        net11956), .Q(dbg_02[0]) );
  SDFFQX1 c_buf_reg_3__0_ ( .D(N503), .SIN(dbg_02[7]), .SMC(test_se), .C(
        net11951), .Q(dbg_03[0]) );
  SDFFQX1 c_buf_reg_4__0_ ( .D(N511), .SIN(dbg_03[7]), .SMC(test_se), .C(
        net11946), .Q(dbg_04[0]) );
  SDFFQX1 c_buf_reg_10__6_ ( .D(N565), .SIN(dbg_0a[5]), .SMC(test_se), .C(
        net11916), .Q(dbg_0a[6]) );
  SDFFQX1 c_buf_reg_10__5_ ( .D(N564), .SIN(dbg_0a[4]), .SMC(test_se), .C(
        net11916), .Q(dbg_0a[5]) );
  SDFFQX1 c_buf_reg_10__4_ ( .D(N563), .SIN(dbg_0a[3]), .SMC(test_se), .C(
        net11916), .Q(dbg_0a[4]) );
  SDFFQX1 c_buf_reg_10__3_ ( .D(N562), .SIN(dbg_0a[2]), .SMC(test_se), .C(
        net11916), .Q(dbg_0a[3]) );
  SDFFQX1 c_buf_reg_10__2_ ( .D(N561), .SIN(dbg_0a[1]), .SMC(test_se), .C(
        net11916), .Q(dbg_0a[2]) );
  SDFFQX1 c_buf_reg_10__0_ ( .D(N559), .SIN(dbg_09[7]), .SMC(test_se), .C(
        net11916), .Q(dbg_0a[0]) );
  SDFFQX1 c_buf_reg_9__6_ ( .D(N557), .SIN(dbg_09[5]), .SMC(test_se), .C(
        net11921), .Q(dbg_09[6]) );
  SDFFQX1 c_buf_reg_9__5_ ( .D(N556), .SIN(dbg_09[4]), .SMC(test_se), .C(
        net11921), .Q(dbg_09[5]) );
  SDFFQX1 c_buf_reg_9__4_ ( .D(N555), .SIN(dbg_09[3]), .SMC(test_se), .C(
        net11921), .Q(dbg_09[4]) );
  SDFFQX1 c_buf_reg_9__3_ ( .D(N554), .SIN(dbg_09[2]), .SMC(test_se), .C(
        net11921), .Q(dbg_09[3]) );
  SDFFQX1 c_buf_reg_9__2_ ( .D(N553), .SIN(dbg_09[1]), .SMC(test_se), .C(
        net11921), .Q(dbg_09[2]) );
  SDFFQX1 c_buf_reg_9__0_ ( .D(N551), .SIN(dbg_08[7]), .SMC(test_se), .C(
        net11921), .Q(dbg_09[0]) );
  SDFFQX1 c_buf_reg_8__6_ ( .D(N549), .SIN(dbg_08[5]), .SMC(test_se), .C(
        net11926), .Q(dbg_08[6]) );
  SDFFQX1 c_buf_reg_8__5_ ( .D(N548), .SIN(dbg_08[4]), .SMC(test_se), .C(
        net11926), .Q(dbg_08[5]) );
  SDFFQX1 c_buf_reg_8__4_ ( .D(N547), .SIN(dbg_08[3]), .SMC(test_se), .C(
        net11926), .Q(dbg_08[4]) );
  SDFFQX1 c_buf_reg_8__3_ ( .D(N546), .SIN(dbg_08[2]), .SMC(test_se), .C(
        net11926), .Q(dbg_08[3]) );
  SDFFQX1 c_buf_reg_8__2_ ( .D(N545), .SIN(dbg_08[1]), .SMC(test_se), .C(
        net11926), .Q(dbg_08[2]) );
  SDFFQX1 c_buf_reg_7__6_ ( .D(N541), .SIN(dbg_07[5]), .SMC(test_se), .C(
        net11931), .Q(dbg_07[6]) );
  SDFFQX1 c_buf_reg_7__5_ ( .D(N540), .SIN(dbg_07[4]), .SMC(test_se), .C(
        net11931), .Q(dbg_07[5]) );
  SDFFQX1 c_buf_reg_7__4_ ( .D(N539), .SIN(dbg_07[3]), .SMC(test_se), .C(
        net11931), .Q(dbg_07[4]) );
  SDFFQX1 c_buf_reg_7__3_ ( .D(N538), .SIN(dbg_07[2]), .SMC(test_se), .C(
        net11931), .Q(dbg_07[3]) );
  SDFFQX1 c_buf_reg_7__2_ ( .D(N537), .SIN(dbg_07[1]), .SMC(test_se), .C(
        net11931), .Q(dbg_07[2]) );
  SDFFQX1 c_buf_reg_11__6_ ( .D(N573), .SIN(dbg_0b[5]), .SMC(test_se), .C(
        net11911), .Q(dbg_0b[6]) );
  SDFFQX1 c_buf_reg_11__5_ ( .D(N572), .SIN(dbg_0b[4]), .SMC(test_se), .C(
        net11911), .Q(dbg_0b[5]) );
  SDFFQX1 c_buf_reg_11__4_ ( .D(N571), .SIN(dbg_0b[3]), .SMC(test_se), .C(
        net11911), .Q(dbg_0b[4]) );
  SDFFQX1 c_buf_reg_11__3_ ( .D(N570), .SIN(dbg_0b[2]), .SMC(test_se), .C(
        net11911), .Q(dbg_0b[3]) );
  SDFFQX1 c_buf_reg_11__2_ ( .D(N569), .SIN(dbg_0b[1]), .SMC(test_se), .C(
        net11911), .Q(dbg_0b[2]) );
  SDFFQX1 c_buf_reg_11__0_ ( .D(N567), .SIN(dbg_0a[7]), .SMC(test_se), .C(
        net11911), .Q(dbg_0b[0]) );
  SDFFQX1 c_buf_reg_0__0_ ( .D(N479), .SIN(c_adr[14]), .SMC(test_se), .C(
        net11966), .Q(rd_buf[0]) );
  SDFFQX1 c_buf_reg_0__6_ ( .D(N485), .SIN(rd_buf[5]), .SMC(test_se), .C(
        net11966), .Q(rd_buf[6]) );
  SDFFQX1 c_buf_reg_0__5_ ( .D(N484), .SIN(rd_buf[4]), .SMC(test_se), .C(
        net11966), .Q(rd_buf[5]) );
  SDFFQX1 c_buf_reg_0__3_ ( .D(N482), .SIN(rd_buf[2]), .SMC(test_se), .C(
        net11966), .Q(rd_buf[3]) );
  SDFFQX1 c_buf_reg_3__4_ ( .D(N507), .SIN(dbg_03[3]), .SMC(test_se), .C(
        net11951), .Q(dbg_03[4]) );
  SDFFQX1 c_buf_reg_5__5_ ( .D(N524), .SIN(dbg_05[4]), .SMC(test_se), .C(
        net11941), .Q(dbg_05[5]) );
  SDFFQX1 c_buf_reg_2__5_ ( .D(N500), .SIN(dbg_02[4]), .SMC(test_se), .C(
        net11956), .Q(dbg_02[5]) );
  SDFFQX1 c_buf_reg_2__4_ ( .D(N499), .SIN(dbg_02[3]), .SMC(test_se), .C(
        net11956), .Q(dbg_02[4]) );
  SDFFQX1 c_buf_reg_3__5_ ( .D(N508), .SIN(dbg_03[4]), .SMC(test_se), .C(
        net11951), .Q(dbg_03[5]) );
  SDFFQX1 c_buf_reg_4__5_ ( .D(N516), .SIN(dbg_04[4]), .SMC(test_se), .C(
        net11946), .Q(dbg_04[5]) );
  SDFFQX1 c_buf_reg_1__5_ ( .D(N492), .SIN(dbg_01[4]), .SMC(test_se), .C(
        net11961), .Q(dbg_01[5]) );
  SDFFQX1 c_buf_reg_4__4_ ( .D(N515), .SIN(dbg_04[3]), .SMC(test_se), .C(
        net11946), .Q(dbg_04[4]) );
  SDFFQX1 c_buf_reg_1__4_ ( .D(N491), .SIN(dbg_01[3]), .SMC(test_se), .C(
        net11961), .Q(dbg_01[4]) );
  SDFFQX1 c_buf_reg_4__3_ ( .D(N514), .SIN(dbg_04[2]), .SMC(test_se), .C(
        net11946), .Q(dbg_04[3]) );
  SDFFQX1 c_buf_reg_8__0_ ( .D(N543), .SIN(dbg_07[7]), .SMC(test_se), .C(
        net11926), .Q(dbg_08[0]) );
  SDFFQX1 c_buf_reg_0__4_ ( .D(N483), .SIN(rd_buf[3]), .SMC(test_se), .C(
        net11966), .Q(rd_buf[4]) );
  SDFFQX1 c_buf_reg_6__2_ ( .D(N529), .SIN(dbg_06[1]), .SMC(test_se), .C(
        net11936), .Q(dbg_06[2]) );
  SDFFQX1 adr_p_reg_14_ ( .D(N868), .SIN(adr_p[13]), .SMC(test_se), .C(
        net11846), .Q(adr_p[14]) );
  SDFFQX1 c_buf_reg_0__2_ ( .D(N481), .SIN(rd_buf[1]), .SMC(test_se), .C(
        net11966), .Q(rd_buf[2]) );
  SDFFQX1 c_buf_reg_0__1_ ( .D(N480), .SIN(rd_buf[0]), .SMC(test_se), .C(
        net11966), .Q(rd_buf[1]) );
  SDFFQX1 c_buf_reg_5__6_ ( .D(N525), .SIN(dbg_05[5]), .SMC(test_se), .C(
        net11941), .Q(dbg_05[6]) );
  SDFFQX1 c_buf_reg_2__6_ ( .D(N501), .SIN(dbg_02[5]), .SMC(test_se), .C(
        net11956), .Q(dbg_02[6]) );
  SDFFQX1 c_buf_reg_5__4_ ( .D(N523), .SIN(dbg_05[3]), .SMC(test_se), .C(
        net11941), .Q(dbg_05[4]) );
  SDFFQX1 c_buf_reg_5__3_ ( .D(N522), .SIN(dbg_05[2]), .SMC(test_se), .C(
        net11941), .Q(dbg_05[3]) );
  SDFFQX1 c_buf_reg_2__3_ ( .D(N498), .SIN(dbg_02[2]), .SMC(test_se), .C(
        net11956), .Q(dbg_02[3]) );
  SDFFQX1 c_buf_reg_5__2_ ( .D(N521), .SIN(dbg_05[1]), .SMC(test_se), .C(
        net11941), .Q(dbg_05[2]) );
  SDFFQX1 c_buf_reg_2__2_ ( .D(N497), .SIN(dbg_02[1]), .SMC(test_se), .C(
        net11956), .Q(dbg_02[2]) );
  SDFFQX1 c_buf_reg_5__1_ ( .D(N520), .SIN(dbg_05[0]), .SMC(test_se), .C(
        net11941), .Q(dbg_05[1]) );
  SDFFQX1 c_buf_reg_2__1_ ( .D(N496), .SIN(dbg_02[0]), .SMC(test_se), .C(
        net11956), .Q(dbg_02[1]) );
  SDFFQX1 c_buf_reg_3__6_ ( .D(N509), .SIN(dbg_03[5]), .SMC(test_se), .C(
        net11951), .Q(dbg_03[6]) );
  SDFFQX1 c_buf_reg_3__3_ ( .D(N506), .SIN(dbg_03[2]), .SMC(test_se), .C(
        net11951), .Q(dbg_03[3]) );
  SDFFQX1 c_buf_reg_3__2_ ( .D(N505), .SIN(dbg_03[1]), .SMC(test_se), .C(
        net11951), .Q(dbg_03[2]) );
  SDFFQX1 c_buf_reg_3__1_ ( .D(N504), .SIN(dbg_03[0]), .SMC(test_se), .C(
        net11951), .Q(dbg_03[1]) );
  SDFFQX1 c_buf_reg_4__6_ ( .D(N517), .SIN(dbg_04[5]), .SMC(test_se), .C(
        net11946), .Q(dbg_04[6]) );
  SDFFQX1 c_buf_reg_1__6_ ( .D(N493), .SIN(dbg_01[5]), .SMC(test_se), .C(
        net11961), .Q(dbg_01[6]) );
  SDFFQX1 c_buf_reg_1__3_ ( .D(N490), .SIN(dbg_01[2]), .SMC(test_se), .C(
        net11961), .Q(dbg_01[3]) );
  SDFFQX1 c_buf_reg_4__2_ ( .D(N513), .SIN(dbg_04[1]), .SMC(test_se), .C(
        net11946), .Q(dbg_04[2]) );
  SDFFQX1 c_buf_reg_1__2_ ( .D(N489), .SIN(dbg_01[1]), .SMC(test_se), .C(
        net11961), .Q(dbg_01[2]) );
  SDFFQX1 c_buf_reg_4__1_ ( .D(N512), .SIN(dbg_04[0]), .SMC(test_se), .C(
        net11946), .Q(dbg_04[1]) );
  SDFFQX1 c_buf_reg_1__1_ ( .D(N488), .SIN(dbg_01[0]), .SMC(test_se), .C(
        net11961), .Q(dbg_01[1]) );
  SDFFQX1 c_buf_reg_10__1_ ( .D(N560), .SIN(dbg_0a[0]), .SMC(test_se), .C(
        net11916), .Q(dbg_0a[1]) );
  SDFFQX1 c_buf_reg_6__1_ ( .D(N528), .SIN(dbg_06[0]), .SMC(test_se), .C(
        net11936), .Q(dbg_06[1]) );
  SDFFQX1 c_buf_reg_9__1_ ( .D(N552), .SIN(dbg_09[0]), .SMC(test_se), .C(
        net11921), .Q(dbg_09[1]) );
  SDFFQX1 c_buf_reg_8__1_ ( .D(N544), .SIN(dbg_08[0]), .SMC(test_se), .C(
        net11926), .Q(dbg_08[1]) );
  SDFFQX1 c_buf_reg_7__1_ ( .D(N536), .SIN(dbg_07[0]), .SMC(test_se), .C(
        net11931), .Q(dbg_07[1]) );
  SDFFQX1 c_buf_reg_15__4_ ( .D(N603), .SIN(dbg_0f[3]), .SMC(test_se), .C(
        net11891), .Q(dbg_0f[4]) );
  SDFFQX1 c_buf_reg_14__4_ ( .D(N595), .SIN(dbg_0e[3]), .SMC(test_se), .C(
        net11896), .Q(dbg_0e[4]) );
  SDFFQX1 c_buf_reg_13__4_ ( .D(N587), .SIN(dbg_0d[3]), .SMC(test_se), .C(
        net11901), .Q(dbg_0d[4]) );
  SDFFQX1 c_buf_reg_12__4_ ( .D(N579), .SIN(dbg_0c[3]), .SMC(test_se), .C(
        net11906), .Q(dbg_0c[4]) );
  SDFFQX1 c_buf_reg_11__1_ ( .D(N568), .SIN(dbg_0b[0]), .SMC(test_se), .C(
        net11911), .Q(dbg_0b[1]) );
  SDFFQX1 c_buf_reg_22__6_ ( .D(N661), .SIN(c_buf_22__5_), .SMC(test_se), .C(
        net11856), .Q(c_buf_22__6_) );
  SDFFQX1 c_buf_reg_22__5_ ( .D(N660), .SIN(c_buf_22__4_), .SMC(test_se), .C(
        net11856), .Q(c_buf_22__5_) );
  SDFFQX1 c_buf_reg_22__4_ ( .D(N659), .SIN(c_buf_22__3_), .SMC(test_se), .C(
        net11856), .Q(c_buf_22__4_) );
  SDFFQX1 c_buf_reg_22__3_ ( .D(N658), .SIN(c_buf_22__2_), .SMC(test_se), .C(
        net11856), .Q(c_buf_22__3_) );
  SDFFQX1 c_buf_reg_22__2_ ( .D(N657), .SIN(c_buf_22__1_), .SMC(test_se), .C(
        net11856), .Q(c_buf_22__2_) );
  SDFFQX1 c_buf_reg_21__6_ ( .D(N653), .SIN(c_buf_21__5_), .SMC(test_se), .C(
        net11861), .Q(c_buf_21__6_) );
  SDFFQX1 c_buf_reg_21__5_ ( .D(N652), .SIN(c_buf_21__4_), .SMC(test_se), .C(
        net11861), .Q(c_buf_21__5_) );
  SDFFQX1 c_buf_reg_21__4_ ( .D(N651), .SIN(c_buf_21__3_), .SMC(test_se), .C(
        net11861), .Q(c_buf_21__4_) );
  SDFFQX1 c_buf_reg_21__3_ ( .D(N650), .SIN(c_buf_21__2_), .SMC(test_se), .C(
        net11861), .Q(c_buf_21__3_) );
  SDFFQX1 c_buf_reg_21__2_ ( .D(N649), .SIN(c_buf_21__1_), .SMC(test_se), .C(
        net11861), .Q(c_buf_21__2_) );
  SDFFQX1 c_buf_reg_20__6_ ( .D(N645), .SIN(c_buf_20__5_), .SMC(test_se), .C(
        net11866), .Q(c_buf_20__6_) );
  SDFFQX1 c_buf_reg_20__5_ ( .D(N644), .SIN(c_buf_20__4_), .SMC(test_se), .C(
        net11866), .Q(c_buf_20__5_) );
  SDFFQX1 c_buf_reg_20__4_ ( .D(N643), .SIN(c_buf_20__3_), .SMC(test_se), .C(
        net11866), .Q(c_buf_20__4_) );
  SDFFQX1 c_buf_reg_20__3_ ( .D(N642), .SIN(c_buf_20__2_), .SMC(test_se), .C(
        net11866), .Q(c_buf_20__3_) );
  SDFFQX1 c_buf_reg_20__2_ ( .D(N641), .SIN(c_buf_20__1_), .SMC(test_se), .C(
        net11866), .Q(c_buf_20__2_) );
  SDFFQX1 c_buf_reg_19__6_ ( .D(N637), .SIN(c_buf_19__5_), .SMC(test_se), .C(
        net11871), .Q(c_buf_19__6_) );
  SDFFQX1 c_buf_reg_19__5_ ( .D(N636), .SIN(c_buf_19__4_), .SMC(test_se), .C(
        net11871), .Q(c_buf_19__5_) );
  SDFFQX1 c_buf_reg_19__4_ ( .D(N635), .SIN(c_buf_19__3_), .SMC(test_se), .C(
        net11871), .Q(c_buf_19__4_) );
  SDFFQX1 c_buf_reg_19__3_ ( .D(N634), .SIN(c_buf_19__2_), .SMC(test_se), .C(
        net11871), .Q(c_buf_19__3_) );
  SDFFQX1 c_buf_reg_18__5_ ( .D(N628), .SIN(c_buf_18__4_), .SMC(test_se), .C(
        net11876), .Q(c_buf_18__5_) );
  SDFFQX1 c_buf_reg_18__4_ ( .D(N627), .SIN(c_buf_18__3_), .SMC(test_se), .C(
        net11876), .Q(c_buf_18__4_) );
  SDFFQX1 c_buf_reg_18__3_ ( .D(N626), .SIN(c_buf_18__2_), .SMC(test_se), .C(
        net11876), .Q(c_buf_18__3_) );
  SDFFQX1 c_buf_reg_17__6_ ( .D(N621), .SIN(c_buf_17__5_), .SMC(test_se), .C(
        net11881), .Q(c_buf_17__6_) );
  SDFFQX1 c_buf_reg_17__5_ ( .D(N620), .SIN(c_buf_17__4_), .SMC(test_se), .C(
        net11881), .Q(c_buf_17__5_) );
  SDFFQX1 c_buf_reg_17__4_ ( .D(N619), .SIN(c_buf_17__3_), .SMC(test_se), .C(
        net11881), .Q(c_buf_17__4_) );
  SDFFQX1 c_buf_reg_17__3_ ( .D(N618), .SIN(c_buf_17__2_), .SMC(test_se), .C(
        net11881), .Q(c_buf_17__3_) );
  SDFFQX1 c_buf_reg_16__5_ ( .D(N612), .SIN(c_buf_16__4_), .SMC(test_se), .C(
        net11886), .Q(c_buf_16__5_) );
  SDFFQX1 c_buf_reg_16__4_ ( .D(N611), .SIN(c_buf_16__3_), .SMC(test_se), .C(
        net11886), .Q(c_buf_16__4_) );
  SDFFQX1 c_buf_reg_16__3_ ( .D(N610), .SIN(c_buf_16__2_), .SMC(test_se), .C(
        net11886), .Q(c_buf_16__3_) );
  SDFFQX1 c_buf_reg_15__5_ ( .D(N604), .SIN(dbg_0f[4]), .SMC(test_se), .C(
        net11891), .Q(dbg_0f[5]) );
  SDFFQX1 c_buf_reg_14__6_ ( .D(N597), .SIN(dbg_0e[5]), .SMC(test_se), .C(
        net11896), .Q(dbg_0e[6]) );
  SDFFQX1 c_buf_reg_14__5_ ( .D(N596), .SIN(dbg_0e[4]), .SMC(test_se), .C(
        net11896), .Q(dbg_0e[5]) );
  SDFFQX1 c_buf_reg_14__3_ ( .D(N594), .SIN(dbg_0e[2]), .SMC(test_se), .C(
        net11896), .Q(dbg_0e[3]) );
  SDFFQX1 c_buf_reg_13__5_ ( .D(N588), .SIN(dbg_0d[4]), .SMC(test_se), .C(
        net11901), .Q(dbg_0d[5]) );
  SDFFQX1 c_buf_reg_12__5_ ( .D(N580), .SIN(dbg_0c[4]), .SMC(test_se), .C(
        net11906), .Q(dbg_0c[5]) );
  SDFFQX1 c_buf_reg_23__4_ ( .D(N790), .SIN(wr_buf[3]), .SMC(test_se), .C(
        net11851), .Q(wr_buf[4]) );
  SDFFQX1 c_buf_reg_23__6_ ( .D(N792), .SIN(wr_buf[5]), .SMC(test_se), .C(
        net11851), .Q(wr_buf[6]) );
  SDFFQX1 c_buf_reg_23__2_ ( .D(N788), .SIN(wr_buf[1]), .SMC(test_se), .C(
        net11851), .Q(wr_buf[2]) );
  SDFFQX1 c_buf_reg_23__3_ ( .D(N789), .SIN(wr_buf[2]), .SMC(test_se), .C(
        net11851), .Q(wr_buf[3]) );
  SDFFQX1 c_buf_reg_23__5_ ( .D(N791), .SIN(wr_buf[4]), .SMC(test_se), .C(
        net11851), .Q(wr_buf[5]) );
  SDFFQX1 c_buf_reg_23__0_ ( .D(N786), .SIN(c_buf_22__7_), .SMC(test_se), .C(
        net11851), .Q(wr_buf[0]) );
  SDFFQX1 c_buf_reg_10__7_ ( .D(N566), .SIN(dbg_0a[6]), .SMC(test_se), .C(
        net11916), .Q(dbg_0a[7]) );
  SDFFQX1 c_buf_reg_9__7_ ( .D(N558), .SIN(dbg_09[6]), .SMC(test_se), .C(
        net11921), .Q(dbg_09[7]) );
  SDFFQX1 c_buf_reg_8__7_ ( .D(N550), .SIN(dbg_08[6]), .SMC(test_se), .C(
        net11926), .Q(dbg_08[7]) );
  SDFFQX1 c_buf_reg_7__7_ ( .D(N542), .SIN(dbg_07[6]), .SMC(test_se), .C(
        net11931), .Q(dbg_07[7]) );
  SDFFQX1 c_buf_reg_11__7_ ( .D(N574), .SIN(dbg_0b[6]), .SMC(test_se), .C(
        net11911), .Q(dbg_0b[7]) );
  SDFFQX1 r_twlb_reg_1_ ( .D(n645), .SIN(pmem_twlb[0]), .SMC(test_se), .C(clk), 
        .Q(pmem_twlb[1]) );
  SDFFQX1 r_twlb_reg_0_ ( .D(n646), .SIN(r_rdy), .SMC(test_se), .C(clk), .Q(
        pmem_twlb[0]) );
  SDFFQX1 c_buf_reg_22__1_ ( .D(N656), .SIN(c_buf_22__0_), .SMC(test_se), .C(
        net11856), .Q(c_buf_22__1_) );
  SDFFQX1 c_buf_reg_22__0_ ( .D(N655), .SIN(c_buf_21__7_), .SMC(test_se), .C(
        net11856), .Q(c_buf_22__0_) );
  SDFFQX1 c_buf_reg_21__1_ ( .D(N648), .SIN(c_buf_21__0_), .SMC(test_se), .C(
        net11861), .Q(c_buf_21__1_) );
  SDFFQX1 c_buf_reg_21__0_ ( .D(N647), .SIN(c_buf_20__7_), .SMC(test_se), .C(
        net11861), .Q(c_buf_21__0_) );
  SDFFQX1 c_buf_reg_20__1_ ( .D(N640), .SIN(c_buf_20__0_), .SMC(test_se), .C(
        net11866), .Q(c_buf_20__1_) );
  SDFFQX1 c_buf_reg_20__0_ ( .D(N639), .SIN(c_buf_19__7_), .SMC(test_se), .C(
        net11866), .Q(c_buf_20__0_) );
  SDFFQX1 c_buf_reg_19__2_ ( .D(N633), .SIN(c_buf_19__1_), .SMC(test_se), .C(
        net11871), .Q(c_buf_19__2_) );
  SDFFQX1 c_buf_reg_19__1_ ( .D(N632), .SIN(c_buf_19__0_), .SMC(test_se), .C(
        net11871), .Q(c_buf_19__1_) );
  SDFFQX1 c_buf_reg_19__0_ ( .D(N631), .SIN(c_buf_18__7_), .SMC(test_se), .C(
        net11871), .Q(c_buf_19__0_) );
  SDFFQX1 c_buf_reg_18__6_ ( .D(N629), .SIN(c_buf_18__5_), .SMC(test_se), .C(
        net11876), .Q(c_buf_18__6_) );
  SDFFQX1 c_buf_reg_18__2_ ( .D(N625), .SIN(c_buf_18__1_), .SMC(test_se), .C(
        net11876), .Q(c_buf_18__2_) );
  SDFFQX1 c_buf_reg_18__1_ ( .D(N624), .SIN(c_buf_18__0_), .SMC(test_se), .C(
        net11876), .Q(c_buf_18__1_) );
  SDFFQX1 c_buf_reg_18__0_ ( .D(N623), .SIN(c_buf_17__7_), .SMC(test_se), .C(
        net11876), .Q(c_buf_18__0_) );
  SDFFQX1 c_buf_reg_17__2_ ( .D(N617), .SIN(c_buf_17__1_), .SMC(test_se), .C(
        net11881), .Q(c_buf_17__2_) );
  SDFFQX1 c_buf_reg_17__1_ ( .D(N616), .SIN(c_buf_17__0_), .SMC(test_se), .C(
        net11881), .Q(c_buf_17__1_) );
  SDFFQX1 c_buf_reg_17__0_ ( .D(N615), .SIN(c_buf_16__7_), .SMC(test_se), .C(
        net11881), .Q(c_buf_17__0_) );
  SDFFQX1 c_buf_reg_16__6_ ( .D(N613), .SIN(c_buf_16__5_), .SMC(test_se), .C(
        net11886), .Q(c_buf_16__6_) );
  SDFFQX1 c_buf_reg_16__2_ ( .D(N609), .SIN(c_buf_16__1_), .SMC(test_se), .C(
        net11886), .Q(c_buf_16__2_) );
  SDFFQX1 c_buf_reg_16__1_ ( .D(N608), .SIN(c_buf_16__0_), .SMC(test_se), .C(
        net11886), .Q(c_buf_16__1_) );
  SDFFQX1 c_buf_reg_16__0_ ( .D(N607), .SIN(dbg_0f[7]), .SMC(test_se), .C(
        net11886), .Q(c_buf_16__0_) );
  SDFFQX1 c_buf_reg_15__6_ ( .D(N605), .SIN(dbg_0f[5]), .SMC(test_se), .C(
        net11891), .Q(dbg_0f[6]) );
  SDFFQX1 c_buf_reg_15__3_ ( .D(N602), .SIN(dbg_0f[2]), .SMC(test_se), .C(
        net11891), .Q(dbg_0f[3]) );
  SDFFQX1 c_buf_reg_15__2_ ( .D(N601), .SIN(dbg_0f[1]), .SMC(test_se), .C(
        net11891), .Q(dbg_0f[2]) );
  SDFFQX1 c_buf_reg_15__1_ ( .D(N600), .SIN(dbg_0f[0]), .SMC(test_se), .C(
        net11891), .Q(dbg_0f[1]) );
  SDFFQX1 c_buf_reg_15__0_ ( .D(N599), .SIN(dbg_0e[7]), .SMC(test_se), .C(
        net11891), .Q(dbg_0f[0]) );
  SDFFQX1 c_buf_reg_14__2_ ( .D(N593), .SIN(dbg_0e[1]), .SMC(test_se), .C(
        net11896), .Q(dbg_0e[2]) );
  SDFFQX1 c_buf_reg_14__1_ ( .D(N592), .SIN(dbg_0e[0]), .SMC(test_se), .C(
        net11896), .Q(dbg_0e[1]) );
  SDFFQX1 c_buf_reg_14__0_ ( .D(N591), .SIN(dbg_0d[7]), .SMC(test_se), .C(
        net11896), .Q(dbg_0e[0]) );
  SDFFQX1 c_buf_reg_13__6_ ( .D(N589), .SIN(dbg_0d[5]), .SMC(test_se), .C(
        net11901), .Q(dbg_0d[6]) );
  SDFFQX1 c_buf_reg_13__3_ ( .D(N586), .SIN(dbg_0d[2]), .SMC(test_se), .C(
        net11901), .Q(dbg_0d[3]) );
  SDFFQX1 c_buf_reg_13__2_ ( .D(N585), .SIN(dbg_0d[1]), .SMC(test_se), .C(
        net11901), .Q(dbg_0d[2]) );
  SDFFQX1 c_buf_reg_13__1_ ( .D(N584), .SIN(dbg_0d[0]), .SMC(test_se), .C(
        net11901), .Q(dbg_0d[1]) );
  SDFFQX1 c_buf_reg_13__0_ ( .D(N583), .SIN(dbg_0c[7]), .SMC(test_se), .C(
        net11901), .Q(dbg_0d[0]) );
  SDFFQX1 c_buf_reg_12__6_ ( .D(N581), .SIN(dbg_0c[5]), .SMC(test_se), .C(
        net11906), .Q(dbg_0c[6]) );
  SDFFQX1 c_buf_reg_12__3_ ( .D(N578), .SIN(dbg_0c[2]), .SMC(test_se), .C(
        net11906), .Q(dbg_0c[3]) );
  SDFFQX1 c_buf_reg_12__2_ ( .D(N577), .SIN(dbg_0c[1]), .SMC(test_se), .C(
        net11906), .Q(dbg_0c[2]) );
  SDFFQX1 c_buf_reg_12__1_ ( .D(N576), .SIN(dbg_0c[0]), .SMC(test_se), .C(
        net11906), .Q(dbg_0c[1]) );
  SDFFQX1 c_buf_reg_12__0_ ( .D(N575), .SIN(dbg_0b[7]), .SMC(test_se), .C(
        net11906), .Q(dbg_0c[0]) );
  SDFFQX1 c_buf_reg_23__1_ ( .D(N787), .SIN(wr_buf[0]), .SMC(test_se), .C(
        net11851), .Q(wr_buf[1]) );
  SDFFQX1 adr_p_reg_13_ ( .D(N867), .SIN(pmem_a[14]), .SMC(test_se), .C(
        net11846), .Q(adr_p[13]) );
  SDFFQX1 wspp_cnt_reg_4_ ( .D(N799), .SIN(wspp_cnt_3_), .SMC(test_se), .C(
        net11835), .Q(wspp_cnt_4_) );
  SDFFQX2 adr_p_reg_6_ ( .D(N860), .SIN(pmem_a[5]), .SMC(test_se), .C(net11846), .Q(pmem_a[9]) );
  SDFFQX1 c_buf_reg_6__7_ ( .D(N534), .SIN(dbg_06[6]), .SMC(test_se), .C(
        net11936), .Q(dbg_06[7]) );
  SDFFQX1 wspp_cnt_reg_5_ ( .D(N800), .SIN(wspp_cnt_4_), .SMC(test_se), .C(
        net11835), .Q(wspp_cnt_5_) );
  SDFFQX1 wspp_cnt_reg_3_ ( .D(N798), .SIN(wspp_cnt_2_), .SMC(test_se), .C(
        net11835), .Q(wspp_cnt_3_) );
  SDFFQX1 wspp_cnt_reg_6_ ( .D(N801), .SIN(wspp_cnt_5_), .SMC(test_se), .C(
        net11835), .Q(test_so2) );
  SDFFQX1 c_buf_reg_0__7_ ( .D(N486), .SIN(rd_buf[6]), .SMC(test_se), .C(
        net11966), .Q(rd_buf[7]) );
  SDFFQX1 c_buf_reg_5__7_ ( .D(N526), .SIN(dbg_05[6]), .SMC(test_se), .C(
        net11941), .Q(dbg_05[7]) );
  SDFFQX1 c_buf_reg_2__7_ ( .D(N502), .SIN(dbg_02[6]), .SMC(test_se), .C(
        net11956), .Q(dbg_02[7]) );
  SDFFQX1 c_buf_reg_3__7_ ( .D(N510), .SIN(dbg_03[6]), .SMC(test_se), .C(
        net11951), .Q(dbg_03[7]) );
  SDFFQX1 c_buf_reg_4__7_ ( .D(N518), .SIN(dbg_04[6]), .SMC(test_se), .C(
        net11946), .Q(dbg_04[7]) );
  SDFFQX1 c_buf_reg_1__7_ ( .D(N494), .SIN(dbg_01[6]), .SMC(test_se), .C(
        net11961), .Q(dbg_01[7]) );
  SDFFQX1 c_buf_reg_22__7_ ( .D(N662), .SIN(c_buf_22__6_), .SMC(test_se), .C(
        net11856), .Q(c_buf_22__7_) );
  SDFFQX1 c_buf_reg_21__7_ ( .D(N654), .SIN(c_buf_21__6_), .SMC(test_se), .C(
        net11861), .Q(c_buf_21__7_) );
  SDFFQX1 c_buf_reg_20__7_ ( .D(N646), .SIN(c_buf_20__6_), .SMC(test_se), .C(
        net11866), .Q(c_buf_20__7_) );
  SDFFQX1 c_buf_reg_19__7_ ( .D(N638), .SIN(c_buf_19__6_), .SMC(test_se), .C(
        net11871), .Q(c_buf_19__7_) );
  SDFFQX1 c_buf_reg_18__7_ ( .D(N630), .SIN(c_buf_18__6_), .SMC(test_se), .C(
        net11876), .Q(c_buf_18__7_) );
  SDFFQX1 c_buf_reg_17__7_ ( .D(N622), .SIN(c_buf_17__6_), .SMC(test_se), .C(
        net11881), .Q(c_buf_17__7_) );
  SDFFQX1 c_buf_reg_16__7_ ( .D(N614), .SIN(c_buf_16__6_), .SMC(test_se), .C(
        net11886), .Q(c_buf_16__7_) );
  SDFFQX1 c_buf_reg_15__7_ ( .D(N606), .SIN(dbg_0f[6]), .SMC(test_se), .C(
        net11891), .Q(dbg_0f[7]) );
  SDFFQX1 c_buf_reg_14__7_ ( .D(N598), .SIN(dbg_0e[6]), .SMC(test_se), .C(
        net11896), .Q(dbg_0e[7]) );
  SDFFQX1 c_buf_reg_13__7_ ( .D(N590), .SIN(dbg_0d[6]), .SMC(test_se), .C(
        net11901), .Q(dbg_0d[7]) );
  SDFFQX1 c_buf_reg_12__7_ ( .D(N582), .SIN(dbg_0c[6]), .SMC(test_se), .C(
        net11906), .Q(dbg_0c[7]) );
  SDFFQX1 c_buf_reg_23__7_ ( .D(N793), .SIN(wr_buf[6]), .SMC(test_se), .C(
        net11851), .Q(wr_buf[7]) );
  SDFFQX2 adr_p_reg_7_ ( .D(N861), .SIN(pmem_a[9]), .SMC(test_se), .C(net11846), .Q(pmem_a[10]) );
  SDFFQX2 adr_p_reg_9_ ( .D(N863), .SIN(pmem_a[11]), .SMC(test_se), .C(
        net11846), .Q(pmem_a[12]) );
  SDFFQX2 adr_p_reg_11_ ( .D(N865), .SIN(pmem_a[13]), .SMC(test_se), .C(
        net11846), .Q(pmem_a[14]) );
  SDFFQX1 c_adr_reg_3_ ( .D(N829), .SIN(c_adr[2]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[3]) );
  SDFFQX1 cs_ft_reg_2_ ( .D(N823), .SIN(cs_ft[1]), .SMC(test_se), .C(net11981), 
        .Q(cs_ft[2]) );
  SDFFQX1 c_adr_reg_4_ ( .D(N830), .SIN(c_adr[3]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[4]) );
  SDFFNQX1 cs_n_reg ( .D(n643), .SIN(pmem_clk[1]), .SMC(test_se), .XC(clk), 
        .Q(test_so1) );
  SDFFQX1 re_p_reg ( .D(n647), .SIN(pmem_twlb[1]), .SMC(test_se), .C(clk), .Q(
        pmem_re) );
  SDFFQX1 c_adr_reg_2_ ( .D(N828), .SIN(c_adr[1]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[2]) );
  SDFFQX1 cs_ft_reg_3_ ( .D(N824), .SIN(cs_ft[2]), .SMC(test_se), .C(net11981), 
        .Q(cs_ft[3]) );
  SDFFQX1 cs_ft_reg_1_ ( .D(N822), .SIN(cs_ft[0]), .SMC(test_se), .C(net11981), 
        .Q(cs_ft[1]) );
  SDFFQX1 cs_ft_reg_0_ ( .D(N821), .SIN(c_ptr[4]), .SMC(test_se), .C(net11981), 
        .Q(cs_ft[0]) );
  SDFFQX1 c_adr_reg_1_ ( .D(N827), .SIN(c_adr[0]), .SMC(test_se), .C(net11976), 
        .Q(c_adr[1]) );
  SDFFQX1 c_adr_reg_0_ ( .D(N826), .SIN(adr_p[14]), .SMC(test_se), .C(net11976), .Q(c_adr[0]) );
  SDFFQX1 un_hold_reg ( .D(n762), .SIN(pmem_re), .SMC(test_se), .C(clk), .Q(
        un_hold) );
  SDFFQX1 r_rdy_reg ( .D(n648), .SIN(pmem_pgm), .SMC(test_se), .C(clk), .Q(
        r_rdy) );
  SDFFQX1 pgm_p_reg ( .D(n644), .SIN(dummy[1]), .SMC(test_se), .C(net11981), 
        .Q(pmem_pgm) );
  SDFFQX2 adr_p_reg_0_ ( .D(N854), .SIN(pmem_a[8]), .SMC(test_se), .C(net11846), .Q(pmem_a[0]) );
  SDFFQX2 adr_p_reg_8_ ( .D(N862), .SIN(pmem_a[10]), .SMC(test_se), .C(
        net11846), .Q(pmem_a[11]) );
  SDFFQX2 adr_p_reg_10_ ( .D(N864), .SIN(pmem_a[12]), .SMC(test_se), .C(
        net11846), .Q(pmem_a[13]) );
  SDFFQX2 adr_p_reg_12_ ( .D(N866), .SIN(test_si3), .SMC(test_se), .C(net11846), .Q(pmem_a[15]) );
  SDFFQX2 a_bit_reg_1_ ( .D(n937), .SIN(pmem_a[6]), .SMC(test_se), .C(net11841), .Q(pmem_a[7]) );
  AOI222XL U3 ( .A(n151), .B(n150), .C(n1), .D(n149), .E(n154), .F(n155), .Y(
        n157) );
  AO21X1 U4 ( .B(n239), .C(n231), .A(n230), .Y(n425) );
  AO21X1 U5 ( .B(n568), .C(n567), .A(n566), .Y(n647) );
  NOR21XL U6 ( .B(n103), .A(n35), .Y(n641) );
  OA22X1 U7 ( .A(n151), .B(n150), .C(n144), .D(n130), .Y(n1) );
  AOI21X1 U8 ( .B(n681), .C(n680), .A(n679), .Y(n2) );
  INVXL U9 ( .A(n441), .Y(n3) );
  INVXL U10 ( .A(n3), .Y(n4) );
  INVX1 U11 ( .A(n483), .Y(n5) );
  INVX1 U12 ( .A(n483), .Y(n6) );
  INVX1 U13 ( .A(n439), .Y(n7) );
  INVX1 U14 ( .A(n485), .Y(n8) );
  INVX1 U15 ( .A(n485), .Y(n9) );
  INVX1 U16 ( .A(n440), .Y(n10) );
  INVX1 U17 ( .A(n489), .Y(n11) );
  INVX1 U18 ( .A(n489), .Y(n12) );
  INVX1 U19 ( .A(n436), .Y(n13) );
  INVX1 U20 ( .A(n491), .Y(n14) );
  INVX1 U21 ( .A(n491), .Y(n15) );
  AOI21X1 U22 ( .B(n111), .C(n512), .A(n519), .Y(n611) );
  INVX1 U23 ( .A(n611), .Y(n16) );
  INVX1 U24 ( .A(n611), .Y(n17) );
  INVX1 U25 ( .A(n493), .Y(n18) );
  INVX1 U26 ( .A(n493), .Y(n19) );
  BUFX3 U27 ( .A(n432), .Y(n20) );
  AOI21XL U28 ( .B(memaddr_c[6]), .C(n432), .A(n77), .Y(n49) );
  INVX1 U29 ( .A(n481), .Y(n21) );
  INVX1 U30 ( .A(n481), .Y(n22) );
  INVX1 U31 ( .A(n515), .Y(n23) );
  INVX1 U32 ( .A(n694), .Y(n24) );
  INVX1 U33 ( .A(n617), .Y(n25) );
  INVX1 U34 ( .A(n487), .Y(n26) );
  INVX1 U35 ( .A(n487), .Y(n27) );
  NAND21X1 U36 ( .B(pwrdn_rst), .A(n104), .Y(n77) );
  NAND21X1 U37 ( .B(pwrdn_rst), .A(n104), .Y(n686) );
  INVX1 U38 ( .A(n495), .Y(n28) );
  INVX1 U39 ( .A(n495), .Y(n29) );
  INVX1 U40 ( .A(n617), .Y(n573) );
  INVX1 U41 ( .A(n655), .Y(n99) );
  NOR32XL U42 ( .B(n206), .C(n172), .A(n171), .Y(n174) );
  INVX1 U43 ( .A(n98), .Y(n78) );
  INVX1 U44 ( .A(n504), .Y(n98) );
  NOR3XL U45 ( .A(n431), .B(n684), .C(cs_ft[2]), .Y(n30) );
  AOI21XL U46 ( .B(n687), .C(n688), .A(n77), .Y(n642) );
  GEN2XL U47 ( .D(c_adr[8]), .E(n249), .C(n197), .B(n374), .A(n196), .Y(n199)
         );
  GEN3XL U48 ( .F(c_adr[12]), .G(n205), .E(n204), .D(n228), .C(n203), .B(n240), 
        .A(n202), .Y(n210) );
  OR2X1 U49 ( .A(d_psrd), .B(n535), .Y(n528) );
  INVXL U50 ( .A(n507), .Y(n509) );
  NAND21XL U51 ( .B(n619), .A(n618), .Y(n93) );
  INVXL U52 ( .A(n655), .Y(n100) );
  NAND21XL U53 ( .B(n523), .A(n615), .Y(n432) );
  INVXL U54 ( .A(n504), .Y(n97) );
  NAND31XL U55 ( .C(n167), .A(n1), .B(n43), .Y(n177) );
  INVXL U56 ( .A(n206), .Y(n207) );
  NAND21XL U57 ( .B(n551), .A(n523), .Y(n572) );
  AO21XL U58 ( .B(n625), .C(n635), .A(n99), .Y(N881) );
  INVXL U59 ( .A(memaddr_c[1]), .Y(n148) );
  OAI211XL U60 ( .C(n564), .D(n669), .A(n688), .B(n672), .Y(n600) );
  INVXL U61 ( .A(n564), .Y(n565) );
  NAND21XL U62 ( .B(n632), .A(n494), .Y(n495) );
  NAND21XL U63 ( .B(n632), .A(n486), .Y(n487) );
  NAND21XL U64 ( .B(n632), .A(n480), .Y(n481) );
  NAND21XL U65 ( .B(n632), .A(n492), .Y(n493) );
  NAND21XL U66 ( .B(n632), .A(n490), .Y(n491) );
  NAND21XL U67 ( .B(n632), .A(n488), .Y(n489) );
  NAND21XL U68 ( .B(n632), .A(n484), .Y(n485) );
  NAND21XL U69 ( .B(n632), .A(n482), .Y(n483) );
  AOI211XL U70 ( .C(n525), .D(n629), .A(n508), .B(n507), .Y(N845) );
  AOI211XL U71 ( .C(n658), .D(n638), .A(n505), .B(n507), .Y(N844) );
  AND2XL U72 ( .A(n655), .B(n662), .Y(n656) );
  AOI31XL U73 ( .A(n672), .B(n671), .C(n670), .D(n77), .Y(n643) );
  NAND31XL U74 ( .C(n534), .A(n435), .B(n694), .Y(n571) );
  INVXL U75 ( .A(memaddr_c[4]), .Y(n150) );
  INVXL U76 ( .A(memaddr_c[3]), .Y(n130) );
  OAI21BBXL U77 ( .A(N432), .B(n573), .C(n44), .Y(N827) );
  AOI21XL U78 ( .B(memaddr_c[1]), .C(n432), .A(n101), .Y(n44) );
  OAI21BBXL U79 ( .A(N434), .B(n25), .C(n46), .Y(N829) );
  AOI21XL U80 ( .B(memaddr_c[3]), .C(n20), .A(n101), .Y(n46) );
  OAI21BBXL U81 ( .A(N435), .B(n25), .C(n47), .Y(N830) );
  AOI21XL U82 ( .B(memaddr_c[4]), .C(n20), .A(n101), .Y(n47) );
  OAI21BBXL U83 ( .A(N437), .B(n573), .C(n49), .Y(N832) );
  OAI21BBXL U84 ( .A(N438), .B(n573), .C(n50), .Y(N833) );
  OAI21BBXL U85 ( .A(N439), .B(n573), .C(n51), .Y(N834) );
  OAI21BBXL U86 ( .A(N440), .B(n573), .C(n52), .Y(N835) );
  OAI21BBXL U87 ( .A(N441), .B(n573), .C(n53), .Y(N836) );
  OAI21BBXL U88 ( .A(N442), .B(n573), .C(n54), .Y(N837) );
  OAI21BBXL U89 ( .A(N444), .B(n573), .C(n55), .Y(N839) );
  OAI21BBXL U90 ( .A(N443), .B(n573), .C(n56), .Y(N838) );
  OAI21BBXL U91 ( .A(N433), .B(n25), .C(n45), .Y(N828) );
  OAI21BBXL U92 ( .A(N436), .B(n25), .C(n48), .Y(N831) );
  OA22XL U93 ( .A(memaddr_c[1]), .B(n187), .C(memaddr_c[0]), .D(n740), .Y(n186) );
  AO21XL U94 ( .B(n623), .C(n639), .A(n99), .Y(N874) );
  AO21XL U95 ( .B(n623), .C(n640), .A(n99), .Y(N875) );
  AO21XL U96 ( .B(n623), .C(n654), .A(n99), .Y(N876) );
  AO21XL U97 ( .B(n623), .C(n635), .A(n99), .Y(N877) );
  AO21XL U98 ( .B(n625), .C(n639), .A(n99), .Y(N878) );
  AO21XL U99 ( .B(n625), .C(n640), .A(n99), .Y(N879) );
  AO21XL U100 ( .B(n625), .C(n654), .A(n99), .Y(N880) );
  AO21XL U101 ( .B(n627), .C(n639), .A(n99), .Y(N882) );
  INVXL U102 ( .A(n182), .Y(n184) );
  AND2XL U103 ( .A(memaddr_c[4]), .B(n731), .Y(n183) );
  XOR3XL U104 ( .A(memaddr_c[4]), .B(n66), .C(n389), .Y(n414) );
  XOR3XL U105 ( .A(memaddr_c[1]), .B(n358), .C(n357), .Y(n419) );
  OAI211XL U106 ( .C(n356), .D(n355), .A(n354), .B(n348), .Y(n420) );
  XOR3XL U107 ( .A(memaddr_c[3]), .B(n391), .C(n390), .Y(n392) );
  AND2XL U108 ( .A(n221), .B(n220), .Y(n222) );
  NAND32XL U109 ( .B(memaddr_c[6]), .C(n193), .A(n236), .Y(n194) );
  OA21XL U110 ( .B(n436), .C(n581), .A(n591), .Y(n437) );
  INVXL U111 ( .A(n580), .Y(n436) );
  NAND21XL U112 ( .B(d_psrd), .A(n571), .Y(n620) );
  AO21XL U113 ( .B(n78), .C(wr_buf[0]), .A(n503), .Y(N655) );
  AO21XL U114 ( .B(n78), .C(wr_buf[4]), .A(n499), .Y(N659) );
  AO21XL U115 ( .B(n78), .C(c_buf_22__7_), .A(n496), .Y(N654) );
  AO21XL U116 ( .B(n78), .C(wr_buf[7]), .A(n21), .Y(N662) );
  AO21XL U117 ( .B(n78), .C(wr_buf[1]), .A(n502), .Y(N656) );
  AO21XL U118 ( .B(n78), .C(wr_buf[2]), .A(n501), .Y(N657) );
  AO21XL U119 ( .B(n78), .C(wr_buf[3]), .A(n500), .Y(N658) );
  AO21XL U120 ( .B(n78), .C(wr_buf[5]), .A(n498), .Y(N660) );
  AO21XL U121 ( .B(n78), .C(wr_buf[6]), .A(n497), .Y(N661) );
  OAI21BBXL U122 ( .A(N431), .B(n25), .C(n31), .Y(N826) );
  AOI21XL U123 ( .B(memaddr_c[0]), .C(n20), .A(n101), .Y(n31) );
  OAI21BBXL U124 ( .A(N445), .B(n25), .C(n32), .Y(N840) );
  AOI21XL U125 ( .B(memaddr_c[14]), .C(n20), .A(n101), .Y(n32) );
  OAI21BBX1 U126 ( .A(n597), .B(n596), .C(n33), .Y(n646) );
  MUX2IX1 U127 ( .D0(n595), .D1(pmem_twlb[0]), .S(n36), .Y(n33) );
  OAI21BBX1 U128 ( .A(n593), .B(n596), .C(n34), .Y(n645) );
  MUX2IXL U129 ( .D0(n595), .D1(pmem_twlb[1]), .S(n36), .Y(n34) );
  AOI21X1 U130 ( .B(n2), .C(n693), .A(n692), .Y(n35) );
  OAI211XL U131 ( .C(n24), .D(n618), .A(n617), .B(n616), .Y(N825) );
  AND2XL U132 ( .A(n102), .B(n615), .Y(n616) );
  NOR43XL U133 ( .B(n102), .C(r_rdy), .D(n17), .A(n558), .Y(n548) );
  AND3XL U134 ( .A(n534), .B(cs_ft[0]), .C(n564), .Y(n547) );
  OA21XL U135 ( .B(r_pwdn_en), .C(n605), .A(n535), .Y(n546) );
  NOR5XL U136 ( .A(c_ptr[3]), .B(d_psrd), .C(n526), .D(n631), .E(n525), .Y(
        n527) );
  NAND21X1 U137 ( .B(n614), .A(n613), .Y(n618) );
  NAND21X1 U138 ( .B(n99), .A(n507), .Y(n441) );
  NAND32X1 U139 ( .B(n573), .C(n619), .A(n572), .Y(N853) );
  AOI21X1 U140 ( .B(we_twlb), .C(n592), .A(N853), .Y(n36) );
  INVX1 U141 ( .A(n431), .Y(n614) );
  INVX1 U142 ( .A(n572), .Y(n613) );
  INVX1 U143 ( .A(n97), .Y(n83) );
  INVX1 U144 ( .A(n98), .Y(n82) );
  INVX1 U145 ( .A(n98), .Y(n81) );
  INVX1 U146 ( .A(n528), .Y(n80) );
  INVX1 U147 ( .A(n528), .Y(n79) );
  INVX1 U148 ( .A(n97), .Y(n86) );
  INVX1 U149 ( .A(n97), .Y(n85) );
  INVX1 U150 ( .A(n97), .Y(n84) );
  INVX1 U151 ( .A(n97), .Y(n90) );
  INVX1 U152 ( .A(n98), .Y(n89) );
  INVX1 U153 ( .A(n97), .Y(n88) );
  INVX1 U154 ( .A(n97), .Y(n87) );
  INVX1 U155 ( .A(n97), .Y(n95) );
  INVX1 U156 ( .A(n98), .Y(n92) );
  INVX1 U157 ( .A(n97), .Y(n94) );
  INVX1 U158 ( .A(n97), .Y(n91) );
  INVX1 U159 ( .A(n98), .Y(n96) );
  INVX1 U160 ( .A(n567), .Y(n602) );
  NAND21X1 U161 ( .B(n594), .A(n568), .Y(n661) );
  INVX1 U162 ( .A(n291), .Y(n910) );
  INVX1 U163 ( .A(n295), .Y(n905) );
  NAND2X1 U164 ( .A(n364), .B(n368), .Y(n275) );
  INVX1 U165 ( .A(n621), .Y(n630) );
  INVX1 U166 ( .A(n282), .Y(n721) );
  INVX1 U167 ( .A(n578), .Y(n568) );
  NOR2X1 U168 ( .A(n924), .B(n23), .Y(n574) );
  INVX1 U169 ( .A(n686), .Y(n103) );
  NAND43X1 U170 ( .B(n179), .C(n178), .D(n177), .A(n176), .Y(n431) );
  INVX1 U171 ( .A(n141), .Y(n179) );
  NOR43XL U172 ( .B(n293), .C(n175), .D(n174), .A(n173), .Y(n176) );
  NAND32X1 U173 ( .B(n614), .C(n564), .A(n430), .Y(n435) );
  NAND21X1 U174 ( .B(n16), .A(n78), .Y(n617) );
  OAI211X1 U175 ( .C(n16), .D(n571), .A(n609), .B(n570), .Y(n619) );
  AND3X1 U176 ( .A(n103), .B(n583), .C(n615), .Y(n570) );
  INVX1 U177 ( .A(n655), .Y(n652) );
  OR2X1 U178 ( .A(n621), .B(n571), .Y(n507) );
  AO21X1 U179 ( .B(n627), .C(n635), .A(n100), .Y(N885) );
  AO21X1 U180 ( .B(n57), .C(n635), .A(n100), .Y(N889) );
  INVX1 U181 ( .A(n657), .Y(n653) );
  INVX1 U182 ( .A(memaddr_c[10]), .Y(n198) );
  INVX1 U183 ( .A(n175), .Y(n160) );
  NAND21X1 U184 ( .B(n577), .A(n592), .Y(n609) );
  INVX1 U185 ( .A(n542), .Y(n594) );
  INVX1 U186 ( .A(n569), .Y(n592) );
  AO21X1 U187 ( .B(n433), .C(n542), .A(n559), .Y(n567) );
  INVX1 U188 ( .A(n662), .Y(n544) );
  AND2X1 U189 ( .A(n377), .B(n366), .Y(n282) );
  AND2X1 U190 ( .A(n378), .B(n367), .Y(n295) );
  AND2X1 U191 ( .A(n377), .B(n367), .Y(n291) );
  NAND2X1 U192 ( .A(n370), .B(n365), .Y(n273) );
  NAND2X1 U193 ( .A(n370), .B(n366), .Y(n278) );
  NAND2X1 U194 ( .A(n378), .B(n366), .Y(n37) );
  NAND2X1 U195 ( .A(n378), .B(n368), .Y(n38) );
  OAI211X1 U196 ( .C(n664), .D(n663), .A(n662), .B(n661), .Y(N898) );
  AND2X1 U197 ( .A(n660), .B(n659), .Y(n664) );
  NOR2X1 U198 ( .A(n369), .B(n931), .Y(n364) );
  NAND2X1 U199 ( .A(n377), .B(n368), .Y(n288) );
  NAND2X1 U200 ( .A(n376), .B(n366), .Y(n286) );
  NAND2X1 U201 ( .A(n376), .B(n367), .Y(n289) );
  NAND2X1 U202 ( .A(n376), .B(n368), .Y(n285) );
  NAND2X1 U203 ( .A(n376), .B(n365), .Y(n287) );
  NAND2X1 U204 ( .A(n366), .B(n371), .Y(n279) );
  NAND2X1 U205 ( .A(n370), .B(n368), .Y(n276) );
  NAND2X1 U206 ( .A(n364), .B(n367), .Y(n270) );
  NAND2X1 U207 ( .A(n365), .B(n371), .Y(n277) );
  NAND2X1 U208 ( .A(n368), .B(n371), .Y(n280) );
  NAND2X1 U209 ( .A(n367), .B(n371), .Y(n281) );
  NAND2X1 U210 ( .A(n370), .B(n367), .Y(n274) );
  NAND2X1 U211 ( .A(n364), .B(n366), .Y(n271) );
  NAND2X1 U212 ( .A(n364), .B(n365), .Y(n272) );
  NAND2X1 U213 ( .A(n377), .B(n365), .Y(n39) );
  NAND2X1 U214 ( .A(n378), .B(n365), .Y(n40) );
  INVX1 U215 ( .A(n369), .Y(n932) );
  OR2XL U216 ( .A(n686), .B(n16), .Y(n621) );
  NOR2X1 U217 ( .A(n933), .B(n379), .Y(n368) );
  NAND21X1 U218 ( .B(o_ofs_inc), .A(n102), .Y(n559) );
  INVX1 U219 ( .A(n440), .Y(n442) );
  INVX1 U220 ( .A(n579), .Y(n596) );
  NAND21X1 U221 ( .B(n578), .A(n577), .Y(n579) );
  NAND21X1 U222 ( .B(n675), .A(n679), .Y(n690) );
  INVX1 U223 ( .A(n659), .Y(n675) );
  INVX1 U224 ( .A(srst), .Y(n104) );
  XOR2X1 U225 ( .A(n129), .B(n391), .Y(n144) );
  XOR2X1 U226 ( .A(n127), .B(n66), .Y(n151) );
  NOR2X1 U227 ( .A(dw_rst), .B(srst), .Y(n418) );
  INVX1 U228 ( .A(n119), .Y(n153) );
  XOR2X1 U229 ( .A(n132), .B(n386), .Y(n143) );
  INVX1 U230 ( .A(n121), .Y(n120) );
  INVX1 U231 ( .A(n125), .Y(n122) );
  INVX1 U232 ( .A(n123), .Y(n124) );
  INVX1 U233 ( .A(n140), .Y(n139) );
  INVX1 U234 ( .A(n381), .Y(n232) );
  INVX1 U235 ( .A(n242), .Y(n246) );
  INVX1 U236 ( .A(n314), .Y(n334) );
  INVX1 U237 ( .A(n344), .Y(n347) );
  AND3X1 U238 ( .A(o_inst[5]), .B(o_inst[7]), .C(o_inst[6]), .Y(n260) );
  AND3X1 U239 ( .A(o_inst[2]), .B(o_inst[4]), .C(o_inst[3]), .Y(n259) );
  INVX1 U240 ( .A(n612), .Y(n523) );
  INVX1 U241 ( .A(n515), .Y(n925) );
  INVX1 U242 ( .A(n669), .Y(n607) );
  INVX1 U243 ( .A(n660), .Y(n924) );
  INVX1 U244 ( .A(n525), .Y(n505) );
  NAND32X1 U245 ( .B(pmem_csb), .C(o_ofs_inc), .A(n669), .Y(n670) );
  NAND21X1 U246 ( .B(n551), .A(n549), .Y(n564) );
  NAND21X1 U247 ( .B(n528), .A(n630), .Y(n655) );
  NAND32X1 U248 ( .B(n16), .C(n435), .A(n694), .Y(n615) );
  GEN2XL U249 ( .D(n64), .E(n148), .C(n356), .B(n43), .A(n147), .Y(n149) );
  INVX1 U250 ( .A(n143), .Y(n146) );
  INVX1 U251 ( .A(n144), .Y(n145) );
  OAI2B11X1 U252 ( .D(n430), .C(n30), .A(n549), .B(n534), .Y(n535) );
  EORX1 U253 ( .A(n141), .B(n41), .C(memaddr_c[7]), .D(n158), .Y(n161) );
  OAI22X1 U254 ( .A(n157), .B(n171), .C(memaddr_c[6]), .D(n156), .Y(n41) );
  NAND2X1 U255 ( .A(n42), .B(n182), .Y(n185) );
  OAI22XL U256 ( .A(memaddr_c[2]), .B(n732), .C(memaddr_c[3]), .D(n739), .Y(
        n42) );
  INVX1 U257 ( .A(n528), .Y(n504) );
  OAI211X1 U258 ( .C(n208), .D(n581), .A(n170), .B(n172), .Y(n206) );
  OAI222XL U259 ( .A(memaddr_c[13]), .B(n169), .C(n168), .D(n167), .E(
        memaddr_c[12]), .F(n166), .Y(n170) );
  OA222X1 U260 ( .A(memaddr_c[11]), .B(n165), .C(n164), .D(n178), .E(
        memaddr_c[10]), .F(n163), .Y(n168) );
  OA222X1 U261 ( .A(memaddr_c[9]), .B(n162), .C(n161), .D(n160), .E(
        memaddr_c[8]), .F(n159), .Y(n164) );
  OAI32X1 U262 ( .A(n190), .B(memaddr_c[4]), .C(n731), .D(n189), .E(n188), .Y(
        n191) );
  GEN2XL U263 ( .D(memaddr_c[1]), .E(n187), .C(n186), .B(n185), .A(n190), .Y(
        n188) );
  INVX1 U264 ( .A(n220), .Y(n190) );
  INVX1 U265 ( .A(n526), .Y(n551) );
  INVX1 U266 ( .A(n142), .Y(n356) );
  NAND21X1 U267 ( .B(memaddr_c[0]), .A(n65), .Y(n142) );
  OA22X1 U268 ( .A(n143), .B(n136), .C(n64), .D(n148), .Y(n43) );
  NAND21X1 U269 ( .B(n638), .A(n637), .Y(n657) );
  OAI22AX1 U270 ( .D(n156), .C(n245), .A(n155), .B(n154), .Y(n171) );
  INVX1 U271 ( .A(n620), .Y(n632) );
  INVX1 U272 ( .A(memaddr_c[6]), .Y(n245) );
  OAI211X1 U273 ( .C(n658), .D(n657), .A(n663), .B(n656), .Y(N897) );
  INVXL U274 ( .A(memaddr_c[5]), .Y(n155) );
  NAND2X1 U275 ( .A(n158), .B(memaddr_c[7]), .Y(n141) );
  INVX1 U276 ( .A(n481), .Y(n496) );
  INVX1 U277 ( .A(n493), .Y(n502) );
  INVX1 U278 ( .A(n491), .Y(n501) );
  INVX1 U279 ( .A(n489), .Y(n500) );
  INVX1 U280 ( .A(n485), .Y(n498) );
  INVX1 U281 ( .A(n483), .Y(n497) );
  INVX1 U282 ( .A(n495), .Y(n503) );
  INVX1 U283 ( .A(n487), .Y(n499) );
  AOI21XL U284 ( .B(memaddr_c[2]), .C(n20), .A(n101), .Y(n45) );
  AOI21XL U285 ( .B(memaddr_c[5]), .C(n20), .A(n101), .Y(n48) );
  AOI21X1 U286 ( .B(memaddr_c[7]), .C(n432), .A(n77), .Y(n50) );
  AOI21X1 U287 ( .B(memaddr_c[8]), .C(n432), .A(n77), .Y(n51) );
  AOI21X1 U288 ( .B(memaddr_c[9]), .C(n432), .A(n77), .Y(n52) );
  AOI21X1 U289 ( .B(memaddr_c[10]), .C(n432), .A(n77), .Y(n53) );
  AOI21X1 U290 ( .B(memaddr_c[11]), .C(n432), .A(n101), .Y(n54) );
  AOI21X1 U291 ( .B(memaddr_c[13]), .C(n432), .A(n77), .Y(n55) );
  AOI21X1 U292 ( .B(memaddr_c[12]), .C(n432), .A(n77), .Y(n56) );
  AO21X1 U293 ( .B(n627), .C(n640), .A(n100), .Y(N883) );
  AO21X1 U294 ( .B(n627), .C(n654), .A(n100), .Y(N884) );
  AO21X1 U295 ( .B(n57), .C(n639), .A(n100), .Y(N886) );
  AO21X1 U296 ( .B(n57), .C(n640), .A(n100), .Y(N887) );
  AO21X1 U297 ( .B(n57), .C(n654), .A(n100), .Y(N888) );
  AO21X1 U298 ( .B(n636), .C(n639), .A(n100), .Y(N890) );
  AO21X1 U299 ( .B(n636), .C(n640), .A(n100), .Y(N891) );
  AO21X1 U300 ( .B(n636), .C(n654), .A(n100), .Y(N892) );
  AO21X1 U301 ( .B(n636), .C(n635), .A(n652), .Y(N893) );
  AO21X1 U302 ( .B(n653), .C(n639), .A(n652), .Y(N894) );
  AO21X1 U303 ( .B(n640), .C(n653), .A(n652), .Y(N895) );
  AO21X1 U304 ( .B(n654), .C(n653), .A(n652), .Y(N896) );
  INVX1 U305 ( .A(n624), .Y(n625) );
  NAND32X1 U306 ( .B(n638), .C(n628), .A(n629), .Y(n624) );
  INVX1 U307 ( .A(n626), .Y(n627) );
  NAND32X1 U308 ( .B(n629), .C(n628), .A(n638), .Y(n626) );
  NOR3XL U309 ( .A(n629), .B(n638), .C(n628), .Y(n57) );
  NAND2X1 U310 ( .A(n159), .B(memaddr_c[8]), .Y(n175) );
  OA21X1 U311 ( .B(n654), .C(n640), .A(n509), .Y(N843) );
  INVX1 U312 ( .A(memaddr_c[8]), .Y(n249) );
  INVX1 U313 ( .A(memaddr_c[12]), .Y(n205) );
  NAND6XL U314 ( .A(n612), .B(n17), .C(n610), .D(n609), .E(n673), .F(n608), 
        .Y(N820) );
  AOI32X1 U315 ( .A(n607), .B(n606), .C(n605), .D(n667), .E(n920), .Y(n608) );
  AND3X1 U316 ( .A(n925), .B(n602), .C(n601), .Y(n610) );
  INVX1 U317 ( .A(n600), .Y(n601) );
  AO22AXL U318 ( .A(n162), .B(memaddr_c[9]), .C(n163), .D(n198), .Y(n178) );
  AO22AXL U319 ( .A(n165), .B(memaddr_c[11]), .C(n166), .D(n205), .Y(n167) );
  AND2X1 U320 ( .A(n509), .B(n427), .Y(N842) );
  INVX1 U321 ( .A(n375), .Y(n196) );
  NAND6XL U322 ( .A(n426), .B(n425), .C(n424), .D(n423), .E(n422), .F(n421), 
        .Y(n430) );
  MUX2X1 U323 ( .D0(n235), .D1(n314), .S(memaddr_c[10]), .Y(n424) );
  XOR2X1 U324 ( .A(n241), .B(n222), .Y(n426) );
  XOR2X1 U325 ( .A(n246), .B(n238), .Y(n423) );
  NAND2X1 U326 ( .A(n169), .B(memaddr_c[13]), .Y(n172) );
  INVX1 U327 ( .A(memaddr_c[13]), .Y(n231) );
  INVX1 U328 ( .A(memaddr_c[14]), .Y(n581) );
  NOR6XL U329 ( .A(n420), .B(n419), .C(n416), .D(n415), .E(n414), .F(n392), 
        .Y(n421) );
  INVX1 U330 ( .A(n293), .Y(n355) );
  OA21X1 U331 ( .B(n347), .C(n346), .A(n345), .Y(n348) );
  AO21X1 U332 ( .B(n335), .C(n334), .A(n325), .Y(n354) );
  NAND32X1 U333 ( .B(n578), .C(n542), .A(n588), .Y(n662) );
  AO21X1 U334 ( .B(sfr_psr), .C(n538), .A(n549), .Y(n542) );
  NAND21X1 U335 ( .B(n560), .A(n594), .Y(n569) );
  NAND21X1 U336 ( .B(n65), .A(memaddr_c[0]), .Y(n293) );
  XOR2X1 U337 ( .A(memaddr_c[14]), .B(n208), .Y(n173) );
  XNOR2XL U338 ( .A(n58), .B(memaddr_c[12]), .Y(n283) );
  AOI21X1 U339 ( .B(n294), .C(n251), .A(n250), .Y(n58) );
  AND4X1 U340 ( .A(n292), .B(n290), .C(n284), .D(n283), .Y(n422) );
  XOR2X1 U341 ( .A(n245), .B(n244), .Y(n290) );
  XOR2X1 U342 ( .A(n249), .B(n248), .Y(n284) );
  XOR2X1 U343 ( .A(n240), .B(n239), .Y(n292) );
  XNOR2XL U344 ( .A(n381), .B(n59), .Y(n416) );
  NAND2X1 U345 ( .A(n375), .B(n374), .Y(n59) );
  AND2X1 U346 ( .A(n237), .B(n236), .Y(n238) );
  INVX1 U347 ( .A(n345), .Y(n202) );
  AND2X1 U348 ( .A(n372), .B(n931), .Y(n370) );
  NOR3XL U349 ( .A(n372), .B(n931), .C(n932), .Y(n377) );
  NOR3XL U350 ( .A(n373), .B(n372), .C(n932), .Y(n378) );
  INVX1 U351 ( .A(n549), .Y(n606) );
  NAND4X1 U352 ( .A(n262), .B(n263), .C(n264), .D(n265), .Y(o_inst[7]) );
  NOR4XL U353 ( .A(n266), .B(n267), .C(n268), .D(n269), .Y(n265) );
  OA222X1 U354 ( .A(n40), .B(n907), .C(n37), .D(n906), .E(n905), .F(n904), .Y(
        n262) );
  OA222X1 U355 ( .A(n39), .B(n911), .C(n910), .D(n909), .E(n38), .F(n908), .Y(
        n263) );
  XNOR2XL U356 ( .A(n383), .B(n384), .Y(n369) );
  XOR2X1 U357 ( .A(n739), .B(n936), .Y(n384) );
  AO21X1 U358 ( .B(n738), .C(n737), .A(n736), .Y(n383) );
  INVX1 U359 ( .A(n385), .Y(n737) );
  INVX1 U360 ( .A(n733), .Y(n736) );
  NAND21X1 U361 ( .B(n732), .A(n935), .Y(n733) );
  AND2X1 U362 ( .A(n372), .B(n373), .Y(n371) );
  NAND21X1 U363 ( .B(n935), .A(n732), .Y(n738) );
  NOR2X1 U364 ( .A(n373), .B(n369), .Y(n376) );
  INVX1 U365 ( .A(n373), .Y(n931) );
  OR4X1 U366 ( .A(n726), .B(n60), .C(n61), .D(n62), .Y(o_inst[1]) );
  OAI222XL U367 ( .A(n39), .B(n718), .C(n38), .D(n717), .E(n910), .F(n716), 
        .Y(n60) );
  OAI222XL U368 ( .A(n288), .B(n722), .C(n721), .D(n720), .E(n287), .F(n719), 
        .Y(n61) );
  OAI222XL U369 ( .A(n286), .B(n725), .C(n289), .D(n724), .E(n285), .F(n723), 
        .Y(n62) );
  NAND31X1 U370 ( .C(n711), .A(n710), .B(n709), .Y(o_inst[0]) );
  NOR43XL U371 ( .B(n708), .C(n707), .D(n706), .A(n705), .Y(n709) );
  NAND31X1 U372 ( .C(n697), .A(n696), .B(n695), .Y(n711) );
  NOR43XL U373 ( .B(n700), .C(n699), .D(n359), .A(n698), .Y(n710) );
  NOR2X1 U374 ( .A(n934), .B(n933), .Y(n366) );
  NOR2X1 U375 ( .A(n380), .B(n934), .Y(n365) );
  NOR2X1 U376 ( .A(n380), .B(n379), .Y(n367) );
  INVX1 U377 ( .A(n582), .Y(n586) );
  INVX1 U378 ( .A(n934), .Y(n379) );
  INVX1 U379 ( .A(n107), .Y(o_ofs_inc) );
  NAND32X1 U380 ( .B(n511), .C(n111), .A(n513), .Y(n107) );
  INVX1 U381 ( .A(n380), .Y(n933) );
  NOR4XL U382 ( .A(n310), .B(n311), .C(n312), .D(n313), .Y(n309) );
  OAI222XL U383 ( .A(n280), .B(n843), .C(n279), .D(n842), .E(n281), .F(n841), 
        .Y(n310) );
  OAI222XL U384 ( .A(n271), .B(n852), .C(n270), .D(n851), .E(n272), .F(n850), 
        .Y(n313) );
  OAI222XL U385 ( .A(n277), .B(n846), .C(n276), .D(n845), .E(n278), .F(n844), 
        .Y(n311) );
  NOR4XL U386 ( .A(n320), .B(n321), .C(n322), .D(n323), .Y(n319) );
  OAI222XL U387 ( .A(n280), .B(n818), .C(n279), .D(n817), .E(n281), .F(n816), 
        .Y(n320) );
  OAI222XL U388 ( .A(n271), .B(n827), .C(n270), .D(n826), .E(n272), .F(n825), 
        .Y(n323) );
  OAI222XL U389 ( .A(n277), .B(n821), .C(n276), .D(n820), .E(n278), .F(n819), 
        .Y(n321) );
  NOR4XL U390 ( .A(n300), .B(n301), .C(n302), .D(n303), .Y(n299) );
  OAI222XL U391 ( .A(n280), .B(n868), .C(n279), .D(n867), .E(n281), .F(n866), 
        .Y(n300) );
  OAI222XL U392 ( .A(n271), .B(n878), .C(n270), .D(n877), .E(n272), .F(n876), 
        .Y(n303) );
  OAI222XL U393 ( .A(n277), .B(n871), .C(n276), .D(n870), .E(n278), .F(n869), 
        .Y(n301) );
  NOR4XL U394 ( .A(n330), .B(n331), .C(n332), .D(n333), .Y(n329) );
  OAI222XL U395 ( .A(n280), .B(n793), .C(n279), .D(n792), .E(n281), .F(n791), 
        .Y(n330) );
  OAI222XL U396 ( .A(n271), .B(n802), .C(n270), .D(n801), .E(n272), .F(n800), 
        .Y(n333) );
  OAI222XL U397 ( .A(n277), .B(n796), .C(n276), .D(n795), .E(n278), .F(n794), 
        .Y(n331) );
  NOR4XL U398 ( .A(n340), .B(n341), .C(n342), .D(n343), .Y(n339) );
  OAI222XL U399 ( .A(n280), .B(n768), .C(n279), .D(n767), .E(n281), .F(n766), 
        .Y(n340) );
  OAI222XL U400 ( .A(n271), .B(n777), .C(n270), .D(n776), .E(n272), .F(n775), 
        .Y(n343) );
  OAI222XL U401 ( .A(n277), .B(n771), .C(n276), .D(n770), .E(n278), .F(n769), 
        .Y(n341) );
  NOR4XL U402 ( .A(n360), .B(n361), .C(n362), .D(n363), .Y(n359) );
  OAI222XL U403 ( .A(n280), .B(n743), .C(n279), .D(n742), .E(n281), .F(n741), 
        .Y(n360) );
  OAI222XL U404 ( .A(n271), .B(n752), .C(n270), .D(n751), .E(n272), .F(n750), 
        .Y(n363) );
  OAI222XL U405 ( .A(n277), .B(n746), .C(n276), .D(n745), .E(n278), .F(n744), 
        .Y(n361) );
  NAND4X1 U406 ( .A(n306), .B(n307), .C(n308), .D(n309), .Y(o_inst[5]) );
  OA222X1 U407 ( .A(n40), .B(n855), .C(n37), .D(n854), .E(n905), .F(n853), .Y(
        n306) );
  OA222X1 U408 ( .A(n39), .B(n858), .C(n910), .D(n857), .E(n38), .F(n856), .Y(
        n307) );
  NOR43XL U409 ( .B(n865), .C(n864), .D(n863), .A(n862), .Y(n308) );
  NAND4X1 U410 ( .A(n336), .B(n337), .C(n338), .D(n339), .Y(o_inst[2]) );
  OA222X1 U411 ( .A(n40), .B(n780), .C(n37), .D(n779), .E(n905), .F(n778), .Y(
        n336) );
  OA222X1 U412 ( .A(n39), .B(n783), .C(n910), .D(n782), .E(n38), .F(n781), .Y(
        n337) );
  NOR43XL U413 ( .B(n790), .C(n789), .D(n788), .A(n787), .Y(n338) );
  NAND4X1 U414 ( .A(n316), .B(n317), .C(n318), .D(n319), .Y(o_inst[4]) );
  OA222X1 U415 ( .A(n905), .B(n830), .C(n40), .D(n829), .E(n37), .F(n828), .Y(
        n316) );
  OA222X1 U416 ( .A(n39), .B(n833), .C(n38), .D(n832), .E(n910), .F(n831), .Y(
        n317) );
  NOR43XL U417 ( .B(n840), .C(n839), .D(n838), .A(n837), .Y(n318) );
  NAND4X1 U418 ( .A(n296), .B(n297), .C(n298), .D(n299), .Y(o_inst[6]) );
  OA222X1 U419 ( .A(n40), .B(n881), .C(n37), .D(n880), .E(n905), .F(n879), .Y(
        n296) );
  OA222X1 U420 ( .A(n39), .B(n884), .C(n910), .D(n883), .E(n38), .F(n882), .Y(
        n297) );
  NOR43XL U421 ( .B(n891), .C(n890), .D(n889), .A(n888), .Y(n298) );
  NAND4X1 U422 ( .A(n326), .B(n327), .C(n328), .D(n329), .Y(o_inst[3]) );
  OA222X1 U423 ( .A(n40), .B(n805), .C(n37), .D(n804), .E(n905), .F(n803), .Y(
        n326) );
  OA222X1 U424 ( .A(n39), .B(n808), .C(n910), .D(n807), .E(n38), .F(n806), .Y(
        n327) );
  NOR43XL U425 ( .B(n815), .C(n814), .D(n813), .A(n812), .Y(n328) );
  OAI21BBX1 U426 ( .A(n478), .B(n583), .C(n102), .Y(n440) );
  AO21X1 U427 ( .B(n925), .C(n940), .A(n77), .Y(n543) );
  INVX1 U428 ( .A(n434), .Y(n557) );
  NAND21X1 U429 ( .B(n929), .A(n102), .Y(n663) );
  INVX1 U430 ( .A(n439), .Y(n443) );
  INVX1 U431 ( .A(n446), .Y(n447) );
  NAND21X1 U432 ( .B(n512), .A(n510), .Y(n659) );
  NAND32X1 U433 ( .B(n513), .C(n512), .A(n511), .Y(n688) );
  INVX1 U434 ( .A(n475), .Y(n693) );
  AND2X1 U435 ( .A(n102), .B(n668), .Y(N899) );
  OAI22X1 U436 ( .A(n940), .B(n667), .C(n925), .D(n666), .Y(n668) );
  AND2X1 U437 ( .A(n665), .B(n743), .Y(n666) );
  INVX1 U438 ( .A(n940), .Y(n920) );
  INVX1 U439 ( .A(n674), .Y(n679) );
  NAND21X1 U440 ( .B(n920), .A(n673), .Y(n674) );
  INVX1 U441 ( .A(n684), .Y(n691) );
  NAND32X1 U442 ( .B(n511), .C(n512), .A(n513), .Y(n669) );
  NAND21X1 U443 ( .B(n513), .A(n109), .Y(n672) );
  INVX1 U444 ( .A(n588), .Y(n577) );
  INVX1 U445 ( .A(n417), .Y(n532) );
  AND2X1 U446 ( .A(n418), .B(n417), .Y(n63) );
  AO21X1 U447 ( .B(n127), .C(n219), .A(n218), .Y(n152) );
  NAND2X1 U448 ( .A(n152), .B(n223), .Y(n119) );
  AO21X1 U449 ( .B(n132), .C(n215), .A(n214), .Y(n129) );
  AO21X1 U450 ( .B(n129), .C(n217), .A(n216), .Y(n127) );
  OAI221X1 U451 ( .A(n187), .B(n137), .C(n740), .D(n658), .E(n133), .Y(n132)
         );
  AO21X1 U452 ( .B(n125), .C(n305), .A(n124), .Y(n165) );
  AO21X1 U453 ( .B(n123), .C(n251), .A(n139), .Y(n166) );
  NAND21X1 U454 ( .B(n225), .A(n153), .Y(n138) );
  OR2X1 U455 ( .A(n224), .B(n138), .Y(n121) );
  NAND21X1 U456 ( .B(n251), .A(n124), .Y(n140) );
  NAND21X1 U457 ( .B(n305), .A(n122), .Y(n123) );
  NAND21X1 U458 ( .B(n226), .A(n120), .Y(n125) );
  INVX1 U459 ( .A(n128), .Y(n391) );
  NAND21X1 U460 ( .B(n216), .A(n217), .Y(n128) );
  XNOR2XL U461 ( .A(n137), .B(n358), .Y(n64) );
  INVX1 U462 ( .A(n133), .Y(n212) );
  INVX1 U463 ( .A(n135), .Y(n358) );
  NAND21X1 U464 ( .B(n212), .A(n213), .Y(n135) );
  INVX1 U465 ( .A(n131), .Y(n386) );
  NAND21X1 U466 ( .B(n214), .A(n215), .Y(n131) );
  AND2X1 U467 ( .A(n357), .B(n137), .Y(n65) );
  INVX1 U468 ( .A(n126), .Y(n218) );
  AND2X1 U469 ( .A(n219), .B(n126), .Y(n66) );
  NAND21X1 U470 ( .B(n226), .A(n232), .Y(n314) );
  AO21X1 U471 ( .B(n389), .C(n219), .A(n218), .Y(n241) );
  NAND32X1 U472 ( .B(n225), .C(n224), .A(n246), .Y(n381) );
  AO21X1 U473 ( .B(n382), .C(n215), .A(n214), .Y(n390) );
  AO21X1 U474 ( .B(n390), .C(n217), .A(n216), .Y(n389) );
  AO21X1 U475 ( .B(n357), .C(n213), .A(n212), .Y(n382) );
  NAND2X1 U476 ( .A(n241), .B(n223), .Y(n242) );
  INVX1 U477 ( .A(n229), .Y(n250) );
  NAND21X1 U478 ( .B(n233), .A(n232), .Y(n344) );
  NAND21X1 U479 ( .B(n665), .A(hit_ps), .Y(n539) );
  NAND21X1 U480 ( .B(n538), .A(n539), .Y(n605) );
  INVX1 U481 ( .A(n560), .Y(n433) );
  INVX1 U482 ( .A(n115), .Y(n534) );
  NAND32X1 U483 ( .B(n631), .C(n629), .A(n180), .Y(n115) );
  NAND21X1 U484 ( .B(n513), .A(n691), .Y(n612) );
  NAND21X1 U485 ( .B(n694), .A(n523), .Y(n583) );
  NOR21XL U486 ( .B(r_hold_mcu), .A(srst), .Y(n874) );
  NAND21X1 U487 ( .B(n675), .A(n671), .Y(n515) );
  INVX1 U488 ( .A(n929), .Y(n919) );
  INVX1 U489 ( .A(n451), .Y(n472) );
  NAND21X1 U490 ( .B(n693), .A(n682), .Y(n451) );
  NAND21X1 U491 ( .B(n638), .A(n635), .Y(n525) );
  NAND2X1 U492 ( .A(n673), .B(n669), .Y(n558) );
  NAND5XL U493 ( .A(n868), .B(n818), .C(n793), .D(n768), .E(n514), .Y(n660) );
  AND4X1 U494 ( .A(n843), .B(n755), .C(n894), .D(n743), .Y(n514) );
  INVX1 U495 ( .A(n658), .Y(n635) );
  INVX1 U496 ( .A(n599), .Y(n921) );
  INVX1 U497 ( .A(n604), .Y(n667) );
  NAND21X1 U498 ( .B(n939), .A(n923), .Y(n604) );
  INVX1 U499 ( .A(n555), .Y(n927) );
  INVX1 U500 ( .A(n554), .Y(n926) );
  INVX1 U501 ( .A(n506), .Y(n508) );
  NAND21X1 U502 ( .B(n629), .A(n505), .Y(n506) );
  OAI31XL U503 ( .A(n691), .B(n690), .C(n689), .D(n688), .Y(n692) );
  INVX1 U504 ( .A(pmem_clk[0]), .Y(n689) );
  AOI32X1 U505 ( .A(pmem_clk[1]), .B(n685), .C(n684), .D(n2), .E(n683), .Y(
        n687) );
  INVX1 U506 ( .A(n690), .Y(n685) );
  INVX1 U507 ( .A(n682), .Y(n683) );
  NAND32X1 U508 ( .B(n211), .C(n210), .A(n209), .Y(n526) );
  AND3X1 U509 ( .A(n631), .B(n629), .C(n180), .Y(n211) );
  AO21X1 U510 ( .B(n208), .C(n581), .A(n207), .Y(n209) );
  NAND2X1 U511 ( .A(n4), .B(pre_1_adr[14]), .Y(n591) );
  AND3X1 U512 ( .A(wd_twlb[0]), .B(we_twlb), .C(n594), .Y(n597) );
  AND3X1 U513 ( .A(wd_twlb[1]), .B(we_twlb), .C(n594), .Y(n593) );
  OAI211X1 U514 ( .C(pre_1_adr[13]), .D(n591), .A(n590), .B(n589), .Y(n595) );
  AOI33X1 U515 ( .A(n588), .B(n587), .C(n586), .D(sfr_psofs[14]), .E(n585), 
        .F(n584), .Y(n589) );
  NAND32X1 U516 ( .B(memaddr_c[13]), .C(n581), .A(n580), .Y(n590) );
  INVX1 U517 ( .A(sfr_psofs[13]), .Y(n584) );
  OA21X1 U518 ( .B(c_adr[12]), .C(n205), .A(n201), .Y(n204) );
  OAI22X1 U519 ( .A(memaddr_c[11]), .B(n305), .C(n335), .D(n200), .Y(n201) );
  AOI22X1 U520 ( .A(n199), .B(n346), .C(c_adr[10]), .D(n198), .Y(n200) );
  AOI32X1 U521 ( .A(n195), .B(n194), .C(n237), .D(memaddr_c[8]), .E(n224), .Y(
        n197) );
  OAI221X1 U522 ( .A(c_adr[6]), .B(n245), .C(n192), .D(n191), .E(n236), .Y(
        n195) );
  INVX1 U523 ( .A(n221), .Y(n192) );
  OAI32X1 U524 ( .A(d_psrd), .B(n101), .C(n612), .D(n435), .E(n434), .Y(n580)
         );
  NAND21XL U525 ( .B(c_adr[3]), .A(memaddr_c[3]), .Y(n182) );
  NAND21XL U526 ( .B(c_adr[5]), .A(memaddr_c[5]), .Y(n220) );
  AO2222XL U527 ( .A(memaddr[9]), .B(n443), .C(sfr_psofs[9]), .D(n442), .E(
        memaddr_c[9]), .F(n580), .G(pre_1_adr[9]), .H(n4), .Y(N863) );
  AO2222XL U528 ( .A(memaddr[2]), .B(n443), .C(sfr_psofs[2]), .D(n442), .E(
        memaddr_c[2]), .F(n580), .G(pre_1_adr[2]), .H(n441), .Y(N856) );
  AO2222XL U529 ( .A(memaddr[12]), .B(n7), .C(sfr_psofs[12]), .D(n10), .E(
        memaddr_c[12]), .F(n13), .G(pre_1_adr[12]), .H(n441), .Y(N866) );
  AO2222XL U530 ( .A(memaddr[11]), .B(n443), .C(sfr_psofs[11]), .D(n442), .E(
        memaddr_c[11]), .F(n580), .G(pre_1_adr[11]), .H(n4), .Y(N865) );
  AO2222XL U531 ( .A(memaddr[8]), .B(n7), .C(sfr_psofs[8]), .D(n10), .E(
        memaddr_c[8]), .F(n13), .G(pre_1_adr[8]), .H(n4), .Y(N862) );
  AO2222XL U532 ( .A(memaddr[7]), .B(n443), .C(sfr_psofs[7]), .D(n442), .E(
        memaddr_c[7]), .F(n580), .G(pre_1_adr[7]), .H(n441), .Y(N861) );
  AO2222XL U533 ( .A(memaddr[3]), .B(n443), .C(sfr_psofs[3]), .D(n442), .E(
        memaddr_c[3]), .F(n580), .G(pre_1_adr[3]), .H(n4), .Y(N857) );
  AO2222XL U534 ( .A(memaddr[13]), .B(n443), .C(sfr_psofs[13]), .D(n442), .E(
        memaddr_c[13]), .F(n580), .G(pre_1_adr[13]), .H(n441), .Y(N867) );
  AO2222XL U535 ( .A(memaddr[6]), .B(n443), .C(sfr_psofs[6]), .D(n442), .E(
        memaddr_c[6]), .F(n580), .G(pre_1_adr[6]), .H(n441), .Y(N860) );
  AO2222XL U536 ( .A(memaddr[4]), .B(n443), .C(sfr_psofs[4]), .D(n442), .E(
        memaddr_c[4]), .F(n580), .G(pre_1_adr[4]), .H(n4), .Y(N858) );
  AO2222XL U537 ( .A(n7), .B(memaddr[0]), .C(sfr_psofs[0]), .D(n10), .E(
        memaddr_c[0]), .F(n13), .G(pre_1_adr[0]), .H(n441), .Y(N854) );
  AO2222XL U538 ( .A(memaddr[5]), .B(n443), .C(sfr_psofs[5]), .D(n442), .E(
        memaddr_c[5]), .F(n13), .G(pre_1_adr[5]), .H(n441), .Y(N859) );
  AO2222XL U539 ( .A(memaddr[10]), .B(n7), .C(sfr_psofs[10]), .D(n10), .E(
        memaddr_c[10]), .F(n13), .G(pre_1_adr[10]), .H(n4), .Y(N864) );
  AO2222XL U540 ( .A(n443), .B(memaddr[1]), .C(sfr_psofs[1]), .D(n442), .E(
        memaddr_c[1]), .F(n13), .G(pre_1_adr[1]), .H(n4), .Y(N855) );
  INVX1 U541 ( .A(n633), .Y(n637) );
  NAND43X1 U542 ( .B(c_ptr[3]), .C(n632), .D(n631), .A(n630), .Y(n633) );
  OAI211X1 U543 ( .C(n438), .D(n440), .A(n582), .B(n437), .Y(N868) );
  INVX1 U544 ( .A(sfr_psofs[14]), .Y(n438) );
  NAND32X1 U545 ( .B(c_ptr[4]), .C(n621), .A(n620), .Y(n628) );
  NAND21XL U546 ( .B(memaddr_c[5]), .A(c_adr[5]), .Y(n221) );
  NAND21X1 U547 ( .B(c_adr[7]), .A(memaddr_c[7]), .Y(n236) );
  GEN2XL U548 ( .D(n547), .E(n546), .C(d_psrd), .B(n630), .A(n545), .Y(N824)
         );
  NAND21X1 U549 ( .B(n544), .A(n543), .Y(n545) );
  NAND21X1 U550 ( .B(memaddr_c[7]), .A(c_adr[7]), .Y(n237) );
  AO21X1 U551 ( .B(n102), .C(n518), .A(n517), .Y(N823) );
  INVX1 U552 ( .A(n661), .Y(n517) );
  NAND32X1 U553 ( .B(n920), .C(n600), .A(n516), .Y(n518) );
  AOI32X1 U554 ( .A(mcu_psw), .B(n659), .C(n515), .D(n660), .E(n919), .Y(n516)
         );
  AO21X1 U555 ( .B(n86), .C(dbg_0d[7]), .A(n22), .Y(N582) );
  AO21X1 U556 ( .B(n85), .C(dbg_0e[7]), .A(n496), .Y(N590) );
  AO21X1 U557 ( .B(n84), .C(dbg_0f[7]), .A(n21), .Y(N598) );
  AO21X1 U558 ( .B(n83), .C(c_buf_16__7_), .A(n22), .Y(N606) );
  AO21X1 U559 ( .B(n82), .C(c_buf_17__7_), .A(n496), .Y(N614) );
  AO21X1 U560 ( .B(n82), .C(c_buf_18__7_), .A(n21), .Y(N622) );
  AO21X1 U561 ( .B(n81), .C(c_buf_19__7_), .A(n22), .Y(N630) );
  AO21X1 U562 ( .B(n80), .C(c_buf_20__7_), .A(n496), .Y(N638) );
  AO21X1 U563 ( .B(n79), .C(c_buf_21__7_), .A(n21), .Y(N646) );
  AO21X1 U564 ( .B(n86), .C(dbg_0c[7]), .A(n22), .Y(N574) );
  AO21X1 U565 ( .B(n90), .C(dbg_08[7]), .A(n496), .Y(N542) );
  AO21X1 U566 ( .B(n89), .C(dbg_09[7]), .A(n21), .Y(N550) );
  AO21X1 U567 ( .B(n88), .C(dbg_0a[7]), .A(n22), .Y(N558) );
  AO21X1 U568 ( .B(n95), .C(dbg_01[7]), .A(n496), .Y(N486) );
  AO21X1 U569 ( .B(n90), .C(dbg_07[7]), .A(n21), .Y(N534) );
  AO21X1 U570 ( .B(n87), .C(dbg_0b[7]), .A(n22), .Y(N566) );
  AO21X1 U571 ( .B(n94), .C(dbg_02[7]), .A(n496), .Y(N494) );
  AO21X1 U572 ( .B(n92), .C(dbg_05[7]), .A(n21), .Y(N518) );
  AO21X1 U573 ( .B(n96), .C(dbg_04[7]), .A(n22), .Y(N510) );
  AO21X1 U574 ( .B(n94), .C(dbg_03[7]), .A(n496), .Y(N502) );
  AO21X1 U575 ( .B(n91), .C(dbg_06[7]), .A(n21), .Y(N526) );
  AO21X1 U576 ( .B(n86), .C(dbg_0d[0]), .A(n28), .Y(N575) );
  AO21X1 U577 ( .B(n86), .C(dbg_0d[1]), .A(n18), .Y(N576) );
  AO21X1 U578 ( .B(n86), .C(dbg_0d[2]), .A(n14), .Y(N577) );
  AO21X1 U579 ( .B(n86), .C(dbg_0d[3]), .A(n11), .Y(N578) );
  AO21X1 U580 ( .B(n86), .C(dbg_0d[5]), .A(n8), .Y(N580) );
  AO21X1 U581 ( .B(n86), .C(dbg_0d[6]), .A(n5), .Y(N581) );
  AO21X1 U582 ( .B(n86), .C(dbg_0e[0]), .A(n29), .Y(N583) );
  AO21X1 U583 ( .B(n85), .C(dbg_0e[1]), .A(n19), .Y(N584) );
  AO21X1 U584 ( .B(n85), .C(dbg_0e[2]), .A(n15), .Y(N585) );
  AO21X1 U585 ( .B(n85), .C(dbg_0e[3]), .A(n12), .Y(N586) );
  AO21X1 U586 ( .B(n85), .C(dbg_0e[5]), .A(n9), .Y(N588) );
  AO21X1 U587 ( .B(n85), .C(dbg_0e[6]), .A(n6), .Y(N589) );
  AO21X1 U588 ( .B(n85), .C(dbg_0f[0]), .A(n503), .Y(N591) );
  AO21X1 U589 ( .B(n85), .C(dbg_0f[1]), .A(n502), .Y(N592) );
  AO21X1 U590 ( .B(n85), .C(dbg_0f[2]), .A(n501), .Y(N593) );
  AO21X1 U591 ( .B(n84), .C(dbg_0f[3]), .A(n500), .Y(N594) );
  AO21X1 U592 ( .B(n84), .C(dbg_0f[5]), .A(n498), .Y(N596) );
  AO21X1 U593 ( .B(n84), .C(dbg_0f[6]), .A(n497), .Y(N597) );
  AO21X1 U594 ( .B(n84), .C(c_buf_16__0_), .A(n28), .Y(N599) );
  AO21X1 U595 ( .B(n84), .C(c_buf_16__1_), .A(n18), .Y(N600) );
  AO21X1 U596 ( .B(n84), .C(c_buf_16__2_), .A(n14), .Y(N601) );
  AO21X1 U597 ( .B(n84), .C(c_buf_16__3_), .A(n11), .Y(N602) );
  AO21X1 U598 ( .B(n83), .C(c_buf_16__5_), .A(n8), .Y(N604) );
  AO21X1 U599 ( .B(n83), .C(c_buf_16__6_), .A(n5), .Y(N605) );
  AO21X1 U600 ( .B(n83), .C(c_buf_17__0_), .A(n29), .Y(N607) );
  AO21X1 U601 ( .B(n83), .C(c_buf_17__1_), .A(n19), .Y(N608) );
  AO21X1 U602 ( .B(n83), .C(c_buf_17__2_), .A(n15), .Y(N609) );
  AO21X1 U603 ( .B(n83), .C(c_buf_17__3_), .A(n12), .Y(N610) );
  AO21X1 U604 ( .B(n83), .C(c_buf_17__4_), .A(n26), .Y(N611) );
  AO21X1 U605 ( .B(n83), .C(c_buf_17__5_), .A(n9), .Y(N612) );
  AO21X1 U606 ( .B(n83), .C(c_buf_17__6_), .A(n6), .Y(N613) );
  AO21X1 U607 ( .B(n82), .C(c_buf_18__0_), .A(n503), .Y(N615) );
  AO21X1 U608 ( .B(n82), .C(c_buf_18__1_), .A(n502), .Y(N616) );
  AO21X1 U609 ( .B(n82), .C(c_buf_18__2_), .A(n501), .Y(N617) );
  AO21X1 U610 ( .B(n82), .C(c_buf_18__3_), .A(n500), .Y(N618) );
  AO21X1 U611 ( .B(n82), .C(c_buf_18__4_), .A(n27), .Y(N619) );
  AO21X1 U612 ( .B(n82), .C(c_buf_18__5_), .A(n498), .Y(N620) );
  AO21X1 U613 ( .B(n82), .C(c_buf_18__6_), .A(n497), .Y(N621) );
  AO21X1 U614 ( .B(n82), .C(c_buf_19__0_), .A(n28), .Y(N623) );
  AO21X1 U615 ( .B(n81), .C(c_buf_19__1_), .A(n18), .Y(N624) );
  AO21X1 U616 ( .B(n81), .C(c_buf_19__2_), .A(n14), .Y(N625) );
  AO21X1 U617 ( .B(n81), .C(c_buf_19__3_), .A(n11), .Y(N626) );
  AO21X1 U618 ( .B(n81), .C(c_buf_19__4_), .A(n499), .Y(N627) );
  AO21X1 U619 ( .B(n81), .C(c_buf_19__5_), .A(n8), .Y(N628) );
  AO21X1 U620 ( .B(n81), .C(c_buf_19__6_), .A(n5), .Y(N629) );
  AO21X1 U621 ( .B(n81), .C(c_buf_20__0_), .A(n29), .Y(N631) );
  AO21X1 U622 ( .B(n81), .C(c_buf_20__1_), .A(n19), .Y(N632) );
  AO21X1 U623 ( .B(n81), .C(c_buf_20__2_), .A(n15), .Y(N633) );
  AO21X1 U624 ( .B(n80), .C(c_buf_20__3_), .A(n12), .Y(N634) );
  AO21X1 U625 ( .B(n80), .C(c_buf_20__4_), .A(n26), .Y(N635) );
  AO21X1 U626 ( .B(n80), .C(c_buf_20__5_), .A(n9), .Y(N636) );
  AO21X1 U627 ( .B(n80), .C(c_buf_20__6_), .A(n6), .Y(N637) );
  AO21X1 U628 ( .B(n80), .C(c_buf_21__0_), .A(n503), .Y(N639) );
  AO21X1 U629 ( .B(n80), .C(c_buf_21__1_), .A(n502), .Y(N640) );
  AO21X1 U630 ( .B(n80), .C(c_buf_21__2_), .A(n501), .Y(N641) );
  AO21X1 U631 ( .B(n80), .C(c_buf_21__3_), .A(n500), .Y(N642) );
  AO21X1 U632 ( .B(n80), .C(c_buf_21__4_), .A(n27), .Y(N643) );
  AO21X1 U633 ( .B(n79), .C(c_buf_21__5_), .A(n498), .Y(N644) );
  AO21X1 U634 ( .B(n79), .C(c_buf_21__6_), .A(n497), .Y(N645) );
  AO21X1 U635 ( .B(n79), .C(c_buf_22__0_), .A(n28), .Y(N647) );
  AO21X1 U636 ( .B(n79), .C(c_buf_22__1_), .A(n18), .Y(N648) );
  AO21X1 U637 ( .B(n79), .C(c_buf_22__2_), .A(n14), .Y(N649) );
  AO21X1 U638 ( .B(n79), .C(c_buf_22__3_), .A(n11), .Y(N650) );
  AO21X1 U639 ( .B(n79), .C(c_buf_22__4_), .A(n499), .Y(N651) );
  AO21X1 U640 ( .B(n79), .C(c_buf_22__5_), .A(n8), .Y(N652) );
  AO21X1 U641 ( .B(n79), .C(c_buf_22__6_), .A(n5), .Y(N653) );
  AO21X1 U642 ( .B(n87), .C(dbg_0c[0]), .A(n29), .Y(N567) );
  AO21X1 U643 ( .B(n87), .C(dbg_0c[1]), .A(n19), .Y(N568) );
  AO21X1 U644 ( .B(n87), .C(dbg_0c[2]), .A(n15), .Y(N569) );
  AO21X1 U645 ( .B(n87), .C(dbg_0c[3]), .A(n12), .Y(N570) );
  AO21X1 U646 ( .B(n87), .C(dbg_0c[4]), .A(n26), .Y(N571) );
  AO21X1 U647 ( .B(n87), .C(dbg_0c[5]), .A(n9), .Y(N572) );
  AO21X1 U648 ( .B(n87), .C(dbg_0c[6]), .A(n6), .Y(N573) );
  AO21X1 U649 ( .B(n86), .C(dbg_0d[4]), .A(n27), .Y(N579) );
  AO21X1 U650 ( .B(n85), .C(dbg_0e[4]), .A(n499), .Y(N587) );
  AO21X1 U651 ( .B(n84), .C(dbg_0f[4]), .A(n26), .Y(N595) );
  AO21X1 U652 ( .B(n84), .C(c_buf_16__4_), .A(n27), .Y(N603) );
  AO21X1 U653 ( .B(n90), .C(dbg_08[0]), .A(n503), .Y(N535) );
  AO21X1 U654 ( .B(n90), .C(dbg_08[1]), .A(n502), .Y(N536) );
  AO21X1 U655 ( .B(n90), .C(dbg_08[2]), .A(n501), .Y(N537) );
  AO21X1 U656 ( .B(n90), .C(dbg_08[3]), .A(n500), .Y(N538) );
  AO21X1 U657 ( .B(n90), .C(dbg_08[4]), .A(n499), .Y(N539) );
  AO21X1 U658 ( .B(n90), .C(dbg_08[5]), .A(n498), .Y(N540) );
  AO21X1 U659 ( .B(n90), .C(dbg_08[6]), .A(n497), .Y(N541) );
  AO21X1 U660 ( .B(n90), .C(dbg_09[0]), .A(n28), .Y(N543) );
  AO21X1 U661 ( .B(n89), .C(dbg_09[1]), .A(n18), .Y(N544) );
  AO21X1 U662 ( .B(n89), .C(dbg_09[2]), .A(n14), .Y(N545) );
  AO21X1 U663 ( .B(n89), .C(dbg_09[3]), .A(n11), .Y(N546) );
  AO21X1 U664 ( .B(n89), .C(dbg_09[4]), .A(n26), .Y(N547) );
  AO21X1 U665 ( .B(n89), .C(dbg_09[5]), .A(n8), .Y(N548) );
  AO21X1 U666 ( .B(n89), .C(dbg_09[6]), .A(n5), .Y(N549) );
  AO21X1 U667 ( .B(n89), .C(dbg_0a[0]), .A(n29), .Y(N551) );
  AO21X1 U668 ( .B(n89), .C(dbg_0a[1]), .A(n19), .Y(N552) );
  AO21X1 U669 ( .B(n89), .C(dbg_0a[2]), .A(n15), .Y(N553) );
  AO21X1 U670 ( .B(n88), .C(dbg_0a[3]), .A(n12), .Y(N554) );
  AO21X1 U671 ( .B(n88), .C(dbg_0a[4]), .A(n27), .Y(N555) );
  AO21X1 U672 ( .B(n88), .C(dbg_0a[5]), .A(n9), .Y(N556) );
  AO21X1 U673 ( .B(n88), .C(dbg_0a[6]), .A(n6), .Y(N557) );
  AO21X1 U674 ( .B(n96), .C(dbg_01[0]), .A(n503), .Y(N479) );
  AO21X1 U675 ( .B(n96), .C(dbg_01[1]), .A(n502), .Y(N480) );
  AO21X1 U676 ( .B(n96), .C(dbg_01[2]), .A(n501), .Y(N481) );
  AO21X1 U677 ( .B(n96), .C(dbg_01[3]), .A(n500), .Y(N482) );
  AO21X1 U678 ( .B(n95), .C(dbg_01[5]), .A(n498), .Y(N484) );
  AO21X1 U679 ( .B(n95), .C(dbg_01[6]), .A(n497), .Y(N485) );
  AO21X1 U680 ( .B(n91), .C(dbg_07[0]), .A(n28), .Y(N527) );
  AO21X1 U681 ( .B(n91), .C(dbg_07[1]), .A(n18), .Y(N528) );
  AO21X1 U682 ( .B(n91), .C(dbg_07[2]), .A(n14), .Y(N529) );
  AO21X1 U683 ( .B(n91), .C(dbg_07[3]), .A(n11), .Y(N530) );
  AO21X1 U684 ( .B(n91), .C(dbg_07[4]), .A(n499), .Y(N531) );
  AO21X1 U685 ( .B(n91), .C(dbg_07[5]), .A(n8), .Y(N532) );
  AO21X1 U686 ( .B(n91), .C(dbg_07[6]), .A(n5), .Y(N533) );
  AO21X1 U687 ( .B(n88), .C(dbg_0b[0]), .A(n29), .Y(N559) );
  AO21X1 U688 ( .B(n88), .C(dbg_0b[1]), .A(n19), .Y(N560) );
  AO21X1 U689 ( .B(n88), .C(dbg_0b[2]), .A(n15), .Y(N561) );
  AO21X1 U690 ( .B(n88), .C(dbg_0b[3]), .A(n12), .Y(N562) );
  AO21X1 U691 ( .B(n88), .C(dbg_0b[4]), .A(n26), .Y(N563) );
  AO21X1 U692 ( .B(n87), .C(dbg_0b[5]), .A(n9), .Y(N564) );
  AO21X1 U693 ( .B(n87), .C(dbg_0b[6]), .A(n6), .Y(N565) );
  AO21X1 U694 ( .B(n95), .C(dbg_02[0]), .A(n503), .Y(N487) );
  AO21X1 U695 ( .B(n96), .C(dbg_05[0]), .A(n28), .Y(N511) );
  AO21X1 U696 ( .B(n95), .C(dbg_02[1]), .A(n502), .Y(N488) );
  AO21X1 U697 ( .B(n96), .C(dbg_05[1]), .A(n18), .Y(N512) );
  AO21X1 U698 ( .B(n95), .C(dbg_02[2]), .A(n501), .Y(N489) );
  AO21X1 U699 ( .B(n96), .C(dbg_05[2]), .A(n14), .Y(N513) );
  AO21X1 U700 ( .B(n95), .C(dbg_02[3]), .A(n500), .Y(N490) );
  AO21X1 U701 ( .B(n92), .C(dbg_05[3]), .A(n11), .Y(N514) );
  AO21X1 U702 ( .B(n95), .C(dbg_02[4]), .A(n27), .Y(N491) );
  AO21X1 U703 ( .B(n92), .C(dbg_05[4]), .A(n499), .Y(N515) );
  AO21X1 U704 ( .B(n95), .C(dbg_02[5]), .A(n498), .Y(N492) );
  AO21X1 U705 ( .B(n92), .C(dbg_05[5]), .A(n8), .Y(N516) );
  AO21X1 U706 ( .B(n95), .C(dbg_02[6]), .A(n497), .Y(N493) );
  AO21X1 U707 ( .B(n92), .C(dbg_05[6]), .A(n5), .Y(N517) );
  AO21X1 U708 ( .B(n94), .C(dbg_04[0]), .A(n29), .Y(N503) );
  AO21X1 U709 ( .B(n504), .C(dbg_04[1]), .A(n19), .Y(N504) );
  AO21X1 U710 ( .B(n504), .C(dbg_04[2]), .A(n15), .Y(N505) );
  AO21X1 U711 ( .B(n504), .C(dbg_04[3]), .A(n12), .Y(N506) );
  AO21X1 U712 ( .B(n504), .C(dbg_04[5]), .A(n9), .Y(N508) );
  AO21X1 U713 ( .B(n504), .C(dbg_04[6]), .A(n6), .Y(N509) );
  AO21X1 U714 ( .B(n94), .C(dbg_03[0]), .A(n503), .Y(N495) );
  AO21X1 U715 ( .B(n92), .C(dbg_06[0]), .A(n28), .Y(N519) );
  AO21X1 U716 ( .B(n94), .C(dbg_03[1]), .A(n502), .Y(N496) );
  AO21X1 U717 ( .B(n92), .C(dbg_06[1]), .A(n18), .Y(N520) );
  AO21X1 U718 ( .B(n94), .C(dbg_03[2]), .A(n501), .Y(N497) );
  AO21X1 U719 ( .B(n92), .C(dbg_06[2]), .A(n14), .Y(N521) );
  AO21X1 U720 ( .B(n94), .C(dbg_03[3]), .A(n500), .Y(N498) );
  AO21X1 U721 ( .B(n92), .C(dbg_06[3]), .A(n11), .Y(N522) );
  AO21X1 U722 ( .B(n94), .C(dbg_03[4]), .A(n26), .Y(N499) );
  AO21X1 U723 ( .B(n92), .C(dbg_06[4]), .A(n27), .Y(N523) );
  AO21X1 U724 ( .B(n94), .C(dbg_03[5]), .A(n498), .Y(N500) );
  AO21X1 U725 ( .B(n91), .C(dbg_06[5]), .A(n8), .Y(N524) );
  AO21X1 U726 ( .B(n94), .C(dbg_03[6]), .A(n497), .Y(N501) );
  AO21X1 U727 ( .B(n91), .C(dbg_06[6]), .A(n5), .Y(N525) );
  AO21X1 U728 ( .B(n96), .C(dbg_01[4]), .A(n499), .Y(N483) );
  AO21X1 U729 ( .B(n96), .C(dbg_04[4]), .A(n26), .Y(N507) );
  OAI21X1 U730 ( .B(n530), .C(n686), .A(n529), .Y(N822) );
  AND4X1 U731 ( .A(n583), .B(n673), .C(n688), .D(n524), .Y(n530) );
  GEN2XL U732 ( .D(n632), .E(n528), .C(n527), .B(n564), .A(n621), .Y(n529) );
  AOI221XL U733 ( .A(n675), .B(mcu_psw), .C(n924), .D(n919), .E(n613), .Y(n524) );
  INVX1 U734 ( .A(n622), .Y(n623) );
  NAND32X1 U735 ( .B(c_ptr[2]), .C(n628), .A(n629), .Y(n622) );
  INVX1 U736 ( .A(n634), .Y(n636) );
  NAND21X1 U737 ( .B(c_ptr[2]), .A(n637), .Y(n634) );
  NAND21X1 U738 ( .B(memaddr_c[9]), .A(c_adr[9]), .Y(n375) );
  GEN3XL U739 ( .F(n102), .G(n558), .E(n557), .D(n551), .C(n550), .B(n549), 
        .A(n548), .Y(n648) );
  AND2X1 U740 ( .A(n30), .B(n557), .Y(n550) );
  NAND21X1 U741 ( .B(c_adr[9]), .A(memaddr_c[9]), .Y(n374) );
  MUX2IX1 U742 ( .D0(n67), .D1(n68), .S(n607), .Y(n566) );
  NAND2X1 U743 ( .A(pmem_re), .B(n602), .Y(n67) );
  NAND2X1 U744 ( .A(n565), .B(n102), .Y(n68) );
  NOR21XL U745 ( .B(n509), .A(n69), .Y(N846) );
  XNOR2XL U746 ( .A(c_ptr[4]), .B(n508), .Y(n69) );
  NAND21X1 U747 ( .B(c_adr[13]), .A(memaddr_c[13]), .Y(n228) );
  NAND21X1 U748 ( .B(memaddr_c[14]), .A(c_adr[14]), .Y(n345) );
  NAND21X1 U749 ( .B(c_adr[10]), .A(memaddr_c[10]), .Y(n346) );
  MUX2X1 U750 ( .D0(n324), .D1(n315), .S(memaddr_c[11]), .Y(n325) );
  AND2X1 U751 ( .A(c_adr[11]), .B(n314), .Y(n315) );
  AO21X1 U752 ( .B(n314), .C(n305), .A(n304), .Y(n324) );
  INVX1 U753 ( .A(n294), .Y(n304) );
  MUX2IX1 U754 ( .D0(n70), .D1(n228), .S(n250), .Y(n230) );
  XNOR2XL U755 ( .A(n231), .B(c_adr[13]), .Y(n70) );
  INVX1 U756 ( .A(n181), .Y(n335) );
  NAND21X1 U757 ( .B(c_adr[11]), .A(memaddr_c[11]), .Y(n181) );
  AND2X1 U758 ( .A(c_adr[13]), .B(n231), .Y(n203) );
  AND2X1 U759 ( .A(hit_ps_c), .B(mcu_psr_c), .Y(n549) );
  NAND21X1 U760 ( .B(c_adr[14]), .A(memaddr_c[14]), .Y(n240) );
  OAI22X1 U761 ( .A(n101), .B(n583), .C(mcu_psw), .D(n662), .Y(n585) );
  INVX1 U762 ( .A(n255), .Y(o_bkp_hold) );
  INVX1 U763 ( .A(memaddr[12]), .Y(n930) );
  XNOR2XL U764 ( .A(memaddr[7]), .B(bkpt_pc[7]), .Y(n402) );
  XNOR2XL U765 ( .A(memaddr[0]), .B(bkpt_pc[0]), .Y(n411) );
  XOR2X1 U766 ( .A(bkpt_pc[9]), .B(memaddr[9]), .Y(n398) );
  XOR2X1 U767 ( .A(bkpt_pc[8]), .B(memaddr[8]), .Y(n397) );
  XOR2X1 U768 ( .A(bkpt_pc[13]), .B(memaddr[13]), .Y(n405) );
  XNOR2XL U769 ( .A(bkpt_pc[12]), .B(n930), .Y(n406) );
  MUX2X1 U770 ( .D0(n108), .D1(n24), .S(n602), .Y(n649) );
  AND2X1 U771 ( .A(n568), .B(n606), .Y(n108) );
  NAND2X1 U772 ( .A(n393), .B(n394), .Y(n255) );
  NOR4XL U773 ( .A(n395), .B(n396), .C(n397), .D(n398), .Y(n394) );
  NOR4XL U774 ( .A(n403), .B(n404), .C(n405), .D(n406), .Y(n393) );
  NAND32X1 U775 ( .B(n727), .C(un_hold), .A(bkpt_ena), .Y(n396) );
  MUX2X1 U776 ( .D0(n568), .D1(pmem_pgm), .S(n562), .Y(n644) );
  AND2X1 U777 ( .A(n561), .B(n569), .Y(n562) );
  INVX1 U778 ( .A(n559), .Y(n561) );
  NAND4X1 U779 ( .A(n410), .B(n411), .C(n412), .D(n413), .Y(n403) );
  XNOR2XL U780 ( .A(memaddr[10]), .B(bkpt_pc[10]), .Y(n410) );
  XNOR2XL U781 ( .A(memaddr[5]), .B(bkpt_pc[5]), .Y(n412) );
  XNOR2XL U782 ( .A(memaddr[4]), .B(bkpt_pc[4]), .Y(n413) );
  NAND4X1 U783 ( .A(n399), .B(n400), .C(n401), .D(n402), .Y(n395) );
  XNOR2XL U784 ( .A(memaddr[1]), .B(bkpt_pc[1]), .Y(n400) );
  XNOR2XL U785 ( .A(memaddr[3]), .B(bkpt_pc[3]), .Y(n399) );
  XNOR2XL U786 ( .A(memaddr[6]), .B(bkpt_pc[6]), .Y(n401) );
  NAND3X1 U787 ( .A(n407), .B(n408), .C(n409), .Y(n404) );
  XNOR2XL U788 ( .A(memaddr[14]), .B(bkpt_pc[14]), .Y(n407) );
  XNOR2XL U789 ( .A(memaddr[11]), .B(bkpt_pc[11]), .Y(n409) );
  XNOR2XL U790 ( .A(memaddr[2]), .B(bkpt_pc[2]), .Y(n408) );
  NOR43XL U791 ( .B(n918), .C(n917), .D(n916), .A(n915), .Y(n264) );
  NAND21X1 U792 ( .B(n287), .A(dbg_08[7]), .Y(n918) );
  NAND21X1 U793 ( .B(n289), .A(dbg_09[7]), .Y(n916) );
  NAND21X1 U794 ( .B(n288), .A(dbg_07[7]), .Y(n917) );
  NAND31X1 U795 ( .C(n914), .A(n913), .B(n912), .Y(n915) );
  NAND21X1 U796 ( .B(n286), .A(dbg_0a[7]), .Y(n913) );
  NAND21X1 U797 ( .B(n285), .A(dbg_0b[7]), .Y(n912) );
  AND2X1 U798 ( .A(n282), .B(dbg_06[7]), .Y(n914) );
  XNOR2XL U799 ( .A(n387), .B(n388), .Y(n372) );
  XOR2X1 U800 ( .A(n731), .B(memaddr[4]), .Y(n387) );
  AO21X1 U801 ( .B(n734), .C(n738), .A(n736), .Y(n735) );
  OAI222XL U802 ( .A(n274), .B(n900), .C(n273), .D(n899), .E(n275), .F(n898), 
        .Y(n268) );
  INVX1 U803 ( .A(c_buf_17__7_), .Y(n900) );
  INVX1 U804 ( .A(c_buf_16__7_), .Y(n899) );
  INVX1 U805 ( .A(dbg_0f[7]), .Y(n898) );
  OAI222XL U806 ( .A(n277), .B(n897), .C(n276), .D(n896), .E(n278), .F(n895), 
        .Y(n267) );
  INVX1 U807 ( .A(c_buf_20__7_), .Y(n897) );
  INVX1 U808 ( .A(c_buf_19__7_), .Y(n896) );
  INVX1 U809 ( .A(c_buf_18__7_), .Y(n895) );
  INVX1 U810 ( .A(n728), .Y(n922) );
  NAND21X1 U811 ( .B(memaddr[0]), .A(c_adr[0]), .Y(n728) );
  INVX1 U812 ( .A(r_rdy), .Y(n727) );
  INVX1 U813 ( .A(memaddr[2]), .Y(n935) );
  XOR2X1 U814 ( .A(n385), .B(n71), .Y(n373) );
  XNOR2XL U815 ( .A(memaddr[2]), .B(c_adr[2]), .Y(n71) );
  OAI22X1 U816 ( .A(c_adr[1]), .B(n730), .C(n922), .D(n729), .Y(n385) );
  AND2X1 U817 ( .A(c_adr[1]), .B(n730), .Y(n729) );
  INVX1 U818 ( .A(memaddr[1]), .Y(n730) );
  OAI222XL U819 ( .A(n274), .B(n761), .C(n273), .D(n760), .E(n275), .F(n759), 
        .Y(n352) );
  INVX1 U820 ( .A(c_buf_17__1_), .Y(n761) );
  INVX1 U821 ( .A(c_buf_16__1_), .Y(n760) );
  INVX1 U822 ( .A(dbg_0f[1]), .Y(n759) );
  OAI222XL U823 ( .A(n271), .B(n765), .C(n270), .D(n764), .E(n272), .F(n763), 
        .Y(n353) );
  INVX1 U824 ( .A(dbg_0e[1]), .Y(n765) );
  INVX1 U825 ( .A(dbg_0d[1]), .Y(n764) );
  INVX1 U826 ( .A(dbg_0c[1]), .Y(n763) );
  OAI222XL U827 ( .A(n271), .B(n903), .C(n270), .D(n902), .E(n272), .F(n901), 
        .Y(n269) );
  INVX1 U828 ( .A(dbg_0e[7]), .Y(n903) );
  INVX1 U829 ( .A(dbg_0d[7]), .Y(n902) );
  INVX1 U830 ( .A(dbg_0c[7]), .Y(n901) );
  OAI222XL U831 ( .A(n277), .B(n758), .C(n276), .D(n757), .E(n278), .F(n756), 
        .Y(n351) );
  INVX1 U832 ( .A(c_buf_20__1_), .Y(n758) );
  INVX1 U833 ( .A(c_buf_19__1_), .Y(n757) );
  INVX1 U834 ( .A(c_buf_18__1_), .Y(n756) );
  OAI222XL U835 ( .A(n280), .B(n755), .C(n279), .D(n754), .E(n281), .F(n753), 
        .Y(n350) );
  INVX1 U836 ( .A(c_buf_22__1_), .Y(n754) );
  INVX1 U837 ( .A(c_buf_21__1_), .Y(n753) );
  OAI222XL U838 ( .A(n280), .B(n894), .C(n279), .D(n893), .E(n281), .F(n892), 
        .Y(n266) );
  INVX1 U839 ( .A(c_buf_22__7_), .Y(n893) );
  INVX1 U840 ( .A(c_buf_21__7_), .Y(n892) );
  MUX2X1 U841 ( .D0(r_rdy), .D1(o_ofs_inc), .S(mcu_psw), .Y(mempsack) );
  OAI211X1 U842 ( .C(n40), .D(n715), .A(n349), .B(n714), .Y(n726) );
  OA22X1 U843 ( .A(n37), .B(n713), .C(n905), .D(n712), .Y(n714) );
  NOR4XL U844 ( .A(n350), .B(n351), .C(n352), .D(n353), .Y(n349) );
  INVX1 U845 ( .A(dbg_02[1]), .Y(n713) );
  NAND21X1 U846 ( .B(n439), .A(memaddr[14]), .Y(n582) );
  AO21X1 U847 ( .B(memaddr[0]), .C(n740), .A(n922), .Y(n934) );
  NAND21X1 U848 ( .B(n578), .A(mcu_psw), .Y(n439) );
  XOR2X1 U849 ( .A(n72), .B(n922), .Y(n380) );
  XNOR2XL U850 ( .A(n730), .B(c_adr[1]), .Y(n72) );
  NAND21X1 U851 ( .B(cs_ft[0]), .A(cs_ft[1]), .Y(n111) );
  INVX1 U852 ( .A(memaddr[3]), .Y(n936) );
  OAI222XL U853 ( .A(n274), .B(n849), .C(n273), .D(n848), .E(n275), .F(n847), 
        .Y(n312) );
  INVX1 U854 ( .A(c_buf_17__5_), .Y(n849) );
  INVX1 U855 ( .A(c_buf_16__5_), .Y(n848) );
  INVX1 U856 ( .A(dbg_0f[5]), .Y(n847) );
  OAI222XL U857 ( .A(n274), .B(n749), .C(n273), .D(n748), .E(n275), .F(n747), 
        .Y(n362) );
  INVX1 U858 ( .A(c_buf_17__0_), .Y(n749) );
  INVX1 U859 ( .A(c_buf_16__0_), .Y(n748) );
  INVX1 U860 ( .A(dbg_0f[0]), .Y(n747) );
  OAI222XL U861 ( .A(n274), .B(n824), .C(n273), .D(n823), .E(n275), .F(n822), 
        .Y(n322) );
  INVX1 U862 ( .A(c_buf_17__4_), .Y(n824) );
  INVX1 U863 ( .A(c_buf_16__4_), .Y(n823) );
  INVX1 U864 ( .A(dbg_0f[4]), .Y(n822) );
  OAI222XL U865 ( .A(n274), .B(n875), .C(n273), .D(n873), .E(n275), .F(n872), 
        .Y(n302) );
  INVX1 U866 ( .A(c_buf_17__6_), .Y(n875) );
  INVX1 U867 ( .A(c_buf_16__6_), .Y(n873) );
  INVX1 U868 ( .A(dbg_0f[6]), .Y(n872) );
  OAI222XL U869 ( .A(n274), .B(n799), .C(n273), .D(n798), .E(n275), .F(n797), 
        .Y(n332) );
  INVX1 U870 ( .A(c_buf_17__3_), .Y(n799) );
  INVX1 U871 ( .A(c_buf_16__3_), .Y(n798) );
  INVX1 U872 ( .A(dbg_0f[3]), .Y(n797) );
  OAI222XL U873 ( .A(n274), .B(n774), .C(n273), .D(n773), .E(n275), .F(n772), 
        .Y(n342) );
  INVX1 U874 ( .A(c_buf_17__2_), .Y(n774) );
  INVX1 U875 ( .A(c_buf_16__2_), .Y(n773) );
  INVX1 U876 ( .A(dbg_0f[2]), .Y(n772) );
  INVX1 U877 ( .A(cs_ft[3]), .Y(n511) );
  INVX1 U878 ( .A(c_adr[2]), .Y(n732) );
  INVX1 U879 ( .A(test_so1), .Y(pmem_csb) );
  NAND31X1 U880 ( .C(n861), .A(n860), .B(n859), .Y(n862) );
  NAND21X1 U881 ( .B(n286), .A(dbg_0a[5]), .Y(n860) );
  NAND21X1 U882 ( .B(n285), .A(dbg_0b[5]), .Y(n859) );
  AND2X1 U883 ( .A(n282), .B(dbg_06[5]), .Y(n861) );
  NAND31X1 U884 ( .C(n836), .A(n835), .B(n834), .Y(n837) );
  NAND21X1 U885 ( .B(n286), .A(dbg_0a[4]), .Y(n835) );
  NAND21X1 U886 ( .B(n285), .A(dbg_0b[4]), .Y(n834) );
  AND2X1 U887 ( .A(n282), .B(dbg_06[4]), .Y(n836) );
  NAND31X1 U888 ( .C(n811), .A(n810), .B(n809), .Y(n812) );
  NAND21X1 U889 ( .B(n286), .A(dbg_0a[3]), .Y(n810) );
  NAND21X1 U890 ( .B(n285), .A(dbg_0b[3]), .Y(n809) );
  AND2X1 U891 ( .A(n282), .B(dbg_06[3]), .Y(n811) );
  NAND31X1 U892 ( .C(n786), .A(n785), .B(n784), .Y(n787) );
  NAND21X1 U893 ( .B(n286), .A(dbg_0a[2]), .Y(n785) );
  NAND21X1 U894 ( .B(n285), .A(dbg_0b[2]), .Y(n784) );
  AND2X1 U895 ( .A(n282), .B(dbg_06[2]), .Y(n786) );
  NAND21X1 U896 ( .B(d_psrd), .A(n630), .Y(n434) );
  NAND21X1 U897 ( .B(n704), .A(n703), .Y(n705) );
  NOR21XL U898 ( .B(dbg_07[0]), .A(n288), .Y(n704) );
  AOI21BBXL U899 ( .B(n702), .C(n287), .A(n701), .Y(n703) );
  INVX1 U900 ( .A(dbg_08[0]), .Y(n702) );
  NAND21X1 U901 ( .B(n38), .A(dbg_03[0]), .Y(n696) );
  NAND21X1 U902 ( .B(n39), .A(dbg_04[0]), .Y(n695) );
  NAND21X1 U903 ( .B(n37), .A(dbg_02[0]), .Y(n700) );
  NAND21X1 U904 ( .B(n287), .A(dbg_08[5]), .Y(n865) );
  NAND21X1 U905 ( .B(n287), .A(dbg_08[4]), .Y(n840) );
  NAND21X1 U906 ( .B(n287), .A(dbg_08[6]), .Y(n891) );
  NAND21X1 U907 ( .B(n289), .A(dbg_09[0]), .Y(n708) );
  NAND21X1 U908 ( .B(n287), .A(dbg_08[3]), .Y(n815) );
  NAND21X1 U909 ( .B(n287), .A(dbg_08[2]), .Y(n790) );
  NAND21X1 U910 ( .B(n40), .A(rd_buf[0]), .Y(n699) );
  NAND21X1 U911 ( .B(n285), .A(dbg_0b[0]), .Y(n707) );
  NAND21X1 U912 ( .B(n288), .A(dbg_07[5]), .Y(n864) );
  NAND21X1 U913 ( .B(n288), .A(dbg_07[4]), .Y(n839) );
  NAND21X1 U914 ( .B(n288), .A(dbg_07[6]), .Y(n890) );
  NAND21X1 U915 ( .B(n288), .A(dbg_07[3]), .Y(n814) );
  NAND21X1 U916 ( .B(n288), .A(dbg_07[2]), .Y(n789) );
  NAND21X1 U917 ( .B(n289), .A(dbg_09[5]), .Y(n863) );
  NAND21X1 U918 ( .B(n289), .A(dbg_09[4]), .Y(n838) );
  NAND21X1 U919 ( .B(n289), .A(dbg_09[6]), .Y(n889) );
  NAND21X1 U920 ( .B(n286), .A(dbg_0a[0]), .Y(n706) );
  NAND21X1 U921 ( .B(n289), .A(dbg_09[3]), .Y(n813) );
  NAND21X1 U922 ( .B(n289), .A(dbg_09[2]), .Y(n788) );
  INVX1 U923 ( .A(cs_ft[2]), .Y(n513) );
  AND2X1 U924 ( .A(dbg_06[0]), .B(n282), .Y(n701) );
  AND2X1 U925 ( .A(dbg_01[0]), .B(n295), .Y(n698) );
  INVX1 U926 ( .A(c_adr[0]), .Y(n740) );
  NAND31X1 U927 ( .C(n887), .A(n886), .B(n885), .Y(n888) );
  NAND21X1 U928 ( .B(n286), .A(dbg_0a[6]), .Y(n886) );
  NAND21X1 U929 ( .B(n285), .A(dbg_0b[6]), .Y(n885) );
  AND2X1 U930 ( .A(n282), .B(dbg_06[6]), .Y(n887) );
  AND2X1 U931 ( .A(dbg_05[0]), .B(n291), .Y(n697) );
  INVX1 U932 ( .A(c_adr[4]), .Y(n731) );
  INVX1 U933 ( .A(c_adr[3]), .Y(n739) );
  OR2X1 U934 ( .A(pmem_a[10]), .B(pmem_a[11]), .Y(n445) );
  OR2X1 U935 ( .A(pmem_a[12]), .B(pmem_a[13]), .Y(n446) );
  AOI21BBXL U936 ( .B(wspp_cnt_3_), .C(n923), .A(test_so2), .Y(n467) );
  AO21X1 U937 ( .B(n102), .C(n112), .A(n557), .Y(N821) );
  NAND32X1 U938 ( .B(n110), .C(n541), .A(n612), .Y(n112) );
  INVX1 U939 ( .A(n672), .Y(n110) );
  OAI31XL U940 ( .A(n929), .B(wr_buf[0]), .C(n924), .D(n940), .Y(n541) );
  AOI221XL U941 ( .A(n465), .B(test_so2), .C(wspp_cnt_5_), .D(n676), .E(n923), 
        .Y(n677) );
  XNOR2XL U942 ( .A(wspp_cnt_5_), .B(wspp_cnt_3_), .Y(n465) );
  INVX1 U943 ( .A(n603), .Y(n923) );
  NAND43X1 U944 ( .B(wspp_cnt_3_), .C(wspp_cnt_5_), .D(test_so2), .A(n676), 
        .Y(n603) );
  MUX2X1 U945 ( .D0(n450), .D1(n449), .S(adr_p[14]), .Y(n682) );
  NAND5XL U946 ( .A(pmem_a[9]), .B(n450), .C(n73), .D(n448), .E(n447), .Y(n449) );
  INVX1 U947 ( .A(adr_p[13]), .Y(n450) );
  INVX1 U948 ( .A(n445), .Y(n448) );
  NOR21XL U949 ( .B(r_multi), .A(n677), .Y(n681) );
  OA21X1 U950 ( .B(n467), .C(wspp_cnt_4_), .A(n678), .Y(n680) );
  NOR2X1 U951 ( .A(pmem_a[14]), .B(pmem_a[15]), .Y(n73) );
  INVX1 U952 ( .A(rd_buf[7]), .Y(n907) );
  INVX1 U953 ( .A(wr_buf[7]), .Y(n894) );
  INVX1 U954 ( .A(dbg_03[7]), .Y(n908) );
  INVX1 U955 ( .A(dbg_01[7]), .Y(n904) );
  INVX1 U956 ( .A(dbg_05[7]), .Y(n909) );
  INVX1 U957 ( .A(dbg_02[7]), .Y(n906) );
  INVX1 U958 ( .A(dbg_04[7]), .Y(n911) );
  NAND21X1 U959 ( .B(n694), .A(n907), .Y(d_inst[7]) );
  NAND32X1 U960 ( .B(cs_ft[1]), .C(cs_ft[0]), .A(n510), .Y(n940) );
  MUX2X1 U961 ( .D0(sfr_psr), .D1(o_ofs_inc), .S(d_psrd), .Y(sfr_psrack) );
  AO21X1 U962 ( .B(adr_p[14]), .C(n444), .A(adr_p[13]), .Y(n475) );
  NAND43X1 U963 ( .B(pmem_a[9]), .C(n445), .D(n446), .A(n73), .Y(n444) );
  NAND21X1 U964 ( .B(cs_ft[2]), .A(n511), .Y(n519) );
  NAND21X1 U965 ( .B(cs_ft[1]), .A(cs_ft[0]), .Y(n512) );
  INVX1 U966 ( .A(n455), .Y(n510) );
  NAND21X1 U967 ( .B(n511), .A(cs_ft[2]), .Y(n455) );
  OR2X1 U968 ( .A(cs_ft[3]), .B(n111), .Y(n684) );
  NAND32X1 U969 ( .B(n522), .C(n521), .A(n520), .Y(n673) );
  INVX1 U970 ( .A(cs_ft[1]), .Y(n521) );
  INVX1 U971 ( .A(n519), .Y(n520) );
  INVX1 U972 ( .A(cs_ft[0]), .Y(n522) );
  INVX1 U973 ( .A(wspp_cnt_4_), .Y(n676) );
  INVX1 U974 ( .A(wr_buf[1]), .Y(n755) );
  INVX1 U975 ( .A(pmem_re), .Y(n678) );
  INVX1 U976 ( .A(c_buf_20__0_), .Y(n746) );
  INVX1 U977 ( .A(dbg_0e[0]), .Y(n752) );
  INVX1 U978 ( .A(dbg_0e[2]), .Y(n777) );
  INVX1 U979 ( .A(c_buf_19__0_), .Y(n745) );
  INVX1 U980 ( .A(dbg_0d[0]), .Y(n751) );
  INVX1 U981 ( .A(c_buf_22__0_), .Y(n742) );
  INVX1 U982 ( .A(dbg_0d[6]), .Y(n877) );
  INVX1 U983 ( .A(dbg_0d[3]), .Y(n801) );
  INVX1 U984 ( .A(c_buf_19__2_), .Y(n770) );
  INVX1 U985 ( .A(dbg_0d[2]), .Y(n776) );
  INVX1 U986 ( .A(c_buf_18__0_), .Y(n744) );
  INVX1 U987 ( .A(dbg_0c[0]), .Y(n750) );
  INVX1 U988 ( .A(c_buf_21__0_), .Y(n741) );
  INVX1 U989 ( .A(c_buf_18__6_), .Y(n869) );
  INVX1 U990 ( .A(dbg_0c[6]), .Y(n876) );
  INVX1 U991 ( .A(dbg_0c[3]), .Y(n800) );
  INVX1 U992 ( .A(c_buf_18__2_), .Y(n769) );
  INVX1 U993 ( .A(dbg_0c[2]), .Y(n775) );
  NAND21X1 U994 ( .B(n540), .A(n539), .Y(n588) );
  AND4X1 U995 ( .A(sfr_psw), .B(n538), .C(n537), .D(n536), .Y(n540) );
  INVX1 U996 ( .A(dummy[0]), .Y(n536) );
  NAND43X1 U997 ( .B(cs_ft[0]), .C(cs_ft[2]), .D(cs_ft[1]), .A(cs_ft[3]), .Y(
        n671) );
  INVX1 U998 ( .A(n105), .Y(n109) );
  NAND32X1 U999 ( .B(cs_ft[1]), .C(cs_ft[3]), .A(n522), .Y(n105) );
  INVX1 U1000 ( .A(rd_buf[1]), .Y(n715) );
  INVX1 U1001 ( .A(rd_buf[2]), .Y(n780) );
  INVX1 U1002 ( .A(wr_buf[0]), .Y(n743) );
  INVX1 U1003 ( .A(wr_buf[6]), .Y(n868) );
  INVX1 U1004 ( .A(wr_buf[2]), .Y(n768) );
  INVX1 U1005 ( .A(wr_buf[3]), .Y(n793) );
  INVX1 U1006 ( .A(wr_buf[4]), .Y(n818) );
  INVX1 U1007 ( .A(wr_buf[5]), .Y(n843) );
  INVX1 U1008 ( .A(dbg_08[1]), .Y(n719) );
  INVX1 U1009 ( .A(dbg_05[1]), .Y(n716) );
  INVX1 U1010 ( .A(dbg_0b[1]), .Y(n723) );
  INVX1 U1011 ( .A(dbg_05[4]), .Y(n831) );
  INVX1 U1012 ( .A(dbg_03[6]), .Y(n882) );
  INVX1 U1013 ( .A(dbg_01[6]), .Y(n879) );
  INVX1 U1014 ( .A(dbg_03[3]), .Y(n806) );
  INVX1 U1015 ( .A(dbg_01[3]), .Y(n803) );
  INVX1 U1016 ( .A(dbg_03[2]), .Y(n781) );
  INVX1 U1017 ( .A(dbg_01[2]), .Y(n778) );
  INVX1 U1018 ( .A(c_buf_20__5_), .Y(n846) );
  INVX1 U1019 ( .A(dbg_0e[5]), .Y(n852) );
  INVX1 U1020 ( .A(c_buf_20__4_), .Y(n821) );
  INVX1 U1021 ( .A(dbg_0e[4]), .Y(n827) );
  INVX1 U1022 ( .A(c_buf_20__6_), .Y(n871) );
  INVX1 U1023 ( .A(dbg_0e[6]), .Y(n878) );
  INVX1 U1024 ( .A(c_buf_20__3_), .Y(n796) );
  INVX1 U1025 ( .A(dbg_0e[3]), .Y(n802) );
  INVX1 U1026 ( .A(c_buf_20__2_), .Y(n771) );
  INVX1 U1027 ( .A(dbg_06[1]), .Y(n720) );
  INVX1 U1028 ( .A(dbg_03[1]), .Y(n717) );
  INVX1 U1029 ( .A(dbg_09[1]), .Y(n724) );
  INVX1 U1030 ( .A(dbg_05[6]), .Y(n883) );
  INVX1 U1031 ( .A(dbg_02[6]), .Y(n880) );
  INVX1 U1032 ( .A(dbg_05[3]), .Y(n807) );
  INVX1 U1033 ( .A(dbg_02[3]), .Y(n804) );
  INVX1 U1034 ( .A(dbg_05[2]), .Y(n782) );
  INVX1 U1035 ( .A(dbg_02[2]), .Y(n779) );
  INVX1 U1036 ( .A(dbg_07[1]), .Y(n722) );
  INVX1 U1037 ( .A(dbg_04[1]), .Y(n718) );
  INVX1 U1038 ( .A(dbg_0a[1]), .Y(n725) );
  INVX1 U1039 ( .A(dbg_04[6]), .Y(n884) );
  INVX1 U1040 ( .A(dbg_04[2]), .Y(n783) );
  INVX1 U1041 ( .A(c_buf_19__5_), .Y(n845) );
  INVX1 U1042 ( .A(dbg_0d[5]), .Y(n851) );
  INVX1 U1043 ( .A(c_buf_22__5_), .Y(n842) );
  INVX1 U1044 ( .A(c_buf_19__4_), .Y(n820) );
  INVX1 U1045 ( .A(dbg_0d[4]), .Y(n826) );
  INVX1 U1046 ( .A(c_buf_22__4_), .Y(n817) );
  INVX1 U1047 ( .A(c_buf_19__6_), .Y(n870) );
  INVX1 U1048 ( .A(c_buf_22__6_), .Y(n867) );
  INVX1 U1049 ( .A(c_buf_19__3_), .Y(n795) );
  INVX1 U1050 ( .A(c_buf_22__3_), .Y(n792) );
  INVX1 U1051 ( .A(c_buf_22__2_), .Y(n767) );
  INVX1 U1052 ( .A(dbg_01[1]), .Y(n712) );
  INVX1 U1053 ( .A(c_buf_18__5_), .Y(n844) );
  INVX1 U1054 ( .A(dbg_0c[5]), .Y(n850) );
  INVX1 U1055 ( .A(c_buf_21__5_), .Y(n841) );
  INVX1 U1056 ( .A(c_buf_18__4_), .Y(n819) );
  INVX1 U1057 ( .A(dbg_0c[4]), .Y(n825) );
  INVX1 U1058 ( .A(c_buf_21__4_), .Y(n816) );
  INVX1 U1059 ( .A(c_buf_21__6_), .Y(n866) );
  INVX1 U1060 ( .A(c_buf_18__3_), .Y(n794) );
  INVX1 U1061 ( .A(c_buf_21__3_), .Y(n791) );
  INVX1 U1062 ( .A(c_buf_21__2_), .Y(n766) );
  NAND21X1 U1063 ( .B(n694), .A(n780), .Y(d_inst[2]) );
  NAND21X1 U1064 ( .B(n694), .A(n855), .Y(d_inst[5]) );
  NAND21X1 U1065 ( .B(n694), .A(n805), .Y(d_inst[3]) );
  AND2X1 U1066 ( .A(d_psrd), .B(rd_buf[4]), .Y(d_inst[4]) );
  NAND21X1 U1067 ( .B(n694), .A(n881), .Y(d_inst[6]) );
  NAND21X1 U1068 ( .B(n694), .A(n715), .Y(d_inst[1]) );
  AND2X1 U1069 ( .A(d_psrd), .B(rd_buf[0]), .Y(d_inst[0]) );
  INVX1 U1070 ( .A(rd_buf[5]), .Y(n855) );
  INVX1 U1071 ( .A(rd_buf[6]), .Y(n881) );
  INVX1 U1072 ( .A(rd_buf[3]), .Y(n805) );
  INVX1 U1073 ( .A(rd_buf[4]), .Y(n829) );
  INVX1 U1074 ( .A(dbg_03[5]), .Y(n856) );
  INVX1 U1075 ( .A(dbg_01[5]), .Y(n853) );
  INVX1 U1076 ( .A(dbg_02[4]), .Y(n828) );
  INVX1 U1077 ( .A(dbg_05[5]), .Y(n857) );
  INVX1 U1078 ( .A(dbg_02[5]), .Y(n854) );
  INVX1 U1079 ( .A(dbg_03[4]), .Y(n832) );
  INVX1 U1080 ( .A(dbg_04[5]), .Y(n858) );
  INVX1 U1081 ( .A(dbg_04[4]), .Y(n833) );
  INVX1 U1082 ( .A(dbg_01[4]), .Y(n830) );
  INVX1 U1083 ( .A(dbg_04[3]), .Y(n808) );
  MUX2X1 U1084 ( .D0(n531), .D1(n63), .S(dummy[0]), .Y(n651) );
  AND2X1 U1085 ( .A(n532), .B(n537), .Y(n531) );
  MUX2X1 U1086 ( .D0(n533), .D1(n63), .S(dummy[1]), .Y(n650) );
  AND2X1 U1087 ( .A(dummy[0]), .B(n532), .Y(n533) );
  NAND3X1 U1088 ( .A(n418), .B(sfr_psw), .C(dw_ena), .Y(n417) );
  OAI222XL U1089 ( .A(n453), .B(n17), .C(sfr_wdat[7]), .D(n478), .E(
        memdatao[7]), .F(n476), .Y(N793) );
  INVX1 U1090 ( .A(n480), .Y(n453) );
  OAI221X1 U1091 ( .A(n462), .B(n17), .C(sfr_wdat[4]), .D(n478), .E(n461), .Y(
        N790) );
  OA22X1 U1092 ( .A(memdatao[4]), .B(n476), .C(n925), .D(n843), .Y(n461) );
  INVX1 U1093 ( .A(n486), .Y(n462) );
  OAI221X1 U1094 ( .A(n474), .B(n17), .C(sfr_wdat[1]), .D(n478), .E(n473), .Y(
        N787) );
  OA22X1 U1095 ( .A(memdatao[1]), .B(n476), .C(n925), .D(n768), .Y(n473) );
  INVX1 U1096 ( .A(n492), .Y(n474) );
  OAI221X1 U1097 ( .A(n479), .B(n17), .C(sfr_wdat[0]), .D(n478), .E(n477), .Y(
        N786) );
  OA22X1 U1098 ( .A(memdatao[0]), .B(n476), .C(n925), .D(n755), .Y(n477) );
  INVX1 U1099 ( .A(n494), .Y(n479) );
  OAI221X1 U1100 ( .A(n460), .B(n17), .C(sfr_wdat[5]), .D(n478), .E(n459), .Y(
        N791) );
  OA22X1 U1101 ( .A(memdatao[5]), .B(n476), .C(n925), .D(n868), .Y(n459) );
  INVX1 U1102 ( .A(n484), .Y(n460) );
  OAI221X1 U1103 ( .A(n466), .B(n17), .C(sfr_wdat[3]), .D(n478), .E(n464), .Y(
        N789) );
  OA22X1 U1104 ( .A(memdatao[3]), .B(n476), .C(n925), .D(n818), .Y(n464) );
  INVX1 U1105 ( .A(n488), .Y(n466) );
  OAI221X1 U1106 ( .A(n457), .B(n17), .C(sfr_wdat[6]), .D(n478), .E(n456), .Y(
        N792) );
  OA22X1 U1107 ( .A(memdatao[6]), .B(n476), .C(n925), .D(n894), .Y(n456) );
  INVX1 U1108 ( .A(n482), .Y(n457) );
  OAI221X1 U1109 ( .A(n470), .B(n17), .C(sfr_wdat[2]), .D(n478), .E(n469), .Y(
        N788) );
  OA22X1 U1110 ( .A(memdatao[2]), .B(n476), .C(n925), .D(n793), .Y(n469) );
  INVX1 U1111 ( .A(n490), .Y(n470) );
  NAND21X1 U1112 ( .B(n134), .A(c_ptr[0]), .Y(n658) );
  NAND21X1 U1113 ( .B(n187), .A(c_ptr[1]), .Y(n133) );
  OR2X1 U1114 ( .A(n153), .B(n74), .Y(n156) );
  AOI21X1 U1115 ( .B(c_adr[5]), .C(n152), .A(c_adr[6]), .Y(n74) );
  NAND21X1 U1116 ( .B(n740), .A(c_ptr[0]), .Y(n137) );
  XOR2X1 U1117 ( .A(n152), .B(c_adr[5]), .Y(n154) );
  INVX1 U1118 ( .A(c_ptr[1]), .Y(n134) );
  INVX1 U1119 ( .A(c_adr[1]), .Y(n187) );
  XOR2X1 U1120 ( .A(n138), .B(c_adr[8]), .Y(n159) );
  XOR2X1 U1121 ( .A(n121), .B(c_adr[9]), .Y(n162) );
  XOR2X1 U1122 ( .A(n119), .B(c_adr[7]), .Y(n158) );
  OR2X1 U1123 ( .A(n122), .B(n75), .Y(n163) );
  AOI21X1 U1124 ( .B(n120), .C(c_adr[9]), .A(c_adr[10]), .Y(n75) );
  NAND21X1 U1125 ( .B(c_adr[2]), .A(n638), .Y(n215) );
  INVX1 U1126 ( .A(c_ptr[2]), .Y(n638) );
  INVX1 U1127 ( .A(n116), .Y(n214) );
  NAND21X1 U1128 ( .B(n732), .A(c_ptr[2]), .Y(n116) );
  INVX1 U1129 ( .A(n117), .Y(n216) );
  NAND21X1 U1130 ( .B(n739), .A(c_ptr[3]), .Y(n117) );
  NAND21X1 U1131 ( .B(n631), .A(c_adr[4]), .Y(n126) );
  NAND21X1 U1132 ( .B(c_adr[0]), .A(n427), .Y(n357) );
  NAND21X1 U1133 ( .B(c_adr[4]), .A(n631), .Y(n219) );
  XOR2X1 U1134 ( .A(n140), .B(c_adr[13]), .Y(n169) );
  NAND21X1 U1135 ( .B(c_adr[3]), .A(n629), .Y(n217) );
  NAND21X1 U1136 ( .B(c_adr[1]), .A(n134), .Y(n213) );
  XNOR2XL U1137 ( .A(c_adr[14]), .B(n76), .Y(n208) );
  NAND2X1 U1138 ( .A(n139), .B(c_adr[13]), .Y(n76) );
  INVX1 U1139 ( .A(c_ptr[3]), .Y(n629) );
  INVX1 U1140 ( .A(c_ptr[0]), .Y(n427) );
  INVX1 U1141 ( .A(c_ptr[4]), .Y(n631) );
  NAND21X1 U1142 ( .B(n314), .A(c_adr[11]), .Y(n294) );
  NAND21X1 U1143 ( .B(n294), .A(c_adr[12]), .Y(n229) );
  INVX1 U1144 ( .A(n227), .Y(n239) );
  NAND21X1 U1145 ( .B(n229), .A(c_adr[13]), .Y(n227) );
  INVX1 U1146 ( .A(n118), .Y(n223) );
  NAND21X1 U1147 ( .B(n193), .A(c_adr[5]), .Y(n118) );
  INVX1 U1148 ( .A(c_adr[6]), .Y(n193) );
  AND2X1 U1149 ( .A(n247), .B(n381), .Y(n248) );
  AO21X1 U1150 ( .B(n246), .C(c_adr[7]), .A(c_adr[8]), .Y(n247) );
  AO21X1 U1151 ( .B(n344), .C(n234), .A(n334), .Y(n235) );
  INVX1 U1152 ( .A(c_adr[10]), .Y(n234) );
  AND2X1 U1153 ( .A(n243), .B(n242), .Y(n244) );
  AO21X1 U1154 ( .B(c_adr[5]), .C(n241), .A(c_adr[6]), .Y(n243) );
  INVX1 U1155 ( .A(c_adr[7]), .Y(n225) );
  NAND21X1 U1156 ( .B(n233), .A(c_adr[10]), .Y(n226) );
  AND3X1 U1157 ( .A(r_rdy), .B(o_inst[1]), .C(o_inst[0]), .Y(n258) );
  INVX1 U1158 ( .A(c_adr[11]), .Y(n305) );
  INVX1 U1159 ( .A(c_adr[9]), .Y(n233) );
  INVX1 U1160 ( .A(c_adr[8]), .Y(n224) );
  OAI31XL U1161 ( .A(n252), .B(n253), .C(n254), .D(n255), .Y(o_set_hold) );
  NAND43X1 U1162 ( .B(memaddr[5]), .C(memaddr[6]), .D(memaddr[4]), .A(n257), 
        .Y(n253) );
  NAND42X1 U1163 ( .C(memaddr[14]), .D(memaddr[13]), .A(n930), .B(n256), .Y(
        n254) );
  NAND4X1 U1164 ( .A(n258), .B(n259), .C(n260), .D(n261), .Y(n252) );
  INVX1 U1165 ( .A(n106), .Y(n538) );
  NAND5XL U1166 ( .A(d_hold[3]), .B(d_hold[0]), .C(d_hold[1]), .D(d_hold[2]), 
        .E(r_hold_mcu), .Y(n106) );
  INVX1 U1167 ( .A(c_adr[12]), .Y(n251) );
  INVX1 U1168 ( .A(n113), .Y(n639) );
  NAND21X1 U1169 ( .B(c_ptr[1]), .A(n427), .Y(n113) );
  INVX1 U1170 ( .A(n114), .Y(n180) );
  NAND21X1 U1171 ( .B(c_ptr[2]), .A(n639), .Y(n114) );
  NAND21X1 U1172 ( .B(cs_ft[2]), .A(n109), .Y(n560) );
  INVX1 U1173 ( .A(d_psrd), .Y(n694) );
  OAI31XL U1174 ( .A(r_rdy), .B(srst), .C(n563), .D(n928), .Y(n762) );
  INVX1 U1175 ( .A(un_hold), .Y(n563) );
  INVX1 U1176 ( .A(n874), .Y(n928) );
  INVX1 U1177 ( .A(dummy[1]), .Y(n537) );
  NAND21X1 U1178 ( .B(mcu_psw), .A(n515), .Y(n929) );
  NAND21X1 U1179 ( .B(n472), .A(n452), .Y(n480) );
  MUX2X1 U1180 ( .D0(pmem_q1[7]), .D1(pmem_q0[7]), .S(n693), .Y(n452) );
  NAND21X1 U1181 ( .B(n472), .A(n471), .Y(n492) );
  MUX2X1 U1182 ( .D0(pmem_q1[1]), .D1(pmem_q0[1]), .S(n693), .Y(n471) );
  NAND21X1 U1183 ( .B(n472), .A(n458), .Y(n484) );
  MUX2X1 U1184 ( .D0(pmem_q1[5]), .D1(pmem_q0[5]), .S(n693), .Y(n458) );
  NAND21X1 U1185 ( .B(n472), .A(n463), .Y(n488) );
  MUX2X1 U1186 ( .D0(pmem_q1[3]), .D1(pmem_q0[3]), .S(n693), .Y(n463) );
  NAND21X1 U1187 ( .B(n472), .A(n468), .Y(n490) );
  MUX2X1 U1188 ( .D0(pmem_q1[2]), .D1(pmem_q0[2]), .S(n693), .Y(n468) );
  NAND21X1 U1189 ( .B(n472), .A(n454), .Y(n482) );
  MUX2X1 U1190 ( .D0(pmem_q1[6]), .D1(pmem_q0[6]), .S(n693), .Y(n454) );
  OAI22X1 U1191 ( .A(pmem_q0[0]), .B(n475), .C(pmem_q1[0]), .D(n682), .Y(n494)
         );
  OAI22X1 U1192 ( .A(pmem_q0[4]), .B(n475), .C(pmem_q1[4]), .D(n682), .Y(n486)
         );
  INVX1 U1193 ( .A(memaddr[13]), .Y(n587) );
  NOR3XL U1194 ( .A(memaddr[7]), .B(memaddr[9]), .C(memaddr[8]), .Y(n257) );
  NOR3XL U1195 ( .A(memaddr[1]), .B(memaddr[3]), .C(memaddr[2]), .Y(n256) );
  INVX1 U1196 ( .A(mcu_psw), .Y(n665) );
  NOR3XL U1197 ( .A(memaddr[0]), .B(memaddr[11]), .C(memaddr[10]), .Y(n261) );
  NAND21X1 U1198 ( .B(wspp_cnt_2_), .A(n921), .Y(n939) );
  NOR21XL U1199 ( .B(n574), .A(pmem_a[6]), .Y(N757) );
  OR2X1 U1200 ( .A(wspp_cnt_0_), .B(wspp_cnt_1_), .Y(n599) );
  NAND21X1 U1201 ( .B(mcu_psw), .A(n433), .Y(n478) );
  NAND21X1 U1202 ( .B(n560), .A(mcu_psw), .Y(n476) );
  GEN2XL U1203 ( .D(n574), .E(n938), .C(N757), .B(pmem_a[8]), .A(n575), .Y(
        N759) );
  NOR42XL U1204 ( .C(pmem_a[6]), .D(n574), .A(n938), .B(pmem_a[8]), .Y(n575)
         );
  GEN2XL U1205 ( .D(wspp_cnt_0_), .E(wspp_cnt_1_), .C(n921), .B(n920), .A(n919), .Y(N796) );
  GEN2XL U1206 ( .D(wspp_cnt_2_), .E(n599), .C(n598), .B(n920), .A(n919), .Y(
        N797) );
  INVX1 U1207 ( .A(n939), .Y(n598) );
  GEN2XL U1208 ( .D(wspp_cnt_4_), .E(n927), .C(n554), .B(n920), .A(n919), .Y(
        N799) );
  GEN2XL U1209 ( .D(wspp_cnt_5_), .E(n926), .C(n553), .B(n920), .A(n919), .Y(
        N800) );
  INVX1 U1210 ( .A(n576), .Y(n937) );
  AOI32X1 U1211 ( .A(pmem_a[6]), .B(n938), .C(n574), .D(pmem_a[7]), .E(N757), 
        .Y(n576) );
  NOR2X1 U1212 ( .A(n939), .B(wspp_cnt_3_), .Y(n555) );
  NOR2X1 U1213 ( .A(n927), .B(wspp_cnt_4_), .Y(n554) );
  OAI21X1 U1214 ( .B(wspp_cnt_0_), .C(n940), .A(n929), .Y(N795) );
  OAI21X1 U1215 ( .B(n552), .C(n940), .A(n929), .Y(N801) );
  XNOR2XL U1216 ( .A(test_so2), .B(n553), .Y(n552) );
  NOR2X1 U1217 ( .A(n926), .B(wspp_cnt_5_), .Y(n553) );
  NOR21XL U1218 ( .B(n920), .A(n556), .Y(N798) );
  AOI21X1 U1219 ( .B(wspp_cnt_3_), .C(n939), .A(n555), .Y(n556) );
  INVX1 U1220 ( .A(pmem_a[7]), .Y(n938) );
  INVX1 U1221 ( .A(n429), .Y(n640) );
  NAND21X1 U1222 ( .B(c_ptr[1]), .A(c_ptr[0]), .Y(n429) );
  INVX1 U1223 ( .A(n428), .Y(n654) );
  NAND21X1 U1224 ( .B(c_ptr[0]), .A(c_ptr[1]), .Y(n428) );
  AND2X1 U1225 ( .A(d_hold[1]), .B(n104), .Y(N153) );
  AND2X1 U1226 ( .A(d_hold[0]), .B(n104), .Y(N152) );
  AND2X1 U1227 ( .A(d_hold[2]), .B(n104), .Y(N154) );
  NAND21XL U1228 ( .B(n686), .A(n433), .Y(n578) );
  INVXL U1229 ( .A(memaddr_c[2]), .Y(n136) );
  OAI22XL U1230 ( .A(memaddr_c[2]), .B(n146), .C(memaddr_c[3]), .D(n145), .Y(
        n147) );
  GEN2XL U1231 ( .D(memaddr_c[2]), .E(n732), .C(n184), .B(n185), .A(n183), .Y(
        n189) );
  XOR3XL U1232 ( .A(memaddr_c[2]), .B(n386), .C(n382), .Y(n415) );
  INVXL U1233 ( .A(n103), .Y(n101) );
  INVXL U1234 ( .A(n686), .Y(n102) );
  MAJ3X1 U1235 ( .A(n730), .B(c_adr[1]), .C(n922), .Y(n734) );
  MAJ3X1 U1236 ( .A(n936), .B(c_adr[3]), .C(n735), .Y(n388) );
endmodule


module ictlr_a0_DW01_inc_2 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module ictlr_a0_DW01_inc_1 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mcu51_a0 ( bclki2c, pc_ini, slp2wakeup, r_hold_mcu, wdt_slow, wdtov, 
        mdubsy, cs_run, t0_intr, clki2c, clkmdu, clkur0, clktm0, clktm1, 
        clkwdt, i2c_autoack, i2c_con_ens1, clkcpu, clkper, reset, ro, port0i, 
        exint_9, exint, clkcpuen, clkperen, port0o, port0ff, rxd0o, txd0, 
        rxd0i, rxd0oe, scli, sdai, sclo, sdao, waitstaten, mempsack, memack, 
        memdatai, memdatao, memaddr, mempswr, mempsrd, memwr, memrd, 
        memdatao_comb, memaddr_comb, mempswr_comb, mempsrd_comb, memwr_comb, 
        memrd_comb, ramdatai, ramdatao, ramaddr, ramwe, ramoe, dbgpo, sfrack, 
        sfrdatai, sfrdatao, sfraddr, sfrwe, sfroe, esfrm_wrdata, esfrm_addr, 
        esfrm_we, esfrm_oe, esfrm_rddata, test_si2, test_si1, test_so1, 
        test_se );
  input [15:0] pc_ini;
  output [1:0] wdtov;
  input [7:0] port0i;
  input [7:0] exint;
  output [7:0] port0o;
  output [7:0] port0ff;
  input [7:0] memdatai;
  output [7:0] memdatao;
  output [15:0] memaddr;
  output [7:0] memdatao_comb;
  output [15:0] memaddr_comb;
  input [7:0] ramdatai;
  output [7:0] ramdatao;
  output [7:0] ramaddr;
  output [31:0] dbgpo;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  output [6:0] sfraddr;
  input [7:0] esfrm_wrdata;
  input [6:0] esfrm_addr;
  output [7:0] esfrm_rddata;
  input bclki2c, slp2wakeup, r_hold_mcu, wdt_slow, clki2c, clkmdu, clkur0,
         clktm0, clktm1, clkwdt, i2c_autoack, clkcpu, clkper, reset, exint_9,
         rxd0i, scli, sdai, mempsack, memack, sfrack, esfrm_we, esfrm_oe,
         test_si2, test_si1, test_se;
  output mdubsy, cs_run, t0_intr, i2c_con_ens1, ro, clkcpuen, clkperen, rxd0o,
         txd0, rxd0oe, sclo, sdao, waitstaten, mempswr, mempsrd, memwr, memrd,
         mempswr_comb, mempsrd_comb, memwr_comb, memrd_comb, ramwe, ramoe,
         sfrwe, sfroe, test_so1;
  wire   n106, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, t0_tf1, t1_tf1, t0_tr1, t1_tr1, stop_flag, idle_flag, isfrwait,
         sfroe_s, sfroe_mcu51_per, sfrwe_s, sfrwe_mcu51_per, newinstr,
         intcall_int, cpu_resume, rmwinstr, pmw, p2sel, gf0, c, ac, ov, f0, f1,
         p, rsttowdt, rsttosrst, rst, int0ff, int1ff, rxd0ff, sdaiff,
         rsttowdtff, rsttosrstff, resetff, smod, ip0wdts, wdt_tm, bd, ie0, it0,
         ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9, isr_tm,
         i2c_int, i2ccon_o_7, tf1_gate, riti0_gate, iex7_gate, iex2_gate,
         srstflag, int_vect_8b, int_vect_93, int_vect_9b, int_vect_a3, wdts,
         srst, pmuintreq_rev, pmuintreq, t1ov, t0ack, t1ack, isr_irq, int0ack,
         int1ack, iex7ack, iex2ack, iex3ack, iex4ack, iex5ack, iex6ack,
         iex8ack, iex9ack, n11, n113, n112, n111, n110, n109, n108, n107, n62,
         n63, n97, n115, n117, n3, n7, n8, n9, n10, n12, n2, n4, n5, n6, n13,
         n14, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36, n38, n39,
         n40, n41, n42, n44, n46, n47, n48, n49, n57, n60, n61, n64, n66, n67,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5;
  wire   [13:0] timer_1ms;
  wire   [5:0] ien2;
  wire   [6:0] ramsfraddr;
  wire   [4:0] intvect_int;
  wire   [7:0] ckcon;
  wire   [7:0] dph;
  wire   [7:0] dpl;
  wire   [3:0] dps;
  wire   [7:0] p2;
  wire   [5:0] dpc;
  wire   [7:0] sp;
  wire   [7:0] acc_s;
  wire   [7:0] b;
  wire   [1:0] rs;
  wire   [7:0] arcon;
  wire   [7:0] md0;
  wire   [7:0] md1;
  wire   [7:0] md2;
  wire   [7:0] md3;
  wire   [7:0] md4;
  wire   [7:0] md5;
  wire   [3:0] t0_tmod;
  wire   [7:0] tl0;
  wire   [7:0] th0;
  wire   [3:0] t1_tmod;
  wire   [7:0] tl1;
  wire   [7:0] th1;
  wire   [7:0] wdtrel;
  wire   [6:5] t2con;
  wire   [7:0] s0con;
  wire   [7:0] s0buf;
  wire   [7:0] s0rell;
  wire   [7:0] s0relh;
  wire   [7:0] ien0;
  wire   [5:0] ien1;
  wire   [5:0] ip0;
  wire   [5:0] ip1;
  wire   [7:0] i2cdat_o;
  wire   [7:0] i2cadr_o;
  wire   [5:0] i2ccon_o;
  wire   [7:0] i2csta_o;
  wire   [3:0] isreg;

  INVX1 U33 ( .A(n63), .Y(n62) );
  INVX1 U34 ( .A(reset), .Y(n63) );
  INVX8 U52 ( .A(n63), .Y(n3) );
  mcu51_cpu_a0 u_cpu ( .clkcpu(clkcpu), .rst(n67), .mempsack(mempsack), 
        .memack(memack), .memdatai(memdatai), .memaddr(memaddr), .mempsrd(
        mempsrd), .mempswr(mempswr), .memrd(memrd), .memwr(memwr), 
        .memaddr_comb({memaddr_comb[15:2], n106, memaddr_comb[0]}), 
        .mempsrd_comb(mempsrd_comb), .mempswr_comb(mempswr_comb), .memrd_comb(
        memrd_comb), .memwr_comb(memwr_comb), .cpu_hold(r_hold_mcu), 
        .cpu_resume(cpu_resume), .irq(dbgpo[20]), .intvect(intvect_int), 
        .intcall(intcall_int), .retiinstr(dbgpo[21]), .newinstr(newinstr), 
        .rmwinstr(rmwinstr), .waitstaten(waitstaten), .ramdatai(ramdatai), 
        .sfrdatai(esfrm_rddata), .ramsfraddr({SYNOPSYS_UNCONNECTED_1, 
        ramsfraddr}), .ramdatao(memdatao), .ramoe(), .ramwe(), .sfroe(sfroe_s), 
        .sfrwe(sfrwe_s), .sfroe_r(), .sfrwe_r(), .sfroe_comb_s(), 
        .sfrwe_comb_s(), .pc_o(dbgpo[15:0]), .pc_ini(pc_ini), .cs_run(cs_run), 
        .instr(dbgpo[31:24]), .codefetch_s(), .sfrack(sfrack), 
        .ramsfraddr_comb(ramaddr), .ramdatao_comb(ramdatao), .ramoe_comb(ramoe), .ramwe_comb(ramwe), .ckcon(ckcon), .pmw(pmw), .p2sel(p2sel), .gf0(gf0), 
        .stop(stop_flag), .idle(idle_flag), .acc(acc_s), .b(b), .rs(rs), .c(c), 
        .ac(ac), .ov(ov), .p(p), .f0(f0), .f1(f1), .dph(dph), .dpl(dpl), .dps(
        dps), .dpc(dpc), .p2(p2), .sp(sp), .test_si(timer_1ms[13]), .test_so(
        n117), .test_se(test_se) );
  syncneg_a0 u_syncneg ( .clk(clkper), .reset(n62), .rsttowdt(rsttowdt), 
        .rsttosrst(rsttosrst), .rst(rst), .int0(exint[0]), .int1(exint[1]), 
        .port0i(port0i), .rxd0i(rxd0i), .sdai(sdai), .int0ff(int0ff), .int1ff(
        int1ff), .port0ff(port0ff), .t0ff(), .t1ff(), .rxd0ff(rxd0ff), 
        .sdaiff(sdaiff), .rsttowdtff(rsttowdtff), .rsttosrstff(rsttosrstff), 
        .rstff(n97), .resetff(resetff), .test_si(srstflag), .test_se(test_se)
         );
  sfrmux_a0 u_sfrmux ( .isfrwait(isfrwait), .sfraddr({n48, n47, sfraddr[4], 
        n41, n39, n36, n13}), .c(c), .ac(ac), .f0(f0), .rs(rs), .ov(ov), .f1(
        f1), .p(p), .acc(acc_s), .b(b), .dpl(dpl), .dph(dph), .dps(dps), .dpc(
        dpc), .p2(p2), .sp(sp), .smod(smod), .pmw(pmw), .p2sel(p2sel), .gf0(
        gf0), .stop(stop_flag), .idle(idle_flag), .ckcon(ckcon), .port0(port0o), .port0ff(port0ff), .rmwinstr(rmwinstr), .arcon(arcon), .md0(md0), .md1(md1), 
        .md2(md2), .md3(md3), .md4(md4), .md5(md5), .t0_tmod(t0_tmod), 
        .t0_tf0(dbgpo[17]), .t0_tf1(t0_tf1), .t0_tr0(dbgpo[16]), .t0_tr1(
        t0_tr1), .tl0(tl0), .th0(th0), .t1_tmod(t1_tmod), .t1_tf1(t1_tf1), 
        .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1), .wdtrel(wdtrel), .ip0wdts(
        ip0wdts), .wdt_tm(wdt_tm), .t2con({1'b0, t2con, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .s0con(s0con), .s0buf(s0buf), .s0rell(s0rell), .s0relh(s0relh), 
        .bd(bd), .ie0(ie0), .it0(it0), .ie1(ie1), .it1(it1), .iex2(iex2), 
        .iex3(iex3), .iex4(iex4), .iex5(iex5), .iex6(iex6), .iex7(iex7), 
        .iex8(iex8), .iex9(iex9), .iex10(1'b0), .iex11(1'b0), .iex12(1'b0), 
        .ien0({ien0[7], 1'b0, ien0[5:0]}), .ien1(ien1), .ien2(ien2), .ip0(ip0), 
        .ip1(ip1), .isr_tm(isr_tm), .i2c_int(i2c_int), .i2cdat_o(i2cdat_o), 
        .i2cadr_o(i2cadr_o), .i2ccon_o({i2ccon_o_7, i2c_con_ens1, i2ccon_o}), 
        .i2csta_o({i2csta_o[7:3], 1'b0, 1'b0, 1'b0}), .sfrdatai(sfrdatai), 
        .tf1_gate(tf1_gate), .riti0_gate(riti0_gate), .iex7_gate(iex7_gate), 
        .iex2_gate(iex2_gate), .srstflag(srstflag), .int_vect_8b(int_vect_8b), 
        .int_vect_93(int_vect_93), .int_vect_9b(int_vect_9b), .int_vect_a3(
        int_vect_a3), .ext_sfr_sel(), .sfrdatao(esfrm_rddata) );
  pmurstctrl_a0 u_pmurstctrl ( .resetff(resetff), .wdts(wdts), .srst(srst), 
        .pmuintreq(pmuintreq_rev), .stop(stop_flag), .idle(idle_flag), 
        .clkcpu_en(clkcpuen), .clkper_en(clkperen), .cpu_resume(cpu_resume), 
        .rsttowdt(rsttowdt), .rsttosrst(rsttosrst), .rst(rst) );
  wakeupctrl_a0 u_wakeupctrl ( .irq(dbgpo[20]), .int0ff(exint[0]), .int1ff(
        exint[1]), .it0(it0), .it1(it1), .isreg(isreg), .intprior0({ip0[2], 
        ip0[0]}), .intprior1({ip1[2], ip1[0]}), .eal(ien0[7]), .eint0(ien0[0]), 
        .eint1(ien0[2]), .pmuintreq(pmuintreq) );
  mdu_a0 u_mdu ( .clkper(clkmdu), .rst(n67), .mdubsy(mdubsy), .sfrdatai({
        sfrdatao[7:6], n57, sfrdatao[4:0]}), .sfraddr({sfraddr[6], n46, n44, 
        n41, n38, n36, n34}), .sfrwe(n28), .sfroe(sfroe_mcu51_per), .arcon(
        arcon), .md0(md0), .md1(md1), .md2(md2), .md3(md3), .md4(md4), .md5(
        md5), .test_si(isr_tm), .test_so(n115), .test_se(test_se) );
  ports_a0 u_ports ( .clkper(clkper), .rst(dbgpo[22]), .port0(port0o), 
        .sfrdatai({sfrdatao[7], n107, n108, n109, sfrdatao[3:0]}), .sfraddr({
        sfraddr[6], n47, n44, n42, n14, n36, n34}), .sfrwe(n28), .test_si(n115), .test_se(test_se) );
  serial0_a0 u_serial0 ( .t_shift_clk(), .r_shift_clk(), .clkper(clkur0), 
        .rst(dbgpo[22]), .newinstr(newinstr), .rxd0ff(rxd0ff), .t1ov(t1ov), 
        .rxd0o(rxd0o), .rxd0oe(rxd0oe), .txd0(txd0), .sfrdatai({n60, 
        sfrdatao[6], n57, sfrdatao[4], n110, n111, n112, n113}), .sfraddr({
        sfraddr[6], n46, n2, n42, n39, n27, n33}), .sfrwe(n29), .s0con(s0con), 
        .s0buf(s0buf), .s0rell(s0rell), .s0relh(s0relh), .smod(smod), .bd(bd), 
        .test_si(port0o[7]), .test_se(test_se) );
  timer0_a0 u_timer0 ( .clkper(clktm0), .rst(n66), .newinstr(newinstr), .t0ff(
        1'b0), .t0ack(t0ack), .t1ack(t1ack), .int0ff(int0ff), .t0_tf0(
        dbgpo[17]), .t0_tf1(t0_tf1), .sfrdatai({sfrdatao[7:6], n57, 
        sfrdatao[4], n110, sfrdatao[2:0]}), .sfraddr({n49, n46, n2, n42, n38, 
        sfraddr[1], n34}), .sfrwe(n28), .t0_tmod(t0_tmod), .t0_tr0(dbgpo[16]), 
        .t0_tr1(t0_tr1), .tl0(tl0), .th0(th0), .test_si(sdaiff), .test_se(
        test_se) );
  timer1_a0 u_timer1 ( .clkper(clktm1), .rst(n61), .newinstr(newinstr), .t1ff(
        1'b0), .t1ack(t1ack), .int1ff(int1ff), .t1_tf1(t1_tf1), .t1ov(t1ov), 
        .sfrdatai({n60, sfrdatao[6], n57, sfrdatao[4], n110, n111, n112, n113}), .sfraddr({n49, n47, n44, sfraddr[3], n38, n27, n33}), .sfrwe(n29), .t1_tmod(
        t1_tmod), .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1), .test_si(tl0[7]), 
        .test_se(test_se) );
  watchdog_a0 u_watchdog ( .wdt_slow(wdt_slow), .clkwdt(clkwdt), .clkper(
        clkper), .resetff(rsttowdtff), .newinstr(newinstr), .wdts_s(wdtov), 
        .wdts(wdts), .ip0wdts(ip0wdts), .wdt_tm(wdt_tm), .sfrdatai({
        sfrdatao[7:6], n108, n109, sfrdatao[3:0]}), .sfraddr({sfraddr[6:5], 
        n44, sfraddr[3], n39, n27, n33}), .sfrwe(n29), .wdtrel(wdtrel), 
        .test_si(tl1[7]), .test_se(test_se) );
  isr_a0 u_isr ( .clkper(clkper), .rst(n64), .intcall(intcall_int), 
        .retiinstr(dbgpo[21]), .int_vect_03(ie0), .int_vect_0b(dbgpo[17]), 
        .t0ff(1'b0), .int_vect_13(ie1), .int_vect_1b(tf1_gate), .t1ff(1'b0), 
        .int_vect_23(riti0_gate), .i2c_int(i2c_int), .rxd0ff(rxd0ff), 
        .int_vect_43(iex7_gate), .sdaiff(sdaiff), .int_vect_4b(iex2_gate), 
        .int_vect_53(iex3), .int_vect_5b(iex4), .int_vect_63(iex5), 
        .int_vect_6b(iex6), .int_vect_8b(int_vect_8b), .int_vect_93(
        int_vect_93), .int_vect_9b(int_vect_9b), .int_vect_a3(int_vect_a3), 
        .int_vect_ab(1'b0), .irq(isr_irq), .intvect(intvect_int), .int_ack_03(
        int0ack), .int_ack_0b(t0ack), .int_ack_13(int1ack), .int_ack_1b(t1ack), 
        .int_ack_43(iex7ack), .int_ack_4b(iex2ack), .int_ack_53(iex3ack), 
        .int_ack_5b(iex4ack), .int_ack_63(iex5ack), .int_ack_6b(iex6ack), 
        .int_ack_8b(iex8ack), .int_ack_93(iex9ack), .int_ack_9b(), 
        .int_ack_a3(), .int_ack_ab(), .is_reg(isreg), .ip0(ip0), .ip1(ip1), 
        .ien0({ien0[7], SYNOPSYS_UNCONNECTED_2, ien0[5:0]}), .ien1(ien1), 
        .ien2(ien2), .isr_tm(isr_tm), .sfraddr({n49, n46, n2, n42, 
        sfraddr[2:1], n34}), .sfrdatai({sfrdatao[7], n107, n57, sfrdatao[4:0]}), .sfrwe(n29), .test_si(test_si2), .test_se(test_se) );
  extint_a0 u_extint ( .clkper(clkper), .rst(n66), .newinstr(newinstr), 
        .int0ff(int0ff), .int0ack(int0ack), .int1ff(int1ff), .int1ack(int1ack), 
        .int2ff(exint[2]), .iex2ack(iex2ack), .int3ff(exint[3]), .iex3ack(
        iex3ack), .int4ff(exint[4]), .iex4ack(iex4ack), .int5ff(exint[5]), 
        .iex5ack(iex5ack), .int6ff(exint[6]), .iex6ack(iex6ack), .int7ff(
        exint[7]), .iex7ack(iex7ack), .int8ff(n11), .iex8ack(iex8ack), 
        .int9ff(exint_9), .iex9ack(iex9ack), .ie0(ie0), .it0(it0), .ie1(ie1), 
        .it1(it1), .i2fr(t2con[5]), .iex2(iex2), .i3fr(t2con[6]), .iex3(iex3), 
        .iex4(iex4), .iex5(iex5), .iex6(iex6), .iex7(iex7), .iex8(iex8), 
        .iex9(iex9), .iex10(), .iex11(), .iex12(), .sfraddr({n49, n47, n44, 
        n41, n38, n36, n34}), .sfrdatai({n60, n107, n57, n109, n110, n111, 
        n112, n113}), .sfrwe(n28), .test_si(n117), .test_se(test_se) );
  i2c_a0 u_i2c ( .clk(clki2c), .rst(n67), .bclksel(bclki2c), .scli(scli), 
        .sdai(sdai), .sclo(sclo), .sdao(sdao), .intack(i2c_autoack), .si(
        i2c_int), .sfrwe(n28), .sfraddr({n49, n46, n2, n42, sfraddr[2:1], n13}), .sfrdatai({sfrdatao[7], n107, n108, sfrdatao[4:3], n111, sfrdatao[1:0]}), 
        .i2cdat_o(i2cdat_o), .i2cadr_o(i2cadr_o), .i2ccon_o({i2ccon_o_7, 
        i2c_con_ens1, i2ccon_o}), .i2csta_o({i2csta_o[7:3], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5}), .test_si(it1), .test_so(test_so1), .test_se(test_se) );
  softrstctrl_a0 u_softrstctrl ( .clkcpu(clkcpu), .resetff(rsttosrstff), 
        .newinstr(newinstr), .srstreq(srst), .srstflag(srstflag), .sfrdatai({
        n60, n107, n57, n109, sfrdatao[3:0]}), .sfraddr({sfraddr[6], n46, n44, 
        n42, n39, n27, n13}), .sfrwe(n29), .test_si(txd0), .test_se(test_se)
         );
  mcu51_a0_DW01_inc_0 add_268 ( .A(timer_1ms), .SUM({N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7}) );
  SDFFQX1 timer_1ms_reg_9_ ( .D(N30), .SIN(timer_1ms[8]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[9]) );
  SDFFQX1 timer_1ms_reg_13_ ( .D(N34), .SIN(timer_1ms[12]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[13]) );
  SDFFQX1 timer_1ms_reg_12_ ( .D(N33), .SIN(timer_1ms[11]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[12]) );
  SDFFQX1 timer_1ms_reg_8_ ( .D(N29), .SIN(timer_1ms[7]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[8]) );
  SDFFQX1 timer_1ms_reg_10_ ( .D(N31), .SIN(timer_1ms[9]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[10]) );
  SDFFQX1 timer_1ms_reg_6_ ( .D(N27), .SIN(timer_1ms[5]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[6]) );
  SDFFQX1 timer_1ms_reg_11_ ( .D(N32), .SIN(timer_1ms[10]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[11]) );
  SDFFQX1 timer_1ms_reg_7_ ( .D(N28), .SIN(timer_1ms[6]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[7]) );
  SDFFQX1 timer_1ms_reg_5_ ( .D(N26), .SIN(timer_1ms[4]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[5]) );
  SDFFQX1 timer_1ms_reg_4_ ( .D(N25), .SIN(timer_1ms[3]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[4]) );
  SDFFQX1 timer_1ms_reg_3_ ( .D(N24), .SIN(timer_1ms[2]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[3]) );
  SDFFQX1 timer_1ms_reg_2_ ( .D(N23), .SIN(timer_1ms[1]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[2]) );
  SDFFQX1 timer_1ms_reg_1_ ( .D(N22), .SIN(timer_1ms[0]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[1]) );
  SDFFQX1 timer_1ms_reg_0_ ( .D(N21), .SIN(test_si1), .SMC(test_se), .C(clkper), .Q(timer_1ms[0]) );
  MUX2IX2 U3 ( .D0(esfrm_addr[3]), .D1(ramsfraddr[3]), .S(n6), .Y(n72) );
  INVX3 U4 ( .A(isfrwait), .Y(n6) );
  INVXL U5 ( .A(n75), .Y(n49) );
  INVX1 U6 ( .A(n75), .Y(n48) );
  INVX3 U7 ( .A(n75), .Y(sfraddr[6]) );
  MUX2IX2 U8 ( .D0(esfrm_addr[6]), .D1(ramsfraddr[6]), .S(n6), .Y(n75) );
  INVX1 U9 ( .A(n92), .Y(n95) );
  INVX2 U10 ( .A(n26), .Y(n36) );
  MUX2XL U11 ( .D0(esfrm_addr[0]), .D1(ramsfraddr[0]), .S(n6), .Y(n13) );
  INVX1 U12 ( .A(n14), .Y(n40) );
  BUFX1 U13 ( .A(n73), .Y(n25) );
  INVXL U14 ( .A(n25), .Y(n44) );
  INVX1 U15 ( .A(n25), .Y(sfraddr[4]) );
  MUX2X1 U16 ( .D0(esfrm_addr[2]), .D1(ramsfraddr[2]), .S(n5), .Y(n14) );
  INVX1 U17 ( .A(n74), .Y(sfraddr[5]) );
  MUX2IX1 U18 ( .D0(esfrm_addr[5]), .D1(ramsfraddr[5]), .S(n6), .Y(n74) );
  INVX1 U19 ( .A(n72), .Y(n41) );
  INVX1 U20 ( .A(n25), .Y(n2) );
  INVX1 U21 ( .A(n40), .Y(sfraddr[2]) );
  BUFXL U22 ( .A(n5), .Y(n4) );
  NAND21X2 U23 ( .B(esfrm_oe), .A(n93), .Y(isfrwait) );
  INVXL U24 ( .A(n13), .Y(n35) );
  AO21XL U25 ( .B(n95), .C(n94), .A(esfrm_we), .Y(sfrwe) );
  INVXL U26 ( .A(isfrwait), .Y(n5) );
  INVX1 U27 ( .A(n35), .Y(n34) );
  INVX1 U28 ( .A(n35), .Y(n33) );
  INVX1 U29 ( .A(n40), .Y(n39) );
  INVX1 U30 ( .A(esfrm_we), .Y(n93) );
  BUFX3 U31 ( .A(sfrwe_mcu51_per), .Y(n28) );
  BUFX3 U32 ( .A(sfrwe_mcu51_per), .Y(n29) );
  INVX1 U35 ( .A(n40), .Y(n38) );
  BUFX3 U36 ( .A(ramdatao[2]), .Y(memdatao_comb[2]) );
  BUFX3 U37 ( .A(ramdatao[4]), .Y(memdatao_comb[4]) );
  BUFX3 U38 ( .A(ramdatao[5]), .Y(memdatao_comb[5]) );
  BUFX3 U39 ( .A(ramdatao[6]), .Y(memdatao_comb[6]) );
  BUFX3 U40 ( .A(ramdatao[7]), .Y(memdatao_comb[7]) );
  BUFX3 U41 ( .A(n106), .Y(memaddr_comb[1]) );
  INVX1 U42 ( .A(n74), .Y(n47) );
  INVX1 U43 ( .A(n85), .Y(sfrdatao[3]) );
  INVX1 U44 ( .A(n35), .Y(sfraddr[0]) );
  INVX1 U45 ( .A(n69), .Y(dbgpo[22]) );
  INVX1 U46 ( .A(n70), .Y(ro) );
  INVX1 U47 ( .A(n91), .Y(sfrdatao[0]) );
  INVX1 U48 ( .A(n81), .Y(sfrdatao[5]) );
  INVX1 U49 ( .A(n83), .Y(sfrdatao[4]) );
  INVX1 U50 ( .A(n79), .Y(sfrdatao[6]) );
  INVX1 U51 ( .A(n77), .Y(sfrdatao[7]) );
  INVX1 U53 ( .A(n89), .Y(sfrdatao[1]) );
  INVX1 U54 ( .A(n87), .Y(sfrdatao[2]) );
  NAND21XL U55 ( .B(esfrm_oe), .A(n96), .Y(sfroe_mcu51_per) );
  INVXL U56 ( .A(n72), .Y(n42) );
  INVXL U57 ( .A(n72), .Y(sfraddr[3]) );
  INVX1 U58 ( .A(n81), .Y(n57) );
  INVX1 U59 ( .A(n69), .Y(n67) );
  NOR21XL U60 ( .B(N19), .A(n30), .Y(N33) );
  NOR21XL U61 ( .B(N18), .A(n31), .Y(N32) );
  NOR21XL U62 ( .B(N17), .A(n30), .Y(N31) );
  NOR21XL U63 ( .B(N16), .A(n31), .Y(N30) );
  INVX1 U64 ( .A(n70), .Y(n61) );
  INVX1 U65 ( .A(n70), .Y(n64) );
  INVX1 U66 ( .A(n69), .Y(n66) );
  NOR21XL U67 ( .B(N8), .A(n31), .Y(N22) );
  NOR21XL U68 ( .B(N9), .A(n30), .Y(N23) );
  NOR21XL U69 ( .B(N10), .A(n31), .Y(N24) );
  NOR21XL U70 ( .B(N11), .A(n30), .Y(N25) );
  NOR21XL U71 ( .B(N14), .A(n31), .Y(N28) );
  NOR21XL U72 ( .B(N13), .A(n30), .Y(N27) );
  NOR21XL U73 ( .B(N12), .A(n31), .Y(N26) );
  NOR21XL U74 ( .B(N15), .A(n30), .Y(N29) );
  BUFX3 U75 ( .A(n7), .Y(n30) );
  BUFX3 U76 ( .A(n7), .Y(n31) );
  BUFX3 U77 ( .A(ramdatao[0]), .Y(memdatao_comb[0]) );
  BUFX3 U78 ( .A(ramdatao[1]), .Y(memdatao_comb[1]) );
  BUFX3 U79 ( .A(ramdatao[3]), .Y(memdatao_comb[3]) );
  BUFX3 U80 ( .A(rxd0i), .Y(dbgpo[23]) );
  INVX1 U81 ( .A(n77), .Y(n60) );
  OR2X1 U82 ( .A(t0_tf1), .B(t1_tf1), .Y(dbgpo[19]) );
  NAND21X1 U83 ( .B(isfrwait), .A(sfrwe_s), .Y(n92) );
  INVX1 U84 ( .A(n85), .Y(n110) );
  INVX1 U85 ( .A(memdatao[3]), .Y(n84) );
  OR2X1 U86 ( .A(pmuintreq), .B(slp2wakeup), .Y(pmuintreq_rev) );
  NOR21XL U87 ( .B(isr_irq), .A(r_hold_mcu), .Y(dbgpo[20]) );
  OR2X1 U88 ( .A(t0_tr1), .B(t1_tr1), .Y(dbgpo[18]) );
  INVX1 U89 ( .A(n97), .Y(n69) );
  INVX1 U90 ( .A(n97), .Y(n70) );
  INVX1 U91 ( .A(n91), .Y(n113) );
  INVX1 U92 ( .A(memdatao[0]), .Y(n90) );
  AO21XL U93 ( .B(sfroe_s), .C(n94), .A(esfrm_oe), .Y(sfroe) );
  INVX1 U94 ( .A(n79), .Y(n107) );
  INVX1 U95 ( .A(memdatao[6]), .Y(n78) );
  INVX1 U96 ( .A(n81), .Y(n108) );
  INVX1 U97 ( .A(memdatao[5]), .Y(n80) );
  INVX1 U98 ( .A(sfroe_s), .Y(n96) );
  INVX1 U99 ( .A(memdatao[7]), .Y(n76) );
  INVX1 U100 ( .A(n83), .Y(n109) );
  INVX1 U101 ( .A(memdatao[4]), .Y(n82) );
  INVX1 U102 ( .A(n89), .Y(n112) );
  INVX1 U103 ( .A(memdatao[1]), .Y(n88) );
  INVX1 U104 ( .A(n87), .Y(n111) );
  INVX1 U105 ( .A(memdatao[2]), .Y(n86) );
  NOR21XL U106 ( .B(N20), .A(n31), .Y(N34) );
  NAND32X1 U107 ( .B(n11), .C(n3), .A(ien2[1]), .Y(n7) );
  NOR21XL U108 ( .B(N7), .A(n30), .Y(N21) );
  NAND43X1 U109 ( .B(timer_1ms[8]), .C(timer_1ms[5]), .D(timer_1ms[12]), .A(
        timer_1ms[0]), .Y(n10) );
  NOR4XL U110 ( .A(n8), .B(n9), .C(n10), .D(n12), .Y(n11) );
  NAND4X1 U111 ( .A(timer_1ms[4]), .B(timer_1ms[3]), .C(timer_1ms[2]), .D(
        timer_1ms[1]), .Y(n8) );
  NAND3X1 U112 ( .A(timer_1ms[7]), .B(timer_1ms[6]), .C(timer_1ms[9]), .Y(n9)
         );
  NAND3X1 U113 ( .A(timer_1ms[11]), .B(timer_1ms[10]), .C(timer_1ms[13]), .Y(
        n12) );
  AND2X1 U114 ( .A(ien0[0]), .B(dbgpo[17]), .Y(t0_intr) );
  MUX2IXL U115 ( .D0(esfrm_addr[4]), .D1(ramsfraddr[4]), .S(n5), .Y(n73) );
  BUFX3 U116 ( .A(n71), .Y(n26) );
  INVXL U117 ( .A(n71), .Y(sfraddr[1]) );
  INVXL U118 ( .A(n26), .Y(n27) );
  INVXL U119 ( .A(n74), .Y(n46) );
  MUX2AXL U120 ( .D0(esfrm_wrdata[3]), .D1(n84), .S(n4), .Y(n85) );
  MUX2AXL U121 ( .D0(esfrm_wrdata[1]), .D1(n88), .S(n6), .Y(n89) );
  MUX2AXL U122 ( .D0(esfrm_wrdata[2]), .D1(n86), .S(n4), .Y(n87) );
  MUX2AXL U123 ( .D0(esfrm_wrdata[4]), .D1(n82), .S(n6), .Y(n83) );
  MUX2AXL U124 ( .D0(esfrm_wrdata[5]), .D1(n80), .S(n4), .Y(n81) );
  MUX2AXL U125 ( .D0(esfrm_wrdata[6]), .D1(n78), .S(n4), .Y(n79) );
  MUX2AXL U126 ( .D0(esfrm_wrdata[7]), .D1(n76), .S(n6), .Y(n77) );
  MUX2AXL U127 ( .D0(esfrm_wrdata[0]), .D1(n90), .S(n6), .Y(n91) );
  NAND21XL U128 ( .B(n95), .A(n93), .Y(sfrwe_mcu51_per) );
  MUX2IX1 U129 ( .D0(esfrm_addr[1]), .D1(ramsfraddr[1]), .S(n5), .Y(n71) );
  INVX8 U130 ( .A(n3), .Y(n94) );
endmodule


module mcu51_a0_DW01_inc_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;

  wire   [13:2] carry;

  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module softrstctrl_a0 ( clkcpu, resetff, newinstr, srstreq, srstflag, sfrdatai, 
        sfraddr, sfrwe, test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkcpu, resetff, newinstr, sfrwe, test_si, test_se;
  output srstreq, srstflag;
  wire   srst_ff0, srst_ff1, N37, N38, N41, net11998, n24, n25, n26, n27, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n28, n29,
         n30, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [3:0] srst_count;

  SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 clk_gate_srst_count_reg ( .CLK(clkcpu), 
        .EN(N37), .ENCLK(net11998), .TE(test_se) );
  SDFFQX1 srst_ff1_reg ( .D(n24), .SIN(srst_ff0), .SMC(test_se), .C(clkcpu), 
        .Q(srst_ff1) );
  SDFFQX1 srst_count_reg_1_ ( .D(n6), .SIN(srst_count[0]), .SMC(test_se), .C(
        net11998), .Q(srst_count[1]) );
  SDFFQX1 srst_count_reg_3_ ( .D(N41), .SIN(srst_count[2]), .SMC(test_se), .C(
        net11998), .Q(srst_count[3]) );
  SDFFQX1 srst_ff0_reg ( .D(n26), .SIN(srst_count[3]), .SMC(test_se), .C(
        clkcpu), .Q(srst_ff0) );
  SDFFQX1 srst_count_reg_0_ ( .D(N38), .SIN(test_si), .SMC(test_se), .C(
        net11998), .Q(srst_count[0]) );
  SDFFQX1 srst_count_reg_2_ ( .D(n4), .SIN(srst_count[1]), .SMC(test_se), .C(
        net11998), .Q(srst_count[2]) );
  SDFFQX1 srst_r_reg ( .D(n27), .SIN(srst_ff1), .SMC(test_se), .C(clkcpu), .Q(
        srstreq) );
  SDFFQX1 srstflag_reg ( .D(n25), .SIN(srstreq), .SMC(test_se), .C(clkcpu), 
        .Q(srstflag) );
  INVX1 U3 ( .A(n15), .Y(n2) );
  NAND42X1 U4 ( .C(sfraddr[3]), .D(n20), .A(sfraddr[0]), .B(n21), .Y(n15) );
  NAND2XL U5 ( .A(sfraddr[2]), .B(sfraddr[1]), .Y(n20) );
  NAND2X1 U6 ( .A(sfrdatai[0]), .B(n2), .Y(n12) );
  INVX1 U7 ( .A(newinstr), .Y(n3) );
  NOR2X1 U8 ( .A(n16), .B(n5), .Y(n22) );
  INVX1 U9 ( .A(n28), .Y(n5) );
  INVX1 U10 ( .A(n16), .Y(n9) );
  NAND2X1 U11 ( .A(n10), .B(n16), .Y(N37) );
  NOR2X1 U12 ( .A(resetff), .B(n18), .Y(n24) );
  AOI22AXL U13 ( .A(srst_ff0), .B(n2), .D(n19), .C(n8), .Y(n18) );
  AOI32X1 U14 ( .A(srst_ff1), .B(n3), .C(n15), .D(srst_ff0), .E(newinstr), .Y(
        n19) );
  NOR2X1 U15 ( .A(resetff), .B(n11), .Y(n27) );
  AOI32X1 U16 ( .A(n12), .B(n13), .C(srstreq), .D(srst_ff1), .E(n1), .Y(n11)
         );
  NAND3X1 U17 ( .A(srst_count[2]), .B(n5), .C(srst_count[3]), .Y(n13) );
  INVX1 U18 ( .A(n12), .Y(n1) );
  NAND2X1 U19 ( .A(n16), .B(n17), .Y(n25) );
  OAI211X1 U20 ( .C(sfrdatai[0]), .D(n15), .A(n10), .B(srstflag), .Y(n17) );
  AOI21X1 U21 ( .B(n12), .C(n14), .A(resetff), .Y(n26) );
  NAND4X1 U22 ( .A(srst_ff0), .B(n15), .C(n3), .D(n8), .Y(n14) );
  GEN2XL U23 ( .D(n9), .E(n7), .C(n22), .B(srst_count[3]), .A(n23), .Y(N41) );
  NOR4XL U24 ( .A(srst_count[3]), .B(n28), .C(n7), .D(n16), .Y(n23) );
  NAND2X1 U25 ( .A(srstreq), .B(n10), .Y(n16) );
  NAND2X1 U26 ( .A(srst_count[1]), .B(srst_count[0]), .Y(n28) );
  INVX1 U27 ( .A(resetff), .Y(n10) );
  INVX1 U28 ( .A(srst_count[2]), .Y(n7) );
  INVX1 U29 ( .A(srstreq), .Y(n8) );
  INVX1 U30 ( .A(n30), .Y(n6) );
  OAI211X1 U31 ( .C(srst_count[0]), .D(srst_count[1]), .A(n9), .B(n28), .Y(n30) );
  INVX1 U32 ( .A(n29), .Y(n4) );
  AOI32X1 U33 ( .A(n9), .B(n7), .C(n5), .D(srst_count[2]), .E(n22), .Y(n29) );
  NOR2X1 U34 ( .A(srst_count[0]), .B(n16), .Y(N38) );
  AND4XL U35 ( .A(sfrwe), .B(sfraddr[6]), .C(sfraddr[5]), .D(sfraddr[4]), .Y(
        n21) );
endmodule


module SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2c_a0 ( clk, rst, bclksel, scli, sdai, sclo, sdao, intack, si, sfrwe, 
        sfraddr, sfrdatai, i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o, test_si, 
        test_so, test_se );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  output [7:0] i2cdat_o;
  output [7:0] i2cadr_o;
  output [7:0] i2ccon_o;
  output [7:0] i2csta_o;
  input clk, rst, bclksel, scli, sdai, intack, sfrwe, test_si, test_se;
  output sclo, sdao, si, test_so;
  wire   scli_ff, N180, sdai_ff, N181, sclo_int, wait_for_setup_r, adrcomp,
         adrcompen, nedetect, ack_bit, bsd7, pedetect, N224, N225, N226, N227,
         N232, N233, N234, sclint, ack, sdaint, bsd7_tmp, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N332, N333, N335, N336, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N406, N407, N408,
         N409, N410, N412, N413, N414, N431, N432, N433, N468, N469, N470,
         N471, N491, N492, N493, N494, N495, busfree, N510, N511, rst_delay,
         clk_count1_ov, N653, N654, N655, N656, N657, clk_count2_ov, N685,
         N686, N687, N688, N689, N690, clkint, clkint_ff, N700, N746, N747,
         N748, N749, N1022, N1023, N1024, N1025, N1026, N1027, N1063, N1064,
         N1065, sclscl, starto_en, N1124, N1125, N1126, net12037, net12043,
         net12048, net12053, net12058, net12063, net12068, net12073, net12078,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n7, n8, n9, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n282, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452;
  wire   [2:0] fsmmod;
  wire   [4:0] fsmsta;
  wire   [3:0] framesync;
  wire   [2:0] fsmdet;
  wire   [2:0] setup_counter_r;
  wire   [2:0] scli_ff_reg0;
  wire   [2:0] sdai_ff_reg0;
  wire   [2:0] indelay;
  wire   [2:0] fsmsync;
  wire   [1:0] bclkcnt;
  wire   [3:0] clk_count1;
  wire   [3:0] clk_count2;

  SNPS_CLOCK_GATE_HIGH_i2c_a0_0 clk_gate_i2ccon_reg ( .CLK(clk), .EN(N224), 
        .ENCLK(net12037), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_8 clk_gate_i2cdat_reg ( .CLK(clk), .EN(N296), 
        .ENCLK(net12043), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_7 clk_gate_setup_counter_r_reg ( .CLK(clk), .EN(
        N332), .ENCLK(net12048), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_6 clk_gate_i2cadr_reg ( .CLK(clk), .EN(N342), 
        .ENCLK(net12053), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_5 clk_gate_indelay_reg ( .CLK(clk), .EN(N468), 
        .ENCLK(net12058), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_4 clk_gate_framesync_reg ( .CLK(clk), .EN(N491), 
        .ENCLK(net12063), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_3 clk_gate_clk_count1_reg ( .CLK(clk), .EN(N653), 
        .ENCLK(net12068), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_2 clk_gate_clk_count2_reg ( .CLK(clk), .EN(N689), 
        .ENCLK(net12073), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_1 clk_gate_fsmsta_reg ( .CLK(clk), .EN(N1022), 
        .ENCLK(net12078), .TE(test_se) );
  SDFFQX1 scli_ff_reg ( .D(N180), .SIN(rst_delay), .SMC(test_se), .C(clk), .Q(
        scli_ff) );
  SDFFQX1 sdai_ff_reg ( .D(N181), .SIN(sclscl), .SMC(test_se), .C(clk), .Q(
        sdai_ff) );
  SDFFQX1 clk_count2_ov_reg ( .D(N690), .SIN(clk_count1[3]), .SMC(test_se), 
        .C(clk), .Q(clk_count2_ov) );
  SDFFQX1 sdai_ff_reg_reg_2_ ( .D(N433), .SIN(sdai_ff_reg0[1]), .SMC(test_se), 
        .C(clk), .Q(sdai_ff_reg0[2]) );
  SDFFQX1 sdai_ff_reg_reg_1_ ( .D(N432), .SIN(sdai_ff_reg0[0]), .SMC(test_se), 
        .C(clk), .Q(sdai_ff_reg0[1]) );
  SDFFQX1 clk_count1_ov_reg ( .D(n505), .SIN(busfree), .SMC(test_se), .C(clk), 
        .Q(clk_count1_ov) );
  SDFFQX1 rst_delay_reg ( .D(n25), .SIN(pedetect), .SMC(test_se), .C(clk), .Q(
        rst_delay) );
  SDFFQX1 ack_bit_reg ( .D(n494), .SIN(test_si), .SMC(test_se), .C(net12037), 
        .Q(ack_bit) );
  SDFFQX1 bsd7_reg ( .D(n491), .SIN(bclkcnt[1]), .SMC(test_se), .C(clk), .Q(
        bsd7) );
  SDFFQX1 clk_count2_reg_3_ ( .D(N688), .SIN(clk_count2[2]), .SMC(test_se), 
        .C(net12073), .Q(clk_count2[3]) );
  SDFFQX1 sdai_ff_reg_reg_0_ ( .D(N431), .SIN(sdai_ff), .SMC(test_se), .C(clk), 
        .Q(sdai_ff_reg0[0]) );
  SDFFQX1 sclscl_reg ( .D(n48), .SIN(sclo_int), .SMC(test_se), .C(clk), .Q(
        sclscl) );
  SDFFQX1 setup_counter_r_reg_2_ ( .D(N335), .SIN(setup_counter_r[1]), .SMC(
        test_se), .C(net12048), .Q(setup_counter_r[2]) );
  SDFFQX1 clk_count2_reg_1_ ( .D(N686), .SIN(clk_count2[0]), .SMC(test_se), 
        .C(net12073), .Q(clk_count2[1]) );
  SDFFQX1 clk_count2_reg_2_ ( .D(N687), .SIN(clk_count2[1]), .SMC(test_se), 
        .C(net12073), .Q(clk_count2[2]) );
  SDFFQX1 bclkcnt_reg_1_ ( .D(N511), .SIN(bclkcnt[0]), .SMC(test_se), .C(clk), 
        .Q(bclkcnt[1]) );
  SDFFQX1 indelay_reg_2_ ( .D(N471), .SIN(indelay[1]), .SMC(test_se), .C(
        net12058), .Q(indelay[2]) );
  SDFFQX1 bclkcnt_reg_0_ ( .D(N510), .SIN(adrcompen), .SMC(test_se), .C(clk), 
        .Q(bclkcnt[0]) );
  SDFFQX1 clkint_ff_reg ( .D(N700), .SIN(clk_count2[3]), .SMC(test_se), .C(clk), .Q(clkint_ff) );
  SDFFQX1 setup_counter_r_reg_0_ ( .D(N333), .SIN(sdao), .SMC(test_se), .C(
        net12048), .Q(setup_counter_r[0]) );
  SDFFQX1 write_data_r_reg ( .D(n500), .SIN(wait_for_setup_r), .SMC(test_se), 
        .C(clk), .Q(test_so) );
  SDFFQX1 clk_count2_reg_0_ ( .D(N685), .SIN(clk_count2_ov), .SMC(test_se), 
        .C(net12073), .Q(clk_count2[0]) );
  SDFFQX1 bsd7_tmp_reg ( .D(n492), .SIN(bsd7), .SMC(test_se), .C(clk), .Q(
        bsd7_tmp) );
  SDFFQX1 busfree_reg ( .D(n506), .SIN(bsd7_tmp), .SMC(test_se), .C(clk), .Q(
        busfree) );
  SDFFQX1 indelay_reg_1_ ( .D(N470), .SIN(indelay[0]), .SMC(test_se), .C(
        net12058), .Q(indelay[1]) );
  SDFFQX1 clkint_reg ( .D(n504), .SIN(clkint_ff), .SMC(test_se), .C(clk), .Q(
        clkint) );
  SDFFQX1 indelay_reg_0_ ( .D(N469), .SIN(i2csta_o[7]), .SMC(test_se), .C(
        net12058), .Q(indelay[0]) );
  SDFFQX1 starto_en_reg ( .D(n490), .SIN(setup_counter_r[2]), .SMC(test_se), 
        .C(clk), .Q(starto_en) );
  SDFFQX1 scli_ff_reg_reg_1_ ( .D(N413), .SIN(scli_ff_reg0[0]), .SMC(test_se), 
        .C(clk), .Q(scli_ff_reg0[1]) );
  SDFFQX1 scli_ff_reg_reg_0_ ( .D(N412), .SIN(scli_ff), .SMC(test_se), .C(clk), 
        .Q(scli_ff_reg0[0]) );
  SDFFQX1 setup_counter_r_reg_1_ ( .D(n40), .SIN(setup_counter_r[0]), .SMC(
        test_se), .C(net12048), .Q(setup_counter_r[1]) );
  SDFFQX1 scli_ff_reg_reg_2_ ( .D(N414), .SIN(scli_ff_reg0[1]), .SMC(test_se), 
        .C(clk), .Q(scli_ff_reg0[2]) );
  SDFFQX1 fsmsync_reg_1_ ( .D(N747), .SIN(fsmsync[0]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[1]) );
  SDFFQX1 fsmsync_reg_0_ ( .D(N746), .SIN(fsmsta[4]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[0]) );
  SDFFQX1 fsmsync_reg_2_ ( .D(N748), .SIN(fsmsync[1]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[2]) );
  SDFFQX1 pedetect_reg ( .D(n497), .SIN(nedetect), .SMC(test_se), .C(clk), .Q(
        pedetect) );
  SDFFQX1 nedetect_reg ( .D(n498), .SIN(indelay[2]), .SMC(test_se), .C(clk), 
        .Q(nedetect) );
  SDFFQX1 sclint_reg ( .D(n499), .SIN(scli_ff_reg0[2]), .SMC(test_se), .C(clk), 
        .Q(sclint) );
  SDFFQX1 clk_count1_reg_2_ ( .D(N656), .SIN(clk_count1[1]), .SMC(test_se), 
        .C(net12068), .Q(clk_count1[2]) );
  SDFFQX1 clk_count1_reg_3_ ( .D(N657), .SIN(clk_count1[2]), .SMC(test_se), 
        .C(net12068), .Q(clk_count1[3]) );
  SDFFQX1 adrcompen_reg ( .D(n496), .SIN(adrcomp), .SMC(test_se), .C(clk), .Q(
        adrcompen) );
  SDFFQX1 adrcomp_reg ( .D(n501), .SIN(ack), .SMC(test_se), .C(clk), .Q(
        adrcomp) );
  SDFFQX1 clk_count1_reg_1_ ( .D(N655), .SIN(clk_count1[0]), .SMC(test_se), 
        .C(net12068), .Q(clk_count1[1]) );
  SDFFQX1 clk_count1_reg_0_ ( .D(N654), .SIN(clk_count1_ov), .SMC(test_se), 
        .C(net12068), .Q(clk_count1[0]) );
  SDFFQX1 ack_reg ( .D(n493), .SIN(ack_bit), .SMC(test_se), .C(clk), .Q(ack)
         );
  SDFFQX1 sdaint_reg ( .D(n507), .SIN(sdai_ff_reg0[2]), .SMC(test_se), .C(clk), 
        .Q(sdaint) );
  SDFFQX1 fsmdet_reg_0_ ( .D(N1063), .SIN(framesync[3]), .SMC(test_se), .C(clk), .Q(fsmdet[0]) );
  SDFFQX1 fsmdet_reg_1_ ( .D(N1064), .SIN(fsmdet[0]), .SMC(test_se), .C(clk), 
        .Q(fsmdet[1]) );
  SDFFQX1 framesync_reg_3_ ( .D(N495), .SIN(framesync[2]), .SMC(test_se), .C(
        net12063), .Q(framesync[3]) );
  SDFFQX1 fsmmod_reg_0_ ( .D(N1124), .SIN(fsmdet[2]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[0]) );
  SDFFQX1 fsmmod_reg_1_ ( .D(N1125), .SIN(fsmmod[0]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[1]) );
  SDFFQX1 fsmdet_reg_2_ ( .D(N1065), .SIN(fsmdet[1]), .SMC(test_se), .C(clk), 
        .Q(fsmdet[2]) );
  SDFFQX1 fsmmod_reg_2_ ( .D(N1126), .SIN(fsmmod[1]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[2]) );
  SDFFQX1 framesync_reg_1_ ( .D(N493), .SIN(framesync[0]), .SMC(test_se), .C(
        net12063), .Q(framesync[1]) );
  SDFFQX1 framesync_reg_2_ ( .D(N494), .SIN(framesync[1]), .SMC(test_se), .C(
        net12063), .Q(framesync[2]) );
  SDFFQX1 framesync_reg_0_ ( .D(N492), .SIN(clkint), .SMC(test_se), .C(
        net12063), .Q(framesync[0]) );
  SDFFQX1 fsmsta_reg_4_ ( .D(N1027), .SIN(n9), .SMC(test_se), .C(net12078), 
        .Q(fsmsta[4]) );
  SDFFQX1 fsmsta_reg_0_ ( .D(N1023), .SIN(fsmmod[2]), .SMC(test_se), .C(
        net12078), .Q(fsmsta[0]) );
  SDFFQX1 fsmsta_reg_2_ ( .D(N1025), .SIN(fsmsta[1]), .SMC(test_se), .C(
        net12078), .Q(fsmsta[2]) );
  SDFFQX1 fsmsta_reg_1_ ( .D(N1024), .SIN(fsmsta[0]), .SMC(test_se), .C(
        net12078), .Q(fsmsta[1]) );
  SDFFQX1 fsmsta_reg_3_ ( .D(N1026), .SIN(fsmsta[2]), .SMC(test_se), .C(
        net12078), .Q(fsmsta[3]) );
  SDFFQX1 i2csta_reg_4_ ( .D(N410), .SIN(i2csta_o[6]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[7]) );
  SDFFQX1 i2csta_reg_3_ ( .D(N409), .SIN(i2csta_o[5]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[6]) );
  SDFFQX1 i2cdat_reg_7_ ( .D(N304), .SIN(i2cdat_o[6]), .SMC(test_se), .C(
        net12043), .Q(i2cdat_o[7]) );
  SDFFQX1 i2cadr_reg_3_ ( .D(N346), .SIN(i2cadr_o[2]), .SMC(test_se), .C(
        net12053), .Q(i2cadr_o[3]) );
  SDFFQX1 i2ccon_reg_5_ ( .D(N232), .SIN(i2ccon_o[4]), .SMC(test_se), .C(
        net12037), .Q(i2ccon_o[5]) );
  SDFFQX1 i2ccon_reg_1_ ( .D(N226), .SIN(i2ccon_o[0]), .SMC(test_se), .C(
        net12037), .Q(i2ccon_o[1]) );
  SDFFQX1 i2cdat_reg_3_ ( .D(N300), .SIN(i2cdat_o[2]), .SMC(test_se), .C(
        net12043), .Q(i2cdat_o[3]) );
  SDFFQX1 i2cdat_reg_6_ ( .D(N303), .SIN(i2cdat_o[5]), .SMC(test_se), .C(
        net12043), .Q(i2cdat_o[6]) );
  SDFFQX1 i2ccon_reg_6_ ( .D(N233), .SIN(i2ccon_o[5]), .SMC(test_se), .C(
        net12037), .Q(i2ccon_o[6]) );
  SDFFQX1 i2cadr_reg_0_ ( .D(N343), .SIN(fsmsync[2]), .SMC(test_se), .C(
        net12053), .Q(i2cadr_o[0]) );
  SDFFQX1 i2ccon_reg_0_ ( .D(N225), .SIN(i2cadr_o[7]), .SMC(test_se), .C(
        net12037), .Q(i2ccon_o[0]) );
  SDFFQX1 i2ccon_reg_7_ ( .D(N234), .SIN(i2ccon_o[6]), .SMC(test_se), .C(
        net12037), .Q(i2ccon_o[7]) );
  SDFFQX1 i2ccon_reg_4_ ( .D(n503), .SIN(si), .SMC(test_se), .C(clk), .Q(
        i2ccon_o[4]) );
  SDFFQX1 i2ccon_reg_3_ ( .D(n495), .SIN(i2ccon_o[2]), .SMC(test_se), .C(clk), 
        .Q(i2ccon_o[3]) );
  SDFFQX1 i2csta_reg_0_ ( .D(N406), .SIN(i2cdat_o[7]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[3]) );
  SDFFQX1 i2csta_reg_1_ ( .D(N407), .SIN(i2csta_o[3]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[4]) );
  SDFFQX1 i2csta_reg_2_ ( .D(N408), .SIN(i2csta_o[4]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[5]) );
  SDFFQX1 i2cadr_reg_4_ ( .D(N347), .SIN(i2cadr_o[3]), .SMC(test_se), .C(
        net12053), .Q(i2cadr_o[4]) );
  SDFFQX1 i2cadr_reg_5_ ( .D(N348), .SIN(i2cadr_o[4]), .SMC(test_se), .C(
        net12053), .Q(i2cadr_o[5]) );
  SDFFQX1 i2cadr_reg_6_ ( .D(N349), .SIN(i2cadr_o[5]), .SMC(test_se), .C(
        net12053), .Q(i2cadr_o[6]) );
  SDFFQX1 i2cadr_reg_7_ ( .D(N350), .SIN(i2cadr_o[6]), .SMC(test_se), .C(
        net12053), .Q(i2cadr_o[7]) );
  SDFFQX1 i2cadr_reg_2_ ( .D(N345), .SIN(i2cadr_o[1]), .SMC(test_se), .C(
        net12053), .Q(i2cadr_o[2]) );
  SDFFQX1 i2cadr_reg_1_ ( .D(N344), .SIN(i2cadr_o[0]), .SMC(test_se), .C(
        net12053), .Q(i2cadr_o[1]) );
  SDFFQX1 i2cdat_reg_5_ ( .D(N302), .SIN(i2cdat_o[4]), .SMC(test_se), .C(
        net12043), .Q(i2cdat_o[5]) );
  SDFFQX1 i2cdat_reg_4_ ( .D(N301), .SIN(i2cdat_o[3]), .SMC(test_se), .C(
        net12043), .Q(i2cdat_o[4]) );
  SDFFQX1 i2ccon_reg_2_ ( .D(N227), .SIN(i2ccon_o[1]), .SMC(test_se), .C(
        net12037), .Q(i2ccon_o[2]) );
  SDFFQX1 i2cdat_reg_1_ ( .D(N298), .SIN(i2cdat_o[0]), .SMC(test_se), .C(
        net12043), .Q(i2cdat_o[1]) );
  SDFFQX1 i2cdat_reg_2_ ( .D(N299), .SIN(i2cdat_o[1]), .SMC(test_se), .C(
        net12043), .Q(i2cdat_o[2]) );
  SDFFQX1 i2cdat_reg_0_ ( .D(N297), .SIN(i2ccon_o[7]), .SMC(test_se), .C(
        net12043), .Q(i2cdat_o[0]) );
  SDFFQX1 sdao_int_reg ( .D(n502), .SIN(sdaint), .SMC(test_se), .C(clk), .Q(
        sdao) );
  SDFFQX1 wait_for_setup_r_reg ( .D(N336), .SIN(starto_en), .SMC(test_se), .C(
        clk), .Q(wait_for_setup_r) );
  SDFFQX1 sclo_int_reg ( .D(N749), .SIN(sclint), .SMC(test_se), .C(clk), .Q(
        sclo_int) );
  INVX1 U3 ( .A(1'b1), .Y(i2csta_o[0]) );
  INVX1 U5 ( .A(1'b1), .Y(i2csta_o[1]) );
  INVX1 U7 ( .A(1'b1), .Y(i2csta_o[2]) );
  BUFX3 U9 ( .A(n441), .Y(n7) );
  INVX1 U10 ( .A(si), .Y(n8) );
  INVX1 U11 ( .A(n437), .Y(n9) );
  INVX1 U12 ( .A(n193), .Y(n10) );
  BUFX3 U13 ( .A(i2ccon_o[3]), .Y(si) );
  INVX1 U14 ( .A(n83), .Y(n12) );
  NAND2X1 U15 ( .A(framesync[3]), .B(n207), .Y(n13) );
  NOR4XL U16 ( .A(n108), .B(n441), .C(fsmsta[0]), .D(fsmsta[3]), .Y(n162) );
  INVX1 U17 ( .A(n27), .Y(n23) );
  INVX1 U18 ( .A(n27), .Y(n24) );
  INVX1 U19 ( .A(n224), .Y(n34) );
  INVX1 U20 ( .A(n135), .Y(n31) );
  NAND2X1 U21 ( .A(n23), .B(n135), .Y(N224) );
  OAI21X1 U22 ( .B(n309), .C(n15), .A(n29), .Y(N343) );
  OAI21X1 U23 ( .B(n18), .C(n309), .A(n24), .Y(N346) );
  OAI21X1 U24 ( .B(n22), .C(n309), .A(n24), .Y(N350) );
  NOR2X1 U25 ( .A(n309), .B(n16), .Y(N344) );
  NOR2X1 U26 ( .A(n309), .B(n20), .Y(N348) );
  NOR2X1 U27 ( .A(n309), .B(n17), .Y(N345) );
  NOR2X1 U28 ( .A(n309), .B(n21), .Y(N349) );
  NOR2X1 U29 ( .A(n19), .B(n309), .Y(N347) );
  NAND2X1 U30 ( .A(n23), .B(n309), .Y(N342) );
  NOR2X1 U31 ( .A(n26), .B(n15), .Y(N225) );
  NOR2X1 U32 ( .A(n27), .B(n22), .Y(N234) );
  NOR2X1 U33 ( .A(n26), .B(n17), .Y(N227) );
  NOR2X1 U34 ( .A(n27), .B(n21), .Y(N233) );
  NOR2X1 U35 ( .A(n26), .B(n16), .Y(N226) );
  NOR2X1 U36 ( .A(n26), .B(n20), .Y(N232) );
  INVX1 U37 ( .A(n28), .Y(n27) );
  INVX1 U38 ( .A(n28), .Y(n26) );
  INVX1 U39 ( .A(n431), .Y(n84) );
  INVX1 U40 ( .A(n29), .Y(n25) );
  NAND21X1 U41 ( .B(sdai), .A(n28), .Y(N181) );
  NAND42X1 U42 ( .C(sfraddr[0]), .D(sfraddr[2]), .A(sfraddr[1]), .B(n311), .Y(
        n224) );
  NOR42XL U43 ( .C(sfraddr[4]), .D(sfraddr[3]), .A(sfraddr[5]), .B(n329), .Y(
        n311) );
  NAND2X1 U44 ( .A(sfrwe), .B(sfraddr[6]), .Y(n329) );
  AOI21X1 U45 ( .B(n224), .C(n228), .A(n318), .Y(n214) );
  NOR2X1 U46 ( .A(n33), .B(n322), .Y(n318) );
  NAND42X1 U47 ( .C(sfraddr[0]), .D(sfraddr[1]), .A(sfraddr[2]), .B(n311), .Y(
        n135) );
  NAND3X1 U48 ( .A(n31), .B(n24), .C(sfrdatai[3]), .Y(n198) );
  NAND4X1 U49 ( .A(sfraddr[0]), .B(sfraddr[1]), .C(n310), .D(n311), .Y(n309)
         );
  NOR2X1 U50 ( .A(sfraddr[2]), .B(n25), .Y(n310) );
  INVX1 U51 ( .A(sfrdatai[4]), .Y(n19) );
  INVX1 U52 ( .A(sfrdatai[5]), .Y(n20) );
  INVX1 U53 ( .A(sfrdatai[6]), .Y(n21) );
  INVX1 U54 ( .A(sfrdatai[1]), .Y(n16) );
  INVX1 U55 ( .A(sfrdatai[2]), .Y(n17) );
  INVX1 U56 ( .A(sfrdatai[7]), .Y(n22) );
  INVX1 U57 ( .A(sfrdatai[0]), .Y(n15) );
  INVX1 U58 ( .A(sfrdatai[3]), .Y(n18) );
  INVX1 U59 ( .A(n324), .Y(n109) );
  NOR32XL U60 ( .B(n84), .C(n433), .A(n157), .Y(n357) );
  NAND2X1 U61 ( .A(n201), .B(n23), .Y(n431) );
  NAND2X1 U62 ( .A(n152), .B(n95), .Y(n376) );
  NOR2X1 U63 ( .A(n86), .B(n210), .Y(n322) );
  INVX1 U64 ( .A(rst), .Y(n28) );
  INVX1 U65 ( .A(n403), .Y(n80) );
  INVX1 U66 ( .A(n228), .Y(n87) );
  AND2X1 U67 ( .A(n385), .B(n386), .Y(n361) );
  NAND41X1 U68 ( .D(n161), .A(n363), .B(n325), .C(n364), .Y(n358) );
  OAI21X1 U69 ( .B(n365), .C(n362), .A(n95), .Y(n363) );
  NAND41X1 U70 ( .D(n357), .A(n75), .B(n403), .C(n430), .Y(N1022) );
  NOR2X1 U71 ( .A(n37), .B(n431), .Y(n430) );
  INVX1 U72 ( .A(rst), .Y(n29) );
  NAND2X1 U73 ( .A(n147), .B(n143), .Y(n145) );
  INVX1 U74 ( .A(n369), .Y(n75) );
  INVX1 U75 ( .A(n132), .Y(n66) );
  INVX1 U76 ( .A(n393), .Y(n96) );
  INVX1 U77 ( .A(n192), .Y(n99) );
  INVX1 U78 ( .A(n251), .Y(n101) );
  NAND2X1 U79 ( .A(n23), .B(n103), .Y(n238) );
  INVX1 U80 ( .A(n308), .Y(n435) );
  INVX1 U81 ( .A(n236), .Y(n282) );
  INVX1 U82 ( .A(n261), .Y(n50) );
  INVX1 U83 ( .A(n231), .Y(n69) );
  INVX1 U84 ( .A(n284), .Y(n35) );
  NAND21X1 U85 ( .B(scli), .A(n28), .Y(N180) );
  OAI21X1 U86 ( .B(n216), .C(n64), .A(n217), .Y(n492) );
  GEN2XL U87 ( .D(n22), .E(n33), .C(n181), .B(n29), .A(n32), .Y(n217) );
  INVX1 U88 ( .A(n216), .Y(n32) );
  OAI21BBX1 U89 ( .A(n34), .B(n215), .C(n218), .Y(n216) );
  OAI22AX1 U90 ( .D(n211), .C(n212), .A(n94), .B(n211), .Y(n493) );
  AND2X1 U91 ( .A(n213), .B(n92), .Y(n212) );
  OAI21X1 U92 ( .B(n214), .C(n78), .A(n213), .Y(n211) );
  NOR2X1 U93 ( .A(n25), .B(n215), .Y(n213) );
  INVX1 U94 ( .A(n226), .Y(n33) );
  OAI22AX1 U95 ( .D(n223), .C(n322), .A(n224), .B(n87), .Y(n320) );
  NOR2X1 U96 ( .A(n319), .B(n320), .Y(n317) );
  OAI32X1 U97 ( .A(n135), .B(n27), .C(n30), .D(n447), .E(n136), .Y(n503) );
  INVX1 U98 ( .A(n136), .Y(n30) );
  OAI221X1 U99 ( .A(n31), .B(n137), .C(n135), .D(n19), .E(n29), .Y(n136) );
  AOI21BBXL U100 ( .B(n123), .C(n122), .A(n119), .Y(n137) );
  AOI21X1 U101 ( .B(n319), .C(n34), .A(n320), .Y(n179) );
  OAI22X1 U102 ( .A(n317), .B(n18), .C(n214), .D(n443), .Y(N300) );
  OAI22X1 U103 ( .A(n317), .B(n16), .C(n214), .D(n449), .Y(N298) );
  OAI22X1 U104 ( .A(n317), .B(n17), .C(n214), .D(n450), .Y(N299) );
  OAI22X1 U105 ( .A(n317), .B(n15), .C(n214), .D(n94), .Y(N297) );
  AOI22X1 U106 ( .A(n86), .B(n223), .C(n215), .D(n224), .Y(n222) );
  NOR2X1 U107 ( .A(n440), .B(n441), .Y(n159) );
  OAI221X1 U108 ( .A(n374), .B(n377), .C(n393), .D(n302), .E(n407), .Y(n392)
         );
  AOI222XL U109 ( .A(n408), .B(n193), .C(n434), .D(n160), .E(n409), .F(n410), 
        .Y(n407) );
  INVX1 U110 ( .A(n303), .Y(n434) );
  OAI221X1 U111 ( .A(n13), .B(n384), .C(n10), .D(n296), .E(n383), .Y(n410) );
  INVX1 U112 ( .A(n193), .Y(n95) );
  NAND2X1 U113 ( .A(n398), .B(n159), .Y(n324) );
  NAND2X1 U114 ( .A(n328), .B(n441), .Y(n296) );
  NAND2X1 U115 ( .A(n109), .B(n437), .Y(n383) );
  NOR21XL U116 ( .B(n323), .A(n150), .Y(n228) );
  NAND42X1 U117 ( .C(n336), .D(n251), .A(n151), .B(n100), .Y(n164) );
  NAND42X1 U118 ( .C(n423), .D(n399), .A(n364), .B(n424), .Y(n406) );
  NAND4X1 U119 ( .A(n328), .B(n159), .C(n93), .D(n13), .Y(n424) );
  OAI22X1 U120 ( .A(n385), .B(n393), .C(n386), .D(n394), .Y(n423) );
  OAI211X1 U121 ( .C(n305), .D(n436), .A(n324), .B(n325), .Y(n150) );
  NOR2X1 U122 ( .A(n193), .B(n452), .Y(n393) );
  NOR4XL U123 ( .A(n431), .B(n78), .C(n157), .D(n433), .Y(n369) );
  NOR2X1 U124 ( .A(n102), .B(n105), .Y(n251) );
  AND2X1 U125 ( .A(n323), .B(n150), .Y(n210) );
  NOR2X1 U126 ( .A(n26), .B(n194), .Y(n121) );
  AOI21X1 U127 ( .B(n194), .C(n342), .A(n420), .Y(n201) );
  NAND4X1 U128 ( .A(n84), .B(n205), .C(n202), .D(n157), .Y(n403) );
  OAI21X1 U129 ( .B(n387), .C(n75), .A(n388), .Y(N1025) );
  OAI21BBX1 U130 ( .A(n166), .B(n94), .C(n357), .Y(n388) );
  NOR4XL U131 ( .A(n389), .B(n390), .C(n391), .D(n392), .Y(n387) );
  NOR2X1 U132 ( .A(n95), .B(n380), .Y(n391) );
  NOR2X1 U133 ( .A(n181), .B(n38), .Y(n215) );
  NAND3X1 U134 ( .A(n295), .B(n110), .C(n306), .Y(n384) );
  INVX1 U135 ( .A(n315), .Y(n41) );
  NAND2X1 U136 ( .A(n194), .B(n446), .Y(n180) );
  INVX1 U137 ( .A(n233), .Y(n446) );
  NAND3X1 U138 ( .A(n160), .B(n110), .C(n295), .Y(n325) );
  INVX1 U139 ( .A(n366), .Y(n37) );
  OAI211X1 U140 ( .C(n418), .D(n75), .A(n367), .B(n419), .Y(N1023) );
  NOR2X1 U141 ( .A(n420), .B(n37), .Y(n419) );
  NOR4XL U142 ( .A(n421), .B(n406), .C(n422), .D(n359), .Y(n418) );
  AOI21X1 U143 ( .B(n411), .C(n383), .A(n393), .Y(n422) );
  INVX1 U144 ( .A(n181), .Y(n86) );
  NAND2X1 U145 ( .A(n379), .B(n383), .Y(n408) );
  INVX1 U146 ( .A(n194), .Y(n85) );
  INVX1 U147 ( .A(n428), .Y(n106) );
  OAI211X1 U148 ( .C(n108), .D(n429), .A(n378), .B(n400), .Y(n428) );
  NAND2X1 U149 ( .A(n441), .B(n437), .Y(n429) );
  INVX1 U150 ( .A(n154), .Y(n100) );
  INVX1 U151 ( .A(n326), .Y(n111) );
  INVX1 U152 ( .A(n398), .Y(n108) );
  NOR21XL U153 ( .B(n151), .A(n152), .Y(n147) );
  NOR2X1 U154 ( .A(n276), .B(n25), .Y(n125) );
  INVX1 U155 ( .A(n206), .Y(n97) );
  NOR2X1 U156 ( .A(n72), .B(n67), .Y(n132) );
  OAI21X1 U157 ( .B(n149), .C(n95), .A(n150), .Y(n143) );
  NOR2X1 U158 ( .A(n447), .B(n164), .Y(n192) );
  AND3X1 U159 ( .A(n380), .B(n325), .C(n384), .Y(n411) );
  NAND2X1 U160 ( .A(n85), .B(n138), .Y(n157) );
  OAI31XL U161 ( .A(n376), .B(n94), .C(n107), .D(n282), .Y(n359) );
  OAI22X1 U162 ( .A(n393), .B(n386), .C(n374), .D(n378), .Y(n390) );
  NOR2X1 U163 ( .A(n77), .B(n79), .Y(n152) );
  AND2X1 U164 ( .A(n382), .B(n92), .Y(n399) );
  AOI21X1 U165 ( .B(n94), .C(n357), .A(n27), .Y(n367) );
  NOR3XL U166 ( .A(n78), .B(n162), .C(n376), .Y(n433) );
  AOI211X1 U167 ( .C(n107), .D(n164), .A(n165), .B(n77), .Y(n163) );
  OAI21X1 U168 ( .B(n166), .C(n94), .A(n167), .Y(n165) );
  OAI22X1 U169 ( .A(n166), .B(n448), .C(n168), .D(n169), .Y(n167) );
  NAND3X1 U170 ( .A(n170), .B(n171), .C(n172), .Y(n169) );
  OAI22AX1 U171 ( .D(n139), .C(n140), .A(n139), .B(n452), .Y(n502) );
  NOR32XL U172 ( .B(n446), .C(n141), .A(n142), .Y(n140) );
  NAND4X1 U173 ( .A(n446), .B(n141), .C(n148), .D(n147), .Y(n139) );
  AOI21X1 U174 ( .B(n79), .C(n153), .A(n154), .Y(n141) );
  NOR3XL U175 ( .A(n193), .B(n94), .C(n296), .Y(n382) );
  OAI31XL U176 ( .A(n78), .B(n186), .C(n182), .D(n187), .Y(n497) );
  NAND4X1 U177 ( .A(n23), .B(n83), .C(n183), .D(n188), .Y(n187) );
  NOR3XL U178 ( .A(n46), .B(n53), .C(n52), .Y(n188) );
  OAI31XL U179 ( .A(n42), .B(n313), .C(n41), .D(n312), .Y(N335) );
  AOI211X1 U180 ( .C(n50), .D(n55), .A(n260), .B(n263), .Y(N687) );
  AOI211X1 U181 ( .C(n54), .D(n51), .A(n260), .B(n261), .Y(N686) );
  AOI211X1 U182 ( .C(n72), .D(n67), .A(n267), .B(n132), .Y(N655) );
  NAND2X1 U183 ( .A(n306), .B(n159), .Y(n385) );
  NAND2X1 U184 ( .A(n425), .B(n441), .Y(n386) );
  NAND2X1 U185 ( .A(n95), .B(n452), .Y(n394) );
  NAND2X1 U186 ( .A(n377), .B(n378), .Y(n362) );
  NAND2X1 U187 ( .A(n52), .B(n29), .Y(N414) );
  NAND2X1 U188 ( .A(n53), .B(n23), .Y(N413) );
  NAND2X1 U189 ( .A(n379), .B(n380), .Y(n365) );
  NAND2X1 U190 ( .A(n41), .B(n312), .Y(N336) );
  NAND2X1 U191 ( .A(n23), .B(n118), .Y(n506) );
  OAI21X1 U192 ( .B(n119), .C(n120), .A(n121), .Y(n118) );
  OAI31XL U193 ( .A(n83), .B(n122), .C(n123), .D(n65), .Y(n120) );
  NAND2X1 U194 ( .A(n125), .B(n73), .Y(N700) );
  INVX1 U195 ( .A(n305), .Y(n113) );
  INVX1 U196 ( .A(n162), .Y(n107) );
  INVX1 U197 ( .A(n287), .Y(n98) );
  INVX1 U198 ( .A(n306), .Y(n436) );
  NOR2X1 U199 ( .A(n38), .B(n25), .Y(n300) );
  NAND21X1 U200 ( .B(n242), .A(n71), .Y(n240) );
  NOR2X1 U201 ( .A(n51), .B(n54), .Y(n261) );
  NOR2X1 U202 ( .A(n70), .B(n82), .Y(n231) );
  NOR2X1 U203 ( .A(n435), .B(n305), .Y(n236) );
  NOR2X1 U204 ( .A(n437), .B(n442), .Y(n308) );
  NOR2X1 U205 ( .A(n293), .B(n95), .Y(n284) );
  NOR2X1 U206 ( .A(n113), .B(n442), .Y(n161) );
  NOR2X1 U207 ( .A(n55), .B(n50), .Y(n263) );
  AOI21X1 U208 ( .B(n49), .C(n81), .A(n69), .Y(n257) );
  AOI21X1 U209 ( .B(n132), .C(n62), .A(n63), .Y(n126) );
  INVX1 U210 ( .A(n183), .Y(n45) );
  NAND2X1 U211 ( .A(n159), .B(n160), .Y(n364) );
  NOR2X1 U212 ( .A(n81), .B(n70), .Y(n244) );
  OAI21AX1 U213 ( .B(n83), .C(n45), .A(n182), .Y(n499) );
  INVX1 U214 ( .A(n409), .Y(n93) );
  INVX1 U215 ( .A(n297), .Y(n68) );
  NAND4X1 U216 ( .A(n300), .B(n301), .C(n302), .D(n438), .Y(N410) );
  NAND2X1 U217 ( .A(n161), .B(n7), .Y(n301) );
  NAND2X1 U218 ( .A(n122), .B(n61), .Y(n338) );
  INVX1 U219 ( .A(n253), .Y(n61) );
  INVX1 U220 ( .A(n243), .Y(n71) );
  INVX1 U221 ( .A(n160), .Y(n438) );
  NOR2X1 U222 ( .A(n299), .B(n68), .Y(N470) );
  XNOR2XL U223 ( .A(n56), .B(n57), .Y(n299) );
  INVX1 U224 ( .A(n245), .Y(n49) );
  NAND2X1 U225 ( .A(n297), .B(n49), .Y(N468) );
  INVX1 U226 ( .A(n153), .Y(n103) );
  INVX1 U227 ( .A(n122), .Y(n60) );
  INVX1 U228 ( .A(n339), .Y(n59) );
  INVX1 U229 ( .A(n258), .Y(n39) );
  INVX1 U230 ( .A(n295), .Y(n439) );
  NOR2X1 U231 ( .A(n91), .B(n90), .Y(n351) );
  NAND4X1 U232 ( .A(n291), .B(n121), .C(n293), .D(n97), .Y(N491) );
  INVX1 U233 ( .A(n133), .Y(n62) );
  NOR2X1 U234 ( .A(wait_for_setup_r), .B(n451), .Y(sclo) );
  INVX1 U235 ( .A(sclo_int), .Y(n451) );
  AO22AXL U236 ( .A(n219), .B(n220), .C(bsd7), .D(n220), .Y(n491) );
  OAI211X1 U237 ( .C(n227), .D(n181), .A(n24), .B(n221), .Y(n219) );
  NAND3X1 U238 ( .A(n221), .B(n218), .C(n222), .Y(n220) );
  NOR2X1 U239 ( .A(n210), .B(n228), .Y(n221) );
  NOR2X1 U240 ( .A(i2ccon_o[3]), .B(n34), .Y(n226) );
  AND3X1 U241 ( .A(n180), .B(n225), .C(n24), .Y(n218) );
  NAND4X1 U242 ( .A(n226), .B(n86), .C(nedetect), .D(n78), .Y(n225) );
  AOI221XL U243 ( .A(i2cdat_o[7]), .B(n226), .C(sfrdatai[7]), .D(n223), .E(
        n229), .Y(n227) );
  AOI21X1 U244 ( .B(n83), .C(n64), .A(n38), .Y(n229) );
  NOR2X1 U245 ( .A(n224), .B(i2ccon_o[3]), .Y(n223) );
  OAI21X1 U246 ( .B(intack), .C(N224), .A(n198), .Y(n199) );
  OAI22AX1 U247 ( .D(i2cdat_o[4]), .C(n214), .A(n317), .B(n20), .Y(N302) );
  OAI22AX1 U248 ( .D(i2cdat_o[3]), .C(n214), .A(n317), .B(n19), .Y(N301) );
  OAI22AX1 U249 ( .D(i2cdat_o[5]), .C(n214), .A(n317), .B(n21), .Y(N303) );
  OAI22AX1 U250 ( .D(i2cdat_o[6]), .C(n214), .A(n317), .B(n22), .Y(N304) );
  OAI21X1 U251 ( .B(n177), .C(n178), .A(n179), .Y(n500) );
  NAND3X1 U252 ( .A(n446), .B(n31), .C(test_so), .Y(n178) );
  NAND4X1 U253 ( .A(n180), .B(n87), .C(n33), .D(n181), .Y(n177) );
  ENOX1 U254 ( .A(n38), .B(n195), .C(n195), .D(n196), .Y(n495) );
  OAI21X1 U255 ( .B(n197), .C(N224), .A(n198), .Y(n196) );
  NAND2X1 U256 ( .A(n199), .B(n197), .Y(n195) );
  OAI21BBX1 U257 ( .A(n200), .B(n201), .C(i2ccon_o[6]), .Y(n197) );
  NAND3X1 U258 ( .A(n321), .B(n24), .C(n179), .Y(N296) );
  OAI21X1 U259 ( .B(n318), .C(n228), .A(pedetect), .Y(n321) );
  ENOX1 U260 ( .A(n208), .B(n209), .C(n208), .D(ack_bit), .Y(n494) );
  NOR2X1 U261 ( .A(n25), .B(sfrdatai[2]), .Y(n209) );
  AOI31X1 U262 ( .A(n210), .B(n31), .C(si), .D(n27), .Y(n208) );
  NAND2X1 U263 ( .A(framesync[3]), .B(n207), .Y(n193) );
  NOR3XL U264 ( .A(fsmsta[3]), .B(fsmsta[4]), .C(fsmsta[2]), .Y(n328) );
  INVX1 U265 ( .A(fsmsta[1]), .Y(n441) );
  NOR2X1 U266 ( .A(n110), .B(fsmsta[4]), .Y(n398) );
  NOR3XL U267 ( .A(framesync[1]), .B(framesync[2]), .C(framesync[0]), .Y(n207)
         );
  INVX1 U268 ( .A(fsmsta[2]), .Y(n110) );
  OAI221X1 U269 ( .A(n401), .B(n75), .C(n79), .D(n366), .E(n402), .Y(N1024) );
  AOI31X1 U270 ( .A(n166), .B(n94), .C(n357), .D(n80), .Y(n402) );
  NOR4XL U271 ( .A(n404), .B(n405), .C(n392), .D(n406), .Y(n401) );
  ENOX1 U272 ( .A(n411), .B(n96), .C(n408), .D(sdao), .Y(n405) );
  INVX1 U273 ( .A(fsmsta[0]), .Y(n440) );
  OAI211X1 U274 ( .C(n258), .D(n432), .A(n157), .B(n84), .Y(n366) );
  NOR32XL U275 ( .B(n207), .C(n38), .A(framesync[3]), .Y(n432) );
  OAI31XL U276 ( .A(n327), .B(fsmsta[3]), .C(n159), .D(n112), .Y(n326) );
  INVX1 U277 ( .A(n328), .Y(n112) );
  OAI21X1 U278 ( .B(fsmsta[4]), .C(n441), .A(fsmsta[2]), .Y(n327) );
  AOI22AXL U279 ( .A(n42), .B(n313), .D(n316), .C(n184), .Y(n315) );
  NOR2X1 U280 ( .A(n25), .B(test_so), .Y(n316) );
  NOR3XL U281 ( .A(n88), .B(fsmdet[2]), .C(n90), .Y(n194) );
  NOR2X1 U282 ( .A(n442), .B(fsmsta[3]), .Y(n160) );
  NOR2X1 U283 ( .A(n440), .B(fsmsta[1]), .Y(n295) );
  NOR2X1 U284 ( .A(n437), .B(fsmsta[4]), .Y(n306) );
  NOR3XL U285 ( .A(n104), .B(fsmmod[2]), .C(n102), .Y(n154) );
  NAND3X1 U286 ( .A(i2ccon_o[6]), .B(n326), .C(n121), .Y(n181) );
  INVX1 U287 ( .A(fsmsta[3]), .Y(n437) );
  AND3X1 U288 ( .A(n121), .B(i2ccon_o[6]), .C(n111), .Y(n323) );
  AOI21X1 U289 ( .B(n104), .C(fsmmod[2]), .A(n342), .Y(n151) );
  OAI221X1 U290 ( .A(n322), .B(n38), .C(n25), .D(i2ccon_o[6]), .E(n180), .Y(
        n319) );
  OAI21X1 U291 ( .B(framesync[3]), .C(n207), .A(n13), .Y(n205) );
  NAND2X1 U292 ( .A(n159), .B(fsmsta[2]), .Y(n303) );
  AOI221XL U293 ( .A(n365), .B(n193), .C(n374), .D(n362), .E(n375), .Y(n373)
         );
  OAI22X1 U294 ( .A(ack), .B(n376), .C(n437), .D(n113), .Y(n375) );
  NOR3XL U295 ( .A(n108), .B(fsmsta[0]), .C(n437), .Y(n425) );
  NAND2X1 U296 ( .A(i2ccon_o[6]), .B(n23), .Y(n233) );
  OAI21X1 U297 ( .B(n394), .C(n379), .A(n426), .Y(n421) );
  AOI33X1 U298 ( .A(sdaint), .B(n427), .C(n95), .D(n93), .E(n13), .F(n295), 
        .Y(n426) );
  OAI211X1 U299 ( .C(ack), .D(n296), .A(n377), .B(n106), .Y(n427) );
  NOR3XL U300 ( .A(fsmmod[0]), .B(fsmmod[2]), .C(n102), .Y(n336) );
  NAND2X1 U301 ( .A(sclint), .B(n23), .Y(n184) );
  NOR3XL U302 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(n104), .Y(n342) );
  INVX1 U303 ( .A(fsmsta[4]), .Y(n442) );
  NOR3XL U304 ( .A(n85), .B(fsmmod[0]), .C(n101), .Y(n420) );
  NAND3X1 U305 ( .A(n160), .B(n441), .C(fsmsta[2]), .Y(n378) );
  NAND2X1 U306 ( .A(n425), .B(fsmsta[1]), .Y(n379) );
  AOI32X1 U307 ( .A(pedetect), .B(n202), .C(n95), .D(n203), .E(n157), .Y(n200)
         );
  ENOX1 U308 ( .A(n204), .B(n79), .C(n202), .D(n205), .Y(n203) );
  NOR2X1 U309 ( .A(n206), .B(n207), .Y(n204) );
  INVX1 U310 ( .A(fsmmod[0]), .Y(n104) );
  OR2X1 U311 ( .A(n164), .B(adrcomp), .Y(n202) );
  INVX1 U312 ( .A(fsmmod[1]), .Y(n102) );
  OAI211X1 U313 ( .C(adrcomp), .D(n366), .A(n367), .B(n368), .Y(N1026) );
  AOI21X1 U314 ( .B(n369), .C(n370), .A(n80), .Y(n368) );
  NAND4X1 U315 ( .A(n371), .B(n282), .C(n372), .D(n373), .Y(n370) );
  OAI21BBX1 U316 ( .A(n384), .B(n361), .C(n96), .Y(n371) );
  NAND2X1 U317 ( .A(n328), .B(fsmsta[1]), .Y(n400) );
  INVX1 U318 ( .A(fsmmod[2]), .Y(n105) );
  INVX1 U319 ( .A(fsmdet[1]), .Y(n90) );
  NOR2X1 U320 ( .A(n41), .B(setup_counter_r[0]), .Y(N333) );
  INVX1 U321 ( .A(fsmdet[0]), .Y(n88) );
  INVX1 U322 ( .A(n314), .Y(n40) );
  AOI32X1 U323 ( .A(setup_counter_r[1]), .B(n315), .C(setup_counter_r[0]), .D(
        n44), .E(N333), .Y(n314) );
  INVX1 U324 ( .A(setup_counter_r[1]), .Y(n44) );
  NOR21XL U325 ( .B(framesync[3]), .A(n146), .Y(n206) );
  GEN2XL U326 ( .D(framesync[3]), .E(n283), .C(n149), .B(n284), .A(n285), .Y(
        N495) );
  AO2222XL U327 ( .A(n95), .B(n412), .C(n162), .D(n413), .E(n414), .F(n193), 
        .G(n415), .H(n305), .Y(n404) );
  AOI31X1 U328 ( .A(n438), .B(n436), .C(n435), .D(n441), .Y(n415) );
  OAI22X1 U329 ( .A(ack), .B(n296), .C(n417), .D(n378), .Y(n412) );
  OAI21X1 U330 ( .B(n106), .C(n93), .A(n400), .Y(n414) );
  NAND32X1 U331 ( .B(framesync[1]), .C(framesync[2]), .A(framesync[0]), .Y(
        n146) );
  INVX1 U332 ( .A(n273), .Y(n63) );
  OAI211X1 U333 ( .C(i2ccon_o[1]), .D(n274), .A(clk_count1[3]), .B(n275), .Y(
        n273) );
  AOI211X1 U334 ( .C(n72), .D(n67), .A(n133), .B(n445), .Y(n274) );
  AOI31X1 U335 ( .A(n133), .B(n445), .C(n66), .D(n272), .Y(n275) );
  OA21X1 U336 ( .B(n12), .C(n8), .A(n138), .Y(n291) );
  XNOR2XL U337 ( .A(i2cdat_o[2]), .B(i2cadr_o[3]), .Y(n176) );
  NOR2X1 U338 ( .A(n97), .B(i2ccon_o[3]), .Y(n258) );
  NOR2X1 U339 ( .A(fsmsta[2]), .B(fsmsta[0]), .Y(n305) );
  XNOR2XL U340 ( .A(i2cdat_o[1]), .B(i2cadr_o[2]), .Y(n170) );
  XNOR2XL U341 ( .A(i2cdat_o[0]), .B(i2cadr_o[1]), .Y(n171) );
  XNOR2XL U342 ( .A(i2cdat_o[4]), .B(i2cadr_o[5]), .Y(n172) );
  OAI32X1 U343 ( .A(n143), .B(ack_bit), .C(n76), .D(n144), .E(n145), .Y(n142)
         );
  INVX1 U344 ( .A(n147), .Y(n76) );
  AOI211X1 U345 ( .C(framesync[3]), .D(n146), .A(bsd7), .B(n111), .Y(n144) );
  INVX1 U346 ( .A(i2ccon_o[3]), .Y(n38) );
  NOR2X1 U347 ( .A(n452), .B(sdaint), .Y(n409) );
  NAND2X1 U348 ( .A(clk_count1[3]), .B(clk_count1[2]), .Y(n133) );
  NOR3XL U349 ( .A(n104), .B(fsmmod[1]), .C(n105), .Y(n115) );
  NAND2X1 U350 ( .A(framesync[1]), .B(framesync[0]), .Y(n287) );
  NOR3XL U351 ( .A(clk_count1[1]), .B(clk_count1[2]), .C(clk_count1[0]), .Y(
        n272) );
  AOI22X1 U352 ( .A(n381), .B(n93), .C(n382), .D(sdaint), .Y(n372) );
  OAI21X1 U353 ( .B(n193), .C(n383), .A(n384), .Y(n381) );
  NOR2X1 U354 ( .A(n343), .B(n333), .Y(N1124) );
  AOI221XL U355 ( .A(n115), .B(n334), .C(n342), .D(n58), .E(n345), .Y(n343) );
  OAI21X1 U356 ( .B(n346), .C(n339), .A(n347), .Y(n345) );
  OAI21BBX1 U357 ( .A(n338), .B(sclint), .C(n154), .Y(n347) );
  AOI21AX1 U358 ( .B(nedetect), .C(n149), .A(n145), .Y(n148) );
  NAND2X1 U359 ( .A(fsmdet[2]), .B(n352), .Y(n138) );
  NOR3XL U360 ( .A(i2ccon_o[2]), .B(sdaint), .C(n13), .Y(n374) );
  NAND3X1 U361 ( .A(n398), .B(n295), .C(fsmsta[3]), .Y(n380) );
  NOR2X1 U362 ( .A(n283), .B(framesync[3]), .Y(n149) );
  NAND4X1 U363 ( .A(n450), .B(n443), .C(n449), .D(n416), .Y(n166) );
  NOR4XL U364 ( .A(i2cdat_o[6]), .B(i2cdat_o[5]), .C(i2cdat_o[4]), .D(
        i2cdat_o[3]), .Y(n416) );
  AOI31X1 U365 ( .A(scli_ff_reg0[2]), .B(N414), .C(N413), .D(n45), .Y(n186) );
  OAI211X1 U366 ( .C(n385), .D(n394), .A(n395), .B(n396), .Y(n389) );
  AO21X1 U367 ( .B(n93), .C(n13), .A(n400), .Y(n395) );
  AOI211X1 U368 ( .C(n397), .D(n398), .A(n399), .B(n162), .Y(n396) );
  NOR2X1 U369 ( .A(fsmsta[3]), .B(fsmsta[1]), .Y(n397) );
  NAND2X1 U370 ( .A(clk_count1_ov), .B(n125), .Y(n260) );
  NAND2X1 U371 ( .A(n125), .B(n270), .Y(n267) );
  OAI211X1 U372 ( .C(i2ccon_o[7]), .D(n63), .A(n271), .B(n131), .Y(n270) );
  OAI21X1 U373 ( .B(n133), .C(n67), .A(n129), .Y(n271) );
  AOI33X1 U374 ( .A(n153), .B(n38), .C(starto_en), .D(n336), .E(n296), .F(n258), .Y(n346) );
  NAND3X1 U375 ( .A(n99), .B(n138), .C(i2ccon_o[6]), .Y(n119) );
  OAI22X1 U376 ( .A(n25), .B(n71), .C(n269), .D(n267), .Y(N656) );
  XNOR2XL U377 ( .A(n132), .B(clk_count1[2]), .Y(n269) );
  NOR2X1 U378 ( .A(n88), .B(fsmdet[1]), .Y(n352) );
  NAND3X1 U379 ( .A(nedetect), .B(n97), .C(n291), .Y(n293) );
  OAI211X1 U380 ( .C(n289), .D(n290), .A(n121), .B(n291), .Y(n285) );
  AOI211X1 U381 ( .C(i2ccon_o[5]), .D(n296), .A(i2ccon_o[4]), .B(i2ccon_o[3]), 
        .Y(n289) );
  EORX1 U382 ( .A(n206), .B(n292), .C(n293), .D(n13), .Y(n290) );
  OAI211X1 U383 ( .C(fsmsta[0]), .D(n110), .A(n439), .B(n294), .Y(n292) );
  NAND4X1 U384 ( .A(fsmsta[2]), .B(n160), .C(fsmsta[1]), .D(n440), .Y(n377) );
  INVX1 U385 ( .A(sdao), .Y(n452) );
  OAI31XL U386 ( .A(n448), .B(ack), .C(n166), .D(n74), .Y(n413) );
  INVX1 U387 ( .A(n376), .Y(n74) );
  OAI21X1 U388 ( .B(n183), .C(n184), .A(n185), .Y(n498) );
  NAND42X1 U389 ( .C(n186), .D(n45), .A(nedetect), .B(n29), .Y(n185) );
  GEN2XL U390 ( .D(n82), .E(n70), .C(n231), .B(n232), .A(n233), .Y(N749) );
  OAI211X1 U391 ( .C(n441), .D(n435), .A(si), .B(n234), .Y(n232) );
  AOI211X1 U392 ( .C(n235), .D(n442), .A(sclint), .B(n236), .Y(n234) );
  OAI21X1 U393 ( .B(fsmsta[2]), .C(n159), .A(fsmsta[3]), .Y(n235) );
  OAI21X1 U394 ( .B(rst_delay), .C(n277), .A(n29), .Y(N653) );
  NOR4XL U395 ( .A(n129), .B(n130), .C(n276), .D(n444), .Y(n277) );
  AOI211X1 U396 ( .C(n79), .D(n155), .A(n156), .B(n157), .Y(n501) );
  OAI211X1 U397 ( .C(n158), .D(n38), .A(n99), .B(n29), .Y(n156) );
  NAND4X1 U398 ( .A(nedetect), .B(n149), .C(i2ccon_o[2]), .D(n163), .Y(n155)
         );
  AOI211X1 U399 ( .C(n159), .D(n160), .A(n161), .B(n162), .Y(n158) );
  NAND3X1 U400 ( .A(n99), .B(n138), .C(n278), .Y(n276) );
  AOI21X1 U401 ( .B(n279), .C(n83), .A(n280), .Y(n278) );
  AOI21X1 U402 ( .B(n81), .C(n82), .A(fsmsync[1]), .Y(n280) );
  OAI22X1 U403 ( .A(n115), .B(n65), .C(n451), .D(n123), .Y(n279) );
  AOI21X1 U404 ( .B(fsmsta[3]), .C(fsmsta[1]), .A(n442), .Y(n294) );
  NAND3X1 U405 ( .A(n104), .B(n102), .C(fsmmod[2]), .Y(n123) );
  OAI2B11X1 U406 ( .D(test_so), .C(sclint), .A(n41), .B(n24), .Y(N332) );
  INVX1 U407 ( .A(adrcomp), .Y(n79) );
  OAI211X1 U408 ( .C(n355), .D(n75), .A(n24), .B(n356), .Y(N1027) );
  NOR3XL U409 ( .A(n358), .B(n359), .C(n360), .Y(n355) );
  AOI22X1 U410 ( .A(n357), .B(ack), .C(n84), .D(n157), .Y(n356) );
  ENOX1 U411 ( .A(n361), .B(n96), .C(n93), .D(n362), .Y(n360) );
  NAND2X1 U412 ( .A(n109), .B(fsmsta[3]), .Y(n302) );
  INVX1 U413 ( .A(clk_count1[1]), .Y(n67) );
  OAI21AX1 U414 ( .B(framesync[0]), .C(n35), .A(n285), .Y(N492) );
  NAND2X1 U415 ( .A(framesync[2]), .B(n98), .Y(n283) );
  INVX1 U416 ( .A(clk_count1[0]), .Y(n72) );
  NAND4X1 U417 ( .A(n173), .B(n174), .C(n175), .D(n176), .Y(n168) );
  XNOR2XL U418 ( .A(i2cdat_o[6]), .B(i2cadr_o[7]), .Y(n173) );
  XNOR2XL U419 ( .A(i2cdat_o[5]), .B(i2cadr_o[6]), .Y(n174) );
  XNOR2XL U420 ( .A(i2cdat_o[3]), .B(i2cadr_o[4]), .Y(n175) );
  INVX1 U421 ( .A(i2ccon_o[0]), .Y(n445) );
  INVX1 U422 ( .A(adrcompen), .Y(n77) );
  NAND2X1 U423 ( .A(n134), .B(n125), .Y(n504) );
  XNOR2XL U424 ( .A(clkint), .B(clk_count2_ov), .Y(n134) );
  NOR2X1 U425 ( .A(clk_count1[0]), .B(n267), .Y(N654) );
  NOR2X1 U426 ( .A(n266), .B(n267), .Y(N657) );
  XNOR2XL U427 ( .A(clk_count1[3]), .B(n268), .Y(n266) );
  NOR21XL U428 ( .B(clk_count1[2]), .A(n66), .Y(n268) );
  NOR2X1 U429 ( .A(n264), .B(n260), .Y(N688) );
  XNOR2XL U430 ( .A(clk_count2[3]), .B(n263), .Y(n264) );
  NOR2X1 U431 ( .A(n259), .B(n260), .Y(N690) );
  AOI222XL U432 ( .A(n261), .B(n444), .C(i2ccon_o[7]), .D(n262), .E(
        clk_count2[3]), .F(n263), .Y(n259) );
  OAI21AX1 U433 ( .B(n445), .C(n54), .A(i2ccon_o[1]), .Y(n262) );
  AOI31X1 U434 ( .A(n53), .B(n46), .C(n52), .D(wait_for_setup_r), .Y(n183) );
  GEN2XL U435 ( .D(n297), .E(n56), .C(N469), .B(indelay[2]), .A(n298), .Y(N471) );
  NOR4XL U436 ( .A(indelay[2]), .B(n56), .C(n68), .D(n57), .Y(n298) );
  GEN2XL U437 ( .D(fsmsta[1]), .E(n440), .C(n295), .B(n435), .A(n36), .Y(N407)
         );
  INVX1 U438 ( .A(n300), .Y(n36) );
  AO33X1 U439 ( .A(clk_count1_ov), .B(n24), .C(rst_delay), .D(n124), .E(n43), 
        .F(n125), .Y(n505) );
  INVX1 U440 ( .A(rst_delay), .Y(n43) );
  OAI21X1 U441 ( .B(i2ccon_o[7]), .C(n126), .A(n127), .Y(n124) );
  AOI33X1 U442 ( .A(i2ccon_o[7]), .B(i2ccon_o[1]), .C(n128), .D(n129), .E(n62), 
        .F(clk_count1[1]), .Y(n127) );
  NAND21X1 U443 ( .B(clk_count1[3]), .A(n272), .Y(n131) );
  NOR3XL U444 ( .A(fsmsync[2]), .B(n25), .C(n69), .Y(n297) );
  NOR3XL U445 ( .A(n82), .B(fsmsync[1]), .C(n81), .Y(n243) );
  NOR3XL U446 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(fsmmod[0]), .Y(n153) );
  NOR21XL U447 ( .B(bclkcnt[1]), .A(n14), .Y(n130) );
  XNOR2XL U448 ( .A(bclksel), .B(bclkcnt[0]), .Y(n14) );
  NAND21X1 U449 ( .B(clk_count1_ov), .A(n125), .Y(N689) );
  NAND2X1 U450 ( .A(clkint_ff), .B(n73), .Y(n122) );
  OAI211X1 U451 ( .C(n107), .D(n344), .A(n138), .B(n446), .Y(n333) );
  NAND2X1 U452 ( .A(n95), .B(pedetect), .Y(n344) );
  NOR2X1 U453 ( .A(n73), .B(clkint_ff), .Y(n253) );
  AOI21X1 U454 ( .B(i2ccon_o[0]), .C(i2ccon_o[1]), .A(n444), .Y(n129) );
  NAND3X1 U455 ( .A(indelay[1]), .B(n57), .C(indelay[2]), .Y(n245) );
  NAND3X1 U456 ( .A(n60), .B(n447), .C(i2ccon_o[5]), .Y(n339) );
  AND3X1 U457 ( .A(n130), .B(n131), .C(i2ccon_o[0]), .Y(n128) );
  INVX1 U458 ( .A(sclint), .Y(n83) );
  INVX1 U459 ( .A(fsmsync[0]), .Y(n82) );
  INVX1 U460 ( .A(fsmsync[1]), .Y(n70) );
  INVX1 U461 ( .A(sdaint), .Y(n92) );
  NOR4XL U462 ( .A(n61), .B(n70), .C(fsmsync[0]), .D(fsmsync[2]), .Y(n242) );
  INVX1 U463 ( .A(pedetect), .Y(n78) );
  INVX1 U464 ( .A(ack), .Y(n94) );
  OAI221X1 U465 ( .A(fsmsta[1]), .B(n113), .C(fsmsta[0]), .D(n308), .E(n300), 
        .Y(N406) );
  INVX1 U466 ( .A(fsmsync[2]), .Y(n81) );
  OAI21X1 U467 ( .B(n35), .C(n288), .A(n121), .Y(N493) );
  OAI21X1 U468 ( .B(framesync[1]), .C(framesync[0]), .A(n287), .Y(n288) );
  OAI21X1 U469 ( .B(n286), .C(n35), .A(n121), .Y(N494) );
  XNOR2XL U470 ( .A(n98), .B(framesync[2]), .Y(n286) );
  OAI211X1 U471 ( .C(n9), .D(n303), .A(n300), .B(n304), .Y(N409) );
  AOI32X1 U472 ( .A(n9), .B(n7), .C(n305), .D(n306), .E(n303), .Y(n304) );
  AOI211X1 U473 ( .C(n47), .D(n122), .A(n230), .B(n115), .Y(n490) );
  INVX1 U474 ( .A(starto_en), .Y(n47) );
  OR2X1 U475 ( .A(n184), .B(n65), .Y(n230) );
  INVX1 U476 ( .A(clkint), .Y(n73) );
  AOI21X1 U477 ( .B(sclint), .C(n60), .A(n123), .Y(n335) );
  NOR3XL U478 ( .A(n103), .B(sdaint), .C(i2ccon_o[3]), .Y(n337) );
  INVX1 U479 ( .A(i2ccon_o[4]), .Y(n447) );
  AOI21X1 U480 ( .B(n254), .C(n255), .A(n238), .Y(N746) );
  AOI211X1 U481 ( .C(n244), .D(n92), .A(n256), .B(n257), .Y(n255) );
  AOI222XL U482 ( .A(n243), .B(si), .C(n240), .D(n447), .E(n242), .F(n39), .Y(
        n254) );
  NOR4XL U483 ( .A(sclint), .B(fsmsync[2]), .C(fsmsync[1]), .D(fsmsync[0]), 
        .Y(n256) );
  AOI21X1 U484 ( .B(n190), .C(n191), .A(n192), .Y(n496) );
  OAI211X1 U485 ( .C(n58), .D(n193), .A(n121), .B(adrcompen), .Y(n191) );
  NAND2X1 U486 ( .A(n194), .B(n28), .Y(n190) );
  AOI21X1 U487 ( .B(n353), .C(n354), .A(n184), .Y(N1063) );
  NAND2X1 U488 ( .A(n351), .B(n92), .Y(n354) );
  AOI32X1 U489 ( .A(n89), .B(n88), .C(sdaint), .D(n352), .E(n91), .Y(n353) );
  INVX1 U490 ( .A(n351), .Y(n89) );
  NAND3X1 U491 ( .A(n24), .B(n83), .C(test_so), .Y(n312) );
  OAI21X1 U492 ( .B(n116), .C(n92), .A(n117), .Y(n507) );
  NOR3XL U493 ( .A(sdai_ff_reg0[0]), .B(sdai_ff_reg0[2]), .C(sdai_ff_reg0[1]), 
        .Y(n116) );
  AOI31X1 U494 ( .A(sdai_ff_reg0[1]), .B(sdai_ff_reg0[0]), .C(sdai_ff_reg0[2]), 
        .D(n27), .Y(n117) );
  AOI31X1 U495 ( .A(n246), .B(n247), .C(n248), .D(n238), .Y(N747) );
  OAI211X1 U496 ( .C(n38), .D(n61), .A(n82), .B(fsmsync[1]), .Y(n247) );
  AOI22X1 U497 ( .A(n243), .B(n38), .C(n231), .D(n245), .Y(n248) );
  AOI31X1 U498 ( .A(n70), .B(n81), .C(n249), .D(n244), .Y(n246) );
  AOI31X1 U499 ( .A(n330), .B(n331), .C(n332), .D(n333), .Y(N1126) );
  NAND3X1 U500 ( .A(n336), .B(i2ccon_o[4]), .C(n258), .Y(n331) );
  AOI221XL U501 ( .A(n251), .B(n58), .C(n115), .D(n334), .E(n335), .Y(n332) );
  AOI33X1 U502 ( .A(starto_en), .B(n59), .C(n337), .D(sclint), .E(n338), .F(
        n154), .Y(n330) );
  AOI31X1 U503 ( .A(n100), .B(n101), .C(n340), .D(n333), .Y(N1125) );
  AOI22X1 U504 ( .A(n336), .B(n341), .C(n342), .D(nedetect), .Y(n340) );
  NAND2X1 U505 ( .A(n258), .B(i2ccon_o[4]), .Y(n341) );
  INVX1 U506 ( .A(indelay[0]), .Y(n57) );
  INVX1 U507 ( .A(i2ccon_o[7]), .Y(n444) );
  INVX1 U508 ( .A(scli_ff_reg0[0]), .Y(n53) );
  INVX1 U509 ( .A(scli_ff_reg0[1]), .Y(n52) );
  INVX1 U510 ( .A(clk_count2[0]), .Y(n54) );
  OAI21BBX1 U511 ( .A(n54), .B(n125), .C(n265), .Y(N685) );
  NAND4X1 U512 ( .A(fsmsync[2]), .B(n82), .C(n70), .D(n29), .Y(n265) );
  NOR2X1 U513 ( .A(setup_counter_r[1]), .B(setup_counter_r[0]), .Y(n313) );
  NOR2X1 U514 ( .A(n68), .B(indelay[0]), .Y(N469) );
  INVX1 U515 ( .A(i2cdat_o[0]), .Y(n449) );
  NAND2X1 U516 ( .A(n23), .B(n189), .Y(n182) );
  NAND4X1 U517 ( .A(scli_ff_reg0[2]), .B(scli_ff_reg0[1]), .C(scli_ff_reg0[0]), 
        .D(n183), .Y(n189) );
  INVX1 U518 ( .A(i2cdat_o[2]), .Y(n443) );
  INVX1 U519 ( .A(i2cdat_o[1]), .Y(n450) );
  NAND2X1 U520 ( .A(n82), .B(n250), .Y(n249) );
  OAI211X1 U521 ( .C(n251), .D(n252), .A(sclint), .B(n253), .Y(n250) );
  AOI22X1 U522 ( .A(fsmmod[2]), .B(n104), .C(fsmmod[1]), .D(fsmmod[0]), .Y(
        n252) );
  INVX1 U523 ( .A(scli_ff_reg0[2]), .Y(n46) );
  NOR2X1 U524 ( .A(i2ccon_o[2]), .B(sdaint), .Y(n417) );
  NAND2X1 U525 ( .A(n300), .B(n307), .Y(N408) );
  OAI211X1 U526 ( .C(fsmsta[2]), .D(n159), .A(n435), .B(n303), .Y(n307) );
  NOR2X1 U527 ( .A(n348), .B(n184), .Y(N1065) );
  AOI221XL U528 ( .A(fsmdet[1]), .B(sdaint), .C(fsmdet[2]), .D(n90), .E(n194), 
        .Y(n348) );
  NOR2X1 U529 ( .A(n349), .B(n184), .Y(N1064) );
  AOI221XL U530 ( .A(fsmdet[2]), .B(fsmdet[0]), .C(n350), .D(n92), .E(n351), 
        .Y(n349) );
  OAI21AX1 U531 ( .B(fsmdet[2]), .C(fsmdet[0]), .A(n352), .Y(n350) );
  NOR2X1 U532 ( .A(n237), .B(n238), .Y(N748) );
  AOI221XL U533 ( .A(n239), .B(n83), .C(i2ccon_o[3]), .D(n240), .E(n241), .Y(
        n237) );
  OAI22X1 U534 ( .A(fsmsync[0]), .B(n81), .C(n245), .D(n69), .Y(n239) );
  GEN2XL U535 ( .D(n206), .E(n242), .C(n243), .B(i2ccon_o[4]), .A(n244), .Y(
        n241) );
  INVX1 U539 ( .A(busfree), .Y(n65) );
  INVX1 U540 ( .A(i2cadr_o[0]), .Y(n448) );
  INVX1 U541 ( .A(n114), .Y(n48) );
  OAI211X1 U542 ( .C(sclscl), .D(pedetect), .A(n115), .B(n29), .Y(n114) );
  INVX1 U543 ( .A(bsd7_tmp), .Y(n64) );
  NAND21X1 U544 ( .B(scli_ff), .A(n28), .Y(N412) );
  NAND21X1 U545 ( .B(sdai_ff), .A(n28), .Y(N431) );
  NAND21X1 U546 ( .B(sdai_ff_reg0[0]), .A(n28), .Y(N432) );
  NAND21X1 U547 ( .B(sdai_ff_reg0[1]), .A(n28), .Y(N433) );
  NOR3XL U548 ( .A(n281), .B(n27), .C(n130), .Y(N511) );
  XNOR2XL U549 ( .A(bclkcnt[1]), .B(bclkcnt[0]), .Y(n281) );
  INVX1 U550 ( .A(nedetect), .Y(n58) );
  NOR3XL U551 ( .A(n130), .B(n27), .C(bclkcnt[0]), .Y(N510) );
  INVX1 U552 ( .A(fsmdet[2]), .Y(n91) );
  NAND2X1 U553 ( .A(sclscl), .B(pedetect), .Y(n334) );
  INVX1 U554 ( .A(clk_count2[1]), .Y(n51) );
  INVX1 U555 ( .A(clk_count2[2]), .Y(n55) );
  INVX1 U556 ( .A(setup_counter_r[2]), .Y(n42) );
  INVX1 U557 ( .A(indelay[1]), .Y(n56) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module extint_a0 ( clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, 
        int2ff, iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, 
        int6ff, iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, 
        ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7, 
        iex8, iex9, iex10, iex11, iex12, sfraddr, sfrdatai, sfrwe, test_si, 
        test_se );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, int2ff,
         iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, int6ff,
         iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, sfrwe,
         test_si, test_se;
  output ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12;
  wire   int0_ff1, int0_fall, int0_clr, N23, int1_ff1, int1_fall, int1_clr,
         N51, int2_ff1, iex2_set, N71, int3_ff1, iex3_set, N90, iex4_set,
         int4_ff1, iex5_set, int5_ff1, iex6_set, int6_ff1, iex7_set, int7_ff1,
         iex8_set, int8_ff1, iex9_set, int9_ff1, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n77, n78, n79, n80,
         n81, n82, n83, n84;

  SDFFQX1 int4_ff1_reg ( .D(n19), .SIN(int3_ff1), .SMC(test_se), .C(clkper), 
        .Q(int4_ff1) );
  SDFFQX1 int5_ff1_reg ( .D(n13), .SIN(int4_ff1), .SMC(test_se), .C(clkper), 
        .Q(int5_ff1) );
  SDFFQX1 int6_ff1_reg ( .D(n11), .SIN(int5_ff1), .SMC(test_se), .C(clkper), 
        .Q(int6_ff1) );
  SDFFQX1 int7_ff1_reg ( .D(n12), .SIN(int6_ff1), .SMC(test_se), .C(clkper), 
        .Q(int7_ff1) );
  SDFFQX1 int8_ff1_reg ( .D(n84), .SIN(int7_ff1), .SMC(test_se), .C(clkper), 
        .Q(int8_ff1) );
  SDFFQX1 int9_ff1_reg ( .D(n10), .SIN(int8_ff1), .SMC(test_se), .C(clkper), 
        .Q(int9_ff1) );
  SDFFQX1 iex4_set_reg ( .D(n105), .SIN(iex4), .SMC(test_se), .C(clkper), .Q(
        iex4_set) );
  SDFFQX1 iex5_set_reg ( .D(n103), .SIN(iex5), .SMC(test_se), .C(clkper), .Q(
        iex5_set) );
  SDFFQX1 iex6_set_reg ( .D(n101), .SIN(iex6), .SMC(test_se), .C(clkper), .Q(
        iex6_set) );
  SDFFQX1 iex7_set_reg ( .D(n99), .SIN(iex7), .SMC(test_se), .C(clkper), .Q(
        iex7_set) );
  SDFFQX1 iex8_set_reg ( .D(n97), .SIN(iex8), .SMC(test_se), .C(clkper), .Q(
        iex8_set) );
  SDFFQX1 iex9_set_reg ( .D(n95), .SIN(iex9), .SMC(test_se), .C(clkper), .Q(
        iex9_set) );
  SDFFQX1 int0_ff1_reg ( .D(N23), .SIN(int0_fall), .SMC(test_se), .C(clkper), 
        .Q(int0_ff1) );
  SDFFQX1 iex2_set_reg ( .D(n110), .SIN(iex2), .SMC(test_se), .C(clkper), .Q(
        iex2_set) );
  SDFFQX1 iex3_set_reg ( .D(n107), .SIN(iex3), .SMC(test_se), .C(clkper), .Q(
        iex3_set) );
  SDFFQX1 int0_clr_reg ( .D(n118), .SIN(iex9_set), .SMC(test_se), .C(clkper), 
        .Q(int0_clr) );
  SDFFQX1 int1_clr_reg ( .D(n114), .SIN(int0_ff1), .SMC(test_se), .C(clkper), 
        .Q(int1_clr) );
  SDFFQX1 int2_ff1_reg ( .D(N71), .SIN(int1_ff1), .SMC(test_se), .C(clkper), 
        .Q(int2_ff1) );
  SDFFQX1 int3_ff1_reg ( .D(N90), .SIN(int2_ff1), .SMC(test_se), .C(clkper), 
        .Q(int3_ff1) );
  SDFFQX1 int1_ff1_reg ( .D(N51), .SIN(int1_fall), .SMC(test_se), .C(clkper), 
        .Q(int1_ff1) );
  SDFFQX1 int0_fall_reg ( .D(n116), .SIN(int0_clr), .SMC(test_se), .C(clkper), 
        .Q(int0_fall) );
  SDFFQX1 int1_fall_reg ( .D(n112), .SIN(int1_clr), .SMC(test_se), .C(clkper), 
        .Q(int1_fall) );
  SDFFQX1 iex9_s_reg ( .D(n94), .SIN(iex8_set), .SMC(test_se), .C(clkper), .Q(
        iex9) );
  SDFFQX1 iex8_s_reg ( .D(n96), .SIN(iex7_set), .SMC(test_se), .C(clkper), .Q(
        iex8) );
  SDFFQX1 it0_s_reg ( .D(n117), .SIN(int9_ff1), .SMC(test_se), .C(clkper), .Q(
        it0) );
  SDFFQX1 iex4_s_reg ( .D(n104), .SIN(iex3_set), .SMC(test_se), .C(clkper), 
        .Q(iex4) );
  SDFFQX1 iex6_s_reg ( .D(n100), .SIN(iex5_set), .SMC(test_se), .C(clkper), 
        .Q(iex6) );
  SDFFQX1 i3fr_s_reg ( .D(n108), .SIN(i2fr), .SMC(test_se), .C(clkper), .Q(
        i3fr) );
  SDFFQX1 ie1_s_reg ( .D(n111), .SIN(ie0), .SMC(test_se), .C(clkper), .Q(ie1)
         );
  SDFFQX1 i2fr_s_reg ( .D(n14), .SIN(test_si), .SMC(test_se), .C(clkper), .Q(
        i2fr) );
  SDFFQX1 ie0_s_reg ( .D(n115), .SIN(i3fr), .SMC(test_se), .C(clkper), .Q(ie0)
         );
  SDFFQX1 iex2_s_reg ( .D(n109), .SIN(ie1), .SMC(test_se), .C(clkper), .Q(iex2) );
  SDFFQX1 iex7_s_reg ( .D(n98), .SIN(iex6_set), .SMC(test_se), .C(clkper), .Q(
        iex7) );
  SDFFQX1 iex5_s_reg ( .D(n102), .SIN(iex4_set), .SMC(test_se), .C(clkper), 
        .Q(iex5) );
  SDFFQX1 it1_s_reg ( .D(n113), .SIN(it0), .SMC(test_se), .C(clkper), .Q(it1)
         );
  SDFFQX1 iex3_s_reg ( .D(n106), .SIN(iex2_set), .SMC(test_se), .C(clkper), 
        .Q(iex3) );
  INVX1 U3 ( .A(1'b1), .Y(iex12) );
  INVX1 U5 ( .A(1'b1), .Y(iex11) );
  INVX1 U7 ( .A(1'b1), .Y(iex10) );
  INVX1 U9 ( .A(n34), .Y(n15) );
  INVX1 U10 ( .A(n52), .Y(n16) );
  NAND2X1 U11 ( .A(n75), .B(n9), .Y(n41) );
  NOR2X1 U12 ( .A(n75), .B(n7), .Y(n43) );
  INVX1 U13 ( .A(n46), .Y(n17) );
  INVX1 U14 ( .A(n8), .Y(n7) );
  AOI21X1 U15 ( .B(n68), .C(sfraddr[3]), .A(rst), .Y(n34) );
  AND2X1 U16 ( .A(sfraddr[6]), .B(n63), .Y(n68) );
  NOR42XL U17 ( .C(sfrwe), .D(n76), .A(sfraddr[0]), .B(sfraddr[1]), .Y(n63) );
  NOR3XL U18 ( .A(sfraddr[2]), .B(sfraddr[5]), .C(sfraddr[4]), .Y(n76) );
  NOR32XL U19 ( .B(n63), .C(sfraddr[3]), .A(sfraddr[6]), .Y(n52) );
  NAND21X1 U20 ( .B(sfraddr[3]), .A(n68), .Y(n75) );
  NAND2X1 U21 ( .A(n49), .B(n50), .Y(n46) );
  NOR43XL U22 ( .B(sfraddr[3]), .C(sfrwe), .D(sfraddr[0]), .A(sfraddr[6]), .Y(
        n50) );
  INVX1 U23 ( .A(n53), .Y(n18) );
  INVX1 U24 ( .A(n35), .Y(n12) );
  INVX1 U25 ( .A(rst), .Y(n8) );
  INVX1 U26 ( .A(rst), .Y(n9) );
  INVX1 U27 ( .A(n40), .Y(n84) );
  INVX1 U28 ( .A(n39), .Y(n13) );
  INVX1 U29 ( .A(n36), .Y(n10) );
  INVX1 U30 ( .A(n38), .Y(n19) );
  NOR2X1 U31 ( .A(n7), .B(newinstr), .Y(n53) );
  OAI22X1 U32 ( .A(n7), .B(n77), .C(n18), .D(n29), .Y(n114) );
  OAI22X1 U33 ( .A(rst), .B(n32), .C(n18), .D(n28), .Y(n118) );
  NAND2X1 U34 ( .A(int7ff), .B(n9), .Y(n35) );
  OR2X1 U35 ( .A(int2ff), .B(rst), .Y(N71) );
  INVX1 U36 ( .A(int0ack), .Y(n32) );
  OR2X1 U37 ( .A(int3ff), .B(rst), .Y(N90) );
  INVX1 U38 ( .A(int1ack), .Y(n77) );
  INVX1 U39 ( .A(iex3ack), .Y(n79) );
  INVX1 U40 ( .A(iex2ack), .Y(n78) );
  INVX1 U41 ( .A(n37), .Y(n11) );
  NAND2X1 U42 ( .A(int8ff), .B(n9), .Y(n40) );
  NOR2X1 U43 ( .A(n7), .B(n83), .Y(N23) );
  NOR2X1 U44 ( .A(n7), .B(n82), .Y(N51) );
  NAND2X1 U45 ( .A(int5ff), .B(n9), .Y(n39) );
  OAI32X1 U46 ( .A(n21), .B(iex5ack), .C(n18), .D(int5_ff1), .E(n39), .Y(n103)
         );
  INVX1 U47 ( .A(iex5_set), .Y(n21) );
  NAND2X1 U48 ( .A(int9ff), .B(n8), .Y(n36) );
  NAND2X1 U49 ( .A(int4ff), .B(n8), .Y(n38) );
  OAI32X1 U50 ( .A(n25), .B(iex9ack), .C(n18), .D(int9_ff1), .E(n36), .Y(n95)
         );
  INVX1 U51 ( .A(iex9_set), .Y(n25) );
  OAI32X1 U52 ( .A(n20), .B(iex4ack), .C(n18), .D(int4_ff1), .E(n38), .Y(n105)
         );
  INVX1 U53 ( .A(iex4_set), .Y(n20) );
  OAI21BBX1 U54 ( .A(n34), .B(i3fr), .C(n67), .Y(n108) );
  NAND3X1 U55 ( .A(n15), .B(n9), .C(sfrdatai[6]), .Y(n67) );
  INVX1 U56 ( .A(n33), .Y(n14) );
  AOI32X1 U57 ( .A(sfrdatai[5]), .B(n9), .C(n15), .D(n34), .E(i2fr), .Y(n33)
         );
  NOR2X1 U58 ( .A(n7), .B(n58), .Y(n113) );
  AOI22X1 U59 ( .A(sfrdatai[2]), .B(n52), .C(it1), .D(n16), .Y(n58) );
  NOR2X1 U60 ( .A(n7), .B(n51), .Y(n117) );
  AOI22X1 U61 ( .A(n52), .B(sfrdatai[0]), .C(it0), .D(n16), .Y(n51) );
  NOR2X1 U62 ( .A(n7), .B(n59), .Y(n111) );
  EORX1 U63 ( .A(sfrdatai[3]), .B(n52), .C(n60), .D(n52), .Y(n59) );
  AOI32X1 U64 ( .A(n29), .B(n77), .C(n61), .D(n82), .E(n31), .Y(n60) );
  ENOX1 U65 ( .A(n62), .B(n31), .C(n82), .D(int1_ff1), .Y(n61) );
  AND2X1 U66 ( .A(n54), .B(n9), .Y(n115) );
  ENOX1 U67 ( .A(n52), .B(n55), .C(sfrdatai[1]), .D(n52), .Y(n54) );
  AOI32X1 U68 ( .A(n28), .B(n32), .C(n56), .D(n83), .E(n30), .Y(n55) );
  ENOX1 U69 ( .A(n57), .B(n30), .C(n83), .D(int0_ff1), .Y(n56) );
  AOI21X1 U70 ( .B(n47), .C(n48), .A(rst), .Y(n94) );
  NAND2X1 U71 ( .A(sfrdatai[1]), .B(n17), .Y(n47) );
  OAI211X1 U72 ( .C(iex9), .D(iex9_set), .A(n46), .B(n80), .Y(n48) );
  INVX1 U73 ( .A(iex9ack), .Y(n80) );
  AOI21X1 U74 ( .B(n44), .C(n45), .A(rst), .Y(n96) );
  NAND2X1 U75 ( .A(n17), .B(sfrdatai[0]), .Y(n44) );
  OAI211X1 U76 ( .C(iex8), .D(iex8_set), .A(n46), .B(n81), .Y(n45) );
  INVX1 U77 ( .A(iex8ack), .Y(n81) );
  ENOX1 U78 ( .A(n41), .B(n42), .C(n43), .D(sfrdatai[0]), .Y(n98) );
  OAI21AX1 U79 ( .B(iex7), .C(iex7_set), .A(iex7ack), .Y(n42) );
  ENOX1 U80 ( .A(n41), .B(n72), .C(n43), .D(sfrdatai[3]), .Y(n104) );
  OAI21AX1 U81 ( .B(iex4), .C(iex4_set), .A(iex4ack), .Y(n72) );
  ENOX1 U82 ( .A(n41), .B(n74), .C(sfrdatai[5]), .D(n43), .Y(n100) );
  OAI21AX1 U83 ( .B(iex6), .C(iex6_set), .A(iex6ack), .Y(n74) );
  ENOX1 U84 ( .A(n41), .B(n73), .C(sfrdatai[4]), .D(n43), .Y(n102) );
  OAI21AX1 U85 ( .B(iex5), .C(iex5_set), .A(iex5ack), .Y(n73) );
  ENOX1 U86 ( .A(n41), .B(n71), .C(n43), .D(sfrdatai[2]), .Y(n106) );
  OAI21X1 U87 ( .B(iex3), .C(iex3_set), .A(n79), .Y(n71) );
  ENOX1 U88 ( .A(n41), .B(n66), .C(n43), .D(sfrdatai[1]), .Y(n109) );
  OAI21X1 U89 ( .B(iex2), .C(iex2_set), .A(n78), .Y(n66) );
  AO33X1 U90 ( .A(int1_ff1), .B(n9), .C(n82), .D(int1_fall), .E(n77), .F(n53), 
        .Y(n112) );
  AO33X1 U91 ( .A(int0_ff1), .B(n9), .C(n83), .D(int0_fall), .E(n32), .F(n53), 
        .Y(n116) );
  OAI32X1 U92 ( .A(n24), .B(iex8ack), .C(n18), .D(int8_ff1), .E(n40), .Y(n97)
         );
  INVX1 U93 ( .A(iex8_set), .Y(n24) );
  OAI32X1 U94 ( .A(n23), .B(iex7ack), .C(n18), .D(int7_ff1), .E(n35), .Y(n99)
         );
  INVX1 U95 ( .A(iex7_set), .Y(n23) );
  OAI32X1 U96 ( .A(n22), .B(iex6ack), .C(n18), .D(int6_ff1), .E(n37), .Y(n101)
         );
  INVX1 U97 ( .A(iex6_set), .Y(n22) );
  OAI31XL U98 ( .A(n27), .B(i3fr), .C(N90), .D(n69), .Y(n107) );
  INVX1 U99 ( .A(int3_ff1), .Y(n27) );
  AOI33X1 U100 ( .A(int3ff), .B(i3fr), .C(n70), .D(n53), .E(n79), .F(iex3_set), 
        .Y(n69) );
  NOR2X1 U101 ( .A(n7), .B(int3_ff1), .Y(n70) );
  OAI31XL U102 ( .A(n26), .B(i2fr), .C(N71), .D(n64), .Y(n110) );
  INVX1 U103 ( .A(int2_ff1), .Y(n26) );
  AOI33X1 U104 ( .A(int2ff), .B(i2fr), .C(n65), .D(n53), .E(n78), .F(iex2_set), 
        .Y(n64) );
  NOR2X1 U105 ( .A(n7), .B(int2_ff1), .Y(n65) );
  NAND2X1 U106 ( .A(int6ff), .B(n9), .Y(n37) );
  INVX1 U107 ( .A(int1ff), .Y(n82) );
  INVX1 U111 ( .A(int0ff), .Y(n83) );
  NOR2X1 U112 ( .A(ie1), .B(int1_fall), .Y(n62) );
  NOR2X1 U113 ( .A(ie0), .B(int0_fall), .Y(n57) );
  INVX1 U114 ( .A(it1), .Y(n31) );
  INVX1 U115 ( .A(it0), .Y(n30) );
  INVX1 U116 ( .A(int1_clr), .Y(n29) );
  INVX1 U117 ( .A(int0_clr), .Y(n28) );
  AND4XL U118 ( .A(sfraddr[1]), .B(sfraddr[2]), .C(sfraddr[4]), .D(sfraddr[5]), 
        .Y(n49) );
endmodule


module isr_a0 ( clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, 
        t0ff, int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff, 
        int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b, 
        int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, int_vect_ab, irq, intvect, int_ack_03, int_ack_0b, 
        int_ack_13, int_ack_1b, int_ack_43, int_ack_4b, int_ack_53, int_ack_5b, 
        int_ack_63, int_ack_6b, int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, 
        int_ack_ab, is_reg, ip0, ip1, ien0, ien1, ien2, isr_tm, sfraddr, 
        sfrdatai, sfrwe, test_si, test_se );
  output [4:0] intvect;
  output [3:0] is_reg;
  output [5:0] ip0;
  output [5:0] ip1;
  output [7:0] ien0;
  output [5:0] ien1;
  output [5:0] ien2;
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, t0ff,
         int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff,
         int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b,
         int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b,
         int_vect_a3, int_vect_ab, sfrwe, test_si, test_se;
  output irq, int_ack_03, int_ack_0b, int_ack_13, int_ack_1b, int_ack_43,
         int_ack_4b, int_ack_53, int_ack_5b, int_ack_63, int_ack_6b,
         int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, int_ack_ab, isr_tm;
  wire   N38, N39, N40, N41, N42, N43, N44, N45, N49, N50, N51, N52, N53, N54,
         N55, N58, N59, N60, N61, N62, N63, N64, N67, N68, N69, N70, N71, N72,
         N73, N76, N77, N78, N79, N80, N81, N82, irq_r, N200, N207, N208, N209,
         N210, N211, N212, net12095, net12101, net12106, net12111, net12116,
         net12121, n196, n197, n198, n199, n200, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n201, n202, n203, n204, n205, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n206, n207;

  SNPS_CLOCK_GATE_HIGH_isr_a0_0 clk_gate_ien0_reg_reg ( .CLK(clkper), .EN(N38), 
        .ENCLK(net12095), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_5 clk_gate_ien1_reg_reg ( .CLK(clkper), .EN(N49), 
        .ENCLK(net12101), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_4 clk_gate_ien2_reg_reg ( .CLK(clkper), .EN(N58), 
        .ENCLK(net12106), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_3 clk_gate_ip0_reg_reg ( .CLK(clkper), .EN(N67), 
        .ENCLK(net12111), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_2 clk_gate_ip1_reg_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12116), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_1 clk_gate_intvect_reg_reg ( .CLK(clkper), .EN(
        N207), .ENCLK(net12121), .TE(test_se) );
  SDFFQX1 intvect_reg_reg_0_ ( .D(N208), .SIN(ien2[5]), .SMC(test_se), .C(
        net12121), .Q(intvect[0]) );
  SDFFQX1 intvect_reg_reg_1_ ( .D(N209), .SIN(intvect[0]), .SMC(test_se), .C(
        net12121), .Q(intvect[1]) );
  SDFFQX1 intvect_reg_reg_4_ ( .D(N212), .SIN(intvect[3]), .SMC(test_se), .C(
        net12121), .Q(intvect[4]) );
  SDFFQX1 intvect_reg_reg_3_ ( .D(N211), .SIN(intvect[2]), .SMC(test_se), .C(
        net12121), .Q(intvect[3]) );
  SDFFQX1 intvect_reg_reg_2_ ( .D(N210), .SIN(intvect[1]), .SMC(test_se), .C(
        net12121), .Q(intvect[2]) );
  SDFFQX1 is_reg_s_reg_0_ ( .D(n199), .SIN(irq_r), .SMC(test_se), .C(clkper), 
        .Q(is_reg[0]) );
  SDFFQX1 is_reg_s_reg_1_ ( .D(n196), .SIN(is_reg[0]), .SMC(test_se), .C(
        clkper), .Q(is_reg[1]) );
  SDFFQX1 is_reg_s_reg_2_ ( .D(n197), .SIN(is_reg[1]), .SMC(test_se), .C(
        clkper), .Q(is_reg[2]) );
  SDFFQX1 is_reg_s_reg_3_ ( .D(n198), .SIN(is_reg[2]), .SMC(test_se), .C(
        clkper), .Q(is_reg[3]) );
  SDFFQX1 ien2_reg_reg_5_ ( .D(N64), .SIN(ien2[4]), .SMC(test_se), .C(net12106), .Q(ien2[5]) );
  SDFFQX1 ien2_reg_reg_4_ ( .D(N63), .SIN(ien2[3]), .SMC(test_se), .C(net12106), .Q(ien2[4]) );
  SDFFQX1 ip0_reg_reg_3_ ( .D(N71), .SIN(ip0[2]), .SMC(test_se), .C(net12111), 
        .Q(ip0[3]) );
  SDFFQX1 ip0_reg_reg_1_ ( .D(N69), .SIN(ip0[0]), .SMC(test_se), .C(net12111), 
        .Q(ip0[1]) );
  SDFFQX1 ien2_reg_reg_0_ ( .D(N59), .SIN(ien1[5]), .SMC(test_se), .C(net12106), .Q(ien2[0]) );
  SDFFQX1 ien1_reg_reg_0_ ( .D(N50), .SIN(ien0[7]), .SMC(test_se), .C(net12101), .Q(ien1[0]) );
  SDFFQX1 ien1_reg_reg_3_ ( .D(N53), .SIN(ien1[2]), .SMC(test_se), .C(net12101), .Q(ien1[3]) );
  SDFFQX1 ien0_reg_reg_3_ ( .D(N42), .SIN(ien0[2]), .SMC(test_se), .C(net12095), .Q(ien0[3]) );
  SDFFQX1 ien1_reg_reg_5_ ( .D(N55), .SIN(ien1[4]), .SMC(test_se), .C(net12101), .Q(ien1[5]) );
  SDFFQX1 ien1_reg_reg_1_ ( .D(N51), .SIN(ien1[0]), .SMC(test_se), .C(net12101), .Q(ien1[1]) );
  SDFFQX1 ien1_reg_reg_4_ ( .D(N54), .SIN(ien1[3]), .SMC(test_se), .C(net12101), .Q(ien1[4]) );
  SDFFQX1 ien0_reg_reg_0_ ( .D(N39), .SIN(test_si), .SMC(test_se), .C(net12095), .Q(ien0[0]) );
  SDFFQX1 ip1_reg_reg_5_ ( .D(N82), .SIN(ip1[4]), .SMC(test_se), .C(net12116), 
        .Q(ip1[5]) );
  SDFFQX1 ip0_reg_reg_0_ ( .D(N68), .SIN(intvect[4]), .SMC(test_se), .C(
        net12111), .Q(ip0[0]) );
  SDFFQX1 ip1_reg_reg_4_ ( .D(N81), .SIN(ip1[3]), .SMC(test_se), .C(net12116), 
        .Q(ip1[4]) );
  SDFFQX1 ip1_reg_reg_0_ ( .D(N77), .SIN(ip0[5]), .SMC(test_se), .C(net12116), 
        .Q(ip1[0]) );
  SDFFQX1 ip1_reg_reg_3_ ( .D(N80), .SIN(ip1[2]), .SMC(test_se), .C(net12116), 
        .Q(ip1[3]) );
  SDFFQX1 isr_tm_reg_reg ( .D(n200), .SIN(is_reg[3]), .SMC(test_se), .C(clkper), .Q(isr_tm) );
  SDFFQX1 ip0_reg_reg_2_ ( .D(N70), .SIN(ip0[1]), .SMC(test_se), .C(net12111), 
        .Q(ip0[2]) );
  SDFFQX1 ip1_reg_reg_1_ ( .D(N78), .SIN(ip1[0]), .SMC(test_se), .C(net12116), 
        .Q(ip1[1]) );
  SDFFQX1 ien1_reg_reg_2_ ( .D(N52), .SIN(ien1[1]), .SMC(test_se), .C(net12101), .Q(ien1[2]) );
  SDFFQX1 ien0_reg_reg_1_ ( .D(N40), .SIN(ien0[0]), .SMC(test_se), .C(net12095), .Q(ien0[1]) );
  SDFFQX1 ien0_reg_reg_4_ ( .D(N43), .SIN(ien0[3]), .SMC(test_se), .C(net12095), .Q(ien0[4]) );
  SDFFQX1 ien0_reg_reg_5_ ( .D(N44), .SIN(ien0[4]), .SMC(test_se), .C(net12095), .Q(ien0[5]) );
  SDFFQX1 ien2_reg_reg_2_ ( .D(N61), .SIN(ien2[1]), .SMC(test_se), .C(net12106), .Q(ien2[2]) );
  SDFFQX1 ien2_reg_reg_3_ ( .D(N62), .SIN(ien2[2]), .SMC(test_se), .C(net12106), .Q(ien2[3]) );
  SDFFQX1 ien0_reg_reg_2_ ( .D(N41), .SIN(ien0[1]), .SMC(test_se), .C(net12095), .Q(ien0[2]) );
  SDFFQX1 ien2_reg_reg_1_ ( .D(N60), .SIN(ien2[0]), .SMC(test_se), .C(net12106), .Q(ien2[1]) );
  SDFFQX1 ip1_reg_reg_2_ ( .D(N79), .SIN(ip1[1]), .SMC(test_se), .C(net12116), 
        .Q(ip1[2]) );
  SDFFQX1 ip0_reg_reg_4_ ( .D(N72), .SIN(ip0[3]), .SMC(test_se), .C(net12111), 
        .Q(ip0[4]) );
  SDFFQX1 ip0_reg_reg_5_ ( .D(N73), .SIN(ip0[4]), .SMC(test_se), .C(net12111), 
        .Q(ip0[5]) );
  SDFFQX1 irq_r_reg ( .D(N200), .SIN(ip1[5]), .SMC(test_se), .C(clkper), .Q(
        irq_r) );
  SDFFQX1 ien0_reg_reg_6_ ( .D(N45), .SIN(ien0[5]), .SMC(test_se), .C(net12095), .Q(ien0[7]) );
  INVX1 U3 ( .A(1'b1), .Y(ien0[6]) );
  NAND4XL U5 ( .A(sfraddr[2]), .B(sfraddr[0]), .C(n59), .D(n60), .Y(n58) );
  AOI221XL U6 ( .A(n204), .B(ien0[4]), .C(ien1[4]), .D(int_vect_63), .E(n48), 
        .Y(n172) );
  OAI222XL U7 ( .A(n24), .B(n176), .C(n177), .D(n47), .E(n46), .F(n178), .Y(
        n128) );
  OAI222XL U8 ( .A(n23), .B(n30), .C(n185), .D(n57), .E(n56), .F(n175), .Y(
        n130) );
  INVX1 U9 ( .A(sfraddr[0]), .Y(n3) );
  NAND3X1 U10 ( .A(n3), .B(n4), .C(n91), .Y(n97) );
  NAND3X1 U11 ( .A(sfraddr[0]), .B(n4), .C(n91), .Y(n92) );
  NAND3X1 U12 ( .A(n91), .B(n3), .C(sfraddr[4]), .Y(n96) );
  NAND3X1 U13 ( .A(n91), .B(sfraddr[0]), .C(sfraddr[4]), .Y(n90) );
  NOR2X1 U14 ( .A(n90), .B(n9), .Y(N81) );
  NOR2X1 U15 ( .A(n90), .B(n8), .Y(N80) );
  NOR2X1 U16 ( .A(n90), .B(n6), .Y(N78) );
  NOR2X1 U17 ( .A(n90), .B(n7), .Y(N79) );
  NOR2X1 U18 ( .A(n90), .B(n5), .Y(N77) );
  NOR2X1 U19 ( .A(n9), .B(n93), .Y(N63) );
  NOR2X1 U20 ( .A(n10), .B(n93), .Y(N64) );
  NOR2X1 U21 ( .A(n6), .B(n93), .Y(N60) );
  NOR2X1 U22 ( .A(n8), .B(n93), .Y(N62) );
  NOR2X1 U23 ( .A(n7), .B(n93), .Y(N61) );
  NOR2X1 U24 ( .A(n5), .B(n93), .Y(N59) );
  NOR2X1 U25 ( .A(n10), .B(n90), .Y(N82) );
  NOR2X1 U26 ( .A(n9), .B(n92), .Y(N72) );
  NOR2X1 U27 ( .A(n8), .B(n92), .Y(N71) );
  NOR2X1 U28 ( .A(n10), .B(n92), .Y(N73) );
  NOR2X1 U29 ( .A(n6), .B(n92), .Y(N69) );
  NOR2X1 U30 ( .A(n6), .B(n96), .Y(N51) );
  NOR2X1 U31 ( .A(n10), .B(n96), .Y(N55) );
  NOR2X1 U32 ( .A(n9), .B(n96), .Y(N54) );
  NOR2X1 U33 ( .A(n8), .B(n96), .Y(N53) );
  NOR2X1 U34 ( .A(n7), .B(n92), .Y(N70) );
  NOR2X1 U35 ( .A(n5), .B(n92), .Y(N68) );
  NOR2X1 U36 ( .A(n7), .B(n96), .Y(N52) );
  NOR2X1 U37 ( .A(n5), .B(n96), .Y(N50) );
  NOR2X1 U38 ( .A(n5), .B(n97), .Y(N39) );
  NOR2X1 U39 ( .A(n10), .B(n97), .Y(N44) );
  NOR2X1 U40 ( .A(n6), .B(n97), .Y(N40) );
  NOR2X1 U41 ( .A(n9), .B(n97), .Y(N43) );
  NOR2X1 U42 ( .A(n7), .B(n97), .Y(N41) );
  NOR2X1 U43 ( .A(n8), .B(n97), .Y(N42) );
  NAND2X1 U44 ( .A(n11), .B(n93), .Y(N58) );
  NAND2X1 U45 ( .A(n11), .B(n92), .Y(N67) );
  NAND2X1 U46 ( .A(n11), .B(n97), .Y(N38) );
  NAND2X1 U47 ( .A(n11), .B(n90), .Y(N76) );
  NAND2X1 U48 ( .A(n11), .B(n96), .Y(N49) );
  INVX1 U49 ( .A(n171), .Y(n23) );
  INVX1 U50 ( .A(n70), .Y(n33) );
  NAND2X1 U51 ( .A(n11), .B(n207), .Y(n66) );
  AND2X1 U52 ( .A(sfraddr[1]), .B(sfrwe), .Y(n95) );
  NOR4XL U53 ( .A(sfraddr[6]), .B(sfraddr[2]), .C(sfraddr[1]), .D(rst), .Y(n98) );
  NOR21XL U54 ( .B(sfrdatai[7]), .A(n97), .Y(N45) );
  NAND4X1 U55 ( .A(sfraddr[4]), .B(sfraddr[3]), .C(n94), .D(n60), .Y(n93) );
  NOR2X1 U56 ( .A(sfraddr[2]), .B(sfraddr[0]), .Y(n94) );
  INVX1 U57 ( .A(sfraddr[4]), .Y(n4) );
  NOR21XL U58 ( .B(n99), .A(rst), .Y(N212) );
  NOR3XL U59 ( .A(n176), .B(n24), .C(n188), .Y(n171) );
  NAND3X1 U60 ( .A(n118), .B(n119), .C(n120), .Y(n106) );
  INVX1 U61 ( .A(sfrdatai[5]), .Y(n10) );
  INVX1 U62 ( .A(sfrdatai[1]), .Y(n6) );
  INVX1 U63 ( .A(sfrdatai[4]), .Y(n9) );
  INVX1 U64 ( .A(sfrdatai[0]), .Y(n5) );
  INVX1 U65 ( .A(sfrdatai[2]), .Y(n7) );
  INVX1 U66 ( .A(sfrdatai[3]), .Y(n8) );
  NAND4X1 U67 ( .A(n118), .B(n123), .C(n102), .D(n126), .Y(n99) );
  AOI21AX1 U68 ( .B(n115), .C(n14), .A(n109), .Y(n126) );
  NAND4X1 U69 ( .A(n119), .B(n11), .C(n124), .D(n125), .Y(N207) );
  NOR21XL U70 ( .B(n100), .A(n99), .Y(n125) );
  INVX1 U71 ( .A(n168), .Y(n26) );
  INVX1 U72 ( .A(n108), .Y(n16) );
  INVX1 U73 ( .A(n145), .Y(n14) );
  INVX1 U74 ( .A(n170), .Y(n30) );
  INVX1 U75 ( .A(n165), .Y(n24) );
  AOI31X1 U76 ( .A(n15), .B(n13), .C(n114), .D(rst), .Y(N208) );
  INVX1 U77 ( .A(n113), .Y(n15) );
  AOI211X1 U78 ( .C(n115), .D(n14), .A(n116), .B(n117), .Y(n114) );
  INVX1 U79 ( .A(n106), .Y(n13) );
  AOI31X1 U80 ( .A(n109), .B(n110), .C(n111), .D(rst), .Y(N209) );
  NOR2X1 U81 ( .A(n112), .B(n113), .Y(n111) );
  NOR2X1 U82 ( .A(rst), .B(n100), .Y(N211) );
  INVX1 U83 ( .A(n193), .Y(n25) );
  NOR21XL U84 ( .B(n62), .A(n61), .Y(n70) );
  INVX1 U85 ( .A(intcall), .Y(n207) );
  NAND32X1 U86 ( .B(retiinstr), .C(rst), .A(n61), .Y(n67) );
  INVX1 U87 ( .A(rst), .Y(n11) );
  NAND2X1 U88 ( .A(intcall), .B(n11), .Y(n61) );
  OAI32X1 U89 ( .A(n52), .B(rst), .C(n12), .D(n58), .E(n10), .Y(n200) );
  INVX1 U90 ( .A(n58), .Y(n12) );
  NOR2XL U91 ( .A(sfraddr[4]), .B(sfraddr[3]), .Y(n59) );
  NOR32XL U92 ( .B(n105), .C(n122), .A(n104), .Y(n124) );
  NAND31X1 U93 ( .C(n127), .A(n128), .B(n129), .Y(n109) );
  OAI221X1 U94 ( .A(n20), .B(n141), .C(n140), .D(n138), .E(n17), .Y(n108) );
  INVX1 U95 ( .A(n139), .Y(n17) );
  OAI21X1 U96 ( .B(n172), .C(n57), .A(n186), .Y(n168) );
  NOR3XL U97 ( .A(n44), .B(n161), .C(n150), .Y(n170) );
  AOI211X1 U98 ( .C(n135), .D(n144), .A(n115), .B(n145), .Y(n129) );
  NOR2X1 U99 ( .A(n194), .B(n55), .Y(n187) );
  NOR2X1 U100 ( .A(n189), .B(n158), .Y(n165) );
  NAND3X1 U101 ( .A(n146), .B(n143), .C(n124), .Y(n139) );
  NOR42XL U102 ( .C(n120), .D(n137), .A(n112), .B(n117), .Y(n100) );
  AOI22AXL U103 ( .A(n16), .B(n142), .D(n143), .C(n124), .Y(n137) );
  NAND2X1 U104 ( .A(n121), .B(n107), .Y(n142) );
  OAI21X1 U105 ( .B(n170), .C(n55), .A(n182), .Y(n175) );
  NAND3X1 U106 ( .A(n121), .B(n107), .C(n16), .Y(n145) );
  NAND3X1 U107 ( .A(n162), .B(n152), .C(n138), .Y(n176) );
  AND2X1 U108 ( .A(n184), .B(n194), .Y(n186) );
  AOI31X1 U109 ( .A(n101), .B(n102), .C(n103), .D(rst), .Y(N210) );
  OR2X1 U110 ( .A(n107), .B(n108), .Y(n101) );
  AOI21X1 U111 ( .B(n104), .C(n105), .A(n106), .Y(n103) );
  NAND3X1 U112 ( .A(n144), .B(n135), .C(n14), .Y(n120) );
  INVX1 U113 ( .A(n130), .Y(n22) );
  NAND31X1 U114 ( .C(n153), .A(n141), .B(n127), .Y(n188) );
  OAI221X1 U115 ( .A(n108), .B(n121), .C(n18), .D(n122), .E(n123), .Y(n113) );
  INVX1 U116 ( .A(n105), .Y(n18) );
  OA21X1 U117 ( .B(n22), .C(n148), .A(n131), .Y(n134) );
  NAND2X1 U118 ( .A(n153), .B(n128), .Y(n110) );
  OAI21X1 U119 ( .B(n20), .C(n127), .A(n129), .Y(n132) );
  AOI21X1 U120 ( .B(n133), .C(n44), .A(n132), .Y(n131) );
  AOI21X1 U121 ( .B(n134), .C(n147), .A(n66), .Y(N200) );
  NAND2X1 U122 ( .A(n136), .B(n135), .Y(n147) );
  INVX1 U123 ( .A(n172), .Y(n28) );
  NOR2X1 U124 ( .A(n152), .B(n140), .Y(n116) );
  NAND2X1 U125 ( .A(n150), .B(n133), .Y(n122) );
  NAND21X1 U126 ( .B(n146), .A(n124), .Y(n119) );
  NOR2X1 U127 ( .A(n51), .B(n190), .Y(n193) );
  NOR3XL U128 ( .A(n139), .B(n20), .C(n141), .Y(n112) );
  NOR3XL U129 ( .A(n138), .B(n139), .C(n140), .Y(n117) );
  NAND2X1 U130 ( .A(n161), .B(n133), .Y(n121) );
  INVX1 U131 ( .A(n128), .Y(n20) );
  NAND2X1 U132 ( .A(n155), .B(n154), .Y(n143) );
  NOR2X1 U133 ( .A(n162), .B(n140), .Y(n115) );
  OAI21X1 U134 ( .B(n46), .C(n166), .A(n167), .Y(n180) );
  NAND2X1 U135 ( .A(n88), .B(n36), .Y(n89) );
  OAI22X1 U136 ( .A(n72), .B(n45), .C(n73), .D(n74), .Y(n62) );
  AOI22X1 U137 ( .A(n38), .B(n75), .C(n76), .D(n37), .Y(n74) );
  OAI22X1 U138 ( .A(n39), .B(n57), .C(n79), .D(n51), .Y(n75) );
  OAI222XL U139 ( .A(n77), .B(n50), .C(n78), .D(n47), .E(n79), .F(n49), .Y(n76) );
  OAI32X1 U140 ( .A(n61), .B(n32), .C(n62), .D(n71), .E(n41), .Y(n196) );
  AOI21BBXL U141 ( .B(n66), .C(n65), .A(n70), .Y(n71) );
  AOI211X1 U142 ( .C(n83), .D(n84), .A(int_ack_03), .B(int_ack_43), .Y(n72) );
  OAI22X1 U143 ( .A(n63), .B(n33), .C(n68), .D(n42), .Y(n197) );
  AOI21BX1 U144 ( .C(n66), .B(n69), .A(n70), .Y(n68) );
  NOR2X1 U145 ( .A(n77), .B(n89), .Y(int_ack_1b) );
  OAI22X1 U146 ( .A(n67), .B(n43), .C(n32), .D(n33), .Y(n198) );
  OAI31XL U147 ( .A(n61), .B(n62), .C(n63), .D(n64), .Y(n199) );
  GEN2XL U148 ( .D(n65), .E(n41), .C(n66), .B(n61), .A(n40), .Y(n64) );
  NOR2X1 U149 ( .A(n87), .B(n39), .Y(int_ack_43) );
  NAND2X1 U150 ( .A(n43), .B(n67), .Y(n69) );
  INVX1 U151 ( .A(n63), .Y(n32) );
  INVX1 U152 ( .A(n86), .Y(n38) );
  NOR2X1 U153 ( .A(n78), .B(n35), .Y(int_ack_93) );
  NOR2X1 U154 ( .A(n79), .B(n35), .Y(int_ack_8b) );
  INVX1 U155 ( .A(n83), .Y(n39) );
  INVX1 U156 ( .A(n84), .Y(n35) );
  NOR2X1 U157 ( .A(n77), .B(n87), .Y(int_ack_5b) );
  NOR2X1 U158 ( .A(n79), .B(n89), .Y(int_ack_0b) );
  NOR2X1 U159 ( .A(n78), .B(n89), .Y(int_ack_13) );
  NOR2X1 U160 ( .A(n78), .B(n87), .Y(int_ack_53) );
  NOR2X1 U161 ( .A(n79), .B(n87), .Y(int_ack_4b) );
  NAND31X1 U162 ( .C(n132), .A(n44), .B(n133), .Y(n123) );
  NAND3X1 U163 ( .A(n48), .B(n130), .C(n131), .Y(n102) );
  NAND3X1 U164 ( .A(n134), .B(n135), .C(n136), .Y(n118) );
  NOR3XL U165 ( .A(n85), .B(n39), .C(n86), .Y(int_ack_a3) );
  NOR3XL U166 ( .A(n85), .B(n79), .C(n86), .Y(int_ack_ab) );
  INVX1 U167 ( .A(n203), .Y(n44) );
  NOR2X1 U168 ( .A(n77), .B(n35), .Y(int_ack_9b) );
  INVX1 U169 ( .A(n148), .Y(n48) );
  AND2X1 U170 ( .A(irq_r), .B(ien0[7]), .Y(irq) );
  NOR21XL U171 ( .B(n202), .A(n166), .Y(n183) );
  AOI33X1 U172 ( .A(ip0[1]), .B(n176), .C(ip1[1]), .D(ip0[2]), .E(n188), .F(
        ip1[2]), .Y(n202) );
  NOR21XL U173 ( .B(ien1[0]), .A(n205), .Y(n155) );
  AOI22X1 U174 ( .A(int_vect_43), .B(n52), .C(sdaiff), .D(isr_tm), .Y(n205) );
  OAI211X1 U175 ( .C(n45), .D(n192), .A(n43), .B(ien0[7]), .Y(n166) );
  NOR43XL U176 ( .B(n26), .C(n192), .D(n25), .A(is_reg[1]), .Y(n164) );
  AOI31X1 U177 ( .A(ip0[4]), .B(n29), .C(n183), .D(n186), .Y(n185) );
  INVX1 U178 ( .A(n187), .Y(n29) );
  AO21X1 U179 ( .B(ien0[0]), .C(int_vect_03), .A(n155), .Y(n189) );
  AOI21X1 U180 ( .B(n188), .C(ip0[2]), .A(n178), .Y(n182) );
  OAI21X1 U181 ( .B(n51), .C(n168), .A(n169), .Y(n135) );
  AOI32X1 U182 ( .A(n170), .B(n171), .C(n172), .D(ip0[5]), .E(n173), .Y(n169)
         );
  OAI22X1 U183 ( .A(n51), .B(n160), .C(n174), .D(n175), .Y(n173) );
  NOR2X1 U184 ( .A(n172), .B(n56), .Y(n174) );
  AND3X1 U185 ( .A(ien0[3]), .B(int_vect_1b), .C(n52), .Y(n150) );
  AOI211X1 U186 ( .C(n52), .D(n206), .A(n22), .B(n149), .Y(n104) );
  OAI21X1 U187 ( .B(n52), .C(rxd0ff), .A(ien0[4]), .Y(n149) );
  NAND2X1 U188 ( .A(n201), .B(n183), .Y(n160) );
  AOI31X1 U189 ( .A(ip0[4]), .B(n28), .C(ip1[4]), .D(n187), .Y(n201) );
  OAI211X1 U190 ( .C(n190), .D(n54), .A(n40), .B(n191), .Y(n158) );
  AOI21X1 U191 ( .B(ip0[4]), .C(n28), .A(n175), .Y(n191) );
  AOI221XL U192 ( .A(n176), .B(ip1[1]), .C(n188), .D(ip1[2]), .E(n167), .Y(
        n184) );
  INVX1 U193 ( .A(isr_tm), .Y(n52) );
  NAND2X1 U194 ( .A(int_vect_8b), .B(ien2[1]), .Y(n162) );
  OAI21BBX1 U195 ( .A(n176), .B(ip0[1]), .C(n164), .Y(n178) );
  NAND4X1 U196 ( .A(int_vect_4b), .B(ien1[1]), .C(n162), .D(n52), .Y(n138) );
  NAND3X1 U197 ( .A(n159), .B(n42), .C(n195), .Y(n167) );
  AOI21X1 U198 ( .B(ip1[0]), .C(n189), .A(n160), .Y(n195) );
  NAND2X1 U199 ( .A(ip1[3]), .B(n30), .Y(n194) );
  NAND3X1 U200 ( .A(i2c_int), .B(n135), .C(ien0[5]), .Y(n146) );
  NAND2X1 U201 ( .A(ip0[0]), .B(n189), .Y(n192) );
  AOI32X1 U202 ( .A(ip0[2]), .B(n53), .C(n31), .D(n179), .E(n180), .Y(n177) );
  NAND2X1 U203 ( .A(ip1[1]), .B(n176), .Y(n179) );
  INVX1 U204 ( .A(n166), .Y(n31) );
  ENOX1 U205 ( .A(n206), .B(isr_tm), .C(rxd0ff), .D(isr_tm), .Y(n204) );
  OAI221X1 U206 ( .A(n181), .B(n50), .C(n55), .D(n19), .E(n23), .Y(n133) );
  AOI21X1 U207 ( .B(n183), .C(ip0[3]), .A(n184), .Y(n181) );
  INVX1 U208 ( .A(n182), .Y(n19) );
  AOI221XL U209 ( .A(n163), .B(ip1[1]), .C(ip0[1]), .D(n164), .E(n165), .Y(
        n140) );
  OAI21X1 U210 ( .B(n166), .C(n53), .A(n167), .Y(n163) );
  AND3X1 U211 ( .A(ien1[3]), .B(int_vect_5b), .C(n203), .Y(n161) );
  OAI211X1 U212 ( .C(n156), .D(n45), .A(n157), .B(n158), .Y(n154) );
  AOI33X1 U213 ( .A(n159), .B(n42), .C(n27), .D(ip0[0]), .E(n43), .F(ien0[7]), 
        .Y(n156) );
  NAND4X1 U214 ( .A(n26), .B(ip0[0]), .C(n25), .D(n41), .Y(n157) );
  INVX1 U215 ( .A(n160), .Y(n27) );
  AND2X1 U216 ( .A(int_vect_13), .B(ien0[2]), .Y(n153) );
  NAND2X1 U217 ( .A(int_vect_93), .B(ien2[2]), .Y(n127) );
  NAND3X1 U218 ( .A(ien1[2]), .B(n127), .C(int_vect_53), .Y(n141) );
  NAND3X1 U219 ( .A(ien0[1]), .B(n52), .C(int_vect_0b), .Y(n152) );
  INVX1 U220 ( .A(int_vect_23), .Y(n206) );
  AOI211X1 U221 ( .C(int_vect_03), .D(n151), .A(n21), .B(n116), .Y(n105) );
  AND2X1 U222 ( .A(ien0[0]), .B(n154), .Y(n151) );
  INVX1 U223 ( .A(n110), .Y(n21) );
  NOR32XL U224 ( .B(ien1[5]), .C(int_vect_6b), .A(n136), .Y(n144) );
  AOI211X1 U225 ( .C(i2c_int), .D(ien0[5]), .A(n144), .B(n136), .Y(n190) );
  NAND4X1 U226 ( .A(int_vect_63), .B(ien1[4]), .C(n130), .D(n148), .Y(n107) );
  INVX1 U227 ( .A(is_reg[3]), .Y(n43) );
  INVX1 U228 ( .A(ip0[3]), .Y(n55) );
  NAND2X1 U229 ( .A(n193), .B(ip0[5]), .Y(n159) );
  INVX1 U230 ( .A(ip1[0]), .Y(n45) );
  INVX1 U231 ( .A(ip1[5]), .Y(n51) );
  INVX1 U232 ( .A(is_reg[2]), .Y(n42) );
  INVX1 U233 ( .A(ip1[4]), .Y(n57) );
  INVX1 U234 ( .A(ip0[2]), .Y(n46) );
  INVX1 U235 ( .A(ip0[5]), .Y(n54) );
  INVX1 U236 ( .A(is_reg[1]), .Y(n41) );
  INVX1 U237 ( .A(ip0[4]), .Y(n56) );
  INVX1 U238 ( .A(ip0[1]), .Y(n53) );
  INVX1 U239 ( .A(ip1[2]), .Y(n47) );
  INVX1 U240 ( .A(is_reg[0]), .Y(n40) );
  INVX1 U241 ( .A(ip1[3]), .Y(n50) );
  AO222X1 U242 ( .A(intcall), .B(n73), .C(n38), .D(intvect[1]), .E(n83), .F(
        n34), .Y(int_ack_03) );
  INVX1 U243 ( .A(n89), .Y(n34) );
  NOR3XL U244 ( .A(intvect[2]), .B(intvect[4]), .C(n207), .Y(n88) );
  OAI22AX1 U245 ( .D(ip0[0]), .C(n72), .A(n73), .B(n80), .Y(n63) );
  AOI22X1 U246 ( .A(n38), .B(n81), .C(n82), .D(n37), .Y(n80) );
  OAI22X1 U247 ( .A(n39), .B(n56), .C(n79), .D(n54), .Y(n81) );
  OAI222XL U248 ( .A(n77), .B(n55), .C(n78), .D(n46), .E(n79), .F(n53), .Y(n82) );
  NOR3XL U249 ( .A(n207), .B(intvect[2]), .C(n85), .Y(n84) );
  NAND2X1 U250 ( .A(intvect[2]), .B(intcall), .Y(n86) );
  NAND2X1 U251 ( .A(n88), .B(intvect[3]), .Y(n87) );
  INVX1 U252 ( .A(intvect[3]), .Y(n36) );
  NOR2X1 U253 ( .A(n69), .B(is_reg[2]), .Y(n65) );
  NAND21X1 U254 ( .B(intvect[1]), .A(intvect[0]), .Y(n79) );
  NAND21X1 U255 ( .B(intvect[0]), .A(intvect[1]), .Y(n78) );
  NOR2X1 U256 ( .A(intvect[0]), .B(intvect[1]), .Y(n83) );
  AND2X1 U257 ( .A(intvect[4]), .B(intvect[3]), .Y(n73) );
  NAND2X1 U258 ( .A(intvect[1]), .B(intvect[0]), .Y(n77) );
  NAND2X1 U259 ( .A(intvect[4]), .B(n36), .Y(n85) );
  INVX1 U260 ( .A(ip1[1]), .Y(n49) );
  NOR4XL U261 ( .A(intvect[4]), .B(n36), .C(n79), .D(n86), .Y(int_ack_6b) );
  NOR4XL U262 ( .A(intvect[4]), .B(n36), .C(n39), .D(n86), .Y(int_ack_63) );
  INVX1 U263 ( .A(intvect[2]), .Y(n37) );
  AND2X1 U264 ( .A(int_vect_ab), .B(ien2[5]), .Y(n136) );
  NAND2X1 U265 ( .A(int_vect_a3), .B(ien2[4]), .Y(n148) );
  NAND2X1 U266 ( .A(int_vect_9b), .B(ien2[3]), .Y(n203) );
  AND4XL U268 ( .A(sfraddr[3]), .B(sfrwe), .C(sfraddr[5]), .D(n98), .Y(n91) );
  NOR42XL U269 ( .C(n11), .D(n95), .A(sfraddr[5]), .B(sfraddr[6]), .Y(n60) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module watchdog_a0 ( wdt_slow, clkwdt, clkper, resetff, newinstr, wdts_s, wdts, 
        ip0wdts, wdt_tm, sfrdatai, sfraddr, sfrwe, wdtrel, test_si, test_se );
  output [1:0] wdts_s;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] wdtrel;
  input wdt_slow, clkwdt, clkper, resetff, newinstr, sfrwe, test_si, test_se;
  output wdts, ip0wdts, wdt_tm;
  wire   wdt_tm_sync, wdt_act_sync, wdt_act, wdtrefresh_sync, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N67, N68, N69, N70, N71, pres_2, N112,
         N113, N114, N115, N116, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, wdt_normal, wdt_normal_ff, N212, net12144, net12150,
         net12155, net12160, net12165, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n117, n118;
  wire   [1:0] pres_8;
  wire   [3:0] cycles_reg;
  wire   [3:0] pres_16;
  wire   [6:0] wdth;
  wire   [7:0] wdtl;

  SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 clk_gate_wdtrel_s_reg ( .CLK(clkper), 
        .EN(N26), .ENCLK(net12144), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 clk_gate_cycles_reg_reg ( .CLK(clkwdt), 
        .EN(N67), .ENCLK(net12150), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 clk_gate_pres_16_reg ( .CLK(clkwdt), .EN(
        N112), .ENCLK(net12155), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 clk_gate_wdth_reg ( .CLK(clkwdt), .EN(
        N165), .ENCLK(net12160), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 clk_gate_wdtl_reg ( .CLK(clkwdt), .EN(
        n116), .ENCLK(net12165), .TE(test_se) );
  watchdog_a0_DW01_inc_0 add_278 ( .A(wdtl), .SUM({N144, N143, N142, N141, 
        N140, N139, N138, N137}) );
  watchdog_a0_DW01_inc_1 add_272 ( .A(wdth), .SUM({N136, N135, N134, N133, 
        N132, N131, N130}) );
  SDFFQX1 wdt_act_reg ( .D(n130), .SIN(pres_16[3]), .SMC(test_se), .C(clkper), 
        .Q(wdt_act) );
  SDFFQX1 wdts_reg ( .D(wdts_s[0]), .SIN(wdtrel[7]), .SMC(test_se), .C(clkper), 
        .Q(wdts) );
  SDFFQX1 wdts_s_reg_1_ ( .D(n126), .SIN(wdts_s[0]), .SMC(test_se), .C(
        net12165), .Q(wdts_s[1]) );
  SDFFQX1 wdts_s_reg_0_ ( .D(n132), .SIN(wdts), .SMC(test_se), .C(net12165), 
        .Q(wdts_s[0]) );
  SDFFQX1 wdt_normal_ff_reg ( .D(n115), .SIN(wdt_act_sync), .SMC(test_se), .C(
        clkper), .Q(wdt_normal_ff) );
  SDFFQX1 wdt_normal_reg ( .D(n133), .SIN(wdt_normal_ff), .SMC(test_se), .C(
        clkper), .Q(wdt_normal) );
  SDFFQX1 wdt_act_sync_reg ( .D(wdt_act), .SIN(wdt_act), .SMC(test_se), .C(
        clkwdt), .Q(wdt_act_sync) );
  SDFFQX1 pres_16_reg_3_ ( .D(N116), .SIN(pres_16[2]), .SMC(test_se), .C(
        net12155), .Q(pres_16[3]) );
  SDFFQX1 wdth_reg_6_ ( .D(N172), .SIN(wdth[5]), .SMC(test_se), .C(net12160), 
        .Q(wdth[6]) );
  SDFFQX1 pres_8_reg_1_ ( .D(n128), .SIN(pres_8[0]), .SMC(test_se), .C(
        net12150), .Q(pres_8[1]) );
  SDFFQX1 pres_16_reg_2_ ( .D(N115), .SIN(pres_16[1]), .SMC(test_se), .C(
        net12155), .Q(pres_16[2]) );
  SDFFQX1 pres_2_reg ( .D(n127), .SIN(ip0wdts), .SMC(test_se), .C(net12150), 
        .Q(pres_2) );
  SDFFQX1 pres_8_reg_0_ ( .D(n129), .SIN(pres_2), .SMC(test_se), .C(net12150), 
        .Q(pres_8[0]) );
  SDFFQX1 wdt_tm_sync_reg ( .D(wdt_tm), .SIN(wdt_tm), .SMC(test_se), .C(clkwdt), .Q(wdt_tm_sync) );
  SDFFQX1 pres_16_reg_1_ ( .D(N114), .SIN(pres_16[0]), .SMC(test_se), .C(
        net12155), .Q(pres_16[1]) );
  SDFFQX1 cycles_reg_reg_2_ ( .D(N70), .SIN(cycles_reg[1]), .SMC(test_se), .C(
        net12150), .Q(cycles_reg[2]) );
  SDFFQX1 pres_16_reg_0_ ( .D(N113), .SIN(pres_8[1]), .SMC(test_se), .C(
        net12155), .Q(pres_16[0]) );
  SDFFQX1 wdth_reg_4_ ( .D(N170), .SIN(wdth[3]), .SMC(test_se), .C(net12160), 
        .Q(wdth[4]) );
  SDFFQX1 wdtl_reg_2_ ( .D(N175), .SIN(wdtl[1]), .SMC(test_se), .C(net12165), 
        .Q(wdtl[2]) );
  SDFFQX1 cycles_reg_reg_3_ ( .D(N71), .SIN(cycles_reg[2]), .SMC(test_se), .C(
        net12150), .Q(cycles_reg[3]) );
  SDFFQX1 wdtl_reg_4_ ( .D(N177), .SIN(wdtl[3]), .SMC(test_se), .C(net12165), 
        .Q(wdtl[4]) );
  SDFFQX1 wdtrefresh_reg ( .D(N212), .SIN(wdtl[7]), .SMC(test_se), .C(clkper), 
        .Q(wdtrefresh_sync) );
  SDFFQX1 cycles_reg_reg_1_ ( .D(N69), .SIN(cycles_reg[0]), .SMC(test_se), .C(
        net12150), .Q(cycles_reg[1]) );
  SDFFQX1 cycles_reg_reg_0_ ( .D(N68), .SIN(test_si), .SMC(test_se), .C(
        net12150), .Q(cycles_reg[0]) );
  SDFFQX1 wdth_reg_1_ ( .D(N167), .SIN(wdth[0]), .SMC(test_se), .C(net12160), 
        .Q(wdth[1]) );
  SDFFQX1 wdth_reg_3_ ( .D(N169), .SIN(wdth[2]), .SMC(test_se), .C(net12160), 
        .Q(wdth[3]) );
  SDFFQX1 wdth_reg_2_ ( .D(N168), .SIN(wdth[1]), .SMC(test_se), .C(net12160), 
        .Q(wdth[2]) );
  SDFFQX1 wdtl_reg_6_ ( .D(N179), .SIN(wdtl[5]), .SMC(test_se), .C(net12165), 
        .Q(wdtl[6]) );
  SDFFQX1 wdtl_reg_5_ ( .D(N178), .SIN(wdtl[4]), .SMC(test_se), .C(net12165), 
        .Q(wdtl[5]) );
  SDFFQX1 wdtl_reg_7_ ( .D(N180), .SIN(wdtl[6]), .SMC(test_se), .C(net12165), 
        .Q(wdtl[7]) );
  SDFFQX1 wdth_reg_5_ ( .D(N171), .SIN(wdth[4]), .SMC(test_se), .C(net12160), 
        .Q(wdth[5]) );
  SDFFQX1 wdtl_reg_1_ ( .D(N174), .SIN(wdtl[0]), .SMC(test_se), .C(net12165), 
        .Q(wdtl[1]) );
  SDFFQX1 wdtl_reg_3_ ( .D(N176), .SIN(wdtl[2]), .SMC(test_se), .C(net12165), 
        .Q(wdtl[3]) );
  SDFFQX1 wdth_reg_0_ ( .D(N166), .SIN(wdt_tm_sync), .SMC(test_se), .C(
        net12160), .Q(wdth[0]) );
  SDFFQX1 wdtl_reg_0_ ( .D(N173), .SIN(wdth[6]), .SMC(test_se), .C(net12165), 
        .Q(wdtl[0]) );
  SDFFQX1 wdtrel_s_reg_1_ ( .D(N28), .SIN(wdtrel[0]), .SMC(test_se), .C(
        net12144), .Q(wdtrel[1]) );
  SDFFQX1 wdtrel_s_reg_3_ ( .D(N30), .SIN(wdtrel[2]), .SMC(test_se), .C(
        net12144), .Q(wdtrel[3]) );
  SDFFQX1 wdtrel_s_reg_2_ ( .D(N29), .SIN(wdtrel[1]), .SMC(test_se), .C(
        net12144), .Q(wdtrel[2]) );
  SDFFQX1 ip0wdts_reg ( .D(n131), .SIN(cycles_reg[3]), .SMC(test_se), .C(
        clkper), .Q(ip0wdts) );
  SDFFQX1 wdtrel_s_reg_7_ ( .D(N34), .SIN(wdtrel[6]), .SMC(test_se), .C(
        net12144), .Q(wdtrel[7]) );
  SDFFQX1 wdt_tm_s_reg ( .D(n134), .SIN(wdt_normal), .SMC(test_se), .C(clkper), 
        .Q(wdt_tm) );
  SDFFQX1 wdtrel_s_reg_6_ ( .D(N33), .SIN(wdtrel[5]), .SMC(test_se), .C(
        net12144), .Q(wdtrel[6]) );
  SDFFQX1 wdtrel_s_reg_4_ ( .D(N31), .SIN(wdtrel[3]), .SMC(test_se), .C(
        net12144), .Q(wdtrel[4]) );
  SDFFQX1 wdtrel_s_reg_0_ ( .D(N27), .SIN(wdtrefresh_sync), .SMC(test_se), .C(
        net12144), .Q(wdtrel[0]) );
  SDFFQX1 wdtrel_s_reg_5_ ( .D(N32), .SIN(wdtrel[4]), .SMC(test_se), .C(
        net12144), .Q(wdtrel[5]) );
  NOR2X1 U3 ( .A(n58), .B(wdtrefresh_sync), .Y(n1) );
  INVX1 U4 ( .A(sfraddr[0]), .Y(n2) );
  NAND2X1 U5 ( .A(n33), .B(n2), .Y(n32) );
  INVX1 U6 ( .A(n4), .Y(n3) );
  INVX1 U7 ( .A(n110), .Y(n11) );
  AND4X1 U8 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(n48), .D(n49), .Y(n33) );
  NOR2XL U9 ( .A(sfraddr[2]), .B(sfraddr[1]), .Y(n48) );
  INVX1 U10 ( .A(n25), .Y(n5) );
  NOR21XL U11 ( .B(sfrdatai[4]), .A(n97), .Y(N31) );
  NOR21XL U12 ( .B(sfrdatai[2]), .A(n97), .Y(N29) );
  NOR21XL U13 ( .B(sfrdatai[5]), .A(n97), .Y(N32) );
  NOR21XL U14 ( .B(sfrdatai[0]), .A(n97), .Y(N27) );
  NOR21XL U15 ( .B(sfrdatai[1]), .A(n97), .Y(N28) );
  NOR21XL U16 ( .B(sfrdatai[3]), .A(n97), .Y(N30) );
  NOR21XL U17 ( .B(sfrdatai[7]), .A(n97), .Y(N34) );
  NOR2X1 U18 ( .A(n4), .B(n97), .Y(N33) );
  NAND4X1 U19 ( .A(sfrwe), .B(n2), .C(n99), .D(n100), .Y(n50) );
  NOR3XL U20 ( .A(sfraddr[1]), .B(sfraddr[6]), .C(sfraddr[2]), .Y(n99) );
  AND4X1 U21 ( .A(sfraddr[3]), .B(sfraddr[5]), .C(sfraddr[4]), .D(n3), .Y(n100) );
  INVX1 U22 ( .A(sfrdatai[6]), .Y(n4) );
  NAND2X1 U23 ( .A(n61), .B(n12), .Y(n110) );
  NOR32XL U24 ( .B(n117), .C(n32), .A(newinstr), .Y(n25) );
  NAND2X1 U25 ( .A(n31), .B(n2), .Y(n97) );
  NAND2X1 U26 ( .A(n117), .B(n97), .Y(N26) );
  NOR32XL U27 ( .B(n39), .C(n9), .A(n61), .Y(n60) );
  NOR3XL U28 ( .A(n14), .B(n13), .C(n15), .Y(n61) );
  NAND3X1 U29 ( .A(n66), .B(n67), .C(n68), .Y(n64) );
  AOI211X1 U30 ( .C(n80), .D(n81), .A(n82), .B(n83), .Y(n67) );
  AOI211X1 U31 ( .C(n87), .D(n118), .A(n88), .B(n89), .Y(n66) );
  NOR4XL U32 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(n68) );
  INVX1 U33 ( .A(n57), .Y(n15) );
  NAND2X1 U34 ( .A(n73), .B(n23), .Y(n85) );
  INVX1 U35 ( .A(n102), .Y(n16) );
  NAND2X1 U36 ( .A(n26), .B(n38), .Y(n35) );
  NOR21XL U37 ( .B(N143), .A(n35), .Y(N179) );
  NOR21XL U38 ( .B(N142), .A(n35), .Y(N178) );
  NOR21XL U39 ( .B(N141), .A(n35), .Y(N177) );
  NOR21XL U40 ( .B(N140), .A(n35), .Y(N176) );
  NOR21XL U41 ( .B(N138), .A(n35), .Y(N174) );
  NOR21XL U42 ( .B(N139), .A(n35), .Y(N175) );
  OAI21X1 U43 ( .B(n112), .C(n110), .A(n53), .Y(N115) );
  XNOR2XL U44 ( .A(n111), .B(n20), .Y(n112) );
  ENOX1 U45 ( .A(n22), .B(n28), .C(N135), .D(n26), .Y(N171) );
  ENOX1 U46 ( .A(n23), .B(n28), .C(N134), .D(n1), .Y(N170) );
  NAND2X1 U47 ( .A(n1), .B(n16), .Y(n93) );
  NOR2X1 U48 ( .A(n20), .B(n111), .Y(n105) );
  OAI211X1 U49 ( .C(n38), .D(n101), .A(n28), .B(n117), .Y(N165) );
  NAND21X1 U50 ( .B(n27), .A(n26), .Y(n101) );
  INVX1 U51 ( .A(n58), .Y(n12) );
  OAI2B11X1 U52 ( .D(n1), .C(n27), .A(n28), .B(n117), .Y(n116) );
  INVX1 U53 ( .A(n94), .Y(n17) );
  NAND2X1 U54 ( .A(n117), .B(n58), .Y(N67) );
  OAI32X1 U55 ( .A(n32), .B(resetff), .C(n4), .D(n10), .E(n5), .Y(n133) );
  OAI32X1 U56 ( .A(n10), .B(resetff), .C(n25), .D(n5), .E(n6), .Y(n115) );
  AND4XL U57 ( .A(sfraddr[1]), .B(n49), .C(sfraddr[2]), .D(n98), .Y(n31) );
  NOR3XL U58 ( .A(resetff), .B(sfraddr[5]), .C(sfraddr[3]), .Y(n98) );
  OAI21X1 U59 ( .B(n29), .C(n4), .A(n30), .Y(n134) );
  NAND3X1 U60 ( .A(n29), .B(n117), .C(wdt_tm), .Y(n30) );
  NAND2X1 U61 ( .A(sfraddr[0]), .B(n31), .Y(n29) );
  AOI21X1 U62 ( .B(n45), .C(n46), .A(resetff), .Y(n131) );
  NAND21X1 U63 ( .B(n47), .A(n3), .Y(n45) );
  OAI21X1 U64 ( .B(ip0wdts), .C(wdts_s[0]), .A(n47), .Y(n46) );
  NAND2X1 U65 ( .A(sfraddr[0]), .B(n33), .Y(n47) );
  OAI31XL U66 ( .A(n50), .B(wdts_s[0]), .C(resetff), .D(n51), .Y(n130) );
  OAI21X1 U67 ( .B(wdts_s[0]), .C(n117), .A(wdt_act), .Y(n51) );
  NOR3XL U68 ( .A(n50), .B(resetff), .C(n6), .Y(N212) );
  NOR21XL U69 ( .B(n75), .A(wdtrel[3]), .Y(n73) );
  NOR21XL U70 ( .B(n77), .A(wdtrel[2]), .Y(n75) );
  XNOR2XL U71 ( .A(wdtrel[1]), .B(wdth[0]), .Y(n80) );
  XNOR2XL U72 ( .A(wdtrel[6]), .B(wdth[5]), .Y(n86) );
  XNOR2XL U73 ( .A(n75), .B(n76), .Y(n71) );
  XNOR2XL U74 ( .A(wdtrel[3]), .B(wdth[2]), .Y(n76) );
  XNOR2XL U75 ( .A(n73), .B(n74), .Y(n72) );
  XNOR2XL U76 ( .A(wdtrel[4]), .B(wdth[3]), .Y(n74) );
  XNOR2XL U77 ( .A(n77), .B(n78), .Y(n70) );
  XNOR2XL U78 ( .A(wdtrel[2]), .B(wdth[1]), .Y(n78) );
  XNOR2XL U79 ( .A(wdtl[7]), .B(wdt_slow), .Y(n44) );
  NOR3XL U80 ( .A(n94), .B(cycles_reg[2]), .C(n21), .Y(n102) );
  OAI22BX1 U81 ( .B(n34), .A(n35), .D(wdts_s[0]), .C(n34), .Y(n132) );
  OAI211X1 U82 ( .C(n36), .D(n37), .A(n38), .B(n39), .Y(n34) );
  NAND4X1 U83 ( .A(wdth[6]), .B(wdth[5]), .C(n40), .D(wdth[4]), .Y(n37) );
  NAND41X1 U84 ( .D(n41), .A(wdth[0]), .B(wdth[1]), .C(n42), .Y(n36) );
  NOR2X1 U85 ( .A(n16), .B(wdtrefresh_sync), .Y(n57) );
  NAND2X1 U86 ( .A(cycles_reg[1]), .B(cycles_reg[0]), .Y(n94) );
  OAI32X1 U87 ( .A(n59), .B(resetff), .C(n60), .D(n7), .E(n8), .Y(n127) );
  INVX1 U88 ( .A(pres_2), .Y(n7) );
  AOI21BBXL U89 ( .B(pres_2), .C(wdtrefresh_sync), .A(wdt_tm_sync), .Y(n59) );
  INVX1 U90 ( .A(n60), .Y(n8) );
  OAI21X1 U91 ( .B(n84), .C(n85), .A(n18), .Y(n82) );
  AOI22X1 U92 ( .A(n86), .B(n22), .C(wdtrel[5]), .D(wdth[4]), .Y(n84) );
  OAI22X1 U93 ( .A(n62), .B(n63), .C(n35), .D(n64), .Y(n126) );
  NAND2X1 U94 ( .A(wdts_s[1]), .B(n39), .Y(n63) );
  OAI2B11X1 U95 ( .D(wdtl[2]), .C(n65), .A(n64), .B(n38), .Y(n62) );
  NAND21X1 U96 ( .B(n43), .A(n41), .Y(n65) );
  NAND4X1 U97 ( .A(n106), .B(n107), .C(wdtl[0]), .D(n108), .Y(n43) );
  XNOR2XL U98 ( .A(n118), .B(wdtl[5]), .Y(n106) );
  NOR2X1 U99 ( .A(n18), .B(n19), .Y(n108) );
  XNOR2XL U100 ( .A(n118), .B(wdtl[6]), .Y(n107) );
  NOR3XL U101 ( .A(n43), .B(wdtl[2]), .C(n44), .Y(n42) );
  AOI21AX1 U102 ( .B(n90), .C(n86), .A(n85), .Y(n89) );
  XNOR2XL U103 ( .A(wdtrel[5]), .B(wdth[4]), .Y(n90) );
  OAI211X1 U104 ( .C(wdtl[7]), .D(n80), .A(wdtl[6]), .B(wdtl[4]), .Y(n87) );
  NOR2X1 U105 ( .A(wdtrel[1]), .B(wdtrel[0]), .Y(n77) );
  NAND3X1 U106 ( .A(wdtl[2]), .B(wdtl[0]), .C(n79), .Y(n69) );
  AOI22AXL U107 ( .A(wdtl[3]), .B(wdtl[5]), .D(wdtl[5]), .C(wdtl[6]), .Y(n79)
         );
  INVX1 U108 ( .A(wdtl[3]), .Y(n19) );
  INVX1 U109 ( .A(wdtl[1]), .Y(n18) );
  NAND2X1 U110 ( .A(n53), .B(n113), .Y(N114) );
  OAI211X1 U111 ( .C(pres_16[1]), .D(pres_16[0]), .A(n111), .B(n11), .Y(n113)
         );
  NAND3X1 U112 ( .A(n53), .B(n117), .C(n114), .Y(N112) );
  AOI22X1 U113 ( .A(n11), .B(pres_2), .C(n12), .D(wdtrefresh_sync), .Y(n114)
         );
  NAND42X1 U114 ( .C(n44), .D(n43), .A(wdtl[2]), .B(wdtl[4]), .Y(n38) );
  NAND31X1 U115 ( .C(n52), .A(n53), .B(n54), .Y(n129) );
  NAND4X1 U116 ( .A(n39), .B(pres_8[0]), .C(n15), .D(n9), .Y(n54) );
  XNOR2XL U117 ( .A(wdtl[4]), .B(n118), .Y(n41) );
  NOR21XL U118 ( .B(N137), .A(n35), .Y(N173) );
  NOR21XL U119 ( .B(N144), .A(n35), .Y(N180) );
  NOR2X1 U120 ( .A(n58), .B(wdtrefresh_sync), .Y(n26) );
  AO22AXL U121 ( .A(N136), .B(n1), .C(wdtrel[6]), .D(n28), .Y(N172) );
  INVX1 U122 ( .A(resetff), .Y(n117) );
  NAND2X1 U123 ( .A(wdt_act_sync), .B(n117), .Y(n58) );
  AND2X1 U124 ( .A(wdth[2]), .B(wdth[3]), .Y(n40) );
  NOR3XL U125 ( .A(n58), .B(pres_8[0]), .C(n15), .Y(n52) );
  OAI22X1 U126 ( .A(wdth[4]), .B(n86), .C(n91), .D(n118), .Y(n88) );
  AOI211X1 U127 ( .C(n80), .D(wdtl[4]), .A(n19), .B(wdtl[7]), .Y(n91) );
  OAI21X1 U128 ( .B(pres_16[0]), .C(n110), .A(n53), .Y(N113) );
  OAI21X1 U129 ( .B(n109), .C(n110), .A(n53), .Y(N116) );
  XNOR2XL U130 ( .A(pres_16[3]), .B(n105), .Y(n109) );
  OAI21X1 U131 ( .B(n92), .C(n93), .A(n53), .Y(N71) );
  AOI32X1 U132 ( .A(n17), .B(n21), .C(cycles_reg[2]), .D(cycles_reg[3]), .E(
        n94), .Y(n92) );
  OAI21X1 U133 ( .B(cycles_reg[0]), .C(n93), .A(n53), .Y(N68) );
  NAND2X1 U134 ( .A(pres_16[1]), .B(pres_16[0]), .Y(n111) );
  AOI21X1 U135 ( .B(wdtl[4]), .C(n24), .A(n80), .Y(n83) );
  OAI211X1 U136 ( .C(n55), .D(n14), .A(n56), .B(n53), .Y(n128) );
  NAND4X1 U137 ( .A(n57), .B(n12), .C(pres_8[0]), .D(n14), .Y(n56) );
  AOI31X1 U138 ( .A(n15), .B(n9), .C(n39), .D(n52), .Y(n55) );
  NAND4X1 U139 ( .A(n102), .B(n103), .C(pres_2), .D(n104), .Y(n27) );
  NOR2X1 U140 ( .A(n13), .B(n14), .Y(n104) );
  OAI21BBX1 U141 ( .A(n105), .B(pres_16[3]), .C(wdtrel[7]), .Y(n103) );
  INVX1 U142 ( .A(wdtrel[4]), .Y(n23) );
  INVX1 U143 ( .A(wdtrel[0]), .Y(n24) );
  INVX1 U144 ( .A(wdtrel[5]), .Y(n22) );
  OR2X1 U145 ( .A(wdtl[7]), .B(n24), .Y(n81) );
  INVX1 U146 ( .A(cycles_reg[3]), .Y(n21) );
  AO22AXL U147 ( .A(N132), .B(n26), .C(wdtrel[2]), .D(n28), .Y(N168) );
  AO22AXL U148 ( .A(N133), .B(n1), .C(wdtrel[3]), .D(n28), .Y(N169) );
  AO22AXL U149 ( .A(N131), .B(n26), .C(wdtrel[1]), .D(n28), .Y(N167) );
  NAND2X1 U150 ( .A(wdt_tm_sync), .B(n12), .Y(n53) );
  NOR2X1 U151 ( .A(wdtrefresh_sync), .B(resetff), .Y(n39) );
  NAND2X1 U152 ( .A(wdtrefresh_sync), .B(n117), .Y(n28) );
  OAI21X1 U153 ( .B(n93), .C(n96), .A(n53), .Y(N69) );
  OAI21X1 U154 ( .B(cycles_reg[1]), .C(cycles_reg[0]), .A(n94), .Y(n96) );
  INVX1 U155 ( .A(wdt_tm_sync), .Y(n9) );
  NOR3XL U156 ( .A(n93), .B(wdt_tm_sync), .C(n95), .Y(N70) );
  XNOR2XL U157 ( .A(n17), .B(cycles_reg[2]), .Y(n95) );
  INVX1 U158 ( .A(pres_8[1]), .Y(n14) );
  ENOX1 U159 ( .A(n24), .B(n28), .C(N130), .D(n26), .Y(N166) );
  INVX1 U160 ( .A(pres_8[0]), .Y(n13) );
  INVX1 U161 ( .A(pres_16[2]), .Y(n20) );
  INVX1 U162 ( .A(wdt_normal), .Y(n10) );
  INVX1 U163 ( .A(wdt_normal_ff), .Y(n6) );
  INVX1 U164 ( .A(wdt_slow), .Y(n118) );
  NOR31XL U165 ( .C(sfrwe), .A(sfraddr[4]), .B(sfraddr[6]), .Y(n49) );
endmodule


module watchdog_a0_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module watchdog_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer1_a0 ( clkper, rst, newinstr, t1ff, t1ack, int1ff, t1_tf1, t1ov, 
        sfrdatai, sfraddr, sfrwe, t1_tmod, t1_tr1, tl1, th1, test_si, test_se
 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t1_tmod;
  output [7:0] tl1;
  output [7:0] th1;
  input clkper, rst, newinstr, t1ff, t1ack, int1ff, sfrwe, test_si, test_se;
  output t1_tf1, t1ov, t1_tr1;
  wire   t1clr, th1_ov_ff, tl1_ov_ff, N31, N32, N33, N34, N35, N36, N37, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N95, N97, N98, clk_ov12, N100, net12182,
         net12188, net12193, n54, n55, n56, n57, n58, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n59, n60, n61, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19;
  wire   [1:0] t0_mode;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer1_a0_0 clk_gate_t1_mode_reg ( .CLK(clkper), .EN(
        N31), .ENCLK(net12182), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_2 clk_gate_tl1_s_reg ( .CLK(clkper), .EN(N50), 
        .ENCLK(net12188), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_1 clk_gate_th1_s_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12193), .TE(test_se) );
  timer1_a0_DW01_inc_0 add_278 ( .A(th1), .SUM({N75, N74, N73, N72, N71, N70, 
        N69, N68}) );
  timer1_a0_DW01_inc_1 add_244 ( .A(tl1), .SUM({N49, N48, N47, N46, N45, N44, 
        N43, N42}) );
  SDFFQX1 th1_ov_ff_reg ( .D(n55), .SIN(t1clr), .SMC(test_se), .C(clkper), .Q(
        th1_ov_ff) );
  SDFFQX1 tl1_ov_ff_reg ( .D(n56), .SIN(th1[7]), .SMC(test_se), .C(clkper), 
        .Q(tl1_ov_ff) );
  SDFFQX1 clk_count_reg_3_ ( .D(N98), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 clk_count_reg_2_ ( .D(N97), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 t1clr_reg ( .D(n57), .SIN(t1_tr1), .SMC(test_se), .C(clkper), .Q(
        t1clr) );
  SDFFQX1 clk_count_reg_1_ ( .D(n10), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 clk_count_reg_0_ ( .D(N95), .SIN(test_si), .SMC(test_se), .C(clkper), 
        .Q(clk_count[0]) );
  SDFFQX1 clk_ov12_reg ( .D(N100), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 t0_mode_reg_1_ ( .D(N37), .SIN(t0_mode[0]), .SMC(test_se), .C(
        net12182), .Q(t0_mode[1]) );
  SDFFQX1 t0_mode_reg_0_ ( .D(N36), .SIN(clk_ov12), .SMC(test_se), .C(net12182), .Q(t0_mode[0]) );
  SDFFQX1 t1_ct_reg ( .D(N33), .SIN(t0_mode[1]), .SMC(test_se), .C(net12182), 
        .Q(t1_tmod[2]) );
  SDFFQX1 t1_gate_reg ( .D(N32), .SIN(t1_tmod[2]), .SMC(test_se), .C(net12182), 
        .Q(t1_tmod[3]) );
  SDFFQX1 tl1_s_reg_7_ ( .D(N58), .SIN(tl1[6]), .SMC(test_se), .C(net12188), 
        .Q(tl1[7]) );
  SDFFQX1 tl1_s_reg_5_ ( .D(N56), .SIN(tl1[4]), .SMC(test_se), .C(net12188), 
        .Q(tl1[5]) );
  SDFFQX1 tl1_s_reg_4_ ( .D(N55), .SIN(tl1[3]), .SMC(test_se), .C(net12188), 
        .Q(tl1[4]) );
  SDFFQX1 th1_s_reg_7_ ( .D(N84), .SIN(th1[6]), .SMC(test_se), .C(net12193), 
        .Q(th1[7]) );
  SDFFQX1 tl1_s_reg_6_ ( .D(N57), .SIN(tl1[5]), .SMC(test_se), .C(net12188), 
        .Q(tl1[6]) );
  SDFFQX1 tl1_s_reg_1_ ( .D(N52), .SIN(tl1[0]), .SMC(test_se), .C(net12188), 
        .Q(tl1[1]) );
  SDFFQX1 th1_s_reg_3_ ( .D(N80), .SIN(th1[2]), .SMC(test_se), .C(net12193), 
        .Q(th1[3]) );
  SDFFQX1 th1_s_reg_6_ ( .D(N83), .SIN(th1[5]), .SMC(test_se), .C(net12193), 
        .Q(th1[6]) );
  SDFFQX1 th1_s_reg_5_ ( .D(N82), .SIN(th1[4]), .SMC(test_se), .C(net12193), 
        .Q(th1[5]) );
  SDFFQX1 th1_s_reg_4_ ( .D(N81), .SIN(th1[3]), .SMC(test_se), .C(net12193), 
        .Q(th1[4]) );
  SDFFQX1 tl1_s_reg_3_ ( .D(N54), .SIN(tl1[2]), .SMC(test_se), .C(net12188), 
        .Q(tl1[3]) );
  SDFFQX1 th1_s_reg_2_ ( .D(N79), .SIN(th1[1]), .SMC(test_se), .C(net12193), 
        .Q(th1[2]) );
  SDFFQX1 th1_s_reg_1_ ( .D(N78), .SIN(th1[0]), .SMC(test_se), .C(net12193), 
        .Q(th1[1]) );
  SDFFQX1 tl1_s_reg_0_ ( .D(N51), .SIN(tl1_ov_ff), .SMC(test_se), .C(net12188), 
        .Q(tl1[0]) );
  SDFFQX1 t1_mode_reg_1_ ( .D(N35), .SIN(t1_tmod[0]), .SMC(test_se), .C(
        net12182), .Q(t1_tmod[1]) );
  SDFFQX1 th1_s_reg_0_ ( .D(N77), .SIN(th1_ov_ff), .SMC(test_se), .C(net12193), 
        .Q(th1[0]) );
  SDFFQX1 tl1_s_reg_2_ ( .D(N53), .SIN(tl1[1]), .SMC(test_se), .C(net12188), 
        .Q(tl1[2]) );
  SDFFQX1 t1_mode_reg_0_ ( .D(N34), .SIN(t1_tmod[3]), .SMC(test_se), .C(
        net12182), .Q(t1_tmod[0]) );
  SDFFQX1 t1_tf1_s_reg ( .D(n54), .SIN(t1_tmod[1]), .SMC(test_se), .C(clkper), 
        .Q(t1_tf1) );
  SDFFQX1 t1_tr1_s_reg ( .D(n58), .SIN(t1_tf1), .SMC(test_se), .C(clkper), .Q(
        t1_tr1) );
  INVX1 U3 ( .A(n21), .Y(n8) );
  NAND32X1 U4 ( .B(sfraddr[0]), .C(sfraddr[1]), .A(n29), .Y(n21) );
  NAND3X1 U5 ( .A(sfraddr[0]), .B(n29), .C(sfraddr[1]), .Y(n49) );
  NAND21X1 U6 ( .B(n43), .A(n7), .Y(n41) );
  NOR2X1 U7 ( .A(n4), .B(n60), .Y(N35) );
  NOR2X1 U8 ( .A(n3), .B(n60), .Y(N34) );
  NOR2X1 U9 ( .A(n6), .B(n60), .Y(N32) );
  NOR2X1 U10 ( .A(n5), .B(n60), .Y(N33) );
  NOR2X1 U11 ( .A(n1), .B(n60), .Y(N36) );
  NOR2X1 U12 ( .A(n2), .B(n60), .Y(N37) );
  NAND2X1 U13 ( .A(n7), .B(n60), .Y(N31) );
  NOR43XL U14 ( .B(sfraddr[3]), .C(n61), .D(sfrwe), .A(sfraddr[2]), .Y(n29) );
  NOR3XL U15 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n61) );
  OR4X1 U16 ( .A(n47), .B(n46), .C(n48), .D(rst), .Y(N50) );
  NOR2X1 U17 ( .A(n49), .B(rst), .Y(n47) );
  NAND4X1 U18 ( .A(sfraddr[2]), .B(sfraddr[0]), .C(n44), .D(n45), .Y(n43) );
  NOR4XL U19 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[4]), .D(sfraddr[1]), 
        .Y(n45) );
  AND2X1 U20 ( .A(sfraddr[3]), .B(sfrwe), .Y(n44) );
  INVX1 U21 ( .A(n42), .Y(n9) );
  NAND3X1 U22 ( .A(n41), .B(n7), .C(n42), .Y(N76) );
  NAND42X1 U23 ( .C(sfraddr[1]), .D(rst), .A(sfraddr[0]), .B(n29), .Y(n60) );
  INVX1 U24 ( .A(sfrdatai[4]), .Y(n3) );
  INVX1 U25 ( .A(sfrdatai[5]), .Y(n4) );
  INVX1 U26 ( .A(sfrdatai[0]), .Y(n1) );
  INVX1 U27 ( .A(sfrdatai[1]), .Y(n2) );
  INVX1 U28 ( .A(sfrdatai[7]), .Y(n6) );
  INVX1 U29 ( .A(sfrdatai[6]), .Y(n5) );
  INVX1 U30 ( .A(rst), .Y(n7) );
  INVX1 U31 ( .A(n37), .Y(n11) );
  NOR42XL U32 ( .C(n31), .D(n49), .A(rst), .B(n50), .Y(n48) );
  NOR32XL U33 ( .B(n49), .C(n7), .A(n31), .Y(n46) );
  AO22AXL U34 ( .A(N70), .B(n9), .C(sfrdatai[2]), .D(n41), .Y(N79) );
  AO22AXL U35 ( .A(N71), .B(n9), .C(sfrdatai[3]), .D(n41), .Y(N80) );
  NAND4X1 U36 ( .A(n16), .B(n43), .C(n7), .D(n18), .Y(n42) );
  ENOX1 U37 ( .A(n41), .B(n2), .C(N69), .D(n9), .Y(N78) );
  ENOX1 U38 ( .A(n41), .B(n3), .C(N72), .D(n9), .Y(N81) );
  ENOX1 U39 ( .A(n41), .B(n4), .C(N73), .D(n9), .Y(N82) );
  ENOX1 U40 ( .A(n5), .B(n41), .C(N74), .D(n9), .Y(N83) );
  NAND21X1 U41 ( .B(newinstr), .A(n7), .Y(n22) );
  NAND2X1 U42 ( .A(n24), .B(n31), .Y(t1ov) );
  INVX1 U43 ( .A(n23), .Y(n16) );
  NAND2X1 U44 ( .A(n7), .B(n40), .Y(n37) );
  NAND2X1 U45 ( .A(n11), .B(n38), .Y(n35) );
  INVX1 U46 ( .A(n38), .Y(n12) );
  NOR2X1 U47 ( .A(rst), .B(n40), .Y(N100) );
  AO222X1 U48 ( .A(n46), .B(th1[0]), .C(n47), .D(sfrdatai[0]), .E(N42), .F(n48), .Y(N51) );
  AO222X1 U49 ( .A(n46), .B(th1[4]), .C(n47), .D(sfrdatai[4]), .E(N46), .F(n48), .Y(N55) );
  AO222X1 U50 ( .A(n46), .B(th1[2]), .C(n47), .D(sfrdatai[2]), .E(N44), .F(n48), .Y(N53) );
  AO222X1 U51 ( .A(n46), .B(th1[3]), .C(n47), .D(sfrdatai[3]), .E(N45), .F(n48), .Y(N54) );
  AO222X1 U52 ( .A(n46), .B(th1[1]), .C(n47), .D(sfrdatai[1]), .E(N43), .F(n48), .Y(N52) );
  AO222X1 U53 ( .A(n46), .B(th1[6]), .C(n47), .D(sfrdatai[6]), .E(N48), .F(n48), .Y(N57) );
  AO222X1 U54 ( .A(n46), .B(th1[5]), .C(n47), .D(sfrdatai[5]), .E(N47), .F(n48), .Y(N56) );
  AO222X1 U55 ( .A(n46), .B(th1[7]), .C(n47), .D(sfrdatai[7]), .E(N49), .F(n48), .Y(N58) );
  OR4X1 U56 ( .A(t1ack), .B(t1clr), .C(n8), .D(rst), .Y(n28) );
  OAI22BX1 U57 ( .B(n25), .A(n26), .D(t1_tf1), .C(n25), .Y(n54) );
  AOI31X1 U58 ( .A(n8), .B(n7), .C(sfrdatai[7]), .D(n27), .Y(n26) );
  GEN2XL U59 ( .D(th1_ov_ff), .E(n18), .C(n15), .B(n27), .A(n28), .Y(n25) );
  AOI21X1 U60 ( .B(t0_mode[0]), .C(t0_mode[1]), .A(n28), .Y(n27) );
  NOR2X1 U61 ( .A(rst), .B(n20), .Y(n58) );
  AOI22X1 U62 ( .A(sfrdatai[6]), .B(n8), .C(t1_tr1), .D(n21), .Y(n20) );
  ENOX1 U63 ( .A(n41), .B(n1), .C(N68), .D(n9), .Y(N77) );
  ENOX1 U64 ( .A(n6), .B(n41), .C(N75), .D(n9), .Y(N84) );
  AO22AXL U65 ( .A(t1ack), .B(n7), .C(t1clr), .D(n22), .Y(n57) );
  OAI22AX1 U66 ( .D(tl1_ov_ff), .C(n22), .A(rst), .B(n23), .Y(n56) );
  OAI22AX1 U67 ( .D(th1_ov_ff), .C(n22), .A(rst), .B(n24), .Y(n55) );
  NAND4X1 U68 ( .A(tl1[3]), .B(tl1[2]), .C(tl1[4]), .D(n51), .Y(n23) );
  NOR42XL U69 ( .C(tl1[1]), .D(tl1[0]), .A(n50), .B(n52), .Y(n51) );
  AOI32X1 U70 ( .A(tl1[6]), .B(tl1[5]), .C(tl1[7]), .D(n18), .E(n17), .Y(n52)
         );
  NAND2X1 U71 ( .A(n16), .B(t1_tmod[1]), .Y(n31) );
  OAI211X1 U72 ( .C(n17), .D(n18), .A(clk_ov12), .B(n53), .Y(n50) );
  AOI211X1 U73 ( .C(t1_tmod[3]), .D(n19), .A(t1_tmod[2]), .B(n59), .Y(n53) );
  INVX1 U74 ( .A(int1ff), .Y(n19) );
  AOI21X1 U75 ( .B(t0_mode[1]), .C(t0_mode[0]), .A(t1_tr1), .Y(n59) );
  NAND4X1 U76 ( .A(th1[2]), .B(th1[1]), .C(n32), .D(n33), .Y(n24) );
  NOR32XL U77 ( .B(th1[7]), .C(th1[6]), .A(n34), .Y(n33) );
  AND3X1 U78 ( .A(th1[0]), .B(n18), .C(n16), .Y(n32) );
  NAND3X1 U79 ( .A(th1[4]), .B(th1[3]), .C(th1[5]), .Y(n34) );
  INVX1 U80 ( .A(n30), .Y(n15) );
  AOI31X1 U81 ( .A(tl1_ov_ff), .B(n17), .C(t1_tmod[1]), .D(t1ov), .Y(n30) );
  INVX1 U82 ( .A(t1_tmod[1]), .Y(n18) );
  INVX1 U83 ( .A(t1_tmod[0]), .Y(n17) );
  NAND2X1 U84 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n38) );
  OAI32X1 U85 ( .A(n37), .B(clk_count[2]), .C(n38), .D(n13), .E(n35), .Y(N97)
         );
  OAI21X1 U86 ( .B(n14), .C(n35), .A(n36), .Y(N98) );
  NAND4X1 U87 ( .A(clk_count[2]), .B(n11), .C(n12), .D(n14), .Y(n36) );
  INVX1 U88 ( .A(clk_count[3]), .Y(n14) );
  NAND3X1 U89 ( .A(n12), .B(n13), .C(clk_count[3]), .Y(n40) );
  INVX1 U90 ( .A(clk_count[2]), .Y(n13) );
  NOR2X1 U91 ( .A(clk_count[0]), .B(n37), .Y(N95) );
  INVX1 U92 ( .A(n39), .Y(n10) );
  OAI211X1 U93 ( .C(clk_count[0]), .D(clk_count[1]), .A(n11), .B(n38), .Y(n39)
         );
endmodule


module timer1_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module timer1_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer0_a0 ( clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, t0_tf0, 
        t0_tf1, sfrdatai, sfraddr, sfrwe, t0_tmod, t0_tr0, t0_tr1, tl0, th0, 
        test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t0_tmod;
  output [7:0] tl0;
  output [7:0] th0;
  input clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, sfrwe, test_si,
         test_se;
  output t0_tf0, t0_tf1, t0_tr0, t0_tr1;
  wire   t0clr, th0_ov_ff, tl0_ov_ff, t1clr, N39, N40, N41, N42, N43, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N101, N103, N104, clk_ov12, N106, net12210,
         net12216, net12221, n60, n61, n62, n63, n64, n65, n66, n67, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n68, n69, n70, n71, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n72, n73, n74;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer0_a0_0 clk_gate_t0_ct_reg ( .CLK(clkper), .EN(N39), 
        .ENCLK(net12210), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_2 clk_gate_th0_s_reg ( .CLK(clkper), .EN(N55), 
        .ENCLK(net12216), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_1 clk_gate_tl0_s_reg ( .CLK(clkper), .EN(N79), 
        .ENCLK(net12221), .TE(test_se) );
  timer0_a0_DW01_inc_0 add_347 ( .A(tl0), .SUM({N78, N77, N76, N75, N74, N73, 
        N72, N71}) );
  timer0_a0_DW01_inc_1 add_309 ( .A(th0), .SUM({N54, N53, N52, N51, N50, N49, 
        N48, N47}) );
  SDFFQX1 th0_ov_ff_reg ( .D(n61), .SIN(t1clr), .SMC(test_se), .C(clkper), .Q(
        th0_ov_ff) );
  SDFFQX1 t1clr_reg ( .D(n63), .SIN(t0clr), .SMC(test_se), .C(clkper), .Q(
        t1clr) );
  SDFFQX1 tl0_ov_ff_reg ( .D(n64), .SIN(th0[7]), .SMC(test_se), .C(clkper), 
        .Q(tl0_ov_ff) );
  SDFFQX1 t0clr_reg ( .D(n65), .SIN(t0_tr1), .SMC(test_se), .C(clkper), .Q(
        t0clr) );
  SDFFQX1 clk_count_reg_3_ ( .D(N104), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 clk_count_reg_2_ ( .D(N103), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 clk_count_reg_1_ ( .D(n17), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 clk_count_reg_0_ ( .D(N101), .SIN(test_si), .SMC(test_se), .C(clkper), .Q(clk_count[0]) );
  SDFFQX1 clk_ov12_reg ( .D(N106), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 tl0_s_reg_7_ ( .D(N87), .SIN(tl0[6]), .SMC(test_se), .C(net12221), 
        .Q(tl0[7]) );
  SDFFQX1 tl0_s_reg_5_ ( .D(N85), .SIN(tl0[4]), .SMC(test_se), .C(net12221), 
        .Q(tl0[5]) );
  SDFFQX1 tl0_s_reg_6_ ( .D(N86), .SIN(tl0[5]), .SMC(test_se), .C(net12221), 
        .Q(tl0[6]) );
  SDFFQX1 tl0_s_reg_4_ ( .D(N84), .SIN(tl0[3]), .SMC(test_se), .C(net12221), 
        .Q(tl0[4]) );
  SDFFQX1 tl0_s_reg_1_ ( .D(N81), .SIN(tl0[0]), .SMC(test_se), .C(net12221), 
        .Q(tl0[1]) );
  SDFFQX1 th0_s_reg_7_ ( .D(N63), .SIN(th0[6]), .SMC(test_se), .C(net12216), 
        .Q(th0[7]) );
  SDFFQX1 t0_ct_reg ( .D(N41), .SIN(clk_ov12), .SMC(test_se), .C(net12210), 
        .Q(t0_tmod[2]) );
  SDFFQX1 t0_gate_reg ( .D(N40), .SIN(t0_tmod[2]), .SMC(test_se), .C(net12210), 
        .Q(t0_tmod[3]) );
  SDFFQX1 th0_s_reg_6_ ( .D(N62), .SIN(th0[5]), .SMC(test_se), .C(net12216), 
        .Q(th0[6]) );
  SDFFQX1 th0_s_reg_5_ ( .D(N61), .SIN(th0[4]), .SMC(test_se), .C(net12216), 
        .Q(th0[5]) );
  SDFFQX1 th0_s_reg_4_ ( .D(N60), .SIN(th0[3]), .SMC(test_se), .C(net12216), 
        .Q(th0[4]) );
  SDFFQX1 tl0_s_reg_3_ ( .D(N83), .SIN(tl0[2]), .SMC(test_se), .C(net12221), 
        .Q(tl0[3]) );
  SDFFQX1 th0_s_reg_1_ ( .D(N57), .SIN(th0[0]), .SMC(test_se), .C(net12216), 
        .Q(th0[1]) );
  SDFFQX1 th0_s_reg_3_ ( .D(N59), .SIN(th0[2]), .SMC(test_se), .C(net12216), 
        .Q(th0[3]) );
  SDFFQX1 th0_s_reg_2_ ( .D(N58), .SIN(th0[1]), .SMC(test_se), .C(net12216), 
        .Q(th0[2]) );
  SDFFQX1 t0_mode_reg_0_ ( .D(N42), .SIN(t0_tmod[3]), .SMC(test_se), .C(
        net12210), .Q(t0_tmod[0]) );
  SDFFQX1 tl0_s_reg_0_ ( .D(N80), .SIN(tl0_ov_ff), .SMC(test_se), .C(net12221), 
        .Q(tl0[0]) );
  SDFFQX1 th0_s_reg_0_ ( .D(N56), .SIN(th0_ov_ff), .SMC(test_se), .C(net12216), 
        .Q(th0[0]) );
  SDFFQX1 t0_mode_reg_1_ ( .D(N43), .SIN(t0_tmod[0]), .SMC(test_se), .C(
        net12210), .Q(t0_tmod[1]) );
  SDFFQX1 tl0_s_reg_2_ ( .D(N82), .SIN(tl0[1]), .SMC(test_se), .C(net12221), 
        .Q(tl0[2]) );
  SDFFQX1 t0_tf1_s_reg ( .D(n62), .SIN(t0_tf0), .SMC(test_se), .C(clkper), .Q(
        t0_tf1) );
  SDFFQX1 t0_tr0_s_reg ( .D(n67), .SIN(t0_tf1), .SMC(test_se), .C(clkper), .Q(
        t0_tr0) );
  SDFFQX1 t0_tr1_s_reg ( .D(n66), .SIN(t0_tr0), .SMC(test_se), .C(clkper), .Q(
        t0_tr1) );
  SDFFQX1 t0_tf0_s_reg ( .D(n60), .SIN(t0_tmod[1]), .SMC(test_se), .C(clkper), 
        .Q(t0_tf0) );
  INVX1 U3 ( .A(n31), .Y(n14) );
  INVX1 U4 ( .A(n2), .Y(n1) );
  NOR2X1 U5 ( .A(n29), .B(n11), .Y(n31) );
  NOR2X1 U6 ( .A(n46), .B(n11), .Y(n43) );
  NOR2X1 U7 ( .A(n31), .B(n11), .Y(n24) );
  INVX1 U8 ( .A(sfraddr[0]), .Y(n2) );
  NAND3X1 U9 ( .A(n40), .B(n2), .C(sfraddr[1]), .Y(n46) );
  NAND3X1 U10 ( .A(n2), .B(n3), .C(n40), .Y(n29) );
  OR2X1 U11 ( .A(n49), .B(n12), .Y(n48) );
  NAND4X1 U12 ( .A(n1), .B(n40), .C(n13), .D(n3), .Y(n56) );
  INVX1 U13 ( .A(sfraddr[1]), .Y(n3) );
  NOR2X1 U14 ( .A(n5), .B(n56), .Y(N43) );
  NOR2X1 U15 ( .A(n4), .B(n56), .Y(N42) );
  NOR2X1 U16 ( .A(n6), .B(n56), .Y(N41) );
  NOR2X1 U17 ( .A(n7), .B(n56), .Y(N40) );
  NAND2X1 U18 ( .A(n13), .B(n56), .Y(N39) );
  INVX1 U19 ( .A(n13), .Y(n11) );
  INVX1 U20 ( .A(n13), .Y(n12) );
  NOR43XL U21 ( .B(sfraddr[3]), .C(n57), .D(sfrwe), .A(sfraddr[2]), .Y(n40) );
  NOR3XL U22 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n57) );
  OR4X1 U23 ( .A(n43), .B(n41), .C(n42), .D(n11), .Y(N79) );
  NAND4X1 U24 ( .A(sfraddr[2]), .B(sfrwe), .C(n50), .D(n51), .Y(n49) );
  NOR21XL U25 ( .B(sfraddr[3]), .A(n1), .Y(n50) );
  NOR4XL U26 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[4]), .D(sfraddr[1]), 
        .Y(n51) );
  INVX1 U27 ( .A(n47), .Y(n15) );
  NAND3X1 U28 ( .A(n47), .B(n13), .C(n48), .Y(N55) );
  INVX1 U29 ( .A(sfrdatai[1]), .Y(n5) );
  INVX1 U30 ( .A(sfrdatai[2]), .Y(n6) );
  INVX1 U31 ( .A(sfrdatai[0]), .Y(n4) );
  INVX1 U32 ( .A(sfrdatai[3]), .Y(n7) );
  INVX1 U33 ( .A(sfrdatai[6]), .Y(n10) );
  INVX1 U34 ( .A(sfrdatai[4]), .Y(n8) );
  INVX1 U35 ( .A(sfrdatai[5]), .Y(n9) );
  INVX1 U36 ( .A(rst), .Y(n13) );
  INVX1 U37 ( .A(n69), .Y(n18) );
  NOR43XL U38 ( .B(n44), .C(n45), .D(n46), .A(n11), .Y(n42) );
  NOR32XL U39 ( .B(n46), .C(n13), .A(n45), .Y(n41) );
  NAND3X1 U40 ( .A(n39), .B(n13), .C(n49), .Y(n47) );
  ENOX1 U41 ( .A(n5), .B(n48), .C(N48), .D(n15), .Y(N57) );
  ENOX1 U42 ( .A(n10), .B(n48), .C(N53), .D(n15), .Y(N62) );
  ENOX1 U43 ( .A(n6), .B(n48), .C(N49), .D(n15), .Y(N58) );
  ENOX1 U44 ( .A(n7), .B(n48), .C(N50), .D(n15), .Y(N59) );
  ENOX1 U45 ( .A(n8), .B(n48), .C(N51), .D(n15), .Y(N60) );
  ENOX1 U46 ( .A(n9), .B(n48), .C(N52), .D(n15), .Y(N61) );
  OAI22X1 U47 ( .A(n11), .B(n16), .C(n25), .D(n22), .Y(n65) );
  OAI22X1 U48 ( .A(n11), .B(n26), .C(n25), .D(n20), .Y(n64) );
  OR2X1 U49 ( .A(newinstr), .B(n12), .Y(n25) );
  INVX1 U50 ( .A(t0ack), .Y(n16) );
  NAND2X1 U51 ( .A(n13), .B(n58), .Y(n69) );
  NAND2X1 U52 ( .A(n18), .B(n70), .Y(n59) );
  INVX1 U53 ( .A(n70), .Y(n19) );
  NOR2X1 U54 ( .A(n11), .B(n58), .Y(N106) );
  AO222X1 U55 ( .A(n41), .B(th0[0]), .C(N71), .D(n42), .E(sfrdatai[0]), .F(n43), .Y(N80) );
  AO222X1 U56 ( .A(n41), .B(th0[2]), .C(N73), .D(n42), .E(sfrdatai[2]), .F(n43), .Y(N82) );
  AO222X1 U57 ( .A(n41), .B(th0[4]), .C(N75), .D(n42), .E(n43), .F(sfrdatai[4]), .Y(N84) );
  AO222X1 U58 ( .A(n41), .B(th0[3]), .C(N74), .D(n42), .E(sfrdatai[3]), .F(n43), .Y(N83) );
  AO222X1 U59 ( .A(n41), .B(th0[1]), .C(N72), .D(n42), .E(sfrdatai[1]), .F(n43), .Y(N81) );
  AO222X1 U60 ( .A(n41), .B(th0[6]), .C(N77), .D(n42), .E(n43), .F(sfrdatai[6]), .Y(N86) );
  AO222X1 U61 ( .A(n41), .B(th0[5]), .C(N76), .D(n42), .E(n43), .F(sfrdatai[5]), .Y(N85) );
  AO222X1 U62 ( .A(n41), .B(th0[7]), .C(N78), .D(n42), .E(n43), .F(sfrdatai[7]), .Y(N87) );
  OAI22BX1 U63 ( .B(n27), .A(n28), .D(t0_tf1), .C(n27), .Y(n62) );
  AOI32X1 U64 ( .A(n29), .B(n13), .C(n30), .D(sfrdatai[7]), .E(n31), .Y(n28)
         );
  OAI211X1 U65 ( .C(n74), .D(n32), .A(n24), .B(n30), .Y(n27) );
  NOR2X1 U66 ( .A(t1clr), .B(t1ack), .Y(n30) );
  OAI211X1 U67 ( .C(n14), .D(n9), .A(n33), .B(n34), .Y(n60) );
  NAND4X1 U68 ( .A(t0_tf0), .B(n24), .C(n16), .D(n22), .Y(n33) );
  NAND4X1 U69 ( .A(n16), .B(n22), .C(n13), .D(n35), .Y(n34) );
  AOI31X1 U70 ( .A(n26), .B(n20), .C(t0_tmod[1]), .D(n36), .Y(n35) );
  OAI31XL U71 ( .A(n72), .B(th0_ov_ff), .C(t0_tmod[1]), .D(n29), .Y(n36) );
  INVX1 U72 ( .A(n32), .Y(n72) );
  OAI22BX1 U73 ( .B(N54), .A(n47), .D(sfrdatai[7]), .C(n48), .Y(N63) );
  ENOX1 U74 ( .A(n14), .B(n8), .C(n24), .D(t0_tr0), .Y(n67) );
  ENOX1 U75 ( .A(n14), .B(n10), .C(n24), .D(t0_tr1), .Y(n66) );
  ENOX1 U76 ( .A(n4), .B(n48), .C(N47), .D(n15), .Y(N56) );
  OAI22BX1 U77 ( .B(t1ack), .A(n11), .D(t1clr), .C(n25), .Y(n63) );
  OAI22AX1 U78 ( .D(th0_ov_ff), .C(n25), .A(n11), .B(n32), .Y(n61) );
  NOR43XL U79 ( .B(t0_tr0), .C(n55), .D(clk_ov12), .A(t0_tmod[2]), .Y(n44) );
  NAND21X1 U80 ( .B(int0ff), .A(t0_tmod[3]), .Y(n55) );
  NAND4X1 U81 ( .A(th0[3]), .B(th0[2]), .C(n37), .D(n38), .Y(n32) );
  AND4X1 U82 ( .A(th0[4]), .B(th0[5]), .C(th0[6]), .D(th0[7]), .Y(n38) );
  AND3X1 U83 ( .A(th0[1]), .B(n39), .C(th0[0]), .Y(n37) );
  OAI21X1 U84 ( .B(t0_tmod[1]), .C(n26), .A(n52), .Y(n39) );
  NAND4X1 U85 ( .A(t0_tmod[1]), .B(t0_tmod[0]), .C(clk_ov12), .D(t0_tr1), .Y(
        n52) );
  NAND4X1 U86 ( .A(tl0[3]), .B(tl0[2]), .C(tl0[4]), .D(n53), .Y(n26) );
  NOR43XL U87 ( .B(tl0[1]), .C(tl0[0]), .D(n44), .A(n54), .Y(n53) );
  AOI32X1 U88 ( .A(tl0[6]), .B(tl0[5]), .C(tl0[7]), .D(n74), .E(n73), .Y(n54)
         );
  INVX1 U89 ( .A(t0_tmod[1]), .Y(n74) );
  INVX1 U90 ( .A(t0_tmod[0]), .Y(n73) );
  NAND31X1 U91 ( .C(n26), .A(n73), .B(t0_tmod[1]), .Y(n45) );
  NAND2X1 U92 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n70) );
  OAI32X1 U93 ( .A(n69), .B(clk_count[2]), .C(n70), .D(n21), .E(n59), .Y(N103)
         );
  NAND3X1 U94 ( .A(n19), .B(n21), .C(clk_count[3]), .Y(n58) );
  OAI21X1 U95 ( .B(n23), .C(n59), .A(n68), .Y(N104) );
  NAND4X1 U96 ( .A(clk_count[2]), .B(n18), .C(n19), .D(n23), .Y(n68) );
  INVX1 U97 ( .A(clk_count[3]), .Y(n23) );
  INVX1 U98 ( .A(t0clr), .Y(n22) );
  INVX1 U99 ( .A(clk_count[2]), .Y(n21) );
  NOR2X1 U100 ( .A(clk_count[0]), .B(n69), .Y(N101) );
  INVX1 U101 ( .A(n71), .Y(n17) );
  OAI211X1 U102 ( .C(clk_count[0]), .D(clk_count[1]), .A(n18), .B(n70), .Y(n71) );
  INVX1 U103 ( .A(tl0_ov_ff), .Y(n20) );
endmodule


module timer0_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module timer0_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module serial0_a0 ( t_shift_clk, r_shift_clk, clkper, rst, newinstr, rxd0ff, 
        t1ov, rxd0o, rxd0oe, txd0, sfrdatai, sfraddr, sfrwe, s0con, s0buf, 
        s0rell, s0relh, smod, bd, test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] s0con;
  output [7:0] s0buf;
  output [7:0] s0rell;
  output [7:0] s0relh;
  input clkper, rst, newinstr, rxd0ff, t1ov, sfrwe, test_si, test_se;
  output t_shift_clk, r_shift_clk, rxd0o, rxd0oe, txd0, smod, bd;
  wire   r_clk_ov2, t1ov_ff, N59, ri_tmp, rxd0_val, s0con2_val, s0con2_tmp,
         ti_tmp, N108, N109, N110, N111, N112, N113, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, baud_rate_ov, N142, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N166, N169, N170, N185, N186, N187,
         N188, N190, clk_ov12, N191, r_start, baud_r_count, baud_r2_clk, N207,
         t_baud_ov, t_start, N223, N224, N225, N226, N227, N230, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N281,
         N282, N283, N284, N303, rxd0_fall, rxd0_ff, rxd0_fall_fl,
         receive_11_bits, N306, N307, N324, N325, N326, N327, N333, ri0_fall,
         ri0_ff, N348, N360, N361, N362, N363, N364, N375, N376, N377, N378,
         N379, N380, N381, N382, N424, N425, N426, N427, N428, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, net12249, net12255,
         net12260, net12265, net12270, net12275, net12280, net12285, net12290,
         net12295, net12300, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n245, n27, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n244;
  wire   [3:0] r_baud_count;
  wire   [3:0] r_shift_count;
  wire   [3:0] t_shift_count;
  wire   [9:0] tim_baud;
  wire   [3:0] clk_count;
  wire   [3:0] t_baud_count;
  wire   [10:0] t_shift_reg;
  wire   [1:0] fluctuation_conter;
  wire   [2:0] rxd0_vec;
  wire   [7:0] r_shift_reg;

  MAJ3X1 U329 ( .A(rxd0_vec[1]), .B(rxd0_vec[0]), .C(rxd0_vec[2]), .Y(n173) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_0 clk_gate_s0con_s_reg ( .CLK(clkper), .EN(
        N108), .ENCLK(net12249), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_10 clk_gate_s0rell_s_reg ( .CLK(clkper), 
        .EN(N117), .ENCLK(net12255), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_9 clk_gate_s0relh_s_reg ( .CLK(clkper), .EN(
        N128), .ENCLK(net12260), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_8 clk_gate_tim_baud_reg ( .CLK(clkper), .EN(
        N166), .ENCLK(net12265), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_7 clk_gate_t_baud_count_reg ( .CLK(clkper), 
        .EN(N223), .ENCLK(net12270), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_6 clk_gate_t_shift_reg_reg ( .CLK(clkper), 
        .EN(N257), .ENCLK(net12275), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_5 clk_gate_rxd0_vec_reg ( .CLK(clkper), .EN(
        N324), .ENCLK(net12280), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_4 clk_gate_r_baud_count_reg ( .CLK(clkper), 
        .EN(N360), .ENCLK(net12285), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_3 clk_gate_r_shift_reg_reg ( .CLK(clkper), 
        .EN(n27), .ENCLK(net12290), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_2 clk_gate_r_shift_count_reg ( .CLK(clkper), 
        .EN(N428), .ENCLK(net12295), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_1 clk_gate_s0buf_r_reg ( .CLK(clkper), .EN(
        N471), .ENCLK(net12300), .TE(test_se) );
  serial0_a0_DW01_inc_0 add_584 ( .A(tim_baud), .SUM({N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145}) );
  SDFFQX1 t_shift_reg_reg_10_ ( .D(N268), .SIN(t_shift_reg[9]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[10]) );
  SDFFQX1 r_shift_reg_reg_0_ ( .D(N375), .SIN(r_shift_count[3]), .SMC(test_se), 
        .C(net12290), .Q(r_shift_reg[0]) );
  SDFFQX1 t_shift_reg_reg_1_ ( .D(N259), .SIN(t_shift_reg[0]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[1]) );
  SDFFQX1 ti_tmp_reg ( .D(n242), .SIN(t_start), .SMC(test_se), .C(clkper), .Q(
        ti_tmp) );
  SDFFQX1 ri_tmp_reg ( .D(n238), .SIN(ri0_ff), .SMC(test_se), .C(clkper), .Q(
        ri_tmp) );
  SDFFQX1 t_shift_reg_reg_2_ ( .D(N260), .SIN(t_shift_reg[1]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[2]) );
  SDFFQX1 t_baud_count_reg_3_ ( .D(N227), .SIN(t_baud_count[2]), .SMC(test_se), 
        .C(net12270), .Q(t_baud_count[3]) );
  SDFFQX1 t_shift_reg_reg_0_ ( .D(N258), .SIN(t_shift_count[3]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[0]) );
  SDFFQX1 baud_r_count_reg ( .D(n245), .SIN(baud_r2_clk), .SMC(test_se), .C(
        clkper), .Q(baud_r_count) );
  SDFFQX1 r_shift_reg_reg_7_ ( .D(N382), .SIN(r_shift_reg[6]), .SMC(test_se), 
        .C(net12290), .Q(r_shift_reg[7]) );
  SDFFQX1 r_shift_reg_reg_6_ ( .D(N381), .SIN(r_shift_reg[5]), .SMC(test_se), 
        .C(net12290), .Q(r_shift_reg[6]) );
  SDFFQX1 r_shift_reg_reg_5_ ( .D(N380), .SIN(r_shift_reg[4]), .SMC(test_se), 
        .C(net12290), .Q(r_shift_reg[5]) );
  SDFFQX1 r_shift_reg_reg_4_ ( .D(N379), .SIN(r_shift_reg[3]), .SMC(test_se), 
        .C(net12290), .Q(r_shift_reg[4]) );
  SDFFQX1 r_shift_reg_reg_3_ ( .D(N378), .SIN(r_shift_reg[2]), .SMC(test_se), 
        .C(net12290), .Q(r_shift_reg[3]) );
  SDFFQX1 r_shift_reg_reg_2_ ( .D(N377), .SIN(r_shift_reg[1]), .SMC(test_se), 
        .C(net12290), .Q(r_shift_reg[2]) );
  SDFFQX1 r_shift_reg_reg_1_ ( .D(N376), .SIN(r_shift_reg[0]), .SMC(test_se), 
        .C(net12290), .Q(r_shift_reg[1]) );
  SDFFQX1 fluctuation_conter_reg_1_ ( .D(n233), .SIN(fluctuation_conter[0]), 
        .SMC(test_se), .C(clkper), .Q(fluctuation_conter[1]) );
  SDFFQX1 t_shift_reg_reg_9_ ( .D(N267), .SIN(t_shift_reg[8]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[9]) );
  SDFFQX1 t_shift_reg_reg_8_ ( .D(N266), .SIN(t_shift_reg[7]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[8]) );
  SDFFQX1 t_shift_reg_reg_7_ ( .D(N265), .SIN(t_shift_reg[6]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[7]) );
  SDFFQX1 t_shift_reg_reg_6_ ( .D(N264), .SIN(t_shift_reg[5]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[6]) );
  SDFFQX1 t_shift_reg_reg_5_ ( .D(N263), .SIN(t_shift_reg[4]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[5]) );
  SDFFQX1 t_shift_reg_reg_4_ ( .D(N262), .SIN(t_shift_reg[3]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[4]) );
  SDFFQX1 t_shift_reg_reg_3_ ( .D(N261), .SIN(t_shift_reg[2]), .SMC(test_se), 
        .C(net12275), .Q(t_shift_reg[3]) );
  SDFFQX1 rxd0_vec_reg_2_ ( .D(N327), .SIN(rxd0_vec[1]), .SMC(test_se), .C(
        net12280), .Q(rxd0_vec[2]) );
  SDFFQX1 rxd0_vec_reg_1_ ( .D(N326), .SIN(rxd0_vec[0]), .SMC(test_se), .C(
        net12280), .Q(rxd0_vec[1]) );
  SDFFQX1 rxd0_fall_fl_reg ( .D(n235), .SIN(ri_tmp), .SMC(test_se), .C(clkper), 
        .Q(rxd0_fall_fl) );
  SDFFQX1 rxd0_ff_reg ( .D(N307), .SIN(rxd0_fall), .SMC(test_se), .C(clkper), 
        .Q(rxd0_ff) );
  SDFFQX1 rxd0_vec_reg_0_ ( .D(N325), .SIN(rxd0_val), .SMC(test_se), .C(
        net12280), .Q(rxd0_vec[0]) );
  SDFFQX1 receive_11_bits_reg ( .D(n229), .SIN(r_start), .SMC(test_se), .C(
        clkper), .Q(receive_11_bits) );
  SDFFQX1 t_shift_count_reg_3_ ( .D(N284), .SIN(t_shift_count[2]), .SMC(
        test_se), .C(net12275), .Q(t_shift_count[3]) );
  SDFFQX1 fluctuation_conter_reg_0_ ( .D(n234), .SIN(clk_ov12), .SMC(test_se), 
        .C(clkper), .Q(fluctuation_conter[0]) );
  SDFFQX1 clk_count_reg_3_ ( .D(N188), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 s0con2_val_reg ( .D(n231), .SIN(s0con2_tmp), .SMC(test_se), .C(
        net12280), .Q(s0con2_val) );
  SDFFQX1 s0con2_tmp_reg ( .D(n232), .SIN(s0buf[7]), .SMC(test_se), .C(clkper), 
        .Q(s0con2_tmp) );
  SDFFQX1 clk_count_reg_2_ ( .D(N187), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 ri0_ff_reg ( .D(N348), .SIN(ri0_fall), .SMC(test_se), .C(clkper), 
        .Q(ri0_ff) );
  SDFFQX1 clk_ov12_reg ( .D(N191), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 t_baud_ov_reg ( .D(N230), .SIN(t_baud_count[3]), .SMC(test_se), .C(
        clkper), .Q(t_baud_ov) );
  SDFFQX1 tim_baud_reg_9_ ( .D(n68), .SIN(tim_baud[8]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[9]) );
  SDFFQX1 tim_baud_reg_8_ ( .D(n75), .SIN(tim_baud[7]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[8]) );
  SDFFQX1 tim_baud_reg_4_ ( .D(n71), .SIN(tim_baud[3]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[4]) );
  SDFFQX1 t_shift_count_reg_1_ ( .D(N282), .SIN(t_shift_count[0]), .SMC(
        test_se), .C(net12275), .Q(t_shift_count[1]) );
  SDFFQX1 t_shift_count_reg_2_ ( .D(N283), .SIN(t_shift_count[1]), .SMC(
        test_se), .C(net12275), .Q(t_shift_count[2]) );
  SDFFQX1 t_shift_count_reg_0_ ( .D(N281), .SIN(t_baud_ov), .SMC(test_se), .C(
        net12275), .Q(t_shift_count[0]) );
  SDFFQX1 ri0_fall_reg ( .D(n236), .SIN(receive_11_bits), .SMC(test_se), .C(
        clkper), .Q(ri0_fall) );
  SDFFQX1 rxd0_val_reg ( .D(N333), .SIN(rxd0_ff), .SMC(test_se), .C(clkper), 
        .Q(rxd0_val) );
  SDFFQX1 t_baud_count_reg_1_ ( .D(N225), .SIN(t_baud_count[0]), .SMC(test_se), 
        .C(net12270), .Q(t_baud_count[1]) );
  SDFFQX1 t_baud_count_reg_2_ ( .D(N226), .SIN(t_baud_count[1]), .SMC(test_se), 
        .C(net12270), .Q(t_baud_count[2]) );
  SDFFQX1 clk_count_reg_1_ ( .D(N186), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 t_baud_count_reg_0_ ( .D(N224), .SIN(t1ov_ff), .SMC(test_se), .C(
        net12270), .Q(t_baud_count[0]) );
  SDFFQX1 r_start_reg ( .D(n240), .SIN(r_shift_reg[7]), .SMC(test_se), .C(
        clkper), .Q(r_start) );
  SDFFQX1 clk_count_reg_0_ ( .D(N185), .SIN(bd), .SMC(test_se), .C(clkper), 
        .Q(clk_count[0]) );
  SDFFQX1 rxd0_fall_reg ( .D(N306), .SIN(rxd0_fall_fl), .SMC(test_se), .C(
        clkper), .Q(rxd0_fall) );
  SDFFQX1 baud_r2_clk_reg ( .D(N207), .SIN(test_si), .SMC(test_se), .C(clkper), 
        .Q(baud_r2_clk) );
  SDFFQX1 tim_baud_reg_2_ ( .D(N169), .SIN(tim_baud[1]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[2]) );
  SDFFQX1 tim_baud_reg_7_ ( .D(n74), .SIN(tim_baud[6]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[7]) );
  SDFFQX1 tim_baud_reg_5_ ( .D(n72), .SIN(tim_baud[4]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[5]) );
  SDFFQX1 tim_baud_reg_1_ ( .D(n70), .SIN(tim_baud[0]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[1]) );
  SDFFQX1 tim_baud_reg_6_ ( .D(n73), .SIN(tim_baud[5]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[6]) );
  SDFFQX1 tim_baud_reg_3_ ( .D(N170), .SIN(tim_baud[2]), .SMC(test_se), .C(
        net12265), .Q(tim_baud[3]) );
  SDFFQX1 r_shift_count_reg_1_ ( .D(N425), .SIN(r_shift_count[0]), .SMC(
        test_se), .C(net12295), .Q(r_shift_count[1]) );
  SDFFQX1 r_shift_count_reg_3_ ( .D(N427), .SIN(r_shift_count[2]), .SMC(
        test_se), .C(net12295), .Q(r_shift_count[3]) );
  SDFFQX1 r_baud_count_reg_1_ ( .D(N362), .SIN(r_baud_count[0]), .SMC(test_se), 
        .C(net12285), .Q(r_baud_count[1]) );
  SDFFQX1 r_shift_count_reg_2_ ( .D(N426), .SIN(r_shift_count[1]), .SMC(
        test_se), .C(net12295), .Q(r_shift_count[2]) );
  SDFFQX1 r_shift_count_reg_0_ ( .D(N424), .SIN(r_clk_ov2), .SMC(test_se), .C(
        net12295), .Q(r_shift_count[0]) );
  SDFFQX1 r_baud_count_reg_3_ ( .D(N364), .SIN(r_baud_count[2]), .SMC(test_se), 
        .C(net12285), .Q(r_baud_count[3]) );
  SDFFQX1 r_baud_count_reg_2_ ( .D(N363), .SIN(r_baud_count[1]), .SMC(test_se), 
        .C(net12285), .Q(r_baud_count[2]) );
  SDFFQX1 tim_baud_reg_0_ ( .D(n69), .SIN(ti_tmp), .SMC(test_se), .C(net12265), 
        .Q(tim_baud[0]) );
  SDFFQX1 r_baud_count_reg_0_ ( .D(N361), .SIN(fluctuation_conter[1]), .SMC(
        test_se), .C(net12285), .Q(r_baud_count[0]) );
  SDFFQX1 t1ov_ff_reg ( .D(N59), .SIN(smod), .SMC(test_se), .C(clkper), .Q(
        t1ov_ff) );
  SDFFQX1 baud_rate_ov_reg ( .D(N142), .SIN(baud_r_count), .SMC(test_se), .C(
        clkper), .Q(baud_rate_ov) );
  SDFFQX1 r_clk_ov2_reg ( .D(N190), .SIN(r_baud_count[3]), .SMC(test_se), .C(
        clkper), .Q(r_clk_ov2) );
  SDFFQX1 s0relh_s_reg_3_ ( .D(N132), .SIN(s0relh[2]), .SMC(test_se), .C(
        net12260), .Q(s0relh[3]) );
  SDFFQX1 s0rell_s_reg_3_ ( .D(N121), .SIN(s0rell[2]), .SMC(test_se), .C(
        net12255), .Q(s0rell[3]) );
  SDFFQX1 s0rell_s_reg_7_ ( .D(N125), .SIN(s0rell[6]), .SMC(test_se), .C(
        net12255), .Q(s0rell[7]) );
  SDFFQX1 s0rell_s_reg_6_ ( .D(N124), .SIN(s0rell[5]), .SMC(test_se), .C(
        net12255), .Q(s0rell[6]) );
  SDFFQX1 s0rell_s_reg_0_ ( .D(N118), .SIN(s0relh[7]), .SMC(test_se), .C(
        net12255), .Q(s0rell[0]) );
  SDFFQX1 s0relh_s_reg_0_ ( .D(N129), .SIN(s0con[7]), .SMC(test_se), .C(
        net12260), .Q(s0relh[0]) );
  SDFFQX1 s0buf_r_reg_7_ ( .D(N479), .SIN(s0buf[6]), .SMC(test_se), .C(
        net12300), .Q(s0buf[7]) );
  SDFFQX1 s0buf_r_reg_6_ ( .D(N478), .SIN(s0buf[5]), .SMC(test_se), .C(
        net12300), .Q(s0buf[6]) );
  SDFFQX1 s0buf_r_reg_3_ ( .D(N475), .SIN(s0buf[2]), .SMC(test_se), .C(
        net12300), .Q(s0buf[3]) );
  SDFFQX1 s0buf_r_reg_0_ ( .D(N472), .SIN(rxd0o), .SMC(test_se), .C(net12300), 
        .Q(s0buf[0]) );
  SDFFQX1 s0relh_s_reg_4_ ( .D(N133), .SIN(s0relh[3]), .SMC(test_se), .C(
        net12260), .Q(s0relh[4]) );
  SDFFQX1 s0relh_s_reg_5_ ( .D(N134), .SIN(s0relh[4]), .SMC(test_se), .C(
        net12260), .Q(s0relh[5]) );
  SDFFQX1 s0relh_s_reg_2_ ( .D(N131), .SIN(s0relh[1]), .SMC(test_se), .C(
        net12260), .Q(s0relh[2]) );
  SDFFQX1 s0buf_r_reg_5_ ( .D(N477), .SIN(s0buf[4]), .SMC(test_se), .C(
        net12300), .Q(s0buf[5]) );
  SDFFQX1 s0con_s_reg_3_ ( .D(N109), .SIN(s0con[2]), .SMC(test_se), .C(
        net12249), .Q(s0con[3]) );
  SDFFQX1 s0rell_s_reg_2_ ( .D(N120), .SIN(s0rell[1]), .SMC(test_se), .C(
        net12255), .Q(s0rell[2]) );
  SDFFQX1 s0rell_s_reg_5_ ( .D(N123), .SIN(s0rell[4]), .SMC(test_se), .C(
        net12255), .Q(s0rell[5]) );
  SDFFQX1 s0rell_s_reg_4_ ( .D(N122), .SIN(s0rell[3]), .SMC(test_se), .C(
        net12255), .Q(s0rell[4]) );
  SDFFQX1 s0rell_s_reg_1_ ( .D(N119), .SIN(s0rell[0]), .SMC(test_se), .C(
        net12255), .Q(s0rell[1]) );
  SDFFQX1 s0relh_s_reg_1_ ( .D(N130), .SIN(s0relh[0]), .SMC(test_se), .C(
        net12260), .Q(s0relh[1]) );
  SDFFQX1 s0con_s_reg_5_ ( .D(N111), .SIN(s0con[4]), .SMC(test_se), .C(
        net12249), .Q(s0con[5]) );
  SDFFQX1 smod_s_reg ( .D(n29), .SIN(s0rell[7]), .SMC(test_se), .C(clkper), 
        .Q(smod) );
  SDFFQX1 bd_s_reg ( .D(n30), .SIN(baud_rate_ov), .SMC(test_se), .C(clkper), 
        .Q(bd) );
  SDFFQX1 s0con_s_reg_0_ ( .D(n237), .SIN(s0con2_val), .SMC(test_se), .C(
        clkper), .Q(s0con[0]) );
  SDFFQX1 s0con_s_reg_4_ ( .D(N110), .SIN(s0con[3]), .SMC(test_se), .C(
        net12249), .Q(s0con[4]) );
  SDFFQX1 s0relh_s_reg_7_ ( .D(N136), .SIN(s0relh[6]), .SMC(test_se), .C(
        net12260), .Q(s0relh[7]) );
  SDFFQX1 s0relh_s_reg_6_ ( .D(N135), .SIN(s0relh[5]), .SMC(test_se), .C(
        net12260), .Q(s0relh[6]) );
  SDFFQX1 s0buf_r_reg_2_ ( .D(N474), .SIN(s0buf[1]), .SMC(test_se), .C(
        net12300), .Q(s0buf[2]) );
  SDFFQX1 s0buf_r_reg_1_ ( .D(N473), .SIN(s0buf[0]), .SMC(test_se), .C(
        net12300), .Q(s0buf[1]) );
  SDFFQX1 s0buf_r_reg_4_ ( .D(N476), .SIN(s0buf[3]), .SMC(test_se), .C(
        net12300), .Q(s0buf[4]) );
  SDFFQX1 s0con_s_reg_2_ ( .D(n230), .SIN(s0con[1]), .SMC(test_se), .C(clkper), 
        .Q(s0con[2]) );
  SDFFQX1 s0con_s_reg_1_ ( .D(n241), .SIN(s0con[0]), .SMC(test_se), .C(clkper), 
        .Q(s0con[1]) );
  SDFFQX1 t_start_reg ( .D(n243), .SIN(t_shift_reg[10]), .SMC(test_se), .C(
        clkper), .Q(t_start) );
  SDFFQX1 s0con_s_reg_6_ ( .D(N112), .SIN(s0con[5]), .SMC(test_se), .C(
        net12249), .Q(s0con[6]) );
  SDFFQX1 s0con_s_reg_7_ ( .D(N113), .SIN(s0con[6]), .SMC(test_se), .C(
        net12249), .Q(s0con[7]) );
  SDFFQX1 rxd0o_reg ( .D(N303), .SIN(rxd0_vec[2]), .SMC(test_se), .C(clkper), 
        .Q(rxd0o) );
  SDFFQX1 txd0_reg ( .D(n239), .SIN(tim_baud[9]), .SMC(test_se), .C(clkper), 
        .Q(txd0) );
  BUFX3 U3 ( .A(n84), .Y(n1) );
  BUFX3 U4 ( .A(n83), .Y(n2) );
  NAND2X1 U5 ( .A(n228), .B(n227), .Y(n3) );
  INVXL U6 ( .A(sfraddr[6]), .Y(n8) );
  AOI221XL U7 ( .A(r_start), .B(n114), .C(n3), .D(r_shift_clk), .E(n22), .Y(
        n81) );
  INVX1 U8 ( .A(N108), .Y(n33) );
  INVX1 U9 ( .A(n181), .Y(n36) );
  NOR2X1 U10 ( .A(n193), .B(n21), .Y(n181) );
  NAND2X1 U11 ( .A(n17), .B(n131), .Y(N108) );
  INVX1 U12 ( .A(n183), .Y(n37) );
  NAND2X1 U13 ( .A(n17), .B(n214), .Y(N117) );
  NAND2X1 U14 ( .A(n18), .B(n212), .Y(N128) );
  INVX1 U15 ( .A(n131), .Y(n32) );
  NOR32XL U16 ( .B(n19), .C(sfraddr[1]), .A(n7), .Y(n100) );
  INVX1 U17 ( .A(n23), .Y(n19) );
  INVX1 U18 ( .A(n23), .Y(n17) );
  INVX1 U19 ( .A(n22), .Y(n20) );
  INVX1 U20 ( .A(n24), .Y(n18) );
  NAND4X1 U21 ( .A(n94), .B(n95), .C(n17), .D(n8), .Y(n131) );
  NOR4XL U22 ( .A(n35), .B(n4), .C(sfraddr[0]), .D(sfraddr[2]), .Y(n94) );
  NAND2X1 U23 ( .A(n181), .B(n226), .Y(n183) );
  NAND4X1 U24 ( .A(n95), .B(sfrwe), .C(sfraddr[0]), .D(n194), .Y(n193) );
  NOR3XL U25 ( .A(n4), .B(n7), .C(sfraddr[2]), .Y(n194) );
  INVX1 U26 ( .A(sfrwe), .Y(n35) );
  NAND2X1 U27 ( .A(n213), .B(n5), .Y(n212) );
  NAND2X1 U28 ( .A(n213), .B(n6), .Y(n214) );
  AOI31X1 U29 ( .A(n94), .B(n8), .C(n95), .D(n24), .Y(n107) );
  INVX1 U30 ( .A(n176), .Y(n39) );
  OAI21X1 U31 ( .B(n131), .C(n15), .A(n20), .Y(N112) );
  OAI21X1 U32 ( .B(n15), .C(n214), .A(n20), .Y(N124) );
  OAI21X1 U33 ( .B(n13), .C(n214), .A(n20), .Y(N122) );
  OAI21X1 U34 ( .B(n16), .C(n214), .A(n20), .Y(N125) );
  OAI21X1 U35 ( .B(n9), .C(n214), .A(n25), .Y(N118) );
  OAI21X1 U36 ( .B(n12), .C(n214), .A(n25), .Y(N121) );
  OAI21X1 U37 ( .B(n9), .C(n212), .A(n20), .Y(N129) );
  OAI21X1 U38 ( .B(n10), .C(n212), .A(n20), .Y(N130) );
  NOR2X1 U39 ( .A(n131), .B(n13), .Y(N110) );
  NOR2X1 U40 ( .A(n131), .B(n12), .Y(N109) );
  NOR2X1 U41 ( .A(n131), .B(n14), .Y(N111) );
  NOR2X1 U42 ( .A(n14), .B(n214), .Y(N123) );
  NOR2X1 U43 ( .A(n11), .B(n214), .Y(N120) );
  NOR2X1 U44 ( .A(n10), .B(n214), .Y(N119) );
  NOR2X1 U45 ( .A(n15), .B(n212), .Y(N135) );
  NOR2X1 U46 ( .A(n16), .B(n212), .Y(N136) );
  NOR2X1 U47 ( .A(n11), .B(n212), .Y(N131) );
  NOR2X1 U48 ( .A(n12), .B(n212), .Y(N132) );
  NOR2X1 U49 ( .A(n14), .B(n212), .Y(N134) );
  NOR2X1 U50 ( .A(n13), .B(n212), .Y(N133) );
  NOR2X1 U51 ( .A(n16), .B(n131), .Y(N113) );
  INVX1 U52 ( .A(n8), .Y(n7) );
  NAND3X1 U53 ( .A(n36), .B(n26), .C(n176), .Y(N257) );
  INVX1 U54 ( .A(n6), .Y(n5) );
  NAND21X1 U55 ( .B(n130), .A(n17), .Y(n127) );
  INVX1 U56 ( .A(n26), .Y(n23) );
  INVX1 U57 ( .A(n28), .Y(n21) );
  INVX1 U58 ( .A(n26), .Y(n24) );
  INVX1 U59 ( .A(n28), .Y(n22) );
  AND3X1 U60 ( .A(n100), .B(n94), .C(sfraddr[5]), .Y(n213) );
  NAND3X1 U61 ( .A(n193), .B(n19), .C(t_shift_clk), .Y(n176) );
  NAND2X1 U62 ( .A(n181), .B(n80), .Y(n179) );
  NOR4XL U63 ( .A(sfraddr[5]), .B(n5), .C(sfraddr[3]), .D(n35), .Y(n101) );
  NOR3XL U64 ( .A(sfraddr[1]), .B(sfraddr[5]), .C(n6), .Y(n95) );
  INVX1 U65 ( .A(sfraddr[4]), .Y(n6) );
  INVX1 U66 ( .A(sfraddr[3]), .Y(n4) );
  INVX1 U67 ( .A(sfrdatai[5]), .Y(n14) );
  INVX1 U68 ( .A(sfrdatai[3]), .Y(n12) );
  INVX1 U69 ( .A(sfrdatai[4]), .Y(n13) );
  INVX1 U70 ( .A(sfrdatai[2]), .Y(n11) );
  INVX1 U71 ( .A(sfrdatai[6]), .Y(n15) );
  INVX1 U72 ( .A(sfrdatai[7]), .Y(n16) );
  INVX1 U73 ( .A(sfrdatai[0]), .Y(n9) );
  INVX1 U74 ( .A(sfrdatai[1]), .Y(n10) );
  INVX1 U75 ( .A(n3), .Y(n226) );
  NAND2X1 U76 ( .A(n145), .B(n3), .Y(n130) );
  NAND32X1 U77 ( .B(n114), .C(rst), .A(n145), .Y(n153) );
  NOR21XL U78 ( .B(t1ov), .A(n21), .Y(N59) );
  OAI211X1 U79 ( .C(n60), .D(n153), .A(n129), .B(n25), .Y(N471) );
  INVX1 U80 ( .A(rst), .Y(n26) );
  NOR3XL U81 ( .A(n120), .B(n24), .C(n3), .Y(n166) );
  INVX1 U82 ( .A(rst), .Y(n25) );
  INVX1 U83 ( .A(rst), .Y(n28) );
  NOR2X1 U84 ( .A(n23), .B(n114), .Y(n134) );
  INVX1 U85 ( .A(n140), .Y(n55) );
  NAND3X1 U86 ( .A(n114), .B(n19), .C(n77), .Y(n129) );
  NAND2X1 U87 ( .A(n228), .B(n227), .Y(n80) );
  NOR2X1 U88 ( .A(n80), .B(n225), .Y(rxd0oe) );
  NOR2X1 U89 ( .A(n24), .B(newinstr), .Y(n104) );
  NOR32XL U90 ( .B(r_shift_clk), .C(n221), .A(n138), .Y(n145) );
  AOI21X1 U91 ( .B(n78), .C(n196), .A(N224), .Y(n199) );
  INVX1 U92 ( .A(n117), .Y(n67) );
  NOR3XL U93 ( .A(n115), .B(n117), .C(n217), .Y(r_shift_clk) );
  INVX1 U94 ( .A(n196), .Y(n66) );
  OAI22X1 U95 ( .A(n153), .B(n48), .C(n129), .D(n47), .Y(N473) );
  OAI22X1 U96 ( .A(n153), .B(n46), .C(n129), .D(n45), .Y(N475) );
  OAI22X1 U97 ( .A(n153), .B(n45), .C(n129), .D(n44), .Y(N476) );
  OAI22X1 U98 ( .A(n153), .B(n44), .C(n129), .D(n43), .Y(N477) );
  OAI22X1 U99 ( .A(n153), .B(n47), .C(n129), .D(n46), .Y(N474) );
  OAI22X1 U100 ( .A(n153), .B(n43), .C(n129), .D(n42), .Y(N478) );
  OAI22X1 U101 ( .A(n153), .B(n42), .C(n61), .D(n129), .Y(N479) );
  AOI211X1 U102 ( .C(n215), .D(n78), .A(n66), .B(n79), .Y(N225) );
  OAI21X1 U103 ( .B(n217), .C(n108), .A(n109), .Y(n240) );
  OAI211X1 U104 ( .C(n110), .D(n111), .A(n108), .B(n25), .Y(n109) );
  NAND32X1 U105 ( .B(n110), .C(rst), .A(n112), .Y(n108) );
  AND3X1 U106 ( .A(n226), .B(n120), .C(n217), .Y(n110) );
  NAND2X1 U107 ( .A(n154), .B(n81), .Y(N428) );
  OAI21X1 U108 ( .B(n62), .C(n126), .A(n20), .Y(n204) );
  NAND21X1 U109 ( .B(n204), .A(n126), .Y(n205) );
  INVX1 U110 ( .A(n138), .Y(n77) );
  AOI22AXL U111 ( .A(n226), .B(n120), .D(n159), .C(n3), .Y(n154) );
  NAND2X1 U112 ( .A(n56), .B(n117), .Y(n140) );
  OAI21AX1 U113 ( .B(n166), .C(n159), .A(n164), .Y(n162) );
  OAI32X1 U114 ( .A(n63), .B(n126), .C(n204), .D(n62), .E(n205), .Y(N188) );
  NOR2X1 U115 ( .A(n156), .B(n80), .Y(n114) );
  NOR3XL U116 ( .A(n53), .B(n156), .C(n224), .Y(n120) );
  OAI21X1 U117 ( .B(n117), .C(n244), .A(n20), .Y(N325) );
  AOI211X1 U118 ( .C(n152), .D(n218), .A(n169), .B(n170), .Y(N363) );
  NOR2X1 U119 ( .A(n225), .B(n156), .Y(t_shift_clk) );
  INVX1 U120 ( .A(n139), .Y(n56) );
  INVX1 U121 ( .A(n81), .Y(n27) );
  NAND2X1 U122 ( .A(n18), .B(n200), .Y(N223) );
  NAND3X1 U123 ( .A(n19), .B(n64), .C(n169), .Y(N360) );
  NAND32X1 U124 ( .B(n1), .C(n2), .A(n17), .Y(N166) );
  AOI21AX1 U125 ( .B(n225), .C(n217), .A(n25), .Y(n122) );
  AOI211X1 U126 ( .C(n59), .D(n57), .A(n204), .B(n58), .Y(N186) );
  INVX1 U127 ( .A(n126), .Y(n58) );
  NOR3XL U128 ( .A(n97), .B(n24), .C(n41), .Y(N207) );
  NOR2X1 U129 ( .A(n221), .B(n22), .Y(N348) );
  NAND2X1 U130 ( .A(n61), .B(n17), .Y(N382) );
  NOR2X1 U131 ( .A(n24), .B(n96), .Y(n245) );
  XNOR2XL U132 ( .A(n41), .B(n97), .Y(n96) );
  NAND3X1 U133 ( .A(n226), .B(n40), .C(n122), .Y(N303) );
  NAND2X1 U134 ( .A(n18), .B(n117), .Y(N324) );
  INVX1 U135 ( .A(n198), .Y(n79) );
  NOR43XL U136 ( .B(n63), .C(n57), .D(N190), .A(n62), .Y(N191) );
  NOR3XL U137 ( .A(n208), .B(n24), .C(n203), .Y(N142) );
  NOR2X1 U138 ( .A(n152), .B(n218), .Y(n170) );
  NOR2X1 U139 ( .A(n59), .B(n22), .Y(N190) );
  NAND2X1 U140 ( .A(n18), .B(n47), .Y(N376) );
  NAND2X1 U141 ( .A(n18), .B(n46), .Y(N377) );
  NAND2X1 U142 ( .A(n18), .B(n45), .Y(N378) );
  NAND2X1 U143 ( .A(n18), .B(n44), .Y(N379) );
  NAND2X1 U144 ( .A(n18), .B(n43), .Y(N380) );
  NAND2X1 U145 ( .A(n18), .B(n42), .Y(N381) );
  NAND2X1 U146 ( .A(n18), .B(n48), .Y(N375) );
  NOR2X1 U147 ( .A(n24), .B(n244), .Y(N307) );
  INVX1 U148 ( .A(n143), .Y(n60) );
  INVX1 U149 ( .A(s0con[6]), .Y(n227) );
  INVX1 U150 ( .A(t_start), .Y(n225) );
  INVX1 U151 ( .A(s0con[7]), .Y(n228) );
  AO222X1 U152 ( .A(sfrdatai[1]), .B(n32), .C(n107), .D(ti_tmp), .E(s0con[1]), 
        .F(n33), .Y(n241) );
  OAI211X1 U153 ( .C(n9), .D(n179), .A(n20), .B(n191), .Y(N260) );
  AOI22X1 U154 ( .A(n37), .B(sfrdatai[1]), .C(t_shift_reg[3]), .D(n39), .Y(
        n191) );
  OAI211X1 U155 ( .C(n10), .D(n179), .A(n28), .B(n190), .Y(N261) );
  AOI22X1 U156 ( .A(n37), .B(sfrdatai[2]), .C(t_shift_reg[4]), .D(n39), .Y(
        n190) );
  OAI211X1 U157 ( .C(n179), .D(n14), .A(n28), .B(n186), .Y(N265) );
  AOI22X1 U158 ( .A(n37), .B(sfrdatai[6]), .C(t_shift_reg[8]), .D(n39), .Y(
        n186) );
  OAI211X1 U159 ( .C(n11), .D(n179), .A(n20), .B(n189), .Y(N262) );
  AOI22X1 U160 ( .A(sfrdatai[3]), .B(n37), .C(t_shift_reg[5]), .D(n39), .Y(
        n189) );
  OAI211X1 U161 ( .C(n179), .D(n12), .A(n28), .B(n188), .Y(N263) );
  AOI22X1 U162 ( .A(sfrdatai[4]), .B(n37), .C(t_shift_reg[6]), .D(n39), .Y(
        n188) );
  OAI211X1 U163 ( .C(n179), .D(n13), .A(n28), .B(n187), .Y(N264) );
  AOI22X1 U164 ( .A(sfrdatai[5]), .B(n37), .C(t_shift_reg[7]), .D(n39), .Y(
        n187) );
  OAI211X1 U165 ( .C(n179), .D(n15), .A(n28), .B(n185), .Y(N266) );
  AOI22X1 U166 ( .A(n37), .B(sfrdatai[7]), .C(t_shift_reg[9]), .D(n39), .Y(
        n185) );
  AO222X1 U167 ( .A(n131), .B(N348), .C(n107), .D(ri_tmp), .E(n32), .F(
        sfrdatai[0]), .Y(n237) );
  GEN2XL U168 ( .D(t_shift_count[1]), .E(t_shift_count[0]), .C(n178), .B(n39), 
        .A(n38), .Y(N282) );
  INVX1 U169 ( .A(n179), .Y(n38) );
  INVX1 U170 ( .A(n98), .Y(n29) );
  AOI32X1 U171 ( .A(smod), .B(n19), .C(n99), .D(sfrdatai[7]), .E(n31), .Y(n98)
         );
  INVX1 U172 ( .A(n99), .Y(n31) );
  NAND4XL U173 ( .A(sfraddr[0]), .B(n100), .C(sfraddr[2]), .D(n101), .Y(n99)
         );
  NAND3X1 U174 ( .A(n176), .B(n28), .C(n182), .Y(N268) );
  OAI21X1 U175 ( .B(s0con[3]), .C(n228), .A(n181), .Y(n182) );
  OAI21X1 U176 ( .B(n131), .C(n11), .A(n147), .Y(n230) );
  AOI33X1 U177 ( .A(s0con2_tmp), .B(n107), .C(s0con2_val), .D(n33), .E(n51), 
        .F(s0con[2]), .Y(n147) );
  INVX1 U178 ( .A(s0con2_tmp), .Y(n51) );
  OAI21X1 U179 ( .B(t_shift_count[0]), .C(n176), .A(n180), .Y(N281) );
  OAI21X1 U180 ( .B(s0con[7]), .C(n227), .A(n181), .Y(n180) );
  OAI21X1 U181 ( .B(n175), .C(n176), .A(n36), .Y(N284) );
  XOR2X1 U182 ( .A(n103), .B(t_shift_count[3]), .Y(n175) );
  NAND3X1 U183 ( .A(n183), .B(n19), .C(n184), .Y(N267) );
  AOI22X1 U184 ( .A(t_shift_reg[10]), .B(n39), .C(n181), .D(sfrdatai[7]), .Y(
        n184) );
  OAI2B11X1 U185 ( .D(t_shift_reg[1]), .C(n176), .A(n36), .B(n25), .Y(N258) );
  OAI211X1 U186 ( .C(n9), .D(n183), .A(n28), .B(n192), .Y(N259) );
  NAND2X1 U187 ( .A(t_shift_reg[2]), .B(n39), .Y(n192) );
  INVX1 U188 ( .A(n92), .Y(n30) );
  AOI32X1 U189 ( .A(bd), .B(n19), .C(n93), .D(n34), .E(sfrdatai[7]), .Y(n92)
         );
  INVX1 U190 ( .A(n93), .Y(n34) );
  NAND4X1 U191 ( .A(n7), .B(n94), .C(n95), .D(n17), .Y(n93) );
  ENOX1 U192 ( .A(n127), .B(n142), .C(n142), .D(s0con2_tmp), .Y(n232) );
  ENOX1 U193 ( .A(n127), .B(n143), .C(n130), .D(n104), .Y(n142) );
  AOI21X1 U194 ( .B(n103), .C(n177), .A(n176), .Y(N283) );
  NAND21X1 U195 ( .B(n178), .A(t_shift_count[2]), .Y(n177) );
  NAND2X1 U196 ( .A(n36), .B(n102), .Y(n243) );
  OAI211X1 U197 ( .C(t_shift_count[3]), .D(n103), .A(n28), .B(t_start), .Y(
        n102) );
  OAI211X1 U198 ( .C(n60), .D(n127), .A(n128), .B(n129), .Y(n238) );
  NAND3X1 U199 ( .A(n104), .B(n130), .C(ri_tmp), .Y(n128) );
  OAI21BBX1 U200 ( .A(n104), .B(ti_tmp), .C(n105), .Y(n242) );
  NAND4X1 U201 ( .A(t_shift_clk), .B(n19), .C(t_shift_count[0]), .D(n106), .Y(
        n105) );
  NOR3XL U202 ( .A(t_shift_count[1]), .B(t_shift_count[3]), .C(
        t_shift_count[2]), .Y(n106) );
  ENOX1 U203 ( .A(smod), .B(baud_r2_clk), .C(n97), .D(smod), .Y(n117) );
  AOI31X1 U204 ( .A(t_baud_count[2]), .B(s0relh[6]), .C(n79), .D(n200), .Y(
        n196) );
  OAI32X1 U205 ( .A(n66), .B(t_baud_count[2]), .C(n198), .D(n199), .E(n216), 
        .Y(N226) );
  OAI32X1 U206 ( .A(n50), .B(rst), .C(n144), .D(n61), .E(n127), .Y(n231) );
  INVX1 U207 ( .A(s0con2_val), .Y(n50) );
  NOR4XL U208 ( .A(n146), .B(n138), .C(n115), .D(n217), .Y(n144) );
  NAND3X1 U209 ( .A(n3), .B(n221), .C(n143), .Y(n146) );
  OAI22AX1 U210 ( .D(n201), .C(t1ov_ff), .A(n202), .B(n201), .Y(n97) );
  NOR2X1 U211 ( .A(n227), .B(bd), .Y(n201) );
  AOI221XL U212 ( .A(s0con[6]), .B(n220), .C(n203), .D(n227), .E(n226), .Y(
        n202) );
  NAND3X1 U213 ( .A(t_start), .B(n19), .C(n67), .Y(n200) );
  NOR2X1 U214 ( .A(s0relh[7]), .B(r_clk_ov2), .Y(n203) );
  NOR2X1 U215 ( .A(n66), .B(t_baud_count[0]), .Y(N224) );
  GEN2XL U216 ( .D(n196), .E(n216), .C(n65), .B(t_baud_count[3]), .A(n197), 
        .Y(N227) );
  NOR4XL U217 ( .A(t_baud_count[3]), .B(n198), .C(n216), .D(n66), .Y(n197) );
  INVX1 U218 ( .A(n199), .Y(n65) );
  AOI22X1 U219 ( .A(n113), .B(n80), .C(n77), .D(n114), .Y(n112) );
  OAI32X1 U220 ( .A(n115), .B(n116), .C(n117), .D(n224), .E(n118), .Y(n113) );
  AOI21X1 U221 ( .B(rxd0_val), .C(n119), .A(n77), .Y(n116) );
  OAI22AX1 U222 ( .D(r_shift_reg[0]), .C(n153), .A(n129), .B(n48), .Y(N472) );
  INVX1 U223 ( .A(baud_rate_ov), .Y(n220) );
  NAND43X1 U224 ( .B(r_shift_count[3]), .C(r_shift_count[1]), .D(
        r_shift_count[2]), .A(r_shift_count[0]), .Y(n138) );
  AOI22X1 U225 ( .A(n222), .B(n220), .C(n208), .D(s0relh[7]), .Y(n83) );
  AOI21X1 U226 ( .B(n222), .C(r_clk_ov2), .A(n83), .Y(n84) );
  GEN2XL U227 ( .D(n56), .E(n49), .C(n55), .B(fluctuation_conter[1]), .A(n141), 
        .Y(n233) );
  NOR4XL U228 ( .A(fluctuation_conter[1]), .B(n55), .C(n139), .D(n49), .Y(n141) );
  INVX1 U229 ( .A(n85), .Y(n75) );
  AOI221XL U230 ( .A(s0relh[0]), .B(n83), .C(N153), .D(n84), .E(n23), .Y(n85)
         );
  NAND21X1 U231 ( .B(r_shift_count[2]), .A(n163), .Y(n160) );
  OAI22X1 U232 ( .A(t_baud_ov), .B(n226), .C(clk_ov12), .D(n80), .Y(n156) );
  NAND2X1 U233 ( .A(rxd0_fall_fl), .B(n17), .Y(n139) );
  NOR42XL U234 ( .C(r_shift_count[3]), .D(r_shift_count[1]), .A(
        r_shift_count[0]), .B(r_shift_count[2]), .Y(n119) );
  OAI32X1 U235 ( .A(n204), .B(clk_count[2]), .C(n126), .D(n63), .E(n205), .Y(
        N187) );
  OAI32X1 U236 ( .A(n139), .B(fluctuation_conter[0]), .C(n55), .D(n140), .E(
        n49), .Y(n234) );
  OAI32X1 U237 ( .A(n49), .B(n64), .C(n139), .D(r_baud_count[0]), .E(n169), 
        .Y(N361) );
  OAI32X1 U238 ( .A(n52), .B(n64), .C(n139), .D(n171), .E(n169), .Y(N362) );
  INVX1 U239 ( .A(fluctuation_conter[1]), .Y(n52) );
  AOI21X1 U240 ( .B(r_baud_count[1]), .C(n219), .A(n151), .Y(n171) );
  OAI32X1 U241 ( .A(n159), .B(n24), .C(n226), .D(n164), .E(n165), .Y(N425) );
  AOI21X1 U242 ( .B(r_shift_count[0]), .C(r_shift_count[1]), .A(n163), .Y(n165) );
  NAND4X1 U243 ( .A(r_start), .B(n67), .C(n17), .D(n64), .Y(n169) );
  NOR2X1 U244 ( .A(r_shift_count[0]), .B(r_shift_count[1]), .Y(n163) );
  NAND41X1 U245 ( .D(n209), .A(n210), .B(tim_baud[8]), .C(tim_baud[9]), .Y(
        n208) );
  NAND3X1 U246 ( .A(tim_baud[6]), .B(tim_baud[5]), .C(tim_baud[7]), .Y(n209)
         );
  NOR32XL U247 ( .B(tim_baud[4]), .C(tim_baud[3]), .A(n211), .Y(n210) );
  NAND3X1 U248 ( .A(tim_baud[1]), .B(tim_baud[0]), .C(tim_baud[2]), .Y(n211)
         );
  INVX1 U249 ( .A(r_baud_count[2]), .Y(n218) );
  NOR4XL U250 ( .A(rxd0_fall), .B(receive_11_bits), .C(r_start), .D(n174), .Y(
        N306) );
  AOI31X1 U251 ( .A(n19), .B(n244), .C(rxd0_ff), .D(n56), .Y(n174) );
  NOR2X1 U252 ( .A(n219), .B(r_baud_count[1]), .Y(n151) );
  NOR2X1 U253 ( .A(n160), .B(r_shift_count[3]), .Y(n111) );
  OAI21X1 U254 ( .B(N382), .C(n157), .A(n158), .Y(N427) );
  GEN2XL U255 ( .D(n119), .E(n80), .C(n157), .B(n154), .A(rst), .Y(n158) );
  AOI21X1 U256 ( .B(n160), .C(r_shift_count[3]), .A(n111), .Y(n157) );
  OAI21X1 U257 ( .B(n53), .C(n132), .A(n133), .Y(n236) );
  NAND4X1 U258 ( .A(ri0_ff), .B(n132), .C(n17), .D(n221), .Y(n133) );
  OAI31XL U259 ( .A(n54), .B(s0con[0]), .C(n80), .D(n134), .Y(n132) );
  INVX1 U260 ( .A(ri0_ff), .Y(n54) );
  AOI221XL U261 ( .A(s0relh[6]), .B(n218), .C(n76), .D(n223), .E(n135), .Y(
        n235) );
  AOI22X1 U262 ( .A(n136), .B(n137), .C(n56), .D(n118), .Y(n135) );
  NOR32XL U263 ( .B(rxd0_ff), .C(s0con[6]), .A(n138), .Y(n136) );
  NOR3XL U264 ( .A(n24), .B(s0con[7]), .C(rxd0ff), .Y(n137) );
  NAND2X1 U265 ( .A(n151), .B(n155), .Y(n115) );
  OAI32X1 U266 ( .A(n76), .B(s0relh[6]), .C(r_baud_count[2]), .D(n218), .E(
        n223), .Y(n155) );
  NOR4XL U267 ( .A(n195), .B(n215), .C(n21), .D(n117), .Y(N230) );
  NAND32X1 U268 ( .B(t_baud_count[3]), .C(t_baud_count[2]), .A(n78), .Y(n195)
         );
  AOI21X1 U269 ( .B(n160), .C(n161), .A(n162), .Y(N426) );
  NAND21X1 U270 ( .B(n163), .A(r_shift_count[2]), .Y(n161) );
  INVX1 U271 ( .A(s0relh[6]), .Y(n223) );
  OAI21BBX1 U272 ( .A(n67), .B(rxd0_vec[0]), .C(n25), .Y(N326) );
  OAI21BBX1 U273 ( .A(n67), .B(rxd0_vec[1]), .C(n25), .Y(N327) );
  NOR2X1 U274 ( .A(n167), .B(n166), .Y(n164) );
  AOI211X1 U275 ( .C(n119), .D(rxd0_val), .A(n226), .B(n21), .Y(n167) );
  NAND2X1 U276 ( .A(rxd0_fall), .B(n111), .Y(n118) );
  INVX1 U277 ( .A(r_baud_count[0]), .Y(n219) );
  INVX1 U278 ( .A(r_baud_count[3]), .Y(n76) );
  NOR2X1 U279 ( .A(n168), .B(n169), .Y(N364) );
  XNOR2XL U280 ( .A(r_baud_count[3]), .B(n170), .Y(n168) );
  NOR2X1 U281 ( .A(n21), .B(n207), .Y(N169) );
  AOI22X1 U282 ( .A(N147), .B(n84), .C(s0rell[2]), .D(n2), .Y(n207) );
  NOR2X1 U283 ( .A(n22), .B(n206), .Y(N170) );
  AOI22X1 U284 ( .A(N148), .B(n1), .C(s0rell[3]), .D(n2), .Y(n206) );
  NOR2X1 U285 ( .A(r_shift_count[0]), .B(n162), .Y(N424) );
  INVX1 U286 ( .A(n87), .Y(n73) );
  AOI221XL U287 ( .A(s0rell[6]), .B(n83), .C(N151), .D(n84), .E(n21), .Y(n87)
         );
  INVX1 U288 ( .A(n90), .Y(n70) );
  AOI221XL U289 ( .A(s0rell[1]), .B(n83), .C(N146), .D(n84), .E(n22), .Y(n90)
         );
  INVX1 U290 ( .A(n88), .Y(n72) );
  AOI221XL U291 ( .A(s0rell[5]), .B(n83), .C(N150), .D(n84), .E(n21), .Y(n88)
         );
  INVX1 U292 ( .A(n86), .Y(n74) );
  AOI221XL U293 ( .A(s0rell[7]), .B(n83), .C(N152), .D(n84), .E(n21), .Y(n86)
         );
  INVX1 U294 ( .A(n89), .Y(n71) );
  AOI221XL U295 ( .A(s0rell[4]), .B(n83), .C(N149), .D(n84), .E(n21), .Y(n89)
         );
  INVX1 U296 ( .A(n82), .Y(n68) );
  AOI221XL U297 ( .A(s0relh[1]), .B(n83), .C(N154), .D(n84), .E(n22), .Y(n82)
         );
  INVX1 U298 ( .A(n91), .Y(n69) );
  AOI221XL U299 ( .A(s0rell[0]), .B(n83), .C(N145), .D(n84), .E(n22), .Y(n91)
         );
  NAND2X1 U300 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n126) );
  NAND2X1 U301 ( .A(t_baud_count[1]), .B(t_baud_count[0]), .Y(n198) );
  NAND2X1 U302 ( .A(s0con[5]), .B(n61), .Y(n143) );
  NOR31X1 U303 ( .C(t_shift_count[0]), .A(t_shift_count[2]), .B(
        t_shift_count[1]), .Y(n125) );
  OAI21X1 U304 ( .B(n80), .C(n244), .A(n172), .Y(N333) );
  AOI21X1 U305 ( .B(n173), .C(n3), .A(n22), .Y(n172) );
  AND2X1 U306 ( .A(n148), .B(s0con[7]), .Y(n229) );
  OAI33XL U307 ( .A(n149), .B(n21), .C(n150), .D(n138), .E(n22), .F(n115), .Y(
        n148) );
  OAI31XL U308 ( .A(n152), .B(r_baud_count[2]), .C(n223), .D(receive_11_bits), 
        .Y(n149) );
  NOR43XL U309 ( .B(n223), .C(n76), .D(n151), .A(n218), .Y(n150) );
  INVX1 U310 ( .A(s0con[0]), .Y(n221) );
  INVX1 U311 ( .A(r_start), .Y(n217) );
  INVX1 U312 ( .A(rxd0_val), .Y(n61) );
  OAI211X1 U313 ( .C(n226), .D(n40), .A(n121), .B(n122), .Y(n239) );
  OAI21BBX1 U314 ( .A(n123), .B(n124), .C(n226), .Y(n121) );
  OAI31XL U315 ( .A(clk_count[0]), .B(clk_count[2]), .C(clk_count[1]), .D(
        clk_count[3]), .Y(n124) );
  AOI33X1 U316 ( .A(txd0), .B(t_shift_count[3]), .C(n125), .D(n63), .E(n62), 
        .F(n126), .Y(n123) );
  NAND2X1 U317 ( .A(rxd0_fall), .B(s0con[4]), .Y(n159) );
  INVX1 U318 ( .A(s0con[4]), .Y(n224) );
  NOR2X1 U319 ( .A(clk_count[0]), .B(n204), .Y(N185) );
  INVX1 U320 ( .A(s0relh[7]), .Y(n222) );
  INVX1 U321 ( .A(ri0_fall), .Y(n53) );
  NAND21X1 U322 ( .B(t_shift_count[2]), .A(n178), .Y(n103) );
  NOR2X1 U323 ( .A(t_shift_count[1]), .B(t_shift_count[0]), .Y(n178) );
  INVX1 U324 ( .A(rxd0_fall), .Y(n64) );
  INVX1 U325 ( .A(clk_count[3]), .Y(n62) );
  NAND2X1 U326 ( .A(r_baud_count[1]), .B(r_baud_count[0]), .Y(n152) );
  INVX1 U327 ( .A(t_baud_count[1]), .Y(n78) );
  INVX1 U328 ( .A(rxd0ff), .Y(n244) );
  INVX1 U330 ( .A(fluctuation_conter[0]), .Y(n49) );
  INVX1 U331 ( .A(clk_count[2]), .Y(n63) );
  INVX1 U332 ( .A(t_baud_count[2]), .Y(n216) );
  INVX1 U333 ( .A(clk_count[0]), .Y(n59) );
  INVX1 U334 ( .A(r_shift_reg[1]), .Y(n48) );
  INVX1 U335 ( .A(r_shift_reg[2]), .Y(n47) );
  INVX1 U336 ( .A(r_shift_reg[3]), .Y(n46) );
  INVX1 U337 ( .A(r_shift_reg[4]), .Y(n45) );
  INVX1 U338 ( .A(r_shift_reg[5]), .Y(n44) );
  INVX1 U339 ( .A(r_shift_reg[6]), .Y(n43) );
  INVX1 U340 ( .A(r_shift_reg[7]), .Y(n42) );
  INVX1 U341 ( .A(t_baud_count[0]), .Y(n215) );
  INVX1 U342 ( .A(clk_count[1]), .Y(n57) );
  INVX1 U343 ( .A(baud_r_count), .Y(n41) );
  INVX1 U344 ( .A(t_shift_reg[0]), .Y(n40) );
endmodule


module serial0_a0_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ports_a0 ( clkper, rst, port0, sfrdatai, sfraddr, sfrwe, test_si, 
        test_se );
  output [7:0] port0;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkper, rst, sfrwe, test_si, test_se;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, net12317, n2, n3, n4, n1;

  SNPS_CLOCK_GATE_HIGH_ports_a0 clk_gate_p0_reg ( .CLK(clkper), .EN(N2), 
        .ENCLK(net12317), .TE(test_se) );
  SDFFQX1 p0_reg_7_ ( .D(N10), .SIN(port0[6]), .SMC(test_se), .C(net12317), 
        .Q(port0[7]) );
  SDFFQX1 p0_reg_4_ ( .D(N7), .SIN(port0[3]), .SMC(test_se), .C(net12317), .Q(
        port0[4]) );
  SDFFQX1 p0_reg_6_ ( .D(N9), .SIN(port0[5]), .SMC(test_se), .C(net12317), .Q(
        port0[6]) );
  SDFFQX1 p0_reg_5_ ( .D(N8), .SIN(port0[4]), .SMC(test_se), .C(net12317), .Q(
        port0[5]) );
  SDFFQX1 p0_reg_1_ ( .D(N4), .SIN(port0[0]), .SMC(test_se), .C(net12317), .Q(
        port0[1]) );
  SDFFQX1 p0_reg_0_ ( .D(N3), .SIN(test_si), .SMC(test_se), .C(net12317), .Q(
        port0[0]) );
  SDFFQX1 p0_reg_2_ ( .D(N5), .SIN(port0[1]), .SMC(test_se), .C(net12317), .Q(
        port0[2]) );
  SDFFQX1 p0_reg_3_ ( .D(N6), .SIN(port0[2]), .SMC(test_se), .C(net12317), .Q(
        port0[3]) );
  NAND2X1 U2 ( .A(n1), .B(n2), .Y(N2) );
  NAND42X1 U3 ( .C(sfraddr[3]), .D(sfraddr[2]), .A(n3), .B(n4), .Y(n2) );
  NOR3XL U4 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n3) );
  NOR42XL U5 ( .C(sfrwe), .D(n1), .A(sfraddr[1]), .B(sfraddr[0]), .Y(n4) );
  NOR21XL U6 ( .B(sfrdatai[2]), .A(n2), .Y(N5) );
  NOR21XL U7 ( .B(sfrdatai[0]), .A(n2), .Y(N3) );
  NOR21XL U8 ( .B(sfrdatai[3]), .A(n2), .Y(N6) );
  NOR21XL U9 ( .B(sfrdatai[1]), .A(n2), .Y(N4) );
  NOR21XL U10 ( .B(sfrdatai[4]), .A(n2), .Y(N7) );
  NOR21XL U11 ( .B(sfrdatai[5]), .A(n2), .Y(N8) );
  NOR21XL U12 ( .B(sfrdatai[6]), .A(n2), .Y(N9) );
  NOR21XL U13 ( .B(sfrdatai[7]), .A(n2), .Y(N10) );
  INVX1 U14 ( .A(rst), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ports_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mdu_a0 ( clkper, rst, mdubsy, sfrdatai, sfraddr, sfrwe, sfroe, arcon, 
        md0, md1, md2, md3, md4, md5, test_si, test_so, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] arcon;
  output [7:0] md0;
  output [7:0] md1;
  output [7:0] md2;
  output [7:0] md3;
  output [7:0] md4;
  output [7:0] md5;
  input clkper, rst, sfrwe, sfroe, test_si, test_se;
  output mdubsy, test_so;
  wire   N104, N105, N106, N107, N108, N109, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N332, N333, N334, N335, N336, N337, N338, N339, N340,
         N405, N406, N407, N408, N409, N410, N411, N412, N413, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N566, N567, N568, N569, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N610,
         N674, N675, N676, N677, N678, set_div16, set_div32, N802, N892, N893,
         N894, N895, net12335, net12341, net12346, net12351, net12356,
         net12361, net12366, n408, n409, n410, n411, n412, n413, n414, n137,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n1, n2, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n405, n406, n407, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2;
  wire   [3:0] oper_reg;
  wire   [4:1] counter_st;
  wire   [17:1] sum1;
  wire   [17:1] sum;
  wire   [15:0] norm_reg;
  wire   [1:0] mdu_op;
  wire   [17:1] arg_a;
  wire   [16:1] arg_b;
  wire   [17:0] arg_c;
  wire   [16:1] arg_d;

  SNPS_CLOCK_GATE_HIGH_mdu_a0_0 clk_gate_arcon_s_reg ( .CLK(clkper), .EN(N104), 
        .ENCLK(net12335), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_6 clk_gate_md0_s_reg ( .CLK(clkper), .EN(N190), 
        .ENCLK(net12341), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_5 clk_gate_md1_s_reg ( .CLK(clkper), .EN(N258), 
        .ENCLK(net12346), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_4 clk_gate_md2_s_reg ( .CLK(clkper), .EN(N332), 
        .ENCLK(net12351), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_3 clk_gate_md3_s_reg ( .CLK(clkper), .EN(N405), 
        .ENCLK(net12356), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_2 clk_gate_md4_s_reg ( .CLK(clkper), .EN(N453), 
        .ENCLK(net12361), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_1 clk_gate_md5_s_reg ( .CLK(clkper), .EN(N483), 
        .ENCLK(net12366), .TE(test_se) );
  mdu_a0_DW01_add_0 add_1040 ( .A(arg_c), .B({1'b0, arg_d, n404}), .CI(1'b0), 
        .SUM({sum, SYNOPSYS_UNCONNECTED_1}), .CO() );
  mdu_a0_DW01_add_1 add_961 ( .A({arg_a, n137}), .B({1'b0, arg_b, n404}), .CI(
        1'b0), .SUM({sum1, SYNOPSYS_UNCONNECTED_2}), .CO() );
  SDFFQX1 set_div16_reg ( .D(n414), .SIN(oper_reg[3]), .SMC(test_se), .C(
        clkper), .Q(set_div16) );
  SDFFQX1 setmdef_reg ( .D(N802), .SIN(set_div32), .SMC(test_se), .C(clkper), 
        .Q(test_so) );
  SDFFQX1 set_div32_reg ( .D(n413), .SIN(set_div16), .SMC(test_se), .C(clkper), 
        .Q(set_div32) );
  SDFFQX1 counter_st_reg_0_ ( .D(N674), .SIN(arcon[7]), .SMC(test_se), .C(
        clkper), .Q(N610) );
  SDFFQX1 counter_st_reg_1_ ( .D(N675), .SIN(N610), .SMC(test_se), .C(clkper), 
        .Q(counter_st[1]) );
  SDFFQX1 counter_st_reg_2_ ( .D(N676), .SIN(counter_st[1]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[2]) );
  SDFFQX1 counter_st_reg_4_ ( .D(N678), .SIN(counter_st[3]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[4]) );
  SDFFQX1 counter_st_reg_3_ ( .D(N677), .SIN(counter_st[2]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[3]) );
  SDFFQX1 oper_reg_reg_3_ ( .D(N895), .SIN(oper_reg[2]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[3]) );
  SDFFQX1 oper_reg_reg_0_ ( .D(N892), .SIN(norm_reg[15]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[0]) );
  SDFFQX1 oper_reg_reg_1_ ( .D(N893), .SIN(oper_reg[0]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[1]) );
  SDFFQX1 oper_reg_reg_2_ ( .D(N894), .SIN(oper_reg[1]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[2]) );
  SDFFQX1 norm_reg_reg_15_ ( .D(N581), .SIN(norm_reg[14]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[15]) );
  SDFFQX1 norm_reg_reg_14_ ( .D(N580), .SIN(norm_reg[13]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[14]) );
  SDFFQX1 norm_reg_reg_13_ ( .D(N579), .SIN(norm_reg[12]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[13]) );
  SDFFQX1 norm_reg_reg_12_ ( .D(N578), .SIN(norm_reg[11]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[12]) );
  SDFFQX1 norm_reg_reg_11_ ( .D(N577), .SIN(norm_reg[10]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[11]) );
  SDFFQX1 norm_reg_reg_10_ ( .D(N576), .SIN(norm_reg[9]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[10]) );
  SDFFQX1 norm_reg_reg_9_ ( .D(N575), .SIN(norm_reg[8]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[9]) );
  SDFFQX1 arcon_s_reg_6_ ( .D(n408), .SIN(arcon[5]), .SMC(test_se), .C(clkper), 
        .Q(arcon[6]) );
  SDFFQX1 arcon_s_reg_3_ ( .D(N108), .SIN(arcon[2]), .SMC(test_se), .C(
        net12335), .Q(arcon[3]) );
  SDFFQX1 md1_s_reg_6_ ( .D(N265), .SIN(md1[5]), .SMC(test_se), .C(net12346), 
        .Q(md1[6]) );
  SDFFQX1 arcon_s_reg_1_ ( .D(N106), .SIN(arcon[0]), .SMC(test_se), .C(
        net12335), .Q(arcon[1]) );
  SDFFQX1 norm_reg_reg_8_ ( .D(N574), .SIN(norm_reg[7]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[8]) );
  SDFFQX1 norm_reg_reg_7_ ( .D(N573), .SIN(norm_reg[6]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[7]) );
  SDFFQX1 md1_s_reg_5_ ( .D(N264), .SIN(md1[4]), .SMC(test_se), .C(net12346), 
        .Q(md1[5]) );
  SDFFQX1 md1_s_reg_4_ ( .D(N263), .SIN(md1[3]), .SMC(test_se), .C(net12346), 
        .Q(md1[4]) );
  SDFFQX1 md0_s_reg_6_ ( .D(N197), .SIN(md0[5]), .SMC(test_se), .C(net12341), 
        .Q(md0[6]) );
  SDFFQX1 md0_s_reg_7_ ( .D(N198), .SIN(md0[6]), .SMC(test_se), .C(net12341), 
        .Q(md0[7]) );
  SDFFQX1 md5_s_reg_3_ ( .D(N487), .SIN(md5[2]), .SMC(test_se), .C(net12366), 
        .Q(md5[3]) );
  SDFFQX1 md5_s_reg_2_ ( .D(N486), .SIN(md5[1]), .SMC(test_se), .C(net12366), 
        .Q(md5[2]) );
  SDFFQX1 md5_s_reg_1_ ( .D(N485), .SIN(md5[0]), .SMC(test_se), .C(net12366), 
        .Q(md5[1]) );
  SDFFQX1 md3_s_reg_6_ ( .D(N412), .SIN(md3[5]), .SMC(test_se), .C(net12356), 
        .Q(md3[6]) );
  SDFFQX1 arcon_s_reg_7_ ( .D(n410), .SIN(arcon[6]), .SMC(test_se), .C(clkper), 
        .Q(arcon[7]) );
  SDFFQX1 arcon_s_reg_0_ ( .D(N105), .SIN(test_si), .SMC(test_se), .C(net12335), .Q(arcon[0]) );
  SDFFQX1 arcon_s_reg_2_ ( .D(N107), .SIN(arcon[1]), .SMC(test_se), .C(
        net12335), .Q(arcon[2]) );
  SDFFQX1 arcon_s_reg_4_ ( .D(N109), .SIN(arcon[3]), .SMC(test_se), .C(
        net12335), .Q(arcon[4]) );
  SDFFQX1 md0_s_reg_3_ ( .D(N194), .SIN(md0[2]), .SMC(test_se), .C(net12341), 
        .Q(md0[3]) );
  SDFFQX1 md3_s_reg_5_ ( .D(N411), .SIN(md3[4]), .SMC(test_se), .C(net12356), 
        .Q(md3[5]) );
  SDFFQX1 norm_reg_reg_6_ ( .D(N572), .SIN(norm_reg[5]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[6]) );
  SDFFQX1 arcon_s_reg_5_ ( .D(n409), .SIN(arcon[4]), .SMC(test_se), .C(
        net12335), .Q(arcon[5]) );
  SDFFQX1 md5_s_reg_6_ ( .D(N490), .SIN(md5[5]), .SMC(test_se), .C(net12366), 
        .Q(md5[6]) );
  SDFFQX1 md5_s_reg_7_ ( .D(N491), .SIN(md5[6]), .SMC(test_se), .C(net12366), 
        .Q(md5[7]) );
  SDFFQX1 md5_s_reg_5_ ( .D(N489), .SIN(md5[4]), .SMC(test_se), .C(net12366), 
        .Q(md5[5]) );
  SDFFQX1 md0_s_reg_4_ ( .D(N195), .SIN(md0[3]), .SMC(test_se), .C(net12341), 
        .Q(md0[4]) );
  SDFFQX1 md0_s_reg_5_ ( .D(N196), .SIN(md0[4]), .SMC(test_se), .C(net12341), 
        .Q(md0[5]) );
  SDFFQX1 md1_s_reg_2_ ( .D(N261), .SIN(md1[1]), .SMC(test_se), .C(net12346), 
        .Q(md1[2]) );
  SDFFQX1 md1_s_reg_0_ ( .D(N259), .SIN(md0[7]), .SMC(test_se), .C(net12346), 
        .Q(md1[0]) );
  SDFFQX1 md1_s_reg_1_ ( .D(N260), .SIN(md1[0]), .SMC(test_se), .C(net12346), 
        .Q(md1[1]) );
  SDFFQX1 md1_s_reg_3_ ( .D(N262), .SIN(md1[2]), .SMC(test_se), .C(net12346), 
        .Q(md1[3]) );
  SDFFQX1 md5_s_reg_4_ ( .D(N488), .SIN(md5[3]), .SMC(test_se), .C(net12366), 
        .Q(md5[4]) );
  SDFFQX1 md3_s_reg_1_ ( .D(N407), .SIN(md3[0]), .SMC(test_se), .C(net12356), 
        .Q(md3[1]) );
  SDFFQX1 md3_s_reg_0_ ( .D(N406), .SIN(md2[7]), .SMC(test_se), .C(net12356), 
        .Q(md3[0]) );
  SDFFQX1 md4_s_reg_7_ ( .D(N461), .SIN(md4[6]), .SMC(test_se), .C(net12361), 
        .Q(md4[7]) );
  SDFFQX1 md3_s_reg_3_ ( .D(N409), .SIN(md3[2]), .SMC(test_se), .C(net12356), 
        .Q(md3[3]) );
  SDFFQX1 md2_s_reg_7_ ( .D(N340), .SIN(md2[6]), .SMC(test_se), .C(net12351), 
        .Q(md2[7]) );
  SDFFQX1 md5_s_reg_0_ ( .D(N484), .SIN(md4[7]), .SMC(test_se), .C(net12366), 
        .Q(md5[0]) );
  SDFFQX1 md0_s_reg_2_ ( .D(N193), .SIN(md0[1]), .SMC(test_se), .C(net12341), 
        .Q(md0[2]) );
  SDFFQX1 md0_s_reg_1_ ( .D(N192), .SIN(md0[0]), .SMC(test_se), .C(net12341), 
        .Q(md0[1]) );
  SDFFQX1 norm_reg_reg_5_ ( .D(N571), .SIN(norm_reg[4]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[5]) );
  SDFFQX1 norm_reg_reg_4_ ( .D(N570), .SIN(norm_reg[3]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[4]) );
  SDFFQX1 md2_s_reg_5_ ( .D(N338), .SIN(md2[4]), .SMC(test_se), .C(net12351), 
        .Q(md2[5]) );
  SDFFQX1 md4_s_reg_6_ ( .D(N460), .SIN(md4[5]), .SMC(test_se), .C(net12361), 
        .Q(md4[6]) );
  SDFFQX1 md2_s_reg_6_ ( .D(N339), .SIN(md2[5]), .SMC(test_se), .C(net12351), 
        .Q(md2[6]) );
  SDFFQX1 md3_s_reg_2_ ( .D(N408), .SIN(md3[1]), .SMC(test_se), .C(net12356), 
        .Q(md3[2]) );
  SDFFQX1 md4_s_reg_5_ ( .D(N459), .SIN(md4[4]), .SMC(test_se), .C(net12361), 
        .Q(md4[5]) );
  SDFFQX1 md3_s_reg_4_ ( .D(N410), .SIN(md3[3]), .SMC(test_se), .C(net12356), 
        .Q(md3[4]) );
  SDFFQX1 norm_reg_reg_3_ ( .D(N569), .SIN(norm_reg[2]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[3]) );
  SDFFQX1 md2_s_reg_4_ ( .D(N337), .SIN(md2[3]), .SMC(test_se), .C(net12351), 
        .Q(md2[4]) );
  SDFFQX1 md4_s_reg_4_ ( .D(N458), .SIN(md4[3]), .SMC(test_se), .C(net12361), 
        .Q(md4[4]) );
  SDFFQX1 norm_reg_reg_2_ ( .D(N568), .SIN(norm_reg[1]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[2]) );
  SDFFQX1 norm_reg_reg_1_ ( .D(N567), .SIN(norm_reg[0]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[1]) );
  SDFFQX1 md2_s_reg_3_ ( .D(N336), .SIN(md2[2]), .SMC(test_se), .C(net12351), 
        .Q(md2[3]) );
  SDFFQX1 md2_s_reg_2_ ( .D(N335), .SIN(md2[1]), .SMC(test_se), .C(net12351), 
        .Q(md2[2]) );
  SDFFQX1 md4_s_reg_2_ ( .D(N456), .SIN(md4[1]), .SMC(test_se), .C(net12361), 
        .Q(md4[2]) );
  SDFFQX1 md4_s_reg_3_ ( .D(N457), .SIN(md4[2]), .SMC(test_se), .C(net12361), 
        .Q(md4[3]) );
  SDFFQX1 norm_reg_reg_0_ ( .D(N566), .SIN(mdu_op[1]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[0]) );
  SDFFQX1 md2_s_reg_1_ ( .D(N334), .SIN(md2[0]), .SMC(test_se), .C(net12351), 
        .Q(md2[1]) );
  SDFFQX1 md4_s_reg_1_ ( .D(N455), .SIN(md4[0]), .SMC(test_se), .C(net12361), 
        .Q(md4[1]) );
  SDFFQX1 md0_s_reg_0_ ( .D(N191), .SIN(counter_st[4]), .SMC(test_se), .C(
        net12341), .Q(md0[0]) );
  SDFFQX1 md2_s_reg_0_ ( .D(N333), .SIN(md1[7]), .SMC(test_se), .C(net12351), 
        .Q(md2[0]) );
  SDFFQX1 md1_s_reg_7_ ( .D(N266), .SIN(md1[6]), .SMC(test_se), .C(net12346), 
        .Q(md1[7]) );
  SDFFQX1 md4_s_reg_0_ ( .D(N454), .SIN(md3[7]), .SMC(test_se), .C(net12361), 
        .Q(md4[0]) );
  SDFFQX1 md3_s_reg_7_ ( .D(N413), .SIN(md3[6]), .SMC(test_se), .C(net12356), 
        .Q(md3[7]) );
  SDFFQX1 mdu_op_reg_0_ ( .D(n411), .SIN(md5[7]), .SMC(test_se), .C(clkper), 
        .Q(mdu_op[0]) );
  SDFFQX1 mdu_op_reg_1_ ( .D(n412), .SIN(mdu_op[0]), .SMC(test_se), .C(clkper), 
        .Q(mdu_op[1]) );
  NAND2X1 U5 ( .A(n242), .B(n271), .Y(n1) );
  NAND2X1 U6 ( .A(n271), .B(n53), .Y(n2) );
  INVX1 U7 ( .A(n298), .Y(n5) );
  INVX1 U8 ( .A(n51), .Y(n6) );
  INVX1 U9 ( .A(n66), .Y(n7) );
  NAND2X1 U10 ( .A(n27), .B(n260), .Y(n8) );
  NAND2X1 U11 ( .A(sum1[17]), .B(arg_c[0]), .Y(n9) );
  INVX1 U12 ( .A(n67), .Y(n10) );
  NAND2X1 U13 ( .A(n107), .B(arg_c[0]), .Y(n11) );
  NAND2X1 U14 ( .A(n259), .B(n260), .Y(n12) );
  INVX1 U15 ( .A(n22), .Y(n13) );
  BUFX3 U16 ( .A(n194), .Y(n14) );
  NOR2X1 U17 ( .A(sum1[17]), .B(n26), .Y(n15) );
  INVX1 U18 ( .A(n65), .Y(n16) );
  BUFX3 U19 ( .A(n254), .Y(n17) );
  BUFX3 U20 ( .A(n188), .Y(n18) );
  INVX1 U21 ( .A(n76), .Y(n19) );
  NOR2X1 U22 ( .A(n107), .B(n26), .Y(n20) );
  INVX1 U23 ( .A(n50), .Y(n21) );
  BUFX3 U24 ( .A(n294), .Y(n22) );
  NOR2X1 U25 ( .A(n376), .B(n68), .Y(n23) );
  INVX1 U26 ( .A(n137), .Y(n24) );
  INVX1 U27 ( .A(sum[17]), .Y(n25) );
  INVX1 U28 ( .A(n25), .Y(n26) );
  INVX1 U29 ( .A(n25), .Y(n27) );
  NOR4XL U30 ( .A(n252), .B(n85), .C(n87), .D(n86), .Y(n380) );
  INVX1 U31 ( .A(n168), .Y(n50) );
  NAND2X1 U32 ( .A(n56), .B(n271), .Y(n166) );
  NAND2X1 U33 ( .A(n55), .B(n271), .Y(n168) );
  NAND2X1 U34 ( .A(n271), .B(n53), .Y(n162) );
  NAND2X1 U35 ( .A(n271), .B(n54), .Y(n237) );
  INVX1 U36 ( .A(n37), .Y(n36) );
  INVX1 U37 ( .A(n352), .Y(n54) );
  INVX1 U38 ( .A(n328), .Y(n53) );
  INVX1 U39 ( .A(n336), .Y(n77) );
  INVX1 U40 ( .A(n369), .Y(n79) );
  INVX1 U41 ( .A(n342), .Y(n67) );
  INVX1 U42 ( .A(n32), .Y(n30) );
  INVX1 U43 ( .A(n404), .Y(n35) );
  INVX1 U44 ( .A(n32), .Y(n31) );
  INVX1 U45 ( .A(n404), .Y(n34) );
  NOR2X1 U46 ( .A(n52), .B(n47), .Y(n271) );
  OAI21AX1 U47 ( .B(n164), .C(n228), .A(n229), .Y(n197) );
  NAND2X1 U48 ( .A(n242), .B(n271), .Y(n161) );
  NAND3X1 U49 ( .A(n37), .B(n38), .C(n272), .Y(n352) );
  NAND3X1 U50 ( .A(n272), .B(n38), .C(n36), .Y(n328) );
  NAND2X1 U51 ( .A(n165), .B(n271), .Y(n355) );
  OR2X1 U52 ( .A(n240), .B(n47), .Y(n159) );
  INVX1 U53 ( .A(n228), .Y(n55) );
  INVX1 U54 ( .A(sfraddr[0]), .Y(n37) );
  INVX1 U55 ( .A(n244), .Y(n56) );
  NAND2X1 U56 ( .A(n311), .B(n161), .Y(N405) );
  NAND2X1 U57 ( .A(n311), .B(n162), .Y(N332) );
  INVX1 U58 ( .A(n374), .Y(n78) );
  NOR2X1 U59 ( .A(n23), .B(n77), .Y(n342) );
  NAND2X1 U60 ( .A(n81), .B(n374), .Y(n369) );
  NAND2X1 U61 ( .A(n81), .B(n78), .Y(n336) );
  NAND2X1 U62 ( .A(n259), .B(n260), .Y(n253) );
  INVX1 U63 ( .A(n404), .Y(n33) );
  INVX1 U64 ( .A(n441), .Y(n32) );
  NAND42X1 U65 ( .C(n243), .D(sfraddr[1]), .A(n36), .B(n285), .Y(n240) );
  NOR2X1 U66 ( .A(n38), .B(n52), .Y(n285) );
  INVX1 U67 ( .A(sfrwe), .Y(n52) );
  NOR21XL U68 ( .B(sfraddr[1]), .A(n243), .Y(n272) );
  OAI21X1 U69 ( .B(n164), .C(n352), .A(n49), .Y(n158) );
  OAI21X1 U70 ( .B(n164), .C(n244), .A(n49), .Y(n229) );
  OAI21BX1 U71 ( .C(n242), .B(n164), .A(n49), .Y(n288) );
  OAI21BX1 U72 ( .C(n165), .B(n164), .A(n49), .Y(n357) );
  OAI21X1 U73 ( .B(n164), .C(n328), .A(n49), .Y(n313) );
  AOI21AX1 U74 ( .B(sfrwe), .C(n55), .A(n48), .Y(n403) );
  NOR4XL U75 ( .A(n37), .B(n243), .C(sfraddr[1]), .D(sfraddr[2]), .Y(n165) );
  NAND3X1 U76 ( .A(n272), .B(n37), .C(sfraddr[2]), .Y(n244) );
  NOR4XL U77 ( .A(n38), .B(n243), .C(n36), .D(sfraddr[1]), .Y(n242) );
  NOR2X1 U78 ( .A(n47), .B(sfrwe), .Y(n164) );
  NAND3X1 U79 ( .A(n36), .B(n272), .C(sfraddr[2]), .Y(n228) );
  OAI31XL U80 ( .A(n37), .B(sfraddr[1]), .C(n243), .D(n244), .Y(n241) );
  NAND2X1 U81 ( .A(n240), .B(n49), .Y(n274) );
  NAND2X1 U82 ( .A(n403), .B(n85), .Y(n379) );
  OAI31XL U83 ( .A(n56), .B(n55), .C(n165), .D(sfrwe), .Y(n239) );
  NAND3X1 U84 ( .A(n75), .B(n49), .C(n159), .Y(N453) );
  INVX1 U85 ( .A(sfraddr[2]), .Y(n38) );
  NAND2X1 U86 ( .A(n354), .B(n355), .Y(N190) );
  NAND2X1 U87 ( .A(n354), .B(n237), .Y(N258) );
  NAND3X1 U88 ( .A(n75), .B(n48), .C(n6), .Y(N483) );
  NOR2X1 U89 ( .A(n376), .B(n68), .Y(n299) );
  NAND2X1 U90 ( .A(n82), .B(n80), .Y(n374) );
  NAND2X1 U91 ( .A(n78), .B(n262), .Y(n376) );
  NAND2X1 U92 ( .A(n330), .B(n331), .Y(n289) );
  OR2X1 U93 ( .A(n375), .B(n68), .Y(n331) );
  INVX1 U94 ( .A(n262), .Y(n81) );
  INVX1 U95 ( .A(n372), .Y(n72) );
  NOR3XL U96 ( .A(n82), .B(n47), .C(n262), .Y(n260) );
  INVX1 U97 ( .A(n298), .Y(n69) );
  NOR32XL U98 ( .B(n330), .C(n332), .A(n77), .Y(n311) );
  NOR43XL U99 ( .B(n291), .C(n375), .D(n376), .A(n47), .Y(n332) );
  INVX1 U100 ( .A(n380), .Y(n84) );
  INVX1 U101 ( .A(n48), .Y(n47) );
  INVX1 U102 ( .A(n286), .Y(n75) );
  NOR2X1 U103 ( .A(n107), .B(n26), .Y(n259) );
  NAND2X1 U104 ( .A(n27), .B(n260), .Y(n255) );
  NAND2X1 U105 ( .A(n261), .B(n260), .Y(n254) );
  NAND2X1 U106 ( .A(n107), .B(arg_c[0]), .Y(n190) );
  INVX1 U107 ( .A(n195), .Y(n441) );
  INVX1 U108 ( .A(n404), .Y(n442) );
  INVX1 U109 ( .A(n195), .Y(n137) );
  AOI31X1 U110 ( .A(n1), .B(n2), .C(n234), .D(n235), .Y(N802) );
  AOI21AX1 U111 ( .B(n236), .C(n49), .A(n237), .Y(n234) );
  OAI2B11X1 U112 ( .D(sfroe), .C(n238), .A(n239), .B(n240), .Y(n236) );
  NOR4XL U113 ( .A(n241), .B(n242), .C(n54), .D(n53), .Y(n238) );
  NAND4X1 U114 ( .A(n377), .B(n379), .C(n168), .D(n49), .Y(N104) );
  INVX1 U115 ( .A(sfrdatai[0]), .Y(n39) );
  INVX1 U116 ( .A(sfrdatai[5]), .Y(n44) );
  INVX1 U117 ( .A(sfrdatai[3]), .Y(n42) );
  INVX1 U118 ( .A(sfrdatai[1]), .Y(n40) );
  INVX1 U119 ( .A(sfrdatai[4]), .Y(n43) );
  INVX1 U120 ( .A(sfrdatai[2]), .Y(n41) );
  INVX1 U121 ( .A(sfrdatai[7]), .Y(n46) );
  INVX1 U122 ( .A(sfrdatai[6]), .Y(n45) );
  NOR32XL U123 ( .B(n201), .C(n398), .A(n86), .Y(n396) );
  NAND2X1 U124 ( .A(n396), .B(n397), .Y(n262) );
  NOR3XL U125 ( .A(n333), .B(n80), .C(n262), .Y(n286) );
  AOI31X1 U126 ( .A(n81), .B(n333), .C(n80), .D(n286), .Y(n330) );
  INVX1 U127 ( .A(n257), .Y(n80) );
  INVX1 U128 ( .A(n388), .Y(n64) );
  INVX1 U129 ( .A(n294), .Y(n71) );
  NOR2X1 U130 ( .A(n383), .B(n375), .Y(n372) );
  NOR2X1 U131 ( .A(n383), .B(n376), .Y(n28) );
  INVX1 U132 ( .A(n333), .Y(n82) );
  NAND3X1 U133 ( .A(n257), .B(n262), .C(n82), .Y(n291) );
  NAND3X1 U134 ( .A(n262), .B(n333), .C(n80), .Y(n375) );
  NAND2X1 U135 ( .A(n207), .B(n205), .Y(n252) );
  INVX1 U136 ( .A(n392), .Y(n70) );
  NOR2X1 U137 ( .A(n383), .B(n376), .Y(n29) );
  NOR2X1 U138 ( .A(n383), .B(n376), .Y(n298) );
  INVX1 U139 ( .A(n397), .Y(n85) );
  NOR32XL U140 ( .B(n19), .C(n332), .A(n79), .Y(n354) );
  INVX1 U141 ( .A(n209), .Y(n87) );
  INVX1 U142 ( .A(n383), .Y(n68) );
  INVX1 U143 ( .A(rst), .Y(n48) );
  INVX1 U144 ( .A(n214), .Y(n83) );
  INVX1 U145 ( .A(rst), .Y(n49) );
  INVX1 U146 ( .A(n206), .Y(n61) );
  OAI21X1 U147 ( .B(n446), .C(n444), .A(n404), .Y(n195) );
  OAI22X1 U148 ( .A(n9), .B(n109), .C(n190), .D(n110), .Y(arg_c[17]) );
  NOR2X1 U149 ( .A(sum1[17]), .B(n26), .Y(n261) );
  INVX1 U150 ( .A(sum[15]), .Y(n94) );
  INVX1 U151 ( .A(sum[16]), .Y(n93) );
  NAND2X1 U152 ( .A(sum1[17]), .B(arg_c[0]), .Y(n189) );
  INVX1 U153 ( .A(sum1[17]), .Y(n107) );
  NAND2X1 U154 ( .A(n444), .B(n446), .Y(n404) );
  OAI222XL U155 ( .A(n428), .B(n12), .C(n429), .D(n254), .E(n255), .F(n105), 
        .Y(N569) );
  OAI222XL U156 ( .A(n432), .B(n253), .C(n433), .D(n254), .E(n8), .F(n106), 
        .Y(N568) );
  OAI222XL U157 ( .A(n421), .B(n12), .C(n422), .D(n254), .E(n255), .F(n104), 
        .Y(N570) );
  OAI222XL U158 ( .A(n420), .B(n253), .C(n423), .D(n254), .E(n8), .F(n103), 
        .Y(N571) );
  OAI222XL U159 ( .A(n416), .B(n12), .C(n417), .D(n254), .E(n255), .F(n102), 
        .Y(N572) );
  OAI222XL U160 ( .A(n145), .B(n253), .C(n146), .D(n254), .E(n8), .F(n101), 
        .Y(N573) );
  OAI222XL U161 ( .A(n123), .B(n12), .C(n124), .D(n254), .E(n255), .F(n99), 
        .Y(N575) );
  OAI222XL U162 ( .A(n143), .B(n253), .C(n144), .D(n254), .E(n8), .F(n100), 
        .Y(N574) );
  OAI222XL U163 ( .A(n120), .B(n12), .C(n121), .D(n254), .E(n255), .F(n98), 
        .Y(N576) );
  OAI222XL U164 ( .A(n119), .B(n253), .C(n122), .D(n17), .E(n8), .F(n97), .Y(
        N577) );
  OAI222XL U165 ( .A(n117), .B(n12), .C(n118), .D(n17), .E(n255), .F(n96), .Y(
        N578) );
  OAI222XL U166 ( .A(n115), .B(n253), .C(n116), .D(n17), .E(n8), .F(n95), .Y(
        N579) );
  OAI222XL U167 ( .A(n113), .B(n12), .C(n114), .D(n17), .E(n255), .F(n94), .Y(
        N580) );
  OAI222XL U168 ( .A(n111), .B(n253), .C(n112), .D(n17), .E(n8), .F(n93), .Y(
        N581) );
  OAI22X1 U169 ( .A(n40), .B(n159), .C(n280), .D(n274), .Y(N455) );
  AOI222XL U170 ( .A(sum[2]), .B(n27), .C(n15), .D(n281), .E(n20), .F(sum1[1]), 
        .Y(n280) );
  OAI22X1 U171 ( .A(n192), .B(n440), .C(n443), .D(n439), .Y(n281) );
  OAI22X1 U172 ( .A(n39), .B(n159), .C(n282), .D(n274), .Y(N454) );
  AOI22X1 U173 ( .A(n283), .B(n284), .C(sum[1]), .D(n27), .Y(n282) );
  OAI22X1 U174 ( .A(n192), .B(n140), .C(n443), .D(n130), .Y(n284) );
  OR2X1 U175 ( .A(n259), .B(n261), .Y(n283) );
  OAI21X1 U176 ( .B(n8), .C(n129), .A(n258), .Y(N566) );
  AO222X1 U177 ( .A(n130), .B(n257), .C(n140), .D(n80), .E(n17), .F(n253), .Y(
        n258) );
  INVX1 U178 ( .A(n192), .Y(n443) );
  INVX1 U179 ( .A(n193), .Y(n445) );
  INVX1 U180 ( .A(sum[14]), .Y(n95) );
  INVX1 U181 ( .A(sum[13]), .Y(n96) );
  INVX1 U182 ( .A(sum[12]), .Y(n97) );
  INVX1 U183 ( .A(sum[11]), .Y(n98) );
  INVX1 U184 ( .A(sum[9]), .Y(n100) );
  INVX1 U185 ( .A(sum[10]), .Y(n99) );
  INVX1 U186 ( .A(sum[8]), .Y(n101) );
  INVX1 U187 ( .A(sum[6]), .Y(n103) );
  INVX1 U188 ( .A(sum[7]), .Y(n102) );
  INVX1 U189 ( .A(sum[5]), .Y(n104) );
  INVX1 U190 ( .A(sum[3]), .Y(n106) );
  INVX1 U191 ( .A(sum[4]), .Y(n105) );
  NAND21X1 U192 ( .B(n401), .A(n403), .Y(n377) );
  INVX1 U193 ( .A(sum1[2]), .Y(n432) );
  INVX1 U194 ( .A(sum1[3]), .Y(n428) );
  INVX1 U195 ( .A(sum1[4]), .Y(n421) );
  INVX1 U196 ( .A(sum1[5]), .Y(n420) );
  INVX1 U197 ( .A(sum1[6]), .Y(n416) );
  INVX1 U198 ( .A(sum1[7]), .Y(n145) );
  INVX1 U199 ( .A(sum1[8]), .Y(n143) );
  INVX1 U200 ( .A(sum1[9]), .Y(n123) );
  INVX1 U201 ( .A(sum1[10]), .Y(n120) );
  INVX1 U202 ( .A(sum1[11]), .Y(n119) );
  INVX1 U203 ( .A(sum1[12]), .Y(n117) );
  INVX1 U204 ( .A(sum1[13]), .Y(n115) );
  INVX1 U205 ( .A(sum1[14]), .Y(n113) );
  INVX1 U206 ( .A(sum1[15]), .Y(n111) );
  INVX1 U207 ( .A(sum[2]), .Y(n108) );
  INVX1 U208 ( .A(sum1[16]), .Y(n109) );
  OAI222XL U209 ( .A(n377), .B(n386), .C(n247), .D(n379), .E(n21), .F(n42), 
        .Y(N108) );
  OAI222XL U210 ( .A(n377), .B(n60), .C(n249), .D(n379), .E(n168), .F(n40), 
        .Y(N106) );
  INVX1 U211 ( .A(n391), .Y(n60) );
  OAI222XL U212 ( .A(n377), .B(n378), .C(n245), .D(n379), .E(n168), .F(n43), 
        .Y(N109) );
  OAI222XL U213 ( .A(n168), .B(n39), .C(n250), .D(n379), .E(n59), .F(n377), 
        .Y(N105) );
  OAI222XL U214 ( .A(n377), .B(n389), .C(n248), .D(n379), .E(n168), .F(n41), 
        .Y(N107) );
  OAI32X1 U215 ( .A(n125), .B(n47), .C(n50), .D(n168), .E(n44), .Y(n409) );
  OAI211X1 U216 ( .C(n196), .D(n197), .A(n166), .B(n168), .Y(N895) );
  AOI211X1 U217 ( .C(n86), .D(n198), .A(n199), .B(n200), .Y(n196) );
  OAI32X1 U218 ( .A(n201), .B(n440), .C(n202), .D(n404), .E(n203), .Y(n200) );
  OAI222XL U219 ( .A(n204), .B(n205), .C(n206), .D(n207), .E(n208), .F(n209), 
        .Y(n199) );
  OAI211X1 U220 ( .C(n160), .D(n57), .A(n161), .B(n162), .Y(n413) );
  NOR2X1 U221 ( .A(n163), .B(n164), .Y(n160) );
  NOR4XL U222 ( .A(n47), .B(n55), .C(n165), .D(n56), .Y(n163) );
  AOI31X1 U223 ( .A(n217), .B(n218), .C(n219), .D(n197), .Y(N893) );
  AOI22AXL U224 ( .A(n87), .B(n208), .D(n207), .C(n61), .Y(n218) );
  AOI21X1 U225 ( .B(n223), .C(n213), .A(n224), .Y(n217) );
  AOI221XL U226 ( .A(n83), .B(n125), .C(n89), .D(n445), .E(n220), .Y(n219) );
  INVX1 U227 ( .A(sum1[1]), .Y(n434) );
  NAND2X1 U228 ( .A(n192), .B(n193), .Y(arg_c[0]) );
  INVX1 U229 ( .A(sum[1]), .Y(n129) );
  NOR42XL U230 ( .C(n400), .D(n401), .A(n235), .B(n172), .Y(n398) );
  NOR21XL U231 ( .B(n178), .A(n89), .Y(n400) );
  NAND3X1 U232 ( .A(n205), .B(n182), .C(n396), .Y(n257) );
  AOI31X1 U233 ( .A(n394), .B(n331), .C(n262), .D(n380), .Y(n388) );
  AOI21X1 U234 ( .B(n140), .C(n257), .A(n299), .Y(n394) );
  INVX1 U235 ( .A(n203), .Y(n89) );
  OAI31XL U236 ( .A(n92), .B(n91), .C(n88), .D(mdubsy), .Y(n235) );
  NAND2X1 U237 ( .A(n172), .B(n91), .Y(mdubsy) );
  NAND42X1 U238 ( .C(n252), .D(n223), .A(n398), .B(n201), .Y(n333) );
  OAI21X1 U239 ( .B(n140), .C(n291), .A(n72), .Y(n294) );
  OAI31XL U240 ( .A(n393), .B(n28), .C(n372), .D(n84), .Y(n392) );
  NOR3XL U241 ( .A(n140), .B(n81), .C(n80), .Y(n393) );
  NAND2X1 U242 ( .A(n77), .B(n221), .Y(n292) );
  NAND3X1 U243 ( .A(n88), .B(n91), .C(n402), .Y(n201) );
  NAND2X1 U244 ( .A(n395), .B(n402), .Y(n205) );
  INVX1 U245 ( .A(n339), .Y(n65) );
  NAND2X1 U246 ( .A(n399), .B(n91), .Y(n207) );
  INVX1 U247 ( .A(n181), .Y(n86) );
  NOR2X1 U248 ( .A(n249), .B(n246), .Y(N675) );
  NOR2X1 U249 ( .A(n247), .B(n246), .Y(N677) );
  NOR2X1 U250 ( .A(n245), .B(n246), .Y(N678) );
  NOR2X1 U251 ( .A(n248), .B(n246), .Y(N676) );
  AOI21X1 U252 ( .B(n91), .C(n232), .A(n223), .Y(n397) );
  NOR2X1 U253 ( .A(n250), .B(n246), .Y(N674) );
  NAND2X1 U254 ( .A(n382), .B(n216), .Y(n383) );
  NAND3X1 U255 ( .A(n90), .B(n92), .C(n395), .Y(n209) );
  NAND21X1 U256 ( .B(n201), .A(n202), .Y(n214) );
  NAND2X1 U257 ( .A(n222), .B(n73), .Y(n206) );
  AOI31X1 U258 ( .A(n216), .B(n62), .C(n59), .D(n68), .Y(n213) );
  OAI31XL U259 ( .A(n251), .B(n85), .C(n252), .D(n49), .Y(n246) );
  NAND3X1 U260 ( .A(n201), .B(n181), .C(n209), .Y(n251) );
  OAI21X1 U261 ( .B(n231), .C(n62), .A(n384), .Y(n389) );
  NAND2X1 U262 ( .A(n382), .B(n59), .Y(n384) );
  NAND2X1 U263 ( .A(n205), .B(n221), .Y(n220) );
  INVX1 U264 ( .A(n208), .Y(n58) );
  OAI22X1 U265 ( .A(md4[1]), .B(n35), .C(n438), .D(n194), .Y(arg_b[2]) );
  OAI22X1 U266 ( .A(n433), .B(n195), .C(n30), .D(n436), .Y(arg_a[2]) );
  OAI22X1 U267 ( .A(md4[2]), .B(n35), .C(n430), .D(n194), .Y(arg_b[3]) );
  OAI22X1 U268 ( .A(n429), .B(n195), .C(n30), .D(n431), .Y(arg_a[3]) );
  OAI22X1 U269 ( .A(md4[3]), .B(n35), .C(n425), .D(n194), .Y(arg_b[4]) );
  OAI22X1 U270 ( .A(n422), .B(n195), .C(n30), .D(n427), .Y(arg_a[4]) );
  OAI22X1 U271 ( .A(md4[4]), .B(n35), .C(n424), .D(n194), .Y(arg_b[5]) );
  OAI22X1 U272 ( .A(n423), .B(n195), .C(n30), .D(n426), .Y(arg_a[5]) );
  OAI22X1 U273 ( .A(md4[5]), .B(n35), .C(n418), .D(n194), .Y(arg_b[6]) );
  OAI22X1 U274 ( .A(n417), .B(n195), .C(n31), .D(n419), .Y(arg_a[6]) );
  OAI22X1 U275 ( .A(md4[2]), .B(n33), .C(n188), .D(n430), .Y(arg_d[3]) );
  OAI222XL U276 ( .A(n9), .B(n432), .C(n190), .D(n433), .E(n137), .F(n421), 
        .Y(arg_c[3]) );
  OAI22X1 U277 ( .A(md4[6]), .B(n35), .C(n153), .D(n194), .Y(arg_b[7]) );
  OAI22X1 U278 ( .A(n146), .B(n195), .C(n31), .D(n156), .Y(arg_a[7]) );
  OAI22X1 U279 ( .A(md4[3]), .B(n33), .C(n188), .D(n425), .Y(arg_d[4]) );
  OAI222XL U280 ( .A(n189), .B(n428), .C(n11), .D(n429), .E(n137), .F(n420), 
        .Y(arg_c[4]) );
  OAI22X1 U281 ( .A(md4[7]), .B(n35), .C(n415), .D(n194), .Y(arg_b[8]) );
  OAI22X1 U282 ( .A(n144), .B(n195), .C(n441), .D(n157), .Y(arg_a[8]) );
  OAI22X1 U283 ( .A(md4[4]), .B(n33), .C(n188), .D(n424), .Y(arg_d[5]) );
  OAI222XL U284 ( .A(n9), .B(n421), .C(n190), .D(n422), .E(n137), .F(n416), 
        .Y(arg_c[5]) );
  OAI22X1 U285 ( .A(md5[0]), .B(n34), .C(n139), .D(n194), .Y(arg_b[9]) );
  OAI22X1 U286 ( .A(n124), .B(n195), .C(n441), .D(n135), .Y(arg_a[9]) );
  OAI22X1 U287 ( .A(md4[5]), .B(n33), .C(n188), .D(n418), .Y(arg_d[6]) );
  OAI222XL U288 ( .A(n189), .B(n420), .C(n11), .D(n423), .E(n137), .F(n145), 
        .Y(arg_c[6]) );
  OAI22X1 U289 ( .A(md5[1]), .B(n33), .C(n407), .D(n14), .Y(arg_b[10]) );
  OAI22X1 U290 ( .A(n121), .B(n24), .C(n30), .D(n155), .Y(arg_a[10]) );
  OAI22X1 U291 ( .A(md4[6]), .B(n34), .C(n188), .D(n153), .Y(arg_d[7]) );
  OAI222XL U292 ( .A(n9), .B(n416), .C(n190), .D(n417), .E(n137), .F(n143), 
        .Y(arg_c[7]) );
  OAI22X1 U293 ( .A(md5[2]), .B(n442), .C(n141), .D(n14), .Y(arg_b[11]) );
  OAI22X1 U294 ( .A(n122), .B(n24), .C(n30), .D(n134), .Y(arg_a[11]) );
  OAI22X1 U295 ( .A(md4[7]), .B(n33), .C(n188), .D(n415), .Y(arg_d[8]) );
  OAI222XL U296 ( .A(n189), .B(n145), .C(n11), .D(n146), .E(n137), .F(n123), 
        .Y(arg_c[8]) );
  OAI22X1 U297 ( .A(md5[3]), .B(n442), .C(n152), .D(n14), .Y(arg_b[12]) );
  OAI22X1 U298 ( .A(n118), .B(n24), .C(n30), .D(n406), .Y(arg_a[12]) );
  OAI22X1 U299 ( .A(md5[0]), .B(n34), .C(n188), .D(n139), .Y(arg_d[9]) );
  OAI222XL U300 ( .A(n9), .B(n143), .C(n190), .D(n144), .E(n441), .F(n120), 
        .Y(arg_c[9]) );
  OAI22X1 U301 ( .A(md5[4]), .B(n442), .C(n154), .D(n14), .Y(arg_b[13]) );
  OAI22X1 U302 ( .A(n116), .B(n24), .C(n30), .D(n147), .Y(arg_a[13]) );
  OAI22X1 U303 ( .A(md5[1]), .B(n34), .C(n18), .D(n407), .Y(arg_d[10]) );
  OAI222XL U304 ( .A(n189), .B(n123), .C(n11), .D(n124), .E(n441), .F(n119), 
        .Y(arg_c[10]) );
  ENOX1 U305 ( .A(n114), .B(n24), .C(n24), .D(md3[5]), .Y(arg_a[14]) );
  OAI22X1 U306 ( .A(md5[5]), .B(n442), .C(n405), .D(n14), .Y(arg_b[14]) );
  OAI22X1 U307 ( .A(md5[2]), .B(n34), .C(n18), .D(n141), .Y(arg_d[11]) );
  OAI222XL U308 ( .A(n9), .B(n120), .C(n190), .D(n121), .E(n441), .F(n117), 
        .Y(arg_c[11]) );
  OAI22X1 U309 ( .A(md5[6]), .B(n35), .C(n138), .D(n14), .Y(arg_b[15]) );
  OAI22X1 U310 ( .A(n112), .B(n24), .C(n30), .D(n140), .Y(arg_a[15]) );
  OAI22X1 U311 ( .A(md5[3]), .B(n34), .C(n18), .D(n152), .Y(arg_d[12]) );
  OAI222XL U312 ( .A(n189), .B(n119), .C(n11), .D(n122), .E(n441), .F(n115), 
        .Y(arg_c[12]) );
  OAI22X1 U313 ( .A(md5[4]), .B(n34), .C(n18), .D(n154), .Y(arg_d[13]) );
  OAI222XL U314 ( .A(n9), .B(n117), .C(n190), .D(n118), .E(n441), .F(n113), 
        .Y(arg_c[13]) );
  OAI22X1 U315 ( .A(md5[5]), .B(n34), .C(n18), .D(n405), .Y(arg_d[14]) );
  OAI222XL U316 ( .A(n189), .B(n115), .C(n11), .D(n116), .E(n441), .F(n111), 
        .Y(arg_c[14]) );
  OAI22X1 U317 ( .A(md5[6]), .B(n34), .C(n18), .D(n138), .Y(arg_d[15]) );
  OAI222XL U318 ( .A(n9), .B(n113), .C(n190), .D(n114), .E(n31), .F(n109), .Y(
        arg_c[15]) );
  OAI22X1 U319 ( .A(md4[0]), .B(n35), .C(n437), .D(n194), .Y(arg_b[1]) );
  OAI21X1 U320 ( .B(n31), .C(n435), .A(n191), .Y(arg_a[1]) );
  NOR21XL U321 ( .B(norm_reg[15]), .A(n24), .Y(arg_a[17]) );
  OAI22X1 U322 ( .A(md5[7]), .B(n35), .C(n136), .D(n14), .Y(arg_b[16]) );
  OAI22X1 U323 ( .A(n110), .B(n24), .C(n30), .D(n440), .Y(arg_a[16]) );
  OAI22X1 U324 ( .A(md5[7]), .B(n34), .C(n18), .D(n136), .Y(arg_d[16]) );
  OAI222XL U325 ( .A(n189), .B(n111), .C(n11), .D(n112), .E(n31), .F(n107), 
        .Y(arg_c[16]) );
  NAND2X1 U326 ( .A(md0[0]), .B(n33), .Y(n194) );
  NAND2X1 U327 ( .A(mdu_op[1]), .B(n444), .Y(n192) );
  OAI22X1 U328 ( .A(md4[1]), .B(n33), .C(n188), .D(n438), .Y(arg_d[2]) );
  OAI222XL U329 ( .A(n189), .B(n434), .C(sum1[17]), .D(n191), .E(n137), .F(
        n428), .Y(arg_c[2]) );
  NAND2X1 U330 ( .A(mdu_op[0]), .B(n446), .Y(n193) );
  OAI222XL U331 ( .A(n434), .B(n12), .C(n256), .D(n17), .E(n255), .F(n108), 
        .Y(N567) );
  AOI22X1 U332 ( .A(n80), .B(md3[7]), .C(md1[7]), .D(n257), .Y(n256) );
  AOI22X1 U333 ( .A(n443), .B(md3[7]), .C(n445), .D(md1[7]), .Y(n191) );
  OAI22X1 U334 ( .A(n39), .B(n355), .C(n373), .D(n357), .Y(N191) );
  AOI222XL U335 ( .A(n29), .B(md0[1]), .C(md0[2]), .D(n67), .E(n79), .F(
        sum[17]), .Y(n373) );
  OAI22X1 U336 ( .A(n41), .B(n159), .C(n279), .D(n274), .Y(N456) );
  AOI222XL U337 ( .A(sum[3]), .B(sum[17]), .C(n261), .D(norm_reg[0]), .E(n259), 
        .F(sum1[2]), .Y(n279) );
  OAI22X1 U338 ( .A(n42), .B(n159), .C(n278), .D(n274), .Y(N457) );
  AOI222XL U339 ( .A(sum[4]), .B(n27), .C(n15), .D(norm_reg[1]), .E(n20), .F(
        sum1[3]), .Y(n278) );
  OAI22X1 U340 ( .A(n43), .B(n159), .C(n277), .D(n274), .Y(N458) );
  AOI222XL U341 ( .A(sum[5]), .B(sum[17]), .C(n261), .D(norm_reg[2]), .E(n259), 
        .F(sum1[4]), .Y(n277) );
  OAI22X1 U342 ( .A(n44), .B(n159), .C(n276), .D(n274), .Y(N459) );
  AOI222XL U343 ( .A(sum[6]), .B(n27), .C(n15), .D(norm_reg[3]), .E(n20), .F(
        sum1[5]), .Y(n276) );
  OAI22X1 U344 ( .A(n46), .B(n159), .C(n273), .D(n274), .Y(N461) );
  AOI222XL U345 ( .A(sum[8]), .B(sum[17]), .C(n261), .D(norm_reg[5]), .E(n259), 
        .F(sum1[7]), .Y(n273) );
  OAI22X1 U346 ( .A(n166), .B(n40), .C(n269), .D(n229), .Y(N485) );
  AOI222XL U347 ( .A(sum[10]), .B(n27), .C(n15), .D(norm_reg[7]), .E(n20), .F(
        sum1[9]), .Y(n269) );
  OAI22X1 U348 ( .A(n166), .B(n44), .C(n265), .D(n229), .Y(N489) );
  AOI222XL U349 ( .A(sum[14]), .B(sum[17]), .C(n261), .D(norm_reg[11]), .E(
        n259), .F(sum1[13]), .Y(n265) );
  OAI22X1 U350 ( .A(n166), .B(n43), .C(n266), .D(n229), .Y(N488) );
  AOI222XL U351 ( .A(sum[13]), .B(n27), .C(n15), .D(norm_reg[10]), .E(n20), 
        .F(sum1[12]), .Y(n266) );
  OAI22X1 U352 ( .A(n45), .B(n159), .C(n275), .D(n274), .Y(N460) );
  AOI222XL U353 ( .A(sum[7]), .B(sum[17]), .C(n15), .D(norm_reg[4]), .E(n20), 
        .F(sum1[6]), .Y(n275) );
  OAI22X1 U354 ( .A(n166), .B(n42), .C(n267), .D(n229), .Y(N487) );
  AOI222XL U355 ( .A(sum[12]), .B(sum[17]), .C(n261), .D(norm_reg[9]), .E(n259), .F(sum1[11]), .Y(n267) );
  OAI22X1 U356 ( .A(n166), .B(n41), .C(n268), .D(n229), .Y(N486) );
  AOI222XL U357 ( .A(sum[11]), .B(n27), .C(n15), .D(norm_reg[8]), .E(n20), .F(
        sum1[10]), .Y(n268) );
  OAI22X1 U358 ( .A(n6), .B(n39), .C(n270), .D(n229), .Y(N484) );
  AOI222XL U359 ( .A(sum[9]), .B(sum[17]), .C(n261), .D(norm_reg[6]), .E(n259), 
        .F(sum1[8]), .Y(n270) );
  OAI22X1 U360 ( .A(n6), .B(n45), .C(n264), .D(n229), .Y(N490) );
  AOI222XL U361 ( .A(sum[15]), .B(n27), .C(n15), .D(norm_reg[12]), .E(n20), 
        .F(sum1[14]), .Y(n264) );
  OAI22X1 U362 ( .A(n6), .B(n46), .C(n263), .D(n229), .Y(N491) );
  AOI222XL U363 ( .A(sum[16]), .B(sum[17]), .C(n261), .D(norm_reg[13]), .E(
        n259), .F(sum1[15]), .Y(n263) );
  OAI22X1 U364 ( .A(n44), .B(n161), .C(n297), .D(n288), .Y(N411) );
  AOI221XL U365 ( .A(n28), .B(md3[6]), .C(n299), .D(md3[7]), .E(n300), .Y(n297) );
  OAI222XL U366 ( .A(n296), .B(n406), .C(n71), .D(n147), .E(n94), .F(n292), 
        .Y(n300) );
  OAI22X1 U367 ( .A(n45), .B(n1), .C(n293), .D(n288), .Y(N412) );
  AOI221XL U368 ( .A(md3[5]), .B(n22), .C(md3[4]), .D(n66), .E(n295), .Y(n293)
         );
  INVX1 U369 ( .A(n296), .Y(n66) );
  OAI22X1 U370 ( .A(n440), .B(n69), .C(n93), .D(n19), .Y(n295) );
  INVX1 U371 ( .A(mdu_op[0]), .Y(n444) );
  OAI22X1 U372 ( .A(n46), .B(n161), .C(n287), .D(n288), .Y(N413) );
  AOI221XL U373 ( .A(md3[5]), .B(n289), .C(n76), .D(n26), .E(n290), .Y(n287)
         );
  INVX1 U374 ( .A(n292), .Y(n76) );
  OAI22X1 U375 ( .A(n179), .B(n291), .C(n140), .D(n72), .Y(n290) );
  INVX1 U376 ( .A(mdu_op[1]), .Y(n446) );
  OAI22X1 U377 ( .A(n43), .B(n1), .C(n301), .D(n288), .Y(N410) );
  AOI221XL U378 ( .A(n298), .B(md3[5]), .C(n23), .D(md3[6]), .E(n302), .Y(n301) );
  OAI222XL U379 ( .A(n296), .B(n134), .C(n71), .D(n406), .E(n95), .F(n292), 
        .Y(n302) );
  INVX1 U380 ( .A(md2[0]), .Y(n435) );
  INVX1 U381 ( .A(md4[0]), .Y(n437) );
  OAI22X1 U382 ( .A(n41), .B(n161), .C(n305), .D(n288), .Y(N408) );
  AOI221XL U383 ( .A(n28), .B(md3[3]), .C(n299), .D(md3[4]), .E(n306), .Y(n305) );
  OAI222XL U384 ( .A(n296), .B(n135), .C(n71), .D(n155), .E(n97), .F(n292), 
        .Y(n306) );
  OAI22X1 U385 ( .A(n42), .B(n1), .C(n303), .D(n288), .Y(N409) );
  AOI221XL U386 ( .A(n29), .B(md3[4]), .C(n23), .D(md3[5]), .E(n304), .Y(n303)
         );
  OAI222XL U387 ( .A(n296), .B(n155), .C(n71), .D(n134), .E(n96), .F(n292), 
        .Y(n304) );
  INVX1 U388 ( .A(md2[1]), .Y(n436) );
  INVX1 U389 ( .A(md4[1]), .Y(n438) );
  INVX1 U390 ( .A(norm_reg[0]), .Y(n433) );
  OAI22X1 U391 ( .A(n40), .B(n161), .C(n307), .D(n288), .Y(N407) );
  AOI221XL U392 ( .A(n29), .B(md3[2]), .C(n299), .D(md3[3]), .E(n308), .Y(n307) );
  OAI222XL U393 ( .A(n296), .B(n157), .C(n71), .D(n135), .E(n98), .F(n292), 
        .Y(n308) );
  INVX1 U394 ( .A(md2[3]), .Y(n427) );
  INVX1 U395 ( .A(md2[2]), .Y(n431) );
  INVX1 U396 ( .A(md4[3]), .Y(n425) );
  INVX1 U397 ( .A(md4[2]), .Y(n430) );
  INVX1 U398 ( .A(norm_reg[1]), .Y(n429) );
  INVX1 U399 ( .A(norm_reg[2]), .Y(n422) );
  OAI22X1 U400 ( .A(n46), .B(n162), .C(n312), .D(n313), .Y(N340) );
  AOI221XL U401 ( .A(n29), .B(md3[0]), .C(n299), .D(md3[1]), .E(n314), .Y(n312) );
  OAI222XL U402 ( .A(n296), .B(n419), .C(n71), .D(n156), .E(n100), .F(n292), 
        .Y(n314) );
  OAI22X1 U403 ( .A(n39), .B(n1), .C(n309), .D(n288), .Y(N406) );
  AOI221XL U404 ( .A(n28), .B(md3[1]), .C(n23), .D(md3[2]), .E(n310), .Y(n309)
         );
  OAI222XL U405 ( .A(n296), .B(n156), .C(n71), .D(n157), .E(n99), .F(n292), 
        .Y(n310) );
  INVX1 U406 ( .A(md2[4]), .Y(n426) );
  INVX1 U407 ( .A(md4[4]), .Y(n424) );
  INVX1 U408 ( .A(norm_reg[3]), .Y(n423) );
  OAI22X1 U409 ( .A(n45), .B(n2), .C(n315), .D(n313), .Y(N339) );
  AOI221XL U410 ( .A(n28), .B(md2[7]), .C(n23), .D(md3[0]), .E(n316), .Y(n315)
         );
  OAI222XL U411 ( .A(n296), .B(n426), .C(n71), .D(n419), .E(n101), .F(n292), 
        .Y(n316) );
  INVX1 U412 ( .A(md2[5]), .Y(n419) );
  INVX1 U413 ( .A(md2[6]), .Y(n156) );
  INVX1 U414 ( .A(md4[5]), .Y(n418) );
  INVX1 U415 ( .A(md4[6]), .Y(n153) );
  INVX1 U416 ( .A(norm_reg[4]), .Y(n417) );
  INVX1 U417 ( .A(norm_reg[5]), .Y(n146) );
  OAI22X1 U418 ( .A(n43), .B(n162), .C(n319), .D(n313), .Y(N337) );
  AOI221XL U419 ( .A(n28), .B(md2[5]), .C(n299), .D(md2[6]), .E(n320), .Y(n319) );
  OAI222XL U420 ( .A(n296), .B(n431), .C(n71), .D(n427), .E(n103), .F(n292), 
        .Y(n320) );
  OAI22X1 U421 ( .A(n44), .B(n2), .C(n317), .D(n313), .Y(N338) );
  AOI221XL U422 ( .A(n29), .B(md2[6]), .C(n23), .D(md2[7]), .E(n318), .Y(n317)
         );
  OAI222XL U423 ( .A(n7), .B(n427), .C(n71), .D(n426), .E(n102), .F(n19), .Y(
        n318) );
  INVX1 U424 ( .A(md2[7]), .Y(n157) );
  INVX1 U425 ( .A(md4[7]), .Y(n415) );
  INVX1 U426 ( .A(norm_reg[6]), .Y(n144) );
  OAI22X1 U427 ( .A(n42), .B(n162), .C(n321), .D(n313), .Y(N336) );
  AOI221XL U428 ( .A(n29), .B(md2[4]), .C(n299), .D(md2[5]), .E(n322), .Y(n321) );
  OAI222XL U429 ( .A(n7), .B(n436), .C(n13), .D(n431), .E(n104), .F(n19), .Y(
        n322) );
  INVX1 U430 ( .A(md3[0]), .Y(n135) );
  INVX1 U431 ( .A(md3[1]), .Y(n155) );
  INVX1 U432 ( .A(md5[0]), .Y(n139) );
  INVX1 U433 ( .A(md5[1]), .Y(n407) );
  INVX1 U434 ( .A(norm_reg[7]), .Y(n124) );
  INVX1 U435 ( .A(norm_reg[8]), .Y(n121) );
  OAI22X1 U436 ( .A(n40), .B(n2), .C(n325), .D(n313), .Y(N334) );
  AOI221XL U437 ( .A(n29), .B(md2[2]), .C(n23), .D(md2[3]), .E(n326), .Y(n325)
         );
  OAI222XL U438 ( .A(n7), .B(n439), .C(n13), .D(n435), .E(n106), .F(n19), .Y(
        n326) );
  OAI22X1 U439 ( .A(n41), .B(n162), .C(n323), .D(n313), .Y(N335) );
  AOI221XL U440 ( .A(n28), .B(md2[3]), .C(n299), .D(md2[4]), .E(n324), .Y(n323) );
  OAI222XL U441 ( .A(n7), .B(n435), .C(n13), .D(n436), .E(n105), .F(n19), .Y(
        n324) );
  INVX1 U442 ( .A(md3[2]), .Y(n134) );
  INVX1 U443 ( .A(md5[2]), .Y(n141) );
  INVX1 U444 ( .A(norm_reg[9]), .Y(n122) );
  OAI22X1 U445 ( .A(md4[0]), .B(n33), .C(n188), .D(n437), .Y(arg_d[1]) );
  OAI222XL U446 ( .A(n192), .B(n140), .C(n193), .D(n130), .E(n137), .F(n432), 
        .Y(arg_c[1]) );
  OAI22X1 U447 ( .A(n39), .B(n2), .C(n327), .D(n313), .Y(N333) );
  AOI221XL U448 ( .A(n28), .B(md2[1]), .C(n23), .D(md2[2]), .E(n329), .Y(n327)
         );
  OAI222XL U449 ( .A(n7), .B(n130), .C(n13), .D(n439), .E(n108), .F(n19), .Y(
        n329) );
  OAI22X1 U450 ( .A(n44), .B(n355), .C(n361), .D(n357), .Y(N196) );
  AOI221XL U451 ( .A(md0[4]), .B(n294), .C(md0[3]), .D(n339), .E(n362), .Y(
        n361) );
  OAI22X1 U452 ( .A(n69), .B(n131), .C(n342), .D(n132), .Y(n362) );
  OAI22X1 U453 ( .A(n43), .B(n355), .C(n363), .D(n357), .Y(N195) );
  AOI221XL U454 ( .A(md0[3]), .B(n294), .C(md0[2]), .D(n339), .E(n364), .Y(
        n363) );
  OAI22X1 U455 ( .A(n69), .B(n151), .C(n342), .D(n131), .Y(n364) );
  OAI22X1 U456 ( .A(n42), .B(n355), .C(n365), .D(n357), .Y(N194) );
  AOI221XL U457 ( .A(md0[2]), .B(n22), .C(md0[1]), .D(n339), .E(n366), .Y(n365) );
  OAI22X1 U458 ( .A(n69), .B(n150), .C(n342), .D(n151), .Y(n366) );
  OAI22X1 U459 ( .A(n40), .B(n355), .C(n370), .D(n357), .Y(N192) );
  AOI221XL U460 ( .A(md0[0]), .B(n22), .C(md0[3]), .D(n67), .E(n371), .Y(n370)
         );
  ENOX1 U461 ( .A(n107), .B(n369), .C(n29), .D(md0[2]), .Y(n371) );
  OAI22X1 U462 ( .A(n46), .B(n355), .C(n356), .D(n357), .Y(N198) );
  AOI221XL U463 ( .A(md0[6]), .B(n22), .C(md0[5]), .D(n16), .E(n358), .Y(n356)
         );
  OAI22X1 U464 ( .A(n5), .B(n128), .C(n10), .D(n148), .Y(n358) );
  OAI22X1 U465 ( .A(n45), .B(n355), .C(n359), .D(n357), .Y(N197) );
  AOI221XL U466 ( .A(md0[5]), .B(n22), .C(md0[4]), .D(n16), .E(n360), .Y(n359)
         );
  OAI22X1 U467 ( .A(n5), .B(n132), .C(n10), .D(n128), .Y(n360) );
  OAI22X1 U468 ( .A(n41), .B(n355), .C(n367), .D(n357), .Y(N193) );
  AOI221XL U469 ( .A(md0[1]), .B(n22), .C(md0[0]), .D(n16), .E(n368), .Y(n367)
         );
  ENOX1 U470 ( .A(n10), .B(n150), .C(n29), .D(md0[3]), .Y(n368) );
  OAI22X1 U471 ( .A(n46), .B(n237), .C(n334), .D(n158), .Y(N266) );
  AOI221XL U472 ( .A(n29), .B(md2[0]), .C(n299), .D(md2[1]), .E(n335), .Y(n334) );
  OAI222XL U473 ( .A(n65), .B(n126), .C(n13), .D(n130), .E(n129), .F(n336), 
        .Y(n335) );
  OAI22X1 U474 ( .A(n42), .B(n237), .C(n345), .D(n158), .Y(N262) );
  AOI221XL U475 ( .A(md1[2]), .B(n294), .C(md1[1]), .D(n339), .E(n346), .Y(
        n345) );
  OAI22X1 U476 ( .A(n69), .B(n133), .C(n342), .D(n126), .Y(n346) );
  OAI22X1 U477 ( .A(n40), .B(n237), .C(n349), .D(n158), .Y(N260) );
  AOI221XL U478 ( .A(md1[0]), .B(n294), .C(md0[7]), .D(n339), .E(n350), .Y(
        n349) );
  OAI22X1 U479 ( .A(n69), .B(n127), .C(n342), .D(n149), .Y(n350) );
  OAI22X1 U480 ( .A(n43), .B(n237), .C(n343), .D(n158), .Y(N263) );
  AOI221XL U481 ( .A(md1[3]), .B(n294), .C(md1[2]), .D(n339), .E(n344), .Y(
        n343) );
  OAI22X1 U482 ( .A(n69), .B(n126), .C(n342), .D(n130), .Y(n344) );
  OAI22X1 U483 ( .A(n45), .B(n237), .C(n337), .D(n158), .Y(N265) );
  AOI221XL U484 ( .A(n28), .B(md1[7]), .C(n23), .D(md2[0]), .E(n338), .Y(n337)
         );
  OAI222XL U485 ( .A(n65), .B(n133), .C(n13), .D(n126), .E(n434), .F(n336), 
        .Y(n338) );
  OAI22X1 U486 ( .A(n39), .B(n237), .C(n351), .D(n158), .Y(N259) );
  AOI221XL U487 ( .A(md0[7]), .B(n294), .C(md0[6]), .D(n339), .E(n353), .Y(
        n351) );
  OAI22X1 U488 ( .A(n69), .B(n148), .C(n342), .D(n127), .Y(n353) );
  OAI22X1 U489 ( .A(n41), .B(n237), .C(n347), .D(n158), .Y(N261) );
  AOI221XL U490 ( .A(md1[1]), .B(n294), .C(md1[0]), .D(n339), .E(n348), .Y(
        n347) );
  OAI22X1 U491 ( .A(n69), .B(n149), .C(n342), .D(n133), .Y(n348) );
  OAI22X1 U492 ( .A(n44), .B(n237), .C(n340), .D(n158), .Y(N264) );
  AOI221XL U493 ( .A(md1[4]), .B(n294), .C(md1[3]), .D(n339), .E(n341), .Y(
        n340) );
  OAI22X1 U494 ( .A(n130), .B(n69), .C(n342), .D(n439), .Y(n341) );
  OAI21BX1 U495 ( .C(set_div16), .B(n158), .A(n159), .Y(n414) );
  OAI31XL U496 ( .A(n444), .B(n47), .C(n51), .D(n169), .Y(n411) );
  AOI31X1 U497 ( .A(set_div16), .B(n57), .C(n51), .D(n50), .Y(n169) );
  INVX1 U498 ( .A(n166), .Y(n51) );
  OAI211X1 U499 ( .C(n57), .D(n166), .A(n167), .B(n168), .Y(n412) );
  NAND3X1 U500 ( .A(n166), .B(n48), .C(mdu_op[1]), .Y(n167) );
  OAI211X1 U501 ( .C(n210), .D(n197), .A(n166), .B(n168), .Y(N894) );
  AOI211X1 U502 ( .C(n89), .D(n444), .A(n211), .B(n212), .Y(n210) );
  OAI221X1 U503 ( .A(n181), .B(n198), .C(n61), .D(n207), .E(n214), .Y(n211) );
  ENOX1 U504 ( .A(md3[7]), .B(n201), .C(n85), .D(n213), .Y(n212) );
  AOI31X1 U505 ( .A(n225), .B(n226), .C(n227), .D(n197), .Y(N892) );
  NAND21X1 U506 ( .B(n205), .A(n204), .Y(n226) );
  AOI32X1 U507 ( .A(n232), .B(n91), .C(n213), .D(n83), .E(arcon[5]), .Y(n225)
         );
  AOI221XL U508 ( .A(n87), .B(n58), .C(n89), .D(n192), .E(n224), .Y(n227) );
  INVX1 U509 ( .A(md3[3]), .Y(n406) );
  INVX1 U510 ( .A(md3[4]), .Y(n147) );
  INVX1 U511 ( .A(norm_reg[10]), .Y(n118) );
  INVX1 U512 ( .A(norm_reg[11]), .Y(n116) );
  INVX1 U513 ( .A(md5[3]), .Y(n152) );
  INVX1 U514 ( .A(md5[4]), .Y(n154) );
  INVX1 U515 ( .A(md5[5]), .Y(n405) );
  INVX1 U516 ( .A(norm_reg[12]), .Y(n114) );
  INVX1 U517 ( .A(md3[6]), .Y(n140) );
  AOI211X1 U518 ( .C(sfroe), .D(n55), .A(n170), .B(n47), .Y(n410) );
  NOR2X1 U519 ( .A(arcon[7]), .B(test_so), .Y(n170) );
  INVX1 U520 ( .A(md3[7]), .Y(n440) );
  INVX1 U521 ( .A(md5[7]), .Y(n136) );
  INVX1 U522 ( .A(md5[6]), .Y(n138) );
  INVX1 U523 ( .A(norm_reg[13]), .Y(n112) );
  INVX1 U524 ( .A(norm_reg[14]), .Y(n110) );
  NAND2X1 U525 ( .A(md0[1]), .B(n33), .Y(n188) );
  INVX1 U526 ( .A(md1[6]), .Y(n130) );
  AOI21BBXL U527 ( .B(md3[6]), .C(n291), .A(n289), .Y(n296) );
  AOI221XL U528 ( .A(n378), .B(n70), .C(n380), .D(arcon[4]), .E(n63), .Y(n245)
         );
  INVX1 U529 ( .A(n381), .Y(n63) );
  GEN2XL U530 ( .D(n382), .E(n74), .C(n73), .B(n383), .A(n64), .Y(n381) );
  NAND2X1 U531 ( .A(n399), .B(oper_reg[3]), .Y(n203) );
  NOR3XL U532 ( .A(oper_reg[0]), .B(oper_reg[1]), .C(n92), .Y(n399) );
  NOR3XL U533 ( .A(oper_reg[1]), .B(oper_reg[2]), .C(oper_reg[0]), .Y(n172) );
  NOR2X1 U534 ( .A(n90), .B(oper_reg[2]), .Y(n402) );
  INVX1 U535 ( .A(oper_reg[0]), .Y(n90) );
  INVX1 U536 ( .A(oper_reg[2]), .Y(n92) );
  NAND3X1 U537 ( .A(oper_reg[3]), .B(n88), .C(n402), .Y(n178) );
  OAI211X1 U538 ( .C(md3[6]), .D(n291), .A(n331), .B(n369), .Y(n339) );
  OA222X1 U539 ( .A(counter_st[1]), .B(n64), .C(n391), .D(n392), .E(n84), .F(
        n142), .Y(n249) );
  NAND3X1 U540 ( .A(n395), .B(oper_reg[0]), .C(oper_reg[2]), .Y(n181) );
  AOI222XL U541 ( .A(n389), .B(n70), .C(n390), .D(n388), .E(n380), .F(arcon[2]), .Y(n248) );
  AO21X1 U542 ( .B(counter_st[2]), .C(counter_st[1]), .A(n382), .Y(n390) );
  AOI222XL U543 ( .A(n388), .B(N610), .C(n59), .D(n70), .E(n380), .F(arcon[0]), 
        .Y(n250) );
  AOI222XL U544 ( .A(n386), .B(n70), .C(n387), .D(n388), .E(n380), .F(arcon[3]), .Y(n247) );
  XNOR2XL U545 ( .A(n74), .B(n382), .Y(n387) );
  INVX1 U546 ( .A(oper_reg[3]), .Y(n91) );
  NOR2X1 U547 ( .A(n88), .B(oper_reg[3]), .Y(n395) );
  INVX1 U548 ( .A(oper_reg[1]), .Y(n88) );
  NAND3X1 U549 ( .A(n402), .B(oper_reg[3]), .C(oper_reg[1]), .Y(n401) );
  AND3X1 U550 ( .A(n395), .B(n90), .C(oper_reg[2]), .Y(n223) );
  NOR3XL U551 ( .A(n90), .B(oper_reg[1]), .C(n92), .Y(n232) );
  NAND3X1 U552 ( .A(n90), .B(n92), .C(oper_reg[3]), .Y(n182) );
  NOR2X1 U553 ( .A(counter_st[2]), .B(counter_st[1]), .Y(n382) );
  NOR2X1 U554 ( .A(counter_st[3]), .B(counter_st[4]), .Y(n216) );
  AND3X1 U555 ( .A(n231), .B(n74), .C(counter_st[2]), .Y(n222) );
  NAND2X1 U556 ( .A(n232), .B(oper_reg[3]), .Y(n221) );
  NOR2X1 U557 ( .A(counter_st[1]), .B(N610), .Y(n231) );
  NAND2X1 U558 ( .A(n179), .B(n215), .Y(n198) );
  NAND4X1 U559 ( .A(counter_st[1]), .B(n216), .C(n59), .D(n62), .Y(n215) );
  NAND42X1 U560 ( .C(arcon[0]), .D(arcon[2]), .A(n142), .B(n233), .Y(n202) );
  NOR2X1 U561 ( .A(arcon[4]), .B(arcon[3]), .Y(n233) );
  AOI21X1 U562 ( .B(counter_st[1]), .C(N610), .A(n231), .Y(n391) );
  XNOR2XL U563 ( .A(n384), .B(counter_st[3]), .Y(n386) );
  NAND4X1 U564 ( .A(counter_st[4]), .B(counter_st[1]), .C(n230), .D(n59), .Y(
        n208) );
  NOR2X1 U565 ( .A(counter_st[3]), .B(counter_st[2]), .Y(n230) );
  OAI22AX1 U566 ( .D(n216), .C(n384), .A(n385), .B(n73), .Y(n378) );
  NOR2X1 U567 ( .A(counter_st[3]), .B(n384), .Y(n385) );
  INVX1 U568 ( .A(N610), .Y(n59) );
  OAI31XL U569 ( .A(n201), .B(md3[7]), .C(n202), .D(n181), .Y(n224) );
  NOR2X1 U570 ( .A(md3[6]), .B(md3[5]), .Y(n179) );
  NOR42XL U571 ( .C(n435), .D(n179), .A(md2[1]), .B(n180), .Y(n177) );
  NAND4X1 U572 ( .A(n431), .B(n427), .C(n426), .D(n419), .Y(n180) );
  NOR4XL U573 ( .A(md3[1]), .B(md3[0]), .C(md2[7]), .D(md2[6]), .Y(n175) );
  NOR4XL U574 ( .A(md3[7]), .B(md3[4]), .C(md3[3]), .D(md3[2]), .Y(n176) );
  NOR4XL U575 ( .A(md4[2]), .B(md4[1]), .C(md4[0]), .D(n182), .Y(n183) );
  NAND2X1 U576 ( .A(counter_st[4]), .B(n222), .Y(n204) );
  NOR3XL U577 ( .A(n187), .B(md5[4]), .C(md5[3]), .Y(n186) );
  NAND3X1 U578 ( .A(n138), .B(n136), .C(n405), .Y(n187) );
  INVX1 U579 ( .A(counter_st[2]), .Y(n62) );
  INVX1 U580 ( .A(counter_st[4]), .Y(n73) );
  INVX1 U581 ( .A(counter_st[3]), .Y(n74) );
  INVX1 U582 ( .A(md1[7]), .Y(n439) );
  INVX1 U583 ( .A(arcon[1]), .Y(n142) );
  INVX1 U584 ( .A(md1[5]), .Y(n126) );
  INVX1 U585 ( .A(md1[4]), .Y(n133) );
  NOR2X1 U586 ( .A(n47), .B(n171), .Y(n408) );
  AOI211X1 U587 ( .C(n172), .D(oper_reg[3]), .A(n173), .B(n174), .Y(n171) );
  AO44X1 U588 ( .A(arcon[6]), .B(n181), .C(n182), .D(n178), .E(n183), .F(n184), 
        .G(n185), .H(n186), .Y(n173) );
  AOI31X1 U589 ( .A(n175), .B(n176), .C(n177), .D(n178), .Y(n174) );
  NOR4XL U590 ( .A(md5[2]), .B(md5[1]), .C(md5[0]), .D(md4[7]), .Y(n185) );
  NOR4XL U591 ( .A(md4[6]), .B(md4[5]), .C(md4[4]), .D(md4[3]), .Y(n184) );
  INVX1 U592 ( .A(set_div32), .Y(n57) );
  INVX1 U593 ( .A(md0[4]), .Y(n150) );
  INVX1 U594 ( .A(md1[0]), .Y(n128) );
  INVX1 U595 ( .A(md1[2]), .Y(n127) );
  INVX1 U596 ( .A(md1[1]), .Y(n148) );
  INVX1 U597 ( .A(md1[3]), .Y(n149) );
  INVX1 U598 ( .A(md0[5]), .Y(n151) );
  INVX1 U599 ( .A(md0[6]), .Y(n131) );
  INVX1 U600 ( .A(md0[7]), .Y(n132) );
  INVX1 U601 ( .A(arcon[5]), .Y(n125) );
  NAND41XL U602 ( .D(sfraddr[4]), .A(sfraddr[5]), .B(sfraddr[3]), .C(
        sfraddr[6]), .Y(n243) );
endmodule


module mdu_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
endmodule


module mdu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module wakeupctrl_a0 ( irq, int0ff, int1ff, it0, it1, isreg, intprior0, 
        intprior1, eal, eint0, eint1, pmuintreq );
  input [3:0] isreg;
  input [1:0] intprior0;
  input [1:0] intprior1;
  input irq, int0ff, int1ff, it0, it1, eal, eint0, eint1;
  output pmuintreq;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n1;

  NAND42X1 U1 ( .C(it0), .D(int0ff), .A(eint0), .B(n9), .Y(n3) );
  OAI2B11X1 U2 ( .D(intprior0[0]), .C(n6), .A(n10), .B(n8), .Y(n9) );
  OAI21X1 U3 ( .B(intprior0[0]), .C(n1), .A(intprior1[0]), .Y(n10) );
  AO21X1 U4 ( .B(n2), .C(eal), .A(irq), .Y(pmuintreq) );
  AOI21X1 U5 ( .B(n3), .C(n4), .A(isreg[3]), .Y(n2) );
  NAND42X1 U6 ( .C(it1), .D(int1ff), .A(eint1), .B(n5), .Y(n4) );
  OAI2B11X1 U7 ( .D(intprior0[1]), .C(n6), .A(n7), .B(n8), .Y(n5) );
  OAI21X1 U8 ( .B(intprior0[1]), .C(n1), .A(intprior1[1]), .Y(n7) );
  OR2X1 U9 ( .A(isreg[1]), .B(isreg[2]), .Y(n6) );
  OR2X1 U10 ( .A(isreg[0]), .B(n6), .Y(n8) );
  INVX1 U11 ( .A(isreg[2]), .Y(n1) );
endmodule


module pmurstctrl_a0 ( resetff, wdts, srst, pmuintreq, stop, idle, clkcpu_en, 
        clkper_en, cpu_resume, rsttowdt, rsttosrst, rst );
  input resetff, wdts, srst, pmuintreq, stop, idle;
  output clkcpu_en, clkper_en, cpu_resume, rsttowdt, rsttosrst, rst;
  wire   n2;

  OAI21X1 U1 ( .B(stop), .C(idle), .A(n2), .Y(clkcpu_en) );
  NAND2X1 U2 ( .A(stop), .B(n2), .Y(clkper_en) );
  BUFX3 U3 ( .A(pmuintreq), .Y(cpu_resume) );
  INVX1 U4 ( .A(pmuintreq), .Y(n2) );
  OR2X1 U5 ( .A(srst), .B(resetff), .Y(rsttowdt) );
  OR2X1 U6 ( .A(wdts), .B(rsttowdt), .Y(rst) );
  OR2X1 U7 ( .A(resetff), .B(wdts), .Y(rsttosrst) );
endmodule


module sfrmux_a0 ( isfrwait, sfraddr, c, ac, f0, rs, ov, f1, p, acc, b, dpl, 
        dph, dps, dpc, p2, sp, smod, pmw, p2sel, gf0, stop, idle, ckcon, port0, 
        port0ff, rmwinstr, arcon, md0, md1, md2, md3, md4, md5, t0_tmod, 
        t0_tf0, t0_tf1, t0_tr0, t0_tr1, tl0, th0, t1_tmod, t1_tf1, t1_tr1, tl1, 
        th1, wdtrel, ip0wdts, wdt_tm, t2con, s0con, s0buf, s0rell, s0relh, bd, 
        ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9, 
        iex10, iex11, iex12, ien0, ien1, ien2, ip0, ip1, isr_tm, i2c_int, 
        i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o, sfrdatai, tf1_gate, riti0_gate, 
        iex7_gate, iex2_gate, srstflag, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, ext_sfr_sel, sfrdatao );
  input [6:0] sfraddr;
  input [1:0] rs;
  input [7:0] acc;
  input [7:0] b;
  input [7:0] dpl;
  input [7:0] dph;
  input [3:0] dps;
  input [5:0] dpc;
  input [7:0] p2;
  input [7:0] sp;
  input [7:0] ckcon;
  input [7:0] port0;
  input [7:0] port0ff;
  input [7:0] arcon;
  input [7:0] md0;
  input [7:0] md1;
  input [7:0] md2;
  input [7:0] md3;
  input [7:0] md4;
  input [7:0] md5;
  input [3:0] t0_tmod;
  input [7:0] tl0;
  input [7:0] th0;
  input [3:0] t1_tmod;
  input [7:0] tl1;
  input [7:0] th1;
  input [7:0] wdtrel;
  input [7:0] t2con;
  input [7:0] s0con;
  input [7:0] s0buf;
  input [7:0] s0rell;
  input [7:0] s0relh;
  input [7:0] ien0;
  input [5:0] ien1;
  input [5:0] ien2;
  input [5:0] ip0;
  input [5:0] ip1;
  input [7:0] i2cdat_o;
  input [7:0] i2cadr_o;
  input [7:0] i2ccon_o;
  input [7:0] i2csta_o;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  input isfrwait, c, ac, f0, ov, f1, p, smod, pmw, p2sel, gf0, stop, idle,
         rmwinstr, t0_tf0, t0_tf1, t0_tr0, t0_tr1, t1_tf1, t1_tr1, ip0wdts,
         wdt_tm, bd, ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12, isr_tm, i2c_int, srstflag;
  output tf1_gate, riti0_gate, iex7_gate, iex2_gate, int_vect_8b, int_vect_93,
         int_vect_9b, int_vect_a3, ext_sfr_sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305;

  NAND2XL U2 ( .A(sfrdatai[3]), .B(n21), .Y(n4) );
  NAND2XL U3 ( .A(sfrdatai[4]), .B(n21), .Y(n13) );
  NAND2X1 U4 ( .A(sfrdatai[2]), .B(n21), .Y(n10) );
  NOR5X1 U5 ( .A(n26), .B(n43), .C(n48), .D(n259), .E(n260), .Y(n83) );
  INVX2 U6 ( .A(n42), .Y(n48) );
  NAND6X1 U7 ( .A(n163), .B(n162), .C(n161), .D(n160), .E(n159), .F(n158), .Y(
        sfrdatao[1]) );
  NOR4X2 U8 ( .A(n50), .B(n51), .C(n49), .D(n52), .Y(n158) );
  NAND6X1 U9 ( .A(n148), .B(n147), .C(n146), .D(n145), .E(n144), .F(n143), .Y(
        sfrdatao[0]) );
  NAND21X1 U10 ( .B(n55), .A(sfraddr[2]), .Y(n72) );
  INVX4 U11 ( .A(sfraddr[1]), .Y(n55) );
  NAND6X2 U12 ( .A(n216), .B(n217), .C(n218), .D(n215), .E(n214), .F(n213), 
        .Y(sfrdatao[4]) );
  NOR2X4 U13 ( .A(n6), .B(n1), .Y(n24) );
  NAND2X1 U14 ( .A(n58), .B(n59), .Y(n6) );
  INVX2 U15 ( .A(n73), .Y(n272) );
  INVX1 U16 ( .A(n74), .Y(n261) );
  NAND21XL U17 ( .B(n53), .A(n36), .Y(n74) );
  NOR2XL U18 ( .A(n85), .B(n62), .Y(n20) );
  NAND32X1 U19 ( .B(n38), .C(n54), .A(n56), .Y(n80) );
  AND4X1 U20 ( .A(n292), .B(n291), .C(n290), .D(n289), .Y(n300) );
  NOR5X1 U21 ( .A(n272), .B(n25), .C(n261), .D(n127), .E(n20), .Y(n78) );
  NAND21XL U22 ( .B(sfraddr[0]), .A(n36), .Y(n115) );
  INVX1 U23 ( .A(n91), .Y(n294) );
  NAND32X2 U24 ( .B(sfraddr[0]), .C(sfraddr[1]), .A(n56), .Y(n122) );
  AND3X1 U25 ( .A(n15), .B(n16), .C(n17), .Y(n226) );
  AND3X1 U26 ( .A(n3), .B(n4), .C(n5), .Y(n194) );
  NAND2X1 U27 ( .A(i2cdat_o[3]), .B(n282), .Y(n5) );
  INVX1 U28 ( .A(n85), .Y(n40) );
  NAND42X1 U29 ( .C(n302), .D(n301), .A(n300), .B(n299), .Y(sfrdatao[7]) );
  NAND42X1 U30 ( .C(n258), .D(n257), .A(n256), .B(n255), .Y(sfrdatao[6]) );
  NOR6XL U31 ( .A(n100), .B(n294), .C(n295), .D(n288), .E(n287), .F(n18), .Y(
        n101) );
  NAND6XL U32 ( .A(n134), .B(n135), .C(n137), .D(n136), .E(n138), .F(n69), .Y(
        n104) );
  NAND6XL U33 ( .A(n78), .B(n115), .C(n125), .D(n124), .E(n126), .F(n120), .Y(
        n103) );
  INVX1 U34 ( .A(n123), .Y(n305) );
  AND3X1 U35 ( .A(n37), .B(n24), .C(n55), .Y(n36) );
  OR2X1 U36 ( .A(n57), .B(sfraddr[6]), .Y(n1) );
  AOI222XL U37 ( .A(th0[7]), .B(n269), .C(md2[7]), .D(n35), .E(port0ff[7]), 
        .F(n268), .Y(n2) );
  NAND32X1 U38 ( .B(n96), .C(n86), .A(n54), .Y(n42) );
  INVX1 U39 ( .A(sfraddr[3]), .Y(n57) );
  NAND32X1 U40 ( .B(sfraddr[3]), .C(n93), .A(n61), .Y(n121) );
  OR2X1 U41 ( .A(n61), .B(n86), .Y(n99) );
  NAND2X1 U42 ( .A(i2ccon_o[3]), .B(n284), .Y(n3) );
  INVX1 U43 ( .A(sfraddr[2]), .Y(n56) );
  AND3XL U44 ( .A(sfraddr[6]), .B(sfraddr[2]), .C(n55), .Y(n41) );
  NAND2XL U45 ( .A(port0[7]), .B(n305), .Y(n7) );
  NAND2X1 U46 ( .A(arcon[7]), .B(n270), .Y(n8) );
  AND3X1 U47 ( .A(n7), .B(n8), .C(n2), .Y(n277) );
  NAND2X1 U48 ( .A(i2cdat_o[2]), .B(n282), .Y(n11) );
  NAND6X2 U49 ( .A(n181), .B(n180), .C(n179), .D(n178), .E(n177), .F(n176), 
        .Y(sfrdatao[2]) );
  NAND2XL U50 ( .A(n58), .B(n59), .Y(n93) );
  AOI221XL U51 ( .A(p2[4]), .B(n274), .C(sp[4]), .D(n266), .E(n207), .Y(n215)
         );
  NAND2X1 U52 ( .A(i2ccon_o[2]), .B(n284), .Y(n9) );
  AND3X2 U53 ( .A(n9), .B(n10), .C(n11), .Y(n175) );
  INVXL U54 ( .A(n134), .Y(n275) );
  AND2X2 U55 ( .A(n19), .B(n98), .Y(n18) );
  AOI221XL U56 ( .A(sp[2]), .B(n266), .C(ip0[2]), .D(n242), .E(n165), .Y(n178)
         );
  AOI221XL U57 ( .A(tl1[4]), .B(n298), .C(tl0[4]), .D(n297), .E(n201), .Y(n218) );
  AOI221XL U58 ( .A(i2cadr_o[2]), .B(n294), .C(it1), .D(n295), .E(n167), .Y(
        n173) );
  NAND2X1 U59 ( .A(i2ccon_o[4]), .B(n284), .Y(n12) );
  NAND2X1 U60 ( .A(i2cdat_o[4]), .B(n282), .Y(n14) );
  AND3X2 U61 ( .A(n12), .B(n13), .C(n14), .Y(n206) );
  NOR21X2 U62 ( .B(n22), .A(n304), .Y(n21) );
  INVXL U63 ( .A(n105), .Y(n282) );
  INVX1 U64 ( .A(n137), .Y(n274) );
  NAND21XL U65 ( .B(n88), .A(n87), .Y(n106) );
  NAND32XL U66 ( .B(n121), .C(n72), .A(n53), .Y(n73) );
  AOI221X1 U67 ( .A(i2cdat_o[6]), .B(n282), .C(sfrdatai[6]), .D(n21), .E(n249), 
        .Y(n253) );
  NAND2X1 U68 ( .A(i2ccon_o[5]), .B(n284), .Y(n15) );
  NAND2X1 U69 ( .A(sfrdatai[5]), .B(n21), .Y(n16) );
  NAND2X1 U70 ( .A(i2cdat_o[5]), .B(n282), .Y(n17) );
  INVXL U71 ( .A(n110), .Y(n293) );
  INVX1 U72 ( .A(n99), .Y(n19) );
  INVXL U73 ( .A(n23), .Y(n22) );
  INVX2 U74 ( .A(n82), .Y(n260) );
  INVX1 U75 ( .A(sfraddr[6]), .Y(n61) );
  AOI221XL U76 ( .A(tl1[7]), .B(n298), .C(tl0[7]), .D(n297), .E(n296), .Y(n299) );
  AND4X1 U77 ( .A(n171), .B(n170), .C(n169), .D(n168), .Y(n172) );
  INVXL U78 ( .A(n113), .Y(n298) );
  NAND21X2 U79 ( .B(n80), .A(n24), .Y(n81) );
  NAND31XL U80 ( .C(n59), .A(n40), .B(n58), .Y(n108) );
  INVXL U81 ( .A(n56), .Y(n37) );
  NAND21XL U82 ( .B(n121), .A(n98), .Y(n138) );
  NAND21XL U83 ( .B(n79), .A(n98), .Y(n111) );
  NAND32XL U84 ( .B(n71), .C(n90), .A(n70), .Y(n120) );
  OR2XL U85 ( .A(n6), .B(n85), .Y(n112) );
  NAND32XL U86 ( .B(n61), .C(n90), .A(n95), .Y(n91) );
  INVXL U87 ( .A(n89), .Y(n284) );
  INVXL U88 ( .A(n126), .Y(n262) );
  INVX3 U89 ( .A(n303), .Y(n268) );
  INVXL U90 ( .A(sfraddr[5]), .Y(n59) );
  NAND32X1 U91 ( .B(n84), .C(n80), .A(n61), .Y(n67) );
  INVX3 U92 ( .A(n67), .Y(n267) );
  INVX2 U93 ( .A(n68), .Y(n264) );
  NAND32XL U94 ( .B(n86), .C(n53), .A(n41), .Y(n82) );
  NOR2XL U95 ( .A(n121), .B(n122), .Y(n23) );
  NOR2XL U96 ( .A(n53), .B(n72), .Y(n39) );
  NAND21XL U97 ( .B(sfraddr[5]), .A(sfraddr[4]), .Y(n71) );
  NAND21XL U98 ( .B(n88), .A(n24), .Y(n114) );
  INVXL U99 ( .A(n63), .Y(n70) );
  NAND32XL U100 ( .B(n99), .C(n72), .A(n53), .Y(n124) );
  NAND32XL U101 ( .B(n88), .C(n61), .A(n95), .Y(n105) );
  NAND21XL U102 ( .B(n122), .A(n95), .Y(n128) );
  NAND32XL U103 ( .B(n88), .C(n86), .A(n60), .Y(n107) );
  NAND32XL U104 ( .B(sfraddr[6]), .C(n57), .A(n77), .Y(n79) );
  NAND32XL U105 ( .B(n54), .C(n99), .A(n75), .Y(n125) );
  NAND21XL U106 ( .B(n122), .A(n87), .Y(n135) );
  INVXL U107 ( .A(n64), .Y(n185) );
  INVXL U108 ( .A(n62), .Y(n77) );
  INVXL U109 ( .A(n76), .Y(n127) );
  OA21XL U110 ( .B(t1_tr1), .C(t0_tr1), .A(n295), .Y(n249) );
  INVXL U111 ( .A(n157), .Y(n49) );
  NAND42XL U112 ( .C(n279), .D(n278), .A(n277), .B(n276), .Y(n301) );
  NAND42XL U113 ( .C(n248), .D(n247), .A(n246), .B(n245), .Y(n257) );
  AND2XL U114 ( .A(i2ccon_o[1]), .B(n284), .Y(n27) );
  AOI22XL U115 ( .A(i2ccon_o[6]), .B(n284), .C(s0rell[6]), .D(n283), .Y(n252)
         );
  AOI22XL U116 ( .A(md0[6]), .B(n18), .C(t2con[6]), .D(n288), .Y(n250) );
  AOI22XL U117 ( .A(i2ccon_o[7]), .B(n284), .C(s0rell[7]), .D(n283), .Y(n291)
         );
  AOI22XL U118 ( .A(md0[7]), .B(n18), .C(t2con[7]), .D(n288), .Y(n289) );
  AOI22XL U119 ( .A(i2cadr_o[4]), .B(n294), .C(t0_tr0), .D(n295), .Y(n203) );
  AOI22XL U120 ( .A(i2cadr_o[5]), .B(n294), .C(t0_tf0), .D(n295), .Y(n223) );
  AND4X1 U121 ( .A(n119), .B(n118), .C(n117), .D(n116), .Y(n145) );
  AO222XL U122 ( .A(md0[0]), .B(n18), .C(i2csta_o[0]), .D(n287), .E(t2con[0]), 
        .F(n288), .Y(n109) );
  AOI22XL U123 ( .A(md2[1]), .B(n35), .C(th0[1]), .D(n269), .Y(n153) );
  AO222XL U124 ( .A(md0[3]), .B(n18), .C(i2csta_o[3]), .D(n287), .E(t2con[3]), 
        .F(n288), .Y(n186) );
  AO222XL U125 ( .A(dph[2]), .B(n275), .C(ien1[2]), .D(n227), .E(p2[2]), .F(
        n274), .Y(n165) );
  AOI22XL U126 ( .A(md2[0]), .B(n35), .C(th0[0]), .D(n269), .Y(n116) );
  AO222XL U127 ( .A(dph[1]), .B(n275), .C(ien1[1]), .D(n227), .E(p2[1]), .F(
        n274), .Y(n150) );
  AO222XL U128 ( .A(dph[3]), .B(n275), .C(ien1[3]), .D(n227), .E(p2[3]), .F(
        n274), .Y(n183) );
  INVX1 U129 ( .A(n136), .Y(n242) );
  INVX1 U130 ( .A(n112), .Y(n220) );
  INVX1 U131 ( .A(n111), .Y(n219) );
  INVX1 U132 ( .A(n108), .Y(n286) );
  INVX1 U133 ( .A(n120), .Y(n231) );
  INVX1 U134 ( .A(n138), .Y(n266) );
  OR2X1 U135 ( .A(n121), .B(n90), .Y(n134) );
  NAND21X1 U136 ( .B(n121), .A(n39), .Y(n110) );
  NAND32X1 U137 ( .B(n57), .C(n59), .A(n58), .Y(n86) );
  INVXL U138 ( .A(n80), .Y(n98) );
  INVX1 U139 ( .A(n65), .Y(n265) );
  NAND21XL U140 ( .B(n71), .A(n40), .Y(n65) );
  INVXL U141 ( .A(n115), .Y(n269) );
  NAND6X1 U142 ( .A(n105), .B(n128), .C(n89), .D(n108), .E(n107), .F(n106), 
        .Y(n100) );
  INVX1 U143 ( .A(n79), .Y(n87) );
  INVX1 U144 ( .A(n114), .Y(n297) );
  INVX1 U145 ( .A(n135), .Y(n227) );
  NOR5X1 U146 ( .A(n185), .B(n265), .C(n230), .D(n267), .E(n264), .Y(n69) );
  INVX1 U147 ( .A(n128), .Y(n281) );
  INVX1 U148 ( .A(n41), .Y(n96) );
  INVX1 U149 ( .A(n107), .Y(n283) );
  INVX1 U150 ( .A(n125), .Y(n270) );
  INVX1 U151 ( .A(n124), .Y(n263) );
  INVX1 U152 ( .A(n106), .Y(n285) );
  NAND43X1 U153 ( .B(n122), .C(n59), .D(sfraddr[4]), .A(n70), .Y(n137) );
  NAND32XL U154 ( .B(n34), .C(n72), .A(n53), .Y(n126) );
  INVXL U155 ( .A(n72), .Y(n75) );
  NAND32X1 U156 ( .B(n122), .C(n61), .A(n57), .Y(n85) );
  NAND32XL U157 ( .B(n55), .C(n53), .A(n56), .Y(n90) );
  NAND32XL U158 ( .B(n47), .C(n96), .A(n53), .Y(n89) );
  INVX1 U159 ( .A(n46), .Y(n95) );
  NAND21XL U160 ( .B(n71), .A(sfraddr[3]), .Y(n46) );
  INVX1 U161 ( .A(n94), .Y(n288) );
  NAND43X1 U162 ( .B(n6), .C(n122), .D(n57), .A(sfraddr[6]), .Y(n94) );
  INVX1 U163 ( .A(n97), .Y(n287) );
  NAND32XL U164 ( .B(n96), .C(n53), .A(n95), .Y(n97) );
  INVX1 U165 ( .A(sfraddr[4]), .Y(n58) );
  NAND32XL U166 ( .B(n122), .C(n86), .A(n61), .Y(n68) );
  NAND21XL U167 ( .B(sfraddr[6]), .A(n57), .Y(n63) );
  NOR2XL U168 ( .A(n121), .B(n88), .Y(n25) );
  NAND21XL U169 ( .B(n58), .A(sfraddr[5]), .Y(n62) );
  INVX1 U170 ( .A(n92), .Y(n295) );
  NAND21XL U171 ( .B(n122), .A(n24), .Y(n92) );
  INVX2 U172 ( .A(n66), .Y(n230) );
  NAND32X1 U173 ( .B(n47), .C(n88), .A(n61), .Y(n66) );
  NOR2X2 U174 ( .A(n88), .B(n99), .Y(n26) );
  NAND5XL U175 ( .A(n39), .B(sfraddr[6]), .C(sfraddr[4]), .D(sfraddr[5]), .E(
        n57), .Y(n76) );
  INVX1 U176 ( .A(n129), .Y(n271) );
  NAND21X1 U177 ( .B(sfraddr[6]), .A(n281), .Y(n129) );
  NAND32XL U178 ( .B(n71), .C(n88), .A(n70), .Y(n64) );
  INVX1 U179 ( .A(sfraddr[0]), .Y(n53) );
  NAND21X1 U180 ( .B(n305), .A(n23), .Y(n303) );
  NAND32XL U181 ( .B(n305), .C(n304), .A(n303), .Y(ext_sfr_sel) );
  AO222XL U182 ( .A(ien0[2]), .B(n264), .C(s0buf[2]), .D(n267), .E(ien2[2]), 
        .F(n230), .Y(n166) );
  AO222XL U183 ( .A(ien0[1]), .B(n264), .C(s0buf[1]), .D(n267), .E(ien2[1]), 
        .F(n230), .Y(n151) );
  AO222XL U184 ( .A(ien0[3]), .B(n264), .C(s0buf[3]), .D(n267), .E(ien2[3]), 
        .F(n230), .Y(n184) );
  AO222XL U185 ( .A(s0buf[4]), .B(n267), .C(ip0[4]), .D(n242), .E(ien0[4]), 
        .F(n264), .Y(n208) );
  AO222XL U186 ( .A(s0buf[5]), .B(n267), .C(ip0[5]), .D(n242), .E(ien0[5]), 
        .F(n264), .Y(n229) );
  AO222XL U187 ( .A(md4[4]), .B(n260), .C(t1_tmod[0]), .D(n259), .E(md3[4]), 
        .F(n48), .Y(n202) );
  AND2XL U188 ( .A(bd), .B(sfraddr[6]), .Y(n280) );
  NAND4X1 U189 ( .A(n156), .B(n155), .C(n154), .D(n153), .Y(n52) );
  AOI221XL U190 ( .A(tl0[6]), .B(n297), .C(t1_tmod[2]), .D(n259), .E(n254), 
        .Y(n255) );
  AOI221XL U191 ( .A(wdtrel[2]), .B(n272), .C(dpl[2]), .D(n25), .E(n164), .Y(
        n179) );
  AO2222XL U192 ( .A(md4[7]), .B(n260), .C(t1_tmod[3]), .D(n259), .E(md1[7]), 
        .F(n26), .G(md3[7]), .H(n48), .Y(n302) );
  NAND31X1 U193 ( .C(n27), .A(n44), .B(n45), .Y(n50) );
  AO222XL U194 ( .A(md4[5]), .B(n260), .C(t1_tmod[1]), .D(n259), .E(md3[5]), 
        .F(n48), .Y(n222) );
  AO222X1 U195 ( .A(iex5), .B(n220), .C(ip1[4]), .D(n219), .E(pmw), .F(n293), 
        .Y(n201) );
  AO222XL U196 ( .A(ien1[4]), .B(n227), .C(dpl[4]), .D(n25), .E(dph[4]), .F(
        n275), .Y(n207) );
  AO222XL U197 ( .A(ien1[5]), .B(n227), .C(dpl[5]), .D(n25), .E(dph[5]), .F(
        n275), .Y(n228) );
  AO222X1 U198 ( .A(iex6), .B(n220), .C(ip1[5]), .D(n219), .E(isr_tm), .F(n293), .Y(n221) );
  AO222X1 U199 ( .A(md0[2]), .B(n18), .C(i2csta_o[2]), .D(n287), .E(t2con[2]), 
        .F(n288), .Y(n167) );
  AOI222XL U200 ( .A(s0relh[0]), .B(n285), .C(s0rell[0]), .D(n283), .E(acc[0]), 
        .F(n286), .Y(n147) );
  AOI221XL U201 ( .A(tl1[5]), .B(n298), .C(tl0[5]), .D(n297), .E(n221), .Y(
        n241) );
  AOI221XL U202 ( .A(p2[5]), .B(n274), .C(sp[5]), .D(n266), .E(n228), .Y(n238)
         );
  AOI221XL U203 ( .A(md1[5]), .B(n26), .C(md2[5]), .D(n35), .E(n222), .Y(n240)
         );
  AOI222XL U204 ( .A(md5[1]), .B(n263), .C(arcon[1]), .D(n270), .E(ckcon[1]), 
        .F(n262), .Y(n162) );
  AOI222XL U205 ( .A(dpc[1]), .B(n231), .C(port0ff[1]), .D(n268), .E(port0[1]), 
        .F(n305), .Y(n163) );
  AOI221XL U206 ( .A(sp[1]), .B(n266), .C(ip0[1]), .D(n242), .E(n150), .Y(n160) );
  AOI222XL U207 ( .A(i2csta_o[7]), .B(n287), .C(acc[7]), .D(n286), .E(
        s0relh[7]), .F(n285), .Y(n290) );
  AOI222XL U208 ( .A(md5[3]), .B(n263), .C(arcon[3]), .D(n270), .E(ckcon[3]), 
        .F(n262), .Y(n199) );
  AOI222XL U209 ( .A(dpc[3]), .B(n231), .C(port0ff[3]), .D(n268), .E(port0[3]), 
        .F(n305), .Y(n200) );
  AOI221XL U210 ( .A(sp[3]), .B(n266), .C(ip0[3]), .D(n242), .E(n183), .Y(n197) );
  AND4X1 U211 ( .A(n212), .B(n211), .C(n210), .D(n209), .Y(n213) );
  AND4X1 U212 ( .A(n253), .B(n252), .C(n251), .D(n250), .Y(n256) );
  AOI222XL U213 ( .A(i2csta_o[6]), .B(n287), .C(acc[6]), .D(n286), .E(
        s0relh[6]), .F(n285), .Y(n251) );
  AOI222XL U214 ( .A(s0relh[4]), .B(n285), .C(s0rell[4]), .D(n283), .E(acc[4]), 
        .F(n286), .Y(n205) );
  AOI222XL U215 ( .A(t2con[4]), .B(n288), .C(i2csta_o[4]), .D(n287), .E(md0[4]), .F(n18), .Y(n204) );
  AOI222XL U216 ( .A(s0relh[3]), .B(n285), .C(s0rell[3]), .D(n283), .E(acc[3]), 
        .F(n286), .Y(n193) );
  AND4X1 U217 ( .A(n190), .B(n189), .C(n188), .D(n187), .Y(n191) );
  AOI221XL U218 ( .A(i2cadr_o[3]), .B(n294), .C(ie1), .D(n295), .E(n186), .Y(
        n192) );
  AOI222XL U219 ( .A(s0relh[2]), .B(n285), .C(s0rell[2]), .D(n283), .E(acc[2]), 
        .F(n286), .Y(n174) );
  AOI222XL U220 ( .A(s0relh[5]), .B(n285), .C(s0rell[5]), .D(n283), .E(acc[5]), 
        .F(n286), .Y(n225) );
  AOI222XL U221 ( .A(t2con[5]), .B(n288), .C(i2csta_o[5]), .D(n287), .E(md0[5]), .F(n18), .Y(n224) );
  AOI222XL U222 ( .A(md5[2]), .B(n263), .C(arcon[2]), .D(n270), .E(ckcon[2]), 
        .F(n262), .Y(n180) );
  AOI222XL U223 ( .A(dpc[2]), .B(n231), .C(port0ff[2]), .D(n268), .E(port0[2]), 
        .F(n305), .Y(n181) );
  AND4X1 U224 ( .A(n133), .B(n132), .C(n131), .D(n130), .Y(n144) );
  AOI22XL U225 ( .A(s0con[0]), .B(n271), .C(wdtrel[0]), .D(n272), .Y(n130) );
  AOI222XL U226 ( .A(md5[0]), .B(n263), .C(arcon[0]), .D(n270), .E(ckcon[0]), 
        .F(n262), .Y(n132) );
  AND4X1 U227 ( .A(n235), .B(n234), .C(n233), .D(n232), .Y(n236) );
  AOI22XL U228 ( .A(s0con[5]), .B(n271), .C(wdtrel[5]), .D(n272), .Y(n232) );
  AOI222XL U229 ( .A(ckcon[5]), .B(n262), .C(dpc[5]), .D(n231), .E(arcon[5]), 
        .F(n270), .Y(n234) );
  NAND32XL U230 ( .B(n122), .C(n121), .A(rmwinstr), .Y(n123) );
  AOI221XL U231 ( .A(arcon[6]), .B(n270), .C(ckcon[6]), .D(n262), .E(n243), 
        .Y(n246) );
  AO222X1 U232 ( .A(port0ff[6]), .B(n268), .C(th0[6]), .D(n269), .E(port0[6]), 
        .F(n305), .Y(n243) );
  AOI221XL U233 ( .A(p2[6]), .B(n274), .C(sp[6]), .D(n266), .E(n244), .Y(n245)
         );
  AO222XL U234 ( .A(dpl[6]), .B(n25), .C(wdtrel[6]), .D(n272), .E(dph[6]), .F(
        n275), .Y(n244) );
  AOI221XL U235 ( .A(dph[7]), .B(n275), .C(p2[7]), .D(n274), .E(n273), .Y(n276) );
  AO222XL U236 ( .A(wdtrel[7]), .B(n272), .C(s0con[7]), .D(n271), .E(dpl[7]), 
        .F(n25), .Y(n273) );
  AOI222XL U237 ( .A(md1[1]), .B(n26), .C(md4[1]), .D(n260), .E(md3[1]), .F(
        n48), .Y(n154) );
  AOI222XL U238 ( .A(stop), .B(n293), .C(ip1[1]), .D(n219), .E(iex2), .F(n220), 
        .Y(n156) );
  AOI222XL U239 ( .A(i2ccon_o[0]), .B(n284), .C(sfrdatai[0]), .D(n21), .E(
        i2cdat_o[0]), .F(n282), .Y(n148) );
  AOI222XL U240 ( .A(md1[3]), .B(n26), .C(md4[3]), .D(n260), .E(md3[3]), .F(
        n48), .Y(n188) );
  AOI222XL U241 ( .A(md1[2]), .B(n26), .C(md4[2]), .D(n260), .E(md3[2]), .F(
        n48), .Y(n169) );
  AOI222XL U242 ( .A(gf0), .B(n293), .C(ip1[2]), .D(n219), .E(iex3), .F(n220), 
        .Y(n171) );
  AOI222XL U243 ( .A(dpc[0]), .B(n231), .C(port0ff[0]), .D(n268), .E(port0[0]), 
        .F(n305), .Y(n133) );
  AOI222XL U244 ( .A(port0[4]), .B(n305), .C(th0[4]), .D(n269), .E(port0ff[4]), 
        .F(n268), .Y(n212) );
  AOI222XL U245 ( .A(port0[5]), .B(n305), .C(th0[5]), .D(n269), .E(port0ff[5]), 
        .F(n268), .Y(n235) );
  AOI222XL U246 ( .A(t0_tmod[2]), .B(n259), .C(tl1[2]), .D(n298), .E(tl0[2]), 
        .F(n297), .Y(n170) );
  AOI221X1 U247 ( .A(i2cadr_o[1]), .B(n294), .C(ie0), .D(n295), .E(n152), .Y(
        n157) );
  AO222X1 U248 ( .A(md0[1]), .B(n18), .C(i2csta_o[1]), .D(n287), .E(t2con[1]), 
        .F(n288), .Y(n152) );
  AOI221XL U249 ( .A(i2cadr_o[0]), .B(n294), .C(it0), .D(n295), .E(n109), .Y(
        n146) );
  AOI221XL U250 ( .A(wdtrel[1]), .B(n272), .C(dpl[1]), .D(n25), .E(n149), .Y(
        n161) );
  AOI221XL U251 ( .A(wdtrel[3]), .B(n272), .C(dpl[3]), .D(n25), .E(n182), .Y(
        n198) );
  AO222X1 U252 ( .A(wdt_tm), .B(n293), .C(i2cadr_o[6]), .D(n294), .E(tl1[6]), 
        .F(n298), .Y(n254) );
  AO222X1 U253 ( .A(n295), .B(tf1_gate), .C(i2cadr_o[7]), .D(n294), .E(smod), 
        .F(n293), .Y(n296) );
  AOI222XL U254 ( .A(t0_tmod[1]), .B(n259), .C(tl1[1]), .D(n298), .E(tl0[1]), 
        .F(n297), .Y(n155) );
  AOI222XL U255 ( .A(ien2[0]), .B(n230), .C(s0buf[0]), .D(n267), .E(ien0[0]), 
        .F(n264), .Y(n140) );
  AOI222XL U256 ( .A(ip0[0]), .B(n242), .C(p2[0]), .D(n274), .E(sp[0]), .F(
        n266), .Y(n141) );
  AOI222XL U257 ( .A(md1[0]), .B(n26), .C(md4[0]), .D(n260), .E(md3[0]), .F(
        n48), .Y(n117) );
  AOI222XL U258 ( .A(p2sel), .B(n293), .C(ip1[3]), .D(n219), .E(iex4), .F(n220), .Y(n190) );
  AOI222XL U259 ( .A(idle), .B(n293), .C(ip1[0]), .D(n219), .E(iex7), .F(n220), 
        .Y(n119) );
  AOI222XL U260 ( .A(t0_tmod[3]), .B(n259), .C(tl1[3]), .D(n298), .E(tl0[3]), 
        .F(n297), .Y(n189) );
  AOI222XL U261 ( .A(t0_tmod[0]), .B(n259), .C(tl1[0]), .D(n298), .E(tl0[0]), 
        .F(n297), .Y(n118) );
  AOI222XL U262 ( .A(ckcon[4]), .B(n262), .C(dpc[4]), .D(n231), .E(arcon[4]), 
        .F(n270), .Y(n211) );
  AOI222XL U263 ( .A(dph[0]), .B(n275), .C(dpl[0]), .D(n25), .E(ien1[0]), .F(
        n227), .Y(n142) );
  AOI22XL U264 ( .A(s0con[4]), .B(n271), .C(wdtrel[4]), .D(n272), .Y(n209) );
  OR2X1 U265 ( .A(t1_tf1), .B(t0_tf1), .Y(tf1_gate) );
  BUFX3 U266 ( .A(iex7), .Y(iex7_gate) );
  BUFX3 U267 ( .A(iex8), .Y(int_vect_8b) );
  BUFX3 U268 ( .A(iex2), .Y(iex2_gate) );
  BUFX3 U269 ( .A(iex9), .Y(int_vect_93) );
  OR2X1 U270 ( .A(s0con[1]), .B(s0con[0]), .Y(riti0_gate) );
  BUFX3 U271 ( .A(iex11), .Y(int_vect_a3) );
  BUFX3 U272 ( .A(iex10), .Y(int_vect_9b) );
  AO222XL U273 ( .A(th1[3]), .B(n261), .C(b[3]), .D(n20), .E(s0con[3]), .F(
        n271), .Y(n182) );
  AO222XL U274 ( .A(th1[1]), .B(n261), .C(b[1]), .D(n20), .E(s0con[1]), .F(
        n271), .Y(n149) );
  AO222XL U275 ( .A(th1[2]), .B(n261), .C(b[2]), .D(n20), .E(s0con[2]), .F(
        n271), .Y(n164) );
  NAND32XL U276 ( .B(n6), .C(n57), .A(n61), .Y(n34) );
  NOR2XL U277 ( .A(n99), .B(n90), .Y(n35) );
  NOR2XL U278 ( .A(n99), .B(n90), .Y(n43) );
  NAND6XL U279 ( .A(n112), .B(n111), .C(n110), .D(n114), .E(n113), .F(n83), 
        .Y(n102) );
  AOI221XL U280 ( .A(md1[4]), .B(n26), .C(md2[4]), .D(n35), .E(n202), .Y(n217)
         );
  AO2222XL U281 ( .A(md3[6]), .B(n48), .C(md4[6]), .D(n260), .E(md2[6]), .F(
        n35), .G(md1[6]), .H(n26), .Y(n258) );
  NAND32X2 U282 ( .B(sfraddr[0]), .C(n55), .A(n56), .Y(n88) );
  INVX1 U283 ( .A(sfraddr[0]), .Y(n54) );
  INVX1 U284 ( .A(n55), .Y(n38) );
  AOI22XL U285 ( .A(md2[2]), .B(n35), .C(th0[2]), .D(n269), .Y(n168) );
  AOI22XL U286 ( .A(md2[3]), .B(n35), .C(th0[3]), .D(n269), .Y(n187) );
  INVX4 U287 ( .A(n81), .Y(n259) );
  NAND32XL U288 ( .B(n86), .C(n80), .A(n60), .Y(n136) );
  AOI222XL U289 ( .A(i2cdat_o[7]), .B(n282), .C(n281), .D(n280), .E(
        sfrdatai[7]), .F(n21), .Y(n292) );
  INVXL U290 ( .A(sfraddr[6]), .Y(n60) );
  NAND21XL U291 ( .B(n90), .A(n24), .Y(n113) );
  AO2222XL U292 ( .A(s0buf[7]), .B(n267), .C(sp[7]), .D(n266), .E(c), .F(n265), 
        .G(ien0[7]), .H(n264), .Y(n278) );
  AO2222XL U293 ( .A(s0buf[6]), .B(n267), .C(ip0wdts), .D(n242), .E(ac), .F(
        n265), .G(ien0[6]), .H(n264), .Y(n247) );
  AOI221XL U294 ( .A(ien2[5]), .B(n230), .C(f0), .D(n265), .E(n229), .Y(n237)
         );
  AOI221XL U295 ( .A(ien2[4]), .B(n230), .C(rs[1]), .D(n265), .E(n208), .Y(
        n214) );
  AOI221XL U296 ( .A(dps[3]), .B(n185), .C(rs[0]), .D(n265), .E(n184), .Y(n196) );
  AOI221XL U297 ( .A(dps[2]), .B(n185), .C(ov), .D(n265), .E(n166), .Y(n177)
         );
  AOI221XL U298 ( .A(dps[1]), .B(n185), .C(f1), .D(n265), .E(n151), .Y(n159)
         );
  AOI22XL U299 ( .A(dps[0]), .B(n185), .C(p), .D(n265), .Y(n139) );
  NAND6X1 U300 ( .A(n241), .B(n240), .C(n239), .D(n238), .E(n237), .F(n236), 
        .Y(sfrdatao[5]) );
  NAND6X2 U301 ( .A(n195), .B(n199), .C(n198), .D(n197), .E(n196), .F(n200), 
        .Y(sfrdatao[3]) );
  AND4X1 U302 ( .A(n142), .B(n141), .C(n140), .D(n139), .Y(n143) );
  AO2222XL U303 ( .A(md5[7]), .B(n263), .C(ckcon[7]), .D(n262), .E(th1[7]), 
        .F(n261), .G(b[7]), .H(n20), .Y(n279) );
  AO2222XL U304 ( .A(b[6]), .B(n20), .C(md5[6]), .D(n263), .E(s0con[6]), .F(
        n271), .G(th1[6]), .H(n261), .Y(n248) );
  AOI222XL U305 ( .A(th1[5]), .B(n261), .C(md5[5]), .D(n263), .E(b[5]), .F(n20), .Y(n233) );
  AOI222XL U306 ( .A(th1[4]), .B(n261), .C(md5[4]), .D(n263), .E(b[4]), .F(n20), .Y(n210) );
  AOI222XL U307 ( .A(th1[0]), .B(n261), .C(srstflag), .D(n127), .E(b[0]), .F(
        n20), .Y(n131) );
  NAND2XL U308 ( .A(sfrdatai[1]), .B(n21), .Y(n44) );
  NAND2XL U309 ( .A(i2cdat_o[1]), .B(n282), .Y(n45) );
  NAND21X1 U310 ( .B(n71), .A(sfraddr[3]), .Y(n47) );
  NAND21X1 U311 ( .B(n71), .A(sfraddr[3]), .Y(n84) );
  AO222X1 U312 ( .A(s0relh[1]), .B(n285), .C(s0rell[1]), .D(n283), .E(acc[1]), 
        .F(n286), .Y(n51) );
  AND4X1 U313 ( .A(n194), .B(n193), .C(n192), .D(n191), .Y(n195) );
  AND4X1 U314 ( .A(n206), .B(n205), .C(n204), .D(n203), .Y(n216) );
  AND4X1 U315 ( .A(n226), .B(n225), .C(n224), .D(n223), .Y(n239) );
  AND4X1 U316 ( .A(n175), .B(n174), .C(n173), .D(n172), .Y(n176) );
  NAND43X1 U317 ( .B(n104), .C(n103), .D(n102), .A(n101), .Y(n304) );
endmodule


module syncneg_a0 ( clk, reset, rsttowdt, rsttosrst, rst, int0, int1, port0i, 
        rxd0i, sdai, int0ff, int1ff, port0ff, t0ff, t1ff, rxd0ff, sdaiff, 
        rsttowdtff, rsttosrstff, rstff, resetff, test_si, test_se );
  input [7:0] port0i;
  output [7:0] port0ff;
  input clk, reset, rsttowdt, rsttosrst, rst, int0, int1, rxd0i, sdai, test_si,
         test_se;
  output int0ff, int1ff, t0ff, t1ff, rxd0ff, sdaiff, rsttowdtff, rsttosrstff,
         rstff, resetff;
  wire   reset_ff1, int0_ff1, int1_ff1, rxd0_ff1, sdai_ff1;
  wire   [7:0] p0_ff1;

  SDFFQX1 reset_ff2_reg ( .D(reset_ff1), .SIN(reset_ff1), .SMC(test_se), .C(
        clk), .Q(resetff) );
  SDFFQX1 rsttosrst_ff1_reg ( .D(rsttosrst), .SIN(rstff), .SMC(test_se), .C(
        clk), .Q(rsttosrstff) );
  SDFFQX1 rsttowdt_ff1_reg ( .D(rsttowdt), .SIN(rsttosrstff), .SMC(test_se), 
        .C(clk), .Q(rsttowdtff) );
  SDFFQX1 int0_ff2_reg ( .D(int0_ff1), .SIN(int0_ff1), .SMC(test_se), .C(clk), 
        .Q(int0ff) );
  SDFFQX1 int1_ff2_reg ( .D(int1_ff1), .SIN(int1_ff1), .SMC(test_se), .C(clk), 
        .Q(int1ff) );
  SDFFQX1 rxd0_ff2_reg ( .D(rxd0_ff1), .SIN(rxd0_ff1), .SMC(test_se), .C(clk), 
        .Q(rxd0ff) );
  SDFFQX1 sdai_ff2_reg ( .D(sdai_ff1), .SIN(sdai_ff1), .SMC(test_se), .C(clk), 
        .Q(sdaiff) );
  SDFFQX1 p0_ff2_reg_1_ ( .D(p0_ff1[1]), .SIN(port0ff[0]), .SMC(test_se), .C(
        clk), .Q(port0ff[1]) );
  SDFFQX1 p0_ff2_reg_3_ ( .D(p0_ff1[3]), .SIN(port0ff[2]), .SMC(test_se), .C(
        clk), .Q(port0ff[3]) );
  SDFFQX1 p0_ff2_reg_4_ ( .D(p0_ff1[4]), .SIN(port0ff[3]), .SMC(test_se), .C(
        clk), .Q(port0ff[4]) );
  SDFFQX1 p0_ff2_reg_5_ ( .D(p0_ff1[5]), .SIN(port0ff[4]), .SMC(test_se), .C(
        clk), .Q(port0ff[5]) );
  SDFFQX1 p0_ff2_reg_0_ ( .D(p0_ff1[0]), .SIN(p0_ff1[7]), .SMC(test_se), .C(
        clk), .Q(port0ff[0]) );
  SDFFQX1 p0_ff2_reg_2_ ( .D(p0_ff1[2]), .SIN(port0ff[1]), .SMC(test_se), .C(
        clk), .Q(port0ff[2]) );
  SDFFQX1 p0_ff2_reg_7_ ( .D(p0_ff1[7]), .SIN(port0ff[6]), .SMC(test_se), .C(
        clk), .Q(port0ff[7]) );
  SDFFQX1 p0_ff2_reg_6_ ( .D(p0_ff1[6]), .SIN(port0ff[5]), .SMC(test_se), .C(
        clk), .Q(port0ff[6]) );
  SDFFQX1 rst_ff1_reg ( .D(rst), .SIN(resetff), .SMC(test_se), .C(clk), .Q(
        rstff) );
  SDFFQX1 int0_ff1_reg ( .D(int0), .SIN(test_si), .SMC(test_se), .C(clk), .Q(
        int0_ff1) );
  SDFFQX1 int1_ff1_reg ( .D(int1), .SIN(int0ff), .SMC(test_se), .C(clk), .Q(
        int1_ff1) );
  SDFFQX1 p0_ff1_reg_6_ ( .D(port0i[6]), .SIN(p0_ff1[5]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[6]) );
  SDFFQX1 p0_ff1_reg_5_ ( .D(port0i[5]), .SIN(p0_ff1[4]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[5]) );
  SDFFQX1 p0_ff1_reg_4_ ( .D(port0i[4]), .SIN(p0_ff1[3]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[4]) );
  SDFFQX1 p0_ff1_reg_2_ ( .D(port0i[2]), .SIN(p0_ff1[1]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[2]) );
  SDFFQX1 p0_ff1_reg_1_ ( .D(port0i[1]), .SIN(p0_ff1[0]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[1]) );
  SDFFQX1 p0_ff1_reg_0_ ( .D(port0i[0]), .SIN(int1ff), .SMC(test_se), .C(clk), 
        .Q(p0_ff1[0]) );
  SDFFQX1 rxd0_ff1_reg ( .D(rxd0i), .SIN(rsttowdtff), .SMC(test_se), .C(clk), 
        .Q(rxd0_ff1) );
  SDFFQX1 p0_ff1_reg_7_ ( .D(port0i[7]), .SIN(p0_ff1[6]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[7]) );
  SDFFQX1 p0_ff1_reg_3_ ( .D(port0i[3]), .SIN(p0_ff1[2]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[3]) );
  SDFFQX1 sdai_ff1_reg ( .D(sdai), .SIN(rxd0ff), .SMC(test_se), .C(clk), .Q(
        sdai_ff1) );
  SDFFQX1 reset_ff1_reg ( .D(reset), .SIN(port0ff[7]), .SMC(test_se), .C(clk), 
        .Q(reset_ff1) );
  INVX1 U5 ( .A(1'b1), .Y(t1ff) );
  INVX1 U7 ( .A(1'b1), .Y(t0ff) );
endmodule


module mcu51_cpu_a0 ( clkcpu, rst, mempsack, memack, memdatai, memaddr, 
        mempsrd, mempswr, memrd, memwr, memaddr_comb, mempsrd_comb, 
        mempswr_comb, memrd_comb, memwr_comb, cpu_hold, cpu_resume, irq, 
        intvect, intcall, retiinstr, newinstr, rmwinstr, waitstaten, ramdatai, 
        sfrdatai, ramsfraddr, ramdatao, ramoe, ramwe, sfroe, sfrwe, sfroe_r, 
        sfrwe_r, sfroe_comb_s, sfrwe_comb_s, pc_o, pc_ini, cs_run, instr, 
        codefetch_s, sfrack, ramsfraddr_comb, ramdatao_comb, ramoe_comb, 
        ramwe_comb, ckcon, pmw, p2sel, gf0, stop, idle, acc, b, rs, c, ac, ov, 
        p, f0, f1, dph, dpl, dps, dpc, p2, sp, test_si, test_so, test_se );
  input [7:0] memdatai;
  output [15:0] memaddr;
  output [15:0] memaddr_comb;
  input [4:0] intvect;
  input [7:0] ramdatai;
  input [7:0] sfrdatai;
  output [7:0] ramsfraddr;
  output [7:0] ramdatao;
  output [15:0] pc_o;
  input [15:0] pc_ini;
  output [7:0] instr;
  output [7:0] ramsfraddr_comb;
  output [7:0] ramdatao_comb;
  output [7:0] ckcon;
  output [7:0] acc;
  output [7:0] b;
  output [1:0] rs;
  output [7:0] dph;
  output [7:0] dpl;
  output [3:0] dps;
  output [5:0] dpc;
  output [7:0] p2;
  output [7:0] sp;
  input clkcpu, rst, mempsack, memack, cpu_hold, cpu_resume, irq, sfrack,
         test_si, test_se;
  output mempsrd, mempswr, memrd, memwr, mempsrd_comb, mempswr_comb,
         memrd_comb, memwr_comb, intcall, retiinstr, newinstr, rmwinstr,
         waitstaten, ramoe, ramwe, sfroe, sfrwe, sfroe_r, sfrwe_r,
         sfroe_comb_s, sfrwe_comb_s, cs_run, codefetch_s, ramoe_comb,
         ramwe_comb, pmw, p2sel, gf0, stop, idle, c, ac, ov, p, f0, f1,
         test_so;
  wire   N343, N344, N345, n2510, n2499, n2501, finishmul, finishdiv, N370,
         N371, N372, N480, N481, N482, N483, N484, N485, N486, N487, N488,
         N489, N490, N491, N492, N493, N494, N495, d_hold, idle_r,
         cpu_resume_fff, stop_r, ramsfrwe, N512, N515, N520, pdmode, interrupt,
         N582, N583, N584, N585, N589, N590, phase0_ff, newinstrlock, N670,
         N671, N672, N673, N674, N675, N676, N677, N679, N680, N681, N682,
         N683, N684, N685, N689, accactv, N10562, N10563, N10564, N10565,
         N10566, N10567, N10568, N10569, N10570, N10571, N10572, N10573,
         N10574, N10575, N10576, N10577, N10578, N10581, N10582, N10583,
         N10584, N10585, N10586, N10587, N10588, N10589, N11478, N11479,
         N11480, N11481, N11482, N11483, N11484, N11485, N11486, N11487,
         N11488, N11489, N11491, N11498, N11499, N11500, N11501, N11502,
         N11503, N11504, N11505, N11524, N11525, N11543, N11544, N11555,
         N12469, N12470, N12472, N12477, N12478, N12479, N12480, N12481,
         N12482, N12483, N12484, N12485, N12486, N12487, N12488, N12489,
         N12490, N12491, N12492, N12493, N12494, N12495, N12496, N12497,
         N12498, N12499, N12500, N12501, N12502, N12503, N12504, N12505,
         N12506, N12507, N12508, N12509, N12510, N12511, N12512, N12513,
         N12514, N12515, N12516, N12517, N12518, N12519, N12520, N12521,
         N12522, N12523, N12524, N12525, N12526, N12527, N12528, N12529,
         N12530, N12531, N12532, N12533, N12534, N12535, N12536, N12537,
         N12538, N12539, N12540, N12541, N12542, N12543, N12544, N12545,
         N12546, N12547, N12548, N12549, N12550, N12551, N12552, N12553,
         N12554, N12555, N12556, N12557, N12558, N12559, N12560, N12561,
         N12562, N12563, N12564, N12566, N12567, N12568, N12569, N12570,
         N12571, N12572, N12573, N12575, N12576, N12577, N12578, N12579,
         N12580, N12581, N12582, N12584, N12585, N12586, N12587, N12588,
         N12589, N12590, N12591, N12593, N12594, N12595, N12596, N12597,
         N12598, N12599, N12600, N12602, N12603, N12604, N12605, N12606,
         N12607, N12608, N12609, N12611, N12612, N12613, N12614, N12615,
         N12616, N12617, N12618, N12620, N12621, N12622, N12623, N12624,
         N12625, N12626, N12627, N12629, N12630, N12631, N12632, N12633,
         N12634, N12635, N12636, N12637, N12644, N12651, N12658, N12665,
         N12672, N12679, N12686, N12690, N12691, N12692, N12693, N12694,
         N12695, N12697, N12698, N12699, N12700, N12701, N12702, N12703,
         N12704, N12705, N12706, N12709, N12710, N12711, N12714, N12715,
         N12716, N12717, N12718, N12719, N12720, N12721, N12722, N12723,
         N12724, N12725, N12726, N12727, N12728, N12729, N12730, N12770,
         N12771, N12772, N12773, N12801, N12802, N12803, N12804, N12805,
         N12806, N12807, N12808, N12824, N12825, N12826, N12827, N12828,
         N12829, N12830, N12831, N12841, N12842, N12843, N12844, N12845,
         N12846, N12847, N12848, N12849, N12850, N12851, N12852, N12853,
         N12854, N12855, N12856, N12905, israccess, N12912, waitcnt_1_,
         waitcnt_0_, N12965, N12966, N12967, N12968, N12969, N12970, N12971,
         N12972, N12974, N12975, N12976, N12977, N13014, N13023, N13032,
         N13041, N13050, N13059, N13068, N13077, N13086, N13095, N13104,
         N13113, N13122, N13131, N13140, N13149, N13158, N13167, N13176,
         N13185, N13194, N13203, N13212, N13221, N13230, N13239, N13248,
         N13257, N13266, N13275, N13284, N13293, multemp1_0_, N13324, N13325,
         N13326, N13327, N13328, N13329, N13330, N13331, N13332, N13336,
         N13337, N13338, N13339, N13340, N13341, N13342, N13343, N13345,
         N13346, N13347, N13348, N13349, N13350, N13351, N13352, N13353,
         N13366, N13367, N13368, N13369, N13370, N13371, N13372, N13373,
         cpu_resume_ff1, N13379, N13380, net12389, net12395, net12400,
         net12405, net12410, net12415, net12420, net12425, net12430, net12435,
         net12440, net12445, net12450, net12455, net12460, net12465, net12470,
         net12475, net12480, net12485, net12490, net12495, net12500, net12505,
         net12510, net12515, net12520, net12525, net12530, net12535, net12540,
         net12545, net12550, net12555, net12560, net12565, net12570, net12575,
         net12580, net12585, net12590, net12595, net12600, net12605, net12610,
         net12615, net12620, net12625, net12630, net12635, net12640, net12645,
         net12650, net12655, net12660, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, N14351, N14350, N14349, N14348, N14347, N14346, N14345,
         N14344, N14343, N14342, N14341, N14340, N14339, N14338, N14337,
         N14336, n2503, n2502, n2504, n2508, n2506, n2507, n189, n190, n191,
         n192, n193, n194, n2509, n2505, n2500, n2031, n2032, n2036,
         multemp1_8_, multemp1_7_, multemp1_6_, multemp1_5_, multemp1_4_,
         multemp1_3_, multemp1_2_, multemp1_1_, n108, n127, n129, n206, n443,
         n444, n449, n450, n451, n456, n464, n466, n467, n475, n476, n477,
         n478, n479, n483, n488, n503, n504, n505, n506, n508, n509, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n580, n581, n582, n583, n584, n585, n586, n587, n588, n593,
         n594, n595, n599, n600, n601, n602, n603, n611, n613, n614, n638,
         n643, n648, n653, n664, n665, n672, n678, n684, n685, n690, n691,
         n692, n693, n698, n701, n706, n711, n716, n721, n726, n731, n736,
         n737, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n760, n761, n762, n763,
         n764, n766, n767, n768, n769, n770, n771, n772, n773, n774, n776,
         n777, n779, n780, n781, n783, n784, n785, n786, n788, n789, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n863, n864, n865, n866, n867, n869, n870, n871, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n887, n890, n891, n892, n894, n895, n899, n900, n901, n902, n906,
         n907, n908, n909, n910, n911, n912, n913, n917, n918, n922, n923,
         n927, n928, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n976, n977, n979, n980, n981, n983, n984, n985, n986, n987,
         n988, n989, n990, n992, n994, n996, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1335, n1336, n1337, n1338,
         n1339, n1340, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1370, n1372,
         n1374, n1375, n1376, n1377, n1378, n1379, n1382, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1408, n1409, n1413, n1414, n1415, n1416, n1417,
         n1419, n1420, n1421, n1422, n1423, n1425, n1427, n1428, n1429, n1430,
         n1431, n1435, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1491, n1492,
         n1493, n1494, n1496, n1497, n1498, n1510, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1536, n1546,
         n1548, n1549, n1550, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1564, n1565, n1566, n1567, n1568, n1569, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1618,
         n1620, n1622, n1623, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1639, n1640, n1641, n1644, n1648,
         n1649, n1650, n1651, n1662, n1663, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1689, n1690, n1698, n1702, n1704, n1706,
         n1710, n1722, n1723, n1725, n1726, n1727, n1735, n1736, n1742, n1744,
         n1745, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1989, n1990, n1991, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2033, n2034, n2037, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2144, n2150, n1, n2, n3,
         n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38, n39,
         n40, n42, n43, n44, n46, n48, n49, n50, n51, n53, n55, n57, n59, n61,
         n62, n63, n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n104, n105, n106, n107,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n128, n130, n131, n132, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n164, n165, n166, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n207, n208, n209, n210,
         n211, n212, n213, n214, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n445, n446, n447, n448, n452, n453,
         n454, n455, n457, n458, n459, n460, n461, n462, n463, n465, n468,
         n469, n470, n471, n472, n473, n474, n480, n481, n482, n484, n485,
         n486, n487, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n507, n510, n579, n589, n590, n591,
         n592, n596, n597, n598, n604, n605, n606, n607, n608, n609, n610,
         n612, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n639, n640, n641, n642, n644, n645, n646, n647, n649,
         n650, n651, n652, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n666, n667, n668, n669, n670, n671, n673, n674, n675,
         n676, n677, n679, n680, n681, n682, n683, n686, n687, n688, n689,
         n694, n695, n696, n697, n699, n700, n702, n703, n704, n705, n707,
         n708, n709, n710, n712, n713, n714, n715, n717, n718, n719, n720,
         n722, n723, n724, n725, n727, n728, n729, n730, n732, n733, n734,
         n735, n738, n739, n740, n741, n759, n765, n775, n778, n782, n787,
         n790, n791, n792, n793, n825, n826, n827, n828, n829, n830, n857,
         n858, n859, n860, n861, n862, n868, n872, n886, n888, n889, n893,
         n896, n897, n898, n903, n904, n905, n914, n915, n916, n919, n920,
         n921, n924, n925, n926, n929, n930, n931, n975, n978, n982, n991,
         n993, n995, n997, n1012, n1020, n1126, n1187, n1228, n1334, n1341,
         n1368, n1369, n1371, n1373, n1380, n1381, n1383, n1384, n1385, n1402,
         n1403, n1404, n1405, n1406, n1407, n1410, n1411, n1412, n1418, n1424,
         n1426, n1432, n1433, n1434, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1489, n1490, n1495, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1511, n1534, n1535, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1547, n1551, n1560,
         n1561, n1562, n1563, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1619,
         n1621, n1624, n1637, n1638, n1642, n1643, n1645, n1646, n1647, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1664,
         n1665, n1666, n1686, n1687, n1688, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1699, n1700, n1701, n1703, n1705, n1707, n1708, n1709,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1724, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1737,
         n1738, n1739, n1740, n1741, n1743, n1746, n1754, n1766, n1767, n1779,
         n1856, n1857, n1858, n1859, n1877, n1885, n1886, n1887, n1931, n1932,
         n1933, n1934, n1954, n1955, n1956, n1957, n1988, n1992, n1993, n1994,
         n1995, n2035, n2038, n2053, n2054, n2055, n2056, n2066, n2067, n2093,
         n2121, n2122, n2123, n2124, n2125, n2141, n2142, n2143, n2145, n2146,
         n2147, n2148, n2149, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         SYNOPSYS_UNCONNECTED_1;
  wire   [2:0] state;
  wire   [5:0] phase;
  wire   [15:0] alu_out;
  wire   [15:0] pc_i;
  wire   [7:0] temp;
  wire   [18:0] dec_accop;
  wire   [7:0] dec_cop;
  wire   [3:2] adder_out;
  wire   [9:1] multemp2;
  wire   [7:0] temp2_comb;
  wire   [15:0] dptr_inc;
  wire   [63:0] dpl_reg;
  wire   [63:0] dph_reg;
  wire   [47:0] dpc_tab;
  wire   [255:0] rn_reg;
  wire   [7:0] multempreg;
  wire   [6:0] divtempreg;
  wire   [3:2] add_1_root_add_5140_2_carry;

  FAD1X1 add_1_root_add_5140_2_U1_2 ( .A(N11524), .B(N11543), .CI(
        add_1_root_add_5140_2_carry[2]), .CO(add_1_root_add_5140_2_carry[3]), 
        .SO(adder_out[2]) );
  FAD1X1 add_1_root_add_5140_2_U1_3 ( .A(N11525), .B(N11544), .CI(
        add_1_root_add_5140_2_carry[3]), .CO(N11555), .SO(adder_out[3]) );
  MAJ3X1 U2627 ( .A(n1453), .B(n1454), .C(n1455), .Y(n1401) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 clk_gate_finishmul_reg ( .CLK(clkcpu), 
        .EN(N370), .ENCLK(net12389), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 clk_gate_instr_reg ( .CLK(clkcpu), .EN(
        N685), .ENCLK(net12395), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 clk_gate_bitno_reg ( .CLK(clkcpu), .EN(
        N11491), .ENCLK(net12400), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 clk_gate_dph_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N12556), .ENCLK(net12405), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 clk_gate_dph_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N12547), .ENCLK(net12410), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 clk_gate_dph_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N12538), .ENCLK(net12415), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 clk_gate_dph_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N12529), .ENCLK(net12420), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 clk_gate_dph_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N12520), .ENCLK(net12425), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 clk_gate_dph_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N12511), .ENCLK(net12430), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 clk_gate_dph_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N12502), .ENCLK(net12435), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 clk_gate_dph_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N12493), .ENCLK(net12440), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 clk_gate_dpc_tab_reg_7_ ( .CLK(clkcpu), 
        .EN(N12686), .ENCLK(net12445), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 clk_gate_dpc_tab_reg_6_ ( .CLK(clkcpu), 
        .EN(N12679), .ENCLK(net12450), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 clk_gate_dpc_tab_reg_5_ ( .CLK(clkcpu), 
        .EN(N12672), .ENCLK(net12455), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 clk_gate_dpc_tab_reg_4_ ( .CLK(clkcpu), 
        .EN(N12665), .ENCLK(net12460), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 clk_gate_dpc_tab_reg_3_ ( .CLK(clkcpu), 
        .EN(N12658), .ENCLK(net12465), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 clk_gate_dpc_tab_reg_2_ ( .CLK(clkcpu), 
        .EN(N12651), .ENCLK(net12470), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 clk_gate_dpc_tab_reg_1_ ( .CLK(clkcpu), 
        .EN(N12644), .ENCLK(net12475), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 clk_gate_dpc_tab_reg_0_ ( .CLK(clkcpu), 
        .EN(N12637), .ENCLK(net12480), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 clk_gate_temp_reg ( .CLK(clkcpu), .EN(
        N12722), .ENCLK(net12485), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 clk_gate_waitcnt_reg ( .CLK(clkcpu), 
        .EN(N12977), .ENCLK(net12490), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 clk_gate_rn_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N13293), .ENCLK(net12495), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 clk_gate_rn_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N13284), .ENCLK(net12500), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 clk_gate_rn_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N13275), .ENCLK(net12505), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 clk_gate_rn_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N13266), .ENCLK(net12510), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 clk_gate_rn_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N13257), .ENCLK(net12515), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 clk_gate_rn_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N13248), .ENCLK(net12520), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 clk_gate_rn_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N13239), .ENCLK(net12525), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 clk_gate_rn_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N13230), .ENCLK(net12530), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 clk_gate_rn_reg_reg_8_ ( .CLK(clkcpu), 
        .EN(N13221), .ENCLK(net12535), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 clk_gate_rn_reg_reg_9_ ( .CLK(clkcpu), 
        .EN(N13212), .ENCLK(net12540), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 clk_gate_rn_reg_reg_10_ ( .CLK(clkcpu), 
        .EN(N13203), .ENCLK(net12545), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 clk_gate_rn_reg_reg_11_ ( .CLK(clkcpu), 
        .EN(N13194), .ENCLK(net12550), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 clk_gate_rn_reg_reg_12_ ( .CLK(clkcpu), 
        .EN(N13185), .ENCLK(net12555), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 clk_gate_rn_reg_reg_13_ ( .CLK(clkcpu), 
        .EN(N13176), .ENCLK(net12560), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 clk_gate_rn_reg_reg_14_ ( .CLK(clkcpu), 
        .EN(N13167), .ENCLK(net12565), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 clk_gate_rn_reg_reg_15_ ( .CLK(clkcpu), 
        .EN(N13158), .ENCLK(net12570), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 clk_gate_rn_reg_reg_16_ ( .CLK(clkcpu), 
        .EN(N13149), .ENCLK(net12575), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 clk_gate_rn_reg_reg_17_ ( .CLK(clkcpu), 
        .EN(N13140), .ENCLK(net12580), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 clk_gate_rn_reg_reg_18_ ( .CLK(clkcpu), 
        .EN(N13131), .ENCLK(net12585), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 clk_gate_rn_reg_reg_19_ ( .CLK(clkcpu), 
        .EN(N13122), .ENCLK(net12590), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 clk_gate_rn_reg_reg_20_ ( .CLK(clkcpu), 
        .EN(N13113), .ENCLK(net12595), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 clk_gate_rn_reg_reg_21_ ( .CLK(clkcpu), 
        .EN(N13104), .ENCLK(net12600), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 clk_gate_rn_reg_reg_22_ ( .CLK(clkcpu), 
        .EN(N13095), .ENCLK(net12605), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 clk_gate_rn_reg_reg_23_ ( .CLK(clkcpu), 
        .EN(N13086), .ENCLK(net12610), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 clk_gate_rn_reg_reg_24_ ( .CLK(clkcpu), 
        .EN(N13077), .ENCLK(net12615), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 clk_gate_rn_reg_reg_25_ ( .CLK(clkcpu), 
        .EN(N13068), .ENCLK(net12620), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 clk_gate_rn_reg_reg_26_ ( .CLK(clkcpu), 
        .EN(N13059), .ENCLK(net12625), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 clk_gate_rn_reg_reg_27_ ( .CLK(clkcpu), 
        .EN(N13050), .ENCLK(net12630), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 clk_gate_rn_reg_reg_28_ ( .CLK(clkcpu), 
        .EN(N13041), .ENCLK(net12635), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 clk_gate_rn_reg_reg_29_ ( .CLK(clkcpu), 
        .EN(N13032), .ENCLK(net12640), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 clk_gate_rn_reg_reg_30_ ( .CLK(clkcpu), 
        .EN(N13023), .ENCLK(net12645), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 clk_gate_rn_reg_reg_31_ ( .CLK(clkcpu), 
        .EN(N13014), .ENCLK(net12650), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 clk_gate_multempreg_reg ( .CLK(clkcpu), 
        .EN(N13324), .ENCLK(net12655), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 clk_gate_divtempreg_reg ( .CLK(clkcpu), 
        .EN(N13366), .ENCLK(net12660), .TE(test_se) );
  mcu51_cpu_a0_DW01_add_0 add_5586 ( .A({n2235, n2235, n2235, n2235, n2235, 
        n2235, n2235, n2235, N12831, N12830, N12829, N12828, N12827, N12826, 
        N12825, N12824}), .B({N12856, N12855, N12854, N12853, N12852, N12851, 
        N12850, N12849, N12848, N12847, N12846, N12845, N12844, N12843, N12842, 
        N12841}), .CI(1'b0), .SUM(alu_out), .CO() );
  mcu51_cpu_a0_DW01_sub_0 sub_5969 ( .A({1'b0, n194, n193, n192, n191, n190, 
        n189, n2120, n77}), .B({1'b0, b}), .CI(1'b0), .DIFF({N13353, N13352, 
        N13351, N13350, N13349, N13348, N13347, N13346, N13345}), .CO() );
  mcu51_cpu_a0_DW01_sub_1 sub_5950 ( .A({1'b0, divtempreg, n90}), .B({1'b0, b}), .CI(1'b0), .DIFF({N13343, SYNOPSYS_UNCONNECTED_1, N13342, N13341, N13340, 
        N13339, N13338, N13337, N13336}), .CO() );
  mcu51_cpu_a0_DW01_inc_0 add_5525 ( .A({n108, n129, n127, N12773, N12772, 
        N12771, N12770, n206}), .SUM({N12808, N12807, N12806, N12805, N12804, 
        N12803, N12802, N12801}) );
  mcu51_cpu_a0_DW01_inc_1 add_5286 ( .A({n2128, n2129, n2130, n2131, n2132, 
        n2126, n2133, n2140, n2144, n2134, n2135, n2136, n2127, n2137, n2138, 
        n2139}), .SUM(dptr_inc) );
  mcu51_cpu_a0_DW01_inc_2 r715 ( .A({pc_o[15:11], n235, pc_o[9:0]}), .SUM(pc_i) );
  mcu51_cpu_a0_DW01_add_8 add_5901_aco ( .A({1'b0, multempreg}), .B({1'b0, 
        N14343, N14342, N14341, N14340, N14339, N14338, N14337, N14336}), .CI(
        1'b0), .SUM({multemp1_8_, multemp1_7_, multemp1_6_, multemp1_5_, 
        multemp1_4_, multemp1_3_, multemp1_2_, multemp1_1_, multemp1_0_}), 
        .CO() );
  mcu51_cpu_a0_DW01_add_7 add_5907_aco ( .A({1'b0, multemp1_8_, multemp1_7_, 
        multemp1_6_, multemp1_5_, multemp1_4_, multemp1_3_, multemp1_2_, 
        multemp1_1_}), .B({1'b0, N14351, N14350, N14349, N14348, N14347, 
        N14346, N14345, N14344}), .CI(1'b0), .SUM(multemp2), .CO() );
  SDFFQXL temp_reg_3_ ( .D(N12717), .SIN(temp[2]), .SMC(test_se), .C(net12485), 
        .Q(temp[3]) );
  SDFFQXL temp_reg_4_ ( .D(N12718), .SIN(temp[3]), .SMC(test_se), .C(net12485), 
        .Q(temp[4]) );
  SDFFQX1 pc_reg_2_ ( .D(N482), .SIN(memaddr[1]), .SMC(test_se), .C(net12389), 
        .Q(n2503) );
  SDFFQX1 pc_reg_5_ ( .D(N485), .SIN(n2502), .SMC(test_se), .C(net12389), .Q(
        memaddr[5]) );
  SDFFQX1 pc_reg_6_ ( .D(N486), .SIN(n50), .SMC(test_se), .C(net12389), .Q(
        pc_o[6]) );
  SDFFQX1 pc_reg_7_ ( .D(N487), .SIN(memaddr[6]), .SMC(test_se), .C(net12389), 
        .Q(memaddr[7]) );
  SDFFQX1 pc_reg_8_ ( .D(N488), .SIN(pc_o[7]), .SMC(test_se), .C(net12389), 
        .Q(pc_o[8]) );
  SDFFQX1 pc_reg_9_ ( .D(N489), .SIN(memaddr[8]), .SMC(test_se), .C(net12389), 
        .Q(pc_o[9]) );
  SDFFQX1 pc_reg_11_ ( .D(N491), .SIN(memaddr[10]), .SMC(test_se), .C(net12389), .Q(memaddr[11]) );
  SDFFQX1 pc_reg_12_ ( .D(N492), .SIN(pc_o[11]), .SMC(test_se), .C(net12389), 
        .Q(memaddr[12]) );
  SDFFQX1 pc_reg_13_ ( .D(N493), .SIN(pc_o[12]), .SMC(test_se), .C(net12389), 
        .Q(pc_o[13]) );
  SDFFQX1 pc_reg_14_ ( .D(N494), .SIN(pc_o[13]), .SMC(test_se), .C(net12389), 
        .Q(memaddr[14]) );
  SDFFQX1 pc_reg_15_ ( .D(N495), .SIN(pc_o[14]), .SMC(test_se), .C(net12389), 
        .Q(pc_o[15]) );
  SDFFQX1 cpu_resume_ff1_reg ( .D(N13379), .SIN(ckcon[7]), .SMC(test_se), .C(
        clkcpu), .Q(cpu_resume_ff1) );
  SDFFQX1 newinstrlock_reg ( .D(n1878), .SIN(multempreg[7]), .SMC(test_se), 
        .C(net12389), .Q(newinstrlock) );
  SDFFQX1 phase0_ff_reg ( .D(N689), .SIN(pdmode), .SMC(test_se), .C(net12389), 
        .Q(phase0_ff) );
  SDFFQX1 finishdiv_reg ( .D(N372), .SIN(f1), .SMC(test_se), .C(net12389), .Q(
        finishdiv) );
  SDFFQX1 finishmul_reg ( .D(N371), .SIN(finishdiv), .SMC(test_se), .C(
        net12389), .Q(finishmul) );
  SDFFQX1 multempreg_reg_7_ ( .D(N13332), .SIN(multempreg[6]), .SMC(test_se), 
        .C(net12655), .Q(multempreg[7]) );
  SDFFQX1 multempreg_reg_6_ ( .D(N13331), .SIN(multempreg[5]), .SMC(test_se), 
        .C(net12655), .Q(multempreg[6]) );
  SDFFQX1 multempreg_reg_5_ ( .D(N13330), .SIN(multempreg[4]), .SMC(test_se), 
        .C(net12655), .Q(multempreg[5]) );
  SDFFQX1 multempreg_reg_4_ ( .D(N13329), .SIN(multempreg[3]), .SMC(test_se), 
        .C(net12655), .Q(multempreg[4]) );
  SDFFQX1 cpu_resume_fff_reg ( .D(N13380), .SIN(cpu_resume_ff1), .SMC(test_se), 
        .C(clkcpu), .Q(cpu_resume_fff) );
  SDFFQX1 multempreg_reg_3_ ( .D(N13328), .SIN(multempreg[2]), .SMC(test_se), 
        .C(net12655), .Q(multempreg[3]) );
  SDFFQX1 pdmode_reg ( .D(n2036), .SIN(pc_o[15]), .SMC(test_se), .C(net12389), 
        .Q(pdmode) );
  SDFFQX1 d_hold_reg ( .D(cpu_hold), .SIN(cpu_resume_fff), .SMC(test_se), .C(
        clkcpu), .Q(d_hold) );
  SDFFQX1 multempreg_reg_2_ ( .D(N13327), .SIN(multempreg[1]), .SMC(test_se), 
        .C(net12655), .Q(multempreg[2]) );
  SDFFQX1 stop_r_reg ( .D(N515), .SIN(state[2]), .SMC(test_se), .C(net12389), 
        .Q(stop_r) );
  SDFFQX1 idle_r_reg ( .D(N512), .SIN(gf0), .SMC(test_se), .C(net12389), .Q(
        idle_r) );
  SDFFQX1 israccess_reg ( .D(N12912), .SIN(interrupt), .SMC(test_se), .C(
        net12389), .Q(israccess) );
  SDFFQX1 phase_reg_5_ ( .D(N684), .SIN(phase[4]), .SMC(test_se), .C(net12389), 
        .Q(phase[5]) );
  SDFFQX1 state_reg_2_ ( .D(N590), .SIN(state[1]), .SMC(test_se), .C(net12389), 
        .Q(state[2]) );
  SDFFQX1 state_reg_0_ ( .D(n2181), .SIN(sp[7]), .SMC(test_se), .C(net12389), 
        .Q(state[0]) );
  SDFFQX1 ramoe_r_reg ( .D(N11486), .SIN(ramdatao[7]), .SMC(test_se), .C(
        net12389), .Q(ramoe) );
  SDFFQX1 state_reg_1_ ( .D(N589), .SIN(state[0]), .SMC(test_se), .C(net12389), 
        .Q(state[1]) );
  SDFFQX1 phase_reg_4_ ( .D(N683), .SIN(phase[3]), .SMC(test_se), .C(net12389), 
        .Q(phase[4]) );
  SDFFQX1 phase_reg_3_ ( .D(N682), .SIN(phase[2]), .SMC(test_se), .C(net12389), 
        .Q(phase[3]) );
  SDFFQX1 f0_reg ( .D(n1882), .SIN(dps[3]), .SMC(test_se), .C(net12389), .Q(f0) );
  SDFFQX1 p2_reg_reg_5_ ( .D(N12490), .SIN(p2[4]), .SMC(test_se), .C(net12389), 
        .Q(p2[5]) );
  SDFFQX1 p2_reg_reg_4_ ( .D(N12489), .SIN(p2[3]), .SMC(test_se), .C(net12389), 
        .Q(p2[4]) );
  SDFFQX1 p_reg ( .D(N12905), .SIN(p2sel), .SMC(test_se), .C(net12389), .Q(p)
         );
  SDFFQX1 dpc_tab_reg_3__2_ ( .D(n264), .SIN(dpc_tab[19]), .SMC(test_se), .C(
        net12465), .Q(dpc_tab[20]) );
  SDFFQX1 dpc_tab_reg_7__2_ ( .D(n2191), .SIN(dpc_tab[43]), .SMC(test_se), .C(
        net12445), .Q(dpc_tab[44]) );
  SDFFQX1 dpc_tab_reg_2__2_ ( .D(n267), .SIN(dpc_tab[13]), .SMC(test_se), .C(
        net12470), .Q(dpc_tab[14]) );
  SDFFQX1 dpc_tab_reg_6__2_ ( .D(n267), .SIN(dpc_tab[37]), .SMC(test_se), .C(
        net12450), .Q(dpc_tab[38]) );
  SDFFQX1 rn_reg_reg_7__2_ ( .D(n267), .SIN(rn_reg[193]), .SMC(test_se), .C(
        net12530), .Q(rn_reg[194]) );
  SDFFQX1 rn_reg_reg_7__6_ ( .D(n268), .SIN(rn_reg[197]), .SMC(test_se), .C(
        net12530), .Q(rn_reg[198]) );
  SDFFQX1 rn_reg_reg_23__6_ ( .D(n2207), .SIN(rn_reg[69]), .SMC(test_se), .C(
        net12610), .Q(rn_reg[70]) );
  SDFFQX1 dpc_tab_reg_3__3_ ( .D(N12690), .SIN(dpc_tab[20]), .SMC(test_se), 
        .C(net12465), .Q(dpc_tab[21]) );
  SDFFQX1 dpc_tab_reg_7__3_ ( .D(N12690), .SIN(dpc_tab[44]), .SMC(test_se), 
        .C(net12445), .Q(dpc_tab[45]) );
  SDFFQX1 rn_reg_reg_31__6_ ( .D(n270), .SIN(rn_reg[5]), .SMC(test_se), .C(
        net12650), .Q(rn_reg[6]) );
  SDFFQX1 rn_reg_reg_15__6_ ( .D(n270), .SIN(rn_reg[133]), .SMC(test_se), .C(
        net12570), .Q(rn_reg[134]) );
  SDFFQX1 rn_reg_reg_15__5_ ( .D(n273), .SIN(rn_reg[132]), .SMC(test_se), .C(
        net12570), .Q(rn_reg[133]) );
  SDFFQX1 rn_reg_reg_15__2_ ( .D(n266), .SIN(rn_reg[129]), .SMC(test_se), .C(
        net12570), .Q(rn_reg[130]) );
  SDFFQX1 rn_reg_reg_4__2_ ( .D(n266), .SIN(rn_reg[217]), .SMC(test_se), .C(
        net12515), .Q(rn_reg[218]) );
  SDFFQX1 rn_reg_reg_4__6_ ( .D(n270), .SIN(rn_reg[221]), .SMC(test_se), .C(
        net12515), .Q(rn_reg[222]) );
  SDFFQX1 rn_reg_reg_20__6_ ( .D(n270), .SIN(rn_reg[93]), .SMC(test_se), .C(
        net12595), .Q(rn_reg[94]) );
  SDFFQX1 rn_reg_reg_28__6_ ( .D(n270), .SIN(rn_reg[29]), .SMC(test_se), .C(
        net12635), .Q(rn_reg[30]) );
  SDFFQX1 rn_reg_reg_12__6_ ( .D(n269), .SIN(rn_reg[157]), .SMC(test_se), .C(
        net12555), .Q(rn_reg[158]) );
  SDFFQX1 rn_reg_reg_12__2_ ( .D(n265), .SIN(rn_reg[153]), .SMC(test_se), .C(
        net12555), .Q(rn_reg[154]) );
  SDFFQX1 rn_reg_reg_5__2_ ( .D(n265), .SIN(rn_reg[209]), .SMC(test_se), .C(
        net12520), .Q(rn_reg[210]) );
  SDFFQX1 rn_reg_reg_5__6_ ( .D(n269), .SIN(rn_reg[213]), .SMC(test_se), .C(
        net12520), .Q(rn_reg[214]) );
  SDFFQX1 rn_reg_reg_5__5_ ( .D(n272), .SIN(rn_reg[212]), .SMC(test_se), .C(
        net12520), .Q(rn_reg[213]) );
  SDFFQX1 rn_reg_reg_21__6_ ( .D(n269), .SIN(rn_reg[85]), .SMC(test_se), .C(
        net12600), .Q(rn_reg[86]) );
  SDFFQX1 rn_reg_reg_21__2_ ( .D(n265), .SIN(rn_reg[81]), .SMC(test_se), .C(
        net12600), .Q(rn_reg[82]) );
  SDFFQX1 rn_reg_reg_29__6_ ( .D(n269), .SIN(rn_reg[21]), .SMC(test_se), .C(
        net12640), .Q(rn_reg[22]) );
  SDFFQX1 rn_reg_reg_13__6_ ( .D(n269), .SIN(rn_reg[149]), .SMC(test_se), .C(
        net12560), .Q(rn_reg[150]) );
  SDFFQX1 rn_reg_reg_13__2_ ( .D(n265), .SIN(rn_reg[145]), .SMC(test_se), .C(
        net12560), .Q(rn_reg[146]) );
  SDFFQX1 dpc_tab_reg_2__3_ ( .D(n2221), .SIN(dpc_tab[14]), .SMC(test_se), .C(
        net12470), .Q(dpc_tab[15]) );
  SDFFQX1 dpc_tab_reg_6__3_ ( .D(n2221), .SIN(dpc_tab[38]), .SMC(test_se), .C(
        net12450), .Q(dpc_tab[39]) );
  SDFFQX1 dpc_tab_reg_3__1_ ( .D(n252), .SIN(dpc_tab[18]), .SMC(test_se), .C(
        net12465), .Q(dpc_tab[19]) );
  SDFFQX1 dpc_tab_reg_7__1_ ( .D(n252), .SIN(dpc_tab[42]), .SMC(test_se), .C(
        net12445), .Q(dpc_tab[43]) );
  SDFFQX1 dpc_tab_reg_2__1_ ( .D(n251), .SIN(dpc_tab[12]), .SMC(test_se), .C(
        net12470), .Q(dpc_tab[13]) );
  SDFFQX1 dpc_tab_reg_6__1_ ( .D(n251), .SIN(dpc_tab[36]), .SMC(test_se), .C(
        net12450), .Q(dpc_tab[37]) );
  SDFFQX1 dpc_tab_reg_0__2_ ( .D(n2191), .SIN(dpc_tab[1]), .SMC(test_se), .C(
        net12480), .Q(dpc_tab[2]) );
  SDFFQX1 dpc_tab_reg_4__2_ ( .D(n267), .SIN(dpc_tab[25]), .SMC(test_se), .C(
        net12460), .Q(dpc_tab[26]) );
  SDFFQX1 dpc_tab_reg_1__2_ ( .D(n267), .SIN(dpc_tab[7]), .SMC(test_se), .C(
        net12475), .Q(dpc_tab[8]) );
  SDFFQX1 dpc_tab_reg_5__2_ ( .D(n267), .SIN(dpc_tab[31]), .SMC(test_se), .C(
        net12455), .Q(dpc_tab[32]) );
  SDFFQX1 rn_reg_reg_3__2_ ( .D(n267), .SIN(rn_reg[225]), .SMC(test_se), .C(
        net12510), .Q(rn_reg[226]) );
  SDFFQX1 rn_reg_reg_3__6_ ( .D(n2207), .SIN(rn_reg[229]), .SMC(test_se), .C(
        net12510), .Q(rn_reg[230]) );
  SDFFQX1 rn_reg_reg_3__5_ ( .D(n2214), .SIN(rn_reg[228]), .SMC(test_se), .C(
        net12510), .Q(rn_reg[229]) );
  SDFFQX1 rn_reg_reg_19__6_ ( .D(n2207), .SIN(rn_reg[101]), .SMC(test_se), .C(
        net12590), .Q(rn_reg[102]) );
  SDFFQX1 rn_reg_reg_19__2_ ( .D(n267), .SIN(rn_reg[97]), .SMC(test_se), .C(
        net12590), .Q(rn_reg[98]) );
  SDFFQX1 rn_reg_reg_27__6_ ( .D(n2207), .SIN(rn_reg[37]), .SMC(test_se), .C(
        net12630), .Q(rn_reg[38]) );
  SDFFQX1 rn_reg_reg_27__2_ ( .D(n267), .SIN(rn_reg[33]), .SMC(test_se), .C(
        net12630), .Q(rn_reg[34]) );
  SDFFQX1 rn_reg_reg_11__6_ ( .D(n270), .SIN(rn_reg[165]), .SMC(test_se), .C(
        net12550), .Q(rn_reg[166]) );
  SDFFQX1 rn_reg_reg_11__5_ ( .D(n273), .SIN(rn_reg[164]), .SMC(test_se), .C(
        net12550), .Q(rn_reg[165]) );
  SDFFQX1 rn_reg_reg_11__2_ ( .D(n266), .SIN(rn_reg[161]), .SMC(test_se), .C(
        net12550), .Q(rn_reg[162]) );
  SDFFQX1 rn_reg_reg_0__2_ ( .D(n266), .SIN(rn_reg[249]), .SMC(test_se), .C(
        net12495), .Q(rn_reg[250]) );
  SDFFQX1 rn_reg_reg_0__6_ ( .D(n270), .SIN(rn_reg[253]), .SMC(test_se), .C(
        net12495), .Q(rn_reg[254]) );
  SDFFQX1 rn_reg_reg_0__5_ ( .D(n273), .SIN(rn_reg[252]), .SMC(test_se), .C(
        net12495), .Q(rn_reg[253]) );
  SDFFQX1 rn_reg_reg_16__6_ ( .D(n270), .SIN(rn_reg[125]), .SMC(test_se), .C(
        net12575), .Q(rn_reg[126]) );
  SDFFQX1 rn_reg_reg_16__2_ ( .D(n266), .SIN(rn_reg[121]), .SMC(test_se), .C(
        net12575), .Q(rn_reg[122]) );
  SDFFQX1 dpc_tab_reg_0__3_ ( .D(n2221), .SIN(dpc_tab[2]), .SMC(test_se), .C(
        net12480), .Q(dpc_tab[3]) );
  SDFFQX1 dpc_tab_reg_4__3_ ( .D(n2221), .SIN(dpc_tab[26]), .SMC(test_se), .C(
        net12460), .Q(dpc_tab[27]) );
  SDFFQX1 rn_reg_reg_24__6_ ( .D(n270), .SIN(rn_reg[61]), .SMC(test_se), .C(
        net12615), .Q(rn_reg[62]) );
  SDFFQX1 rn_reg_reg_24__2_ ( .D(n266), .SIN(rn_reg[57]), .SMC(test_se), .C(
        net12615), .Q(rn_reg[58]) );
  SDFFQX1 rn_reg_reg_8__6_ ( .D(n270), .SIN(rn_reg[189]), .SMC(test_se), .C(
        net12535), .Q(rn_reg[190]) );
  SDFFQX1 rn_reg_reg_8__5_ ( .D(n272), .SIN(rn_reg[188]), .SMC(test_se), .C(
        net12535), .Q(rn_reg[189]) );
  SDFFQX1 rn_reg_reg_8__2_ ( .D(n265), .SIN(rn_reg[185]), .SMC(test_se), .C(
        net12535), .Q(rn_reg[186]) );
  SDFFQX1 rn_reg_reg_1__2_ ( .D(n265), .SIN(rn_reg[241]), .SMC(test_se), .C(
        net12500), .Q(rn_reg[242]) );
  SDFFQX1 rn_reg_reg_1__6_ ( .D(n269), .SIN(rn_reg[245]), .SMC(test_se), .C(
        net12500), .Q(rn_reg[246]) );
  SDFFQX1 rn_reg_reg_1__5_ ( .D(n272), .SIN(rn_reg[244]), .SMC(test_se), .C(
        net12500), .Q(rn_reg[245]) );
  SDFFQX1 rn_reg_reg_17__6_ ( .D(n269), .SIN(rn_reg[117]), .SMC(test_se), .C(
        net12580), .Q(rn_reg[118]) );
  SDFFQX1 rn_reg_reg_17__2_ ( .D(n265), .SIN(rn_reg[113]), .SMC(test_se), .C(
        net12580), .Q(rn_reg[114]) );
  SDFFQX1 dpc_tab_reg_1__3_ ( .D(N12690), .SIN(dpc_tab[8]), .SMC(test_se), .C(
        net12475), .Q(dpc_tab[9]) );
  SDFFQX1 dpc_tab_reg_5__0_ ( .D(n257), .SIN(dpc_tab[29]), .SMC(test_se), .C(
        net12455), .Q(dpc_tab[30]) );
  SDFFQX1 rn_reg_reg_26__6_ ( .D(n268), .SIN(rn_reg[45]), .SMC(test_se), .C(
        net12625), .Q(rn_reg[46]) );
  SDFFQX1 rn_reg_reg_26__2_ ( .D(n264), .SIN(rn_reg[41]), .SMC(test_se), .C(
        net12625), .Q(rn_reg[42]) );
  SDFFQX1 rn_reg_reg_10__6_ ( .D(n268), .SIN(rn_reg[173]), .SMC(test_se), .C(
        net12545), .Q(rn_reg[174]) );
  SDFFQX1 rn_reg_reg_10__5_ ( .D(n271), .SIN(rn_reg[172]), .SMC(test_se), .C(
        net12545), .Q(rn_reg[173]) );
  SDFFQX1 rn_reg_reg_10__2_ ( .D(n264), .SIN(rn_reg[169]), .SMC(test_se), .C(
        net12545), .Q(rn_reg[170]) );
  SDFFQX1 dpc_tab_reg_0__1_ ( .D(n252), .SIN(dpc_tab[0]), .SMC(test_se), .C(
        net12480), .Q(dpc_tab[1]) );
  SDFFQX1 dpc_tab_reg_4__1_ ( .D(n252), .SIN(dpc_tab[24]), .SMC(test_se), .C(
        net12460), .Q(dpc_tab[25]) );
  SDFFQX1 dpc_tab_reg_1__1_ ( .D(n251), .SIN(dpc_tab[6]), .SMC(test_se), .C(
        net12475), .Q(dpc_tab[7]) );
  SDFFQX1 dpc_tab_reg_5__3_ ( .D(N12690), .SIN(dpc_tab[32]), .SMC(test_se), 
        .C(net12455), .Q(dpc_tab[33]) );
  SDFFQX1 dpc_tab_reg_5__1_ ( .D(n251), .SIN(dpc_tab[30]), .SMC(test_se), .C(
        net12455), .Q(dpc_tab[31]) );
  SDFFQX1 rn_reg_reg_25__6_ ( .D(n269), .SIN(rn_reg[53]), .SMC(test_se), .C(
        net12620), .Q(rn_reg[54]) );
  SDFFQX1 rn_reg_reg_25__2_ ( .D(n265), .SIN(rn_reg[49]), .SMC(test_se), .C(
        net12620), .Q(rn_reg[50]) );
  SDFFQX1 rn_reg_reg_9__6_ ( .D(n269), .SIN(rn_reg[181]), .SMC(test_se), .C(
        net12540), .Q(rn_reg[182]) );
  SDFFQX1 rn_reg_reg_9__5_ ( .D(n272), .SIN(rn_reg[180]), .SMC(test_se), .C(
        net12540), .Q(rn_reg[181]) );
  SDFFQX1 rn_reg_reg_9__2_ ( .D(n266), .SIN(rn_reg[177]), .SMC(test_se), .C(
        net12540), .Q(rn_reg[178]) );
  SDFFQX1 rn_reg_reg_2__2_ ( .D(n264), .SIN(rn_reg[233]), .SMC(test_se), .C(
        net12505), .Q(rn_reg[234]) );
  SDFFQX1 rn_reg_reg_18__6_ ( .D(n268), .SIN(rn_reg[109]), .SMC(test_se), .C(
        net12585), .Q(rn_reg[110]) );
  SDFFQX1 rn_reg_reg_6__2_ ( .D(n264), .SIN(rn_reg[201]), .SMC(test_se), .C(
        net12525), .Q(rn_reg[202]) );
  SDFFQX1 rn_reg_reg_6__6_ ( .D(n268), .SIN(rn_reg[205]), .SMC(test_se), .C(
        net12525), .Q(rn_reg[206]) );
  SDFFQX1 rn_reg_reg_22__6_ ( .D(n268), .SIN(rn_reg[77]), .SMC(test_se), .C(
        net12605), .Q(rn_reg[78]) );
  SDFFQX1 rn_reg_reg_30__6_ ( .D(n268), .SIN(rn_reg[13]), .SMC(test_se), .C(
        net12645), .Q(rn_reg[14]) );
  SDFFQX1 rn_reg_reg_30__2_ ( .D(n264), .SIN(rn_reg[9]), .SMC(test_se), .C(
        net12645), .Q(rn_reg[10]) );
  SDFFQX1 rn_reg_reg_14__6_ ( .D(n268), .SIN(rn_reg[141]), .SMC(test_se), .C(
        net12565), .Q(rn_reg[142]) );
  SDFFQX1 rn_reg_reg_14__5_ ( .D(n271), .SIN(rn_reg[140]), .SMC(test_se), .C(
        net12565), .Q(rn_reg[141]) );
  SDFFQX1 rn_reg_reg_14__2_ ( .D(n265), .SIN(rn_reg[137]), .SMC(test_se), .C(
        net12565), .Q(rn_reg[138]) );
  SDFFQX1 dec_cop_reg_0_ ( .D(N10582), .SIN(dec_accop[18]), .SMC(test_se), .C(
        net12389), .Q(dec_cop[0]) );
  SDFFQX1 f1_reg ( .D(n1883), .SIN(f0), .SMC(test_se), .C(net12389), .Q(f1) );
  SDFFQX1 ov_reg_reg ( .D(N12711), .SIN(newinstrlock), .SMC(test_se), .C(
        net12389), .Q(ov) );
  SDFFQX1 dpl_reg_reg_3__3_ ( .D(N12596), .SIN(dpl_reg[26]), .SMC(test_se), 
        .C(net12425), .Q(dpl_reg[27]) );
  SDFFQX1 dpl_reg_reg_7__3_ ( .D(N12632), .SIN(dpl_reg[58]), .SMC(test_se), 
        .C(net12405), .Q(dpl_reg[59]) );
  SDFFQX1 dpl_reg_reg_7__2_ ( .D(N12631), .SIN(dpl_reg[57]), .SMC(test_se), 
        .C(net12405), .Q(dpl_reg[58]) );
  SDFFQX1 dph_reg_reg_7__7_ ( .D(N12564), .SIN(dph_reg[62]), .SMC(test_se), 
        .C(net12405), .Q(dph_reg[63]) );
  SDFFQX1 dpl_reg_reg_1__3_ ( .D(N12578), .SIN(dpl_reg[10]), .SMC(test_se), 
        .C(net12435), .Q(dpl_reg[11]) );
  SDFFQX1 dpl_reg_reg_5__3_ ( .D(N12614), .SIN(dpl_reg[42]), .SMC(test_se), 
        .C(net12415), .Q(dpl_reg[43]) );
  SDFFQX1 dpl_reg_reg_2__3_ ( .D(N12587), .SIN(dpl_reg[18]), .SMC(test_se), 
        .C(net12430), .Q(dpl_reg[19]) );
  SDFFQX1 dpl_reg_reg_6__3_ ( .D(N12623), .SIN(dpl_reg[50]), .SMC(test_se), 
        .C(net12410), .Q(dpl_reg[51]) );
  SDFFQX1 dpl_reg_reg_1__2_ ( .D(N12577), .SIN(dpl_reg[9]), .SMC(test_se), .C(
        net12435), .Q(dpl_reg[10]) );
  SDFFQX1 dpl_reg_reg_5__2_ ( .D(N12613), .SIN(dpl_reg[41]), .SMC(test_se), 
        .C(net12415), .Q(dpl_reg[42]) );
  SDFFQX1 dph_reg_reg_5__0_ ( .D(N12539), .SIN(dph_reg[39]), .SMC(test_se), 
        .C(net12415), .Q(dph_reg[40]) );
  SDFFQX1 dph_reg_reg_1__7_ ( .D(N12510), .SIN(dph_reg[14]), .SMC(test_se), 
        .C(net12435), .Q(dph_reg[15]) );
  SDFFQX1 dph_reg_reg_5__7_ ( .D(N12546), .SIN(dph_reg[46]), .SMC(test_se), 
        .C(net12415), .Q(dph_reg[47]) );
  SDFFQX1 dpl_reg_reg_0__3_ ( .D(N12569), .SIN(dpl_reg[2]), .SMC(test_se), .C(
        net12440), .Q(dpl_reg[3]) );
  SDFFQX1 dpl_reg_reg_4__3_ ( .D(N12605), .SIN(dpl_reg[34]), .SMC(test_se), 
        .C(net12420), .Q(dpl_reg[35]) );
  SDFFQX1 dpl_reg_reg_0__2_ ( .D(N12568), .SIN(dpl_reg[1]), .SMC(test_se), .C(
        net12440), .Q(dpl_reg[2]) );
  SDFFQX1 dpl_reg_reg_4__2_ ( .D(N12604), .SIN(dpl_reg[33]), .SMC(test_se), 
        .C(net12420), .Q(dpl_reg[34]) );
  SDFFQX1 dph_reg_reg_4__0_ ( .D(N12530), .SIN(dph_reg[31]), .SMC(test_se), 
        .C(net12420), .Q(dph_reg[32]) );
  SDFFQX1 dph_reg_reg_0__7_ ( .D(N12501), .SIN(dph_reg[6]), .SMC(test_se), .C(
        net12440), .Q(dph_reg[7]) );
  SDFFQX1 dph_reg_reg_4__7_ ( .D(N12537), .SIN(dph_reg[38]), .SMC(test_se), 
        .C(net12420), .Q(dph_reg[39]) );
  SDFFQX1 gf0_reg ( .D(n1881), .SIN(finishmul), .SMC(test_se), .C(net12389), 
        .Q(gf0) );
  SDFFQX1 p2sel_s_reg ( .D(N520), .SIN(p2[7]), .SMC(test_se), .C(net12389), 
        .Q(p2sel) );
  SDFFQX1 p2_reg_reg_7_ ( .D(N12492), .SIN(p2[6]), .SMC(test_se), .C(net12389), 
        .Q(p2[7]) );
  SDFFQX1 p2_reg_reg_3_ ( .D(N12488), .SIN(p2[2]), .SMC(test_se), .C(net12389), 
        .Q(p2[3]) );
  SDFFQX1 p2_reg_reg_6_ ( .D(N12491), .SIN(p2[5]), .SMC(test_se), .C(net12389), 
        .Q(p2[6]) );
  SDFFQX1 idle_s_reg ( .D(n1879), .SIN(idle_r), .SMC(test_se), .C(net12389), 
        .Q(idle) );
  SDFFQX1 stop_s_reg ( .D(n1880), .SIN(stop_r), .SMC(test_se), .C(net12389), 
        .Q(stop) );
  SDFFQX1 p2_reg_reg_0_ ( .D(N12485), .SIN(ov), .SMC(test_se), .C(net12389), 
        .Q(p2[0]) );
  SDFFQX1 dpc_tab_reg_3__5_ ( .D(n2214), .SIN(dpc_tab[22]), .SMC(test_se), .C(
        net12465), .Q(dpc_tab[23]) );
  SDFFQX1 dpc_tab_reg_3__4_ ( .D(N12691), .SIN(dpc_tab[21]), .SMC(test_se), 
        .C(net12465), .Q(dpc_tab[22]) );
  SDFFQX1 dpc_tab_reg_7__5_ ( .D(N12692), .SIN(dpc_tab[46]), .SMC(test_se), 
        .C(net12445), .Q(dpc_tab[47]) );
  SDFFQX1 dpc_tab_reg_7__4_ ( .D(N12691), .SIN(dpc_tab[45]), .SMC(test_se), 
        .C(net12445), .Q(dpc_tab[46]) );
  SDFFQX1 dpc_tab_reg_2__5_ ( .D(n2214), .SIN(dpc_tab[16]), .SMC(test_se), .C(
        net12470), .Q(dpc_tab[17]) );
  SDFFQX1 dpc_tab_reg_2__4_ ( .D(N12691), .SIN(dpc_tab[15]), .SMC(test_se), 
        .C(net12470), .Q(dpc_tab[16]) );
  SDFFQX1 dpc_tab_reg_6__5_ ( .D(N12692), .SIN(dpc_tab[40]), .SMC(test_se), 
        .C(net12450), .Q(dpc_tab[41]) );
  SDFFQX1 dpc_tab_reg_6__4_ ( .D(N12691), .SIN(dpc_tab[39]), .SMC(test_se), 
        .C(net12450), .Q(dpc_tab[40]) );
  SDFFQX1 rn_reg_reg_7__7_ ( .D(n2231), .SIN(rn_reg[198]), .SMC(test_se), .C(
        net12530), .Q(rn_reg[199]) );
  SDFFQX1 rn_reg_reg_7__1_ ( .D(n254), .SIN(rn_reg[192]), .SMC(test_se), .C(
        net12530), .Q(rn_reg[193]) );
  SDFFQX1 rn_reg_reg_7__0_ ( .D(n258), .SIN(rn_reg[207]), .SMC(test_se), .C(
        net12530), .Q(rn_reg[192]) );
  SDFFQX1 rn_reg_reg_7__5_ ( .D(n2214), .SIN(rn_reg[196]), .SMC(test_se), .C(
        net12530), .Q(rn_reg[197]) );
  SDFFQX1 rn_reg_reg_23__7_ ( .D(n2231), .SIN(rn_reg[70]), .SMC(test_se), .C(
        net12610), .Q(rn_reg[71]) );
  SDFFQX1 rn_reg_reg_23__5_ ( .D(n273), .SIN(rn_reg[68]), .SMC(test_se), .C(
        net12610), .Q(rn_reg[69]) );
  SDFFQX1 rn_reg_reg_23__2_ ( .D(n267), .SIN(rn_reg[65]), .SMC(test_se), .C(
        net12610), .Q(rn_reg[66]) );
  SDFFQX1 rn_reg_reg_23__1_ ( .D(n254), .SIN(rn_reg[64]), .SMC(test_se), .C(
        net12610), .Q(rn_reg[65]) );
  SDFFQX1 dpc_tab_reg_3__0_ ( .D(n258), .SIN(dpc_tab[17]), .SMC(test_se), .C(
        net12465), .Q(dpc_tab[18]) );
  SDFFQX1 dpc_tab_reg_7__0_ ( .D(n258), .SIN(dpc_tab[41]), .SMC(test_se), .C(
        net12445), .Q(dpc_tab[42]) );
  SDFFQX1 rn_reg_reg_31__7_ ( .D(n2231), .SIN(rn_reg[6]), .SMC(test_se), .C(
        net12650), .Q(rn_reg[7]) );
  SDFFQX1 rn_reg_reg_31__5_ ( .D(n273), .SIN(rn_reg[4]), .SMC(test_se), .C(
        net12650), .Q(rn_reg[5]) );
  SDFFQX1 rn_reg_reg_31__2_ ( .D(n266), .SIN(rn_reg[1]), .SMC(test_se), .C(
        net12650), .Q(rn_reg[2]) );
  SDFFQX1 rn_reg_reg_31__1_ ( .D(n254), .SIN(rn_reg[0]), .SMC(test_se), .C(
        net12650), .Q(rn_reg[1]) );
  SDFFQX1 rn_reg_reg_15__7_ ( .D(n2231), .SIN(rn_reg[134]), .SMC(test_se), .C(
        net12570), .Q(rn_reg[135]) );
  SDFFQX1 rn_reg_reg_15__1_ ( .D(n254), .SIN(rn_reg[128]), .SMC(test_se), .C(
        net12570), .Q(rn_reg[129]) );
  SDFFQX1 rn_reg_reg_15__0_ ( .D(n258), .SIN(rn_reg[143]), .SMC(test_se), .C(
        net12570), .Q(rn_reg[128]) );
  SDFFQX1 rn_reg_reg_4__7_ ( .D(n2231), .SIN(rn_reg[222]), .SMC(test_se), .C(
        net12515), .Q(rn_reg[223]) );
  SDFFQX1 rn_reg_reg_4__1_ ( .D(n254), .SIN(rn_reg[216]), .SMC(test_se), .C(
        net12515), .Q(rn_reg[217]) );
  SDFFQX1 rn_reg_reg_4__0_ ( .D(n258), .SIN(rn_reg[231]), .SMC(test_se), .C(
        net12515), .Q(rn_reg[216]) );
  SDFFQX1 rn_reg_reg_4__5_ ( .D(n273), .SIN(rn_reg[220]), .SMC(test_se), .C(
        net12515), .Q(rn_reg[221]) );
  SDFFQX1 rn_reg_reg_20__7_ ( .D(n280), .SIN(rn_reg[94]), .SMC(test_se), .C(
        net12595), .Q(rn_reg[95]) );
  SDFFQX1 rn_reg_reg_20__5_ ( .D(n273), .SIN(rn_reg[92]), .SMC(test_se), .C(
        net12595), .Q(rn_reg[93]) );
  SDFFQX1 rn_reg_reg_20__2_ ( .D(n266), .SIN(rn_reg[89]), .SMC(test_se), .C(
        net12595), .Q(rn_reg[90]) );
  SDFFQX1 rn_reg_reg_20__1_ ( .D(n254), .SIN(rn_reg[88]), .SMC(test_se), .C(
        net12595), .Q(rn_reg[89]) );
  SDFFQX1 rn_reg_reg_28__7_ ( .D(n280), .SIN(rn_reg[30]), .SMC(test_se), .C(
        net12635), .Q(rn_reg[31]) );
  SDFFQX1 rn_reg_reg_28__5_ ( .D(n272), .SIN(rn_reg[28]), .SMC(test_se), .C(
        net12635), .Q(rn_reg[29]) );
  SDFFQX1 rn_reg_reg_28__2_ ( .D(n266), .SIN(rn_reg[25]), .SMC(test_se), .C(
        net12635), .Q(rn_reg[26]) );
  SDFFQX1 rn_reg_reg_28__1_ ( .D(n254), .SIN(rn_reg[24]), .SMC(test_se), .C(
        net12635), .Q(rn_reg[25]) );
  SDFFQX1 rn_reg_reg_12__7_ ( .D(n280), .SIN(rn_reg[158]), .SMC(test_se), .C(
        net12555), .Q(rn_reg[159]) );
  SDFFQX1 rn_reg_reg_12__5_ ( .D(n272), .SIN(rn_reg[156]), .SMC(test_se), .C(
        net12555), .Q(rn_reg[157]) );
  SDFFQX1 rn_reg_reg_12__1_ ( .D(n253), .SIN(rn_reg[152]), .SMC(test_se), .C(
        net12555), .Q(rn_reg[153]) );
  SDFFQX1 rn_reg_reg_12__0_ ( .D(n257), .SIN(rn_reg[167]), .SMC(test_se), .C(
        net12555), .Q(rn_reg[152]) );
  SDFFQX1 rn_reg_reg_5__7_ ( .D(n280), .SIN(rn_reg[214]), .SMC(test_se), .C(
        net12520), .Q(rn_reg[215]) );
  SDFFQX1 rn_reg_reg_5__1_ ( .D(n253), .SIN(rn_reg[208]), .SMC(test_se), .C(
        net12520), .Q(rn_reg[209]) );
  SDFFQX1 rn_reg_reg_5__0_ ( .D(n257), .SIN(rn_reg[223]), .SMC(test_se), .C(
        net12520), .Q(rn_reg[208]) );
  SDFFQX1 rn_reg_reg_21__7_ ( .D(n280), .SIN(rn_reg[86]), .SMC(test_se), .C(
        net12600), .Q(rn_reg[87]) );
  SDFFQX1 rn_reg_reg_21__5_ ( .D(n272), .SIN(rn_reg[84]), .SMC(test_se), .C(
        net12600), .Q(rn_reg[85]) );
  SDFFQX1 rn_reg_reg_29__7_ ( .D(n281), .SIN(rn_reg[22]), .SMC(test_se), .C(
        net12640), .Q(rn_reg[23]) );
  SDFFQX1 rn_reg_reg_29__5_ ( .D(n272), .SIN(rn_reg[20]), .SMC(test_se), .C(
        net12640), .Q(rn_reg[21]) );
  SDFFQX1 rn_reg_reg_29__2_ ( .D(n265), .SIN(rn_reg[17]), .SMC(test_se), .C(
        net12640), .Q(rn_reg[18]) );
  SDFFQX1 rn_reg_reg_13__7_ ( .D(n281), .SIN(rn_reg[150]), .SMC(test_se), .C(
        net12560), .Q(rn_reg[151]) );
  SDFFQX1 rn_reg_reg_13__5_ ( .D(n271), .SIN(rn_reg[148]), .SMC(test_se), .C(
        net12560), .Q(rn_reg[149]) );
  SDFFQX1 rn_reg_reg_13__1_ ( .D(n253), .SIN(rn_reg[144]), .SMC(test_se), .C(
        net12560), .Q(rn_reg[145]) );
  SDFFQX1 rn_reg_reg_13__0_ ( .D(n257), .SIN(rn_reg[159]), .SMC(test_se), .C(
        net12560), .Q(rn_reg[144]) );
  SDFFQX1 dpc_tab_reg_2__0_ ( .D(n257), .SIN(dpc_tab[11]), .SMC(test_se), .C(
        net12470), .Q(dpc_tab[12]) );
  SDFFQX1 dpc_tab_reg_6__0_ ( .D(n256), .SIN(dpc_tab[35]), .SMC(test_se), .C(
        net12450), .Q(dpc_tab[36]) );
  SDFFQX1 rn_reg_reg_7__4_ ( .D(n2220), .SIN(rn_reg[195]), .SMC(test_se), .C(
        net12530), .Q(rn_reg[196]) );
  SDFFQX1 rn_reg_reg_23__3_ ( .D(n279), .SIN(rn_reg[66]), .SMC(test_se), .C(
        net12610), .Q(rn_reg[67]) );
  SDFFQX1 rn_reg_reg_23__0_ ( .D(n256), .SIN(rn_reg[79]), .SMC(test_se), .C(
        net12610), .Q(rn_reg[64]) );
  SDFFQX1 rn_reg_reg_31__4_ ( .D(n276), .SIN(rn_reg[3]), .SMC(test_se), .C(
        net12650), .Q(rn_reg[4]) );
  SDFFQX1 rn_reg_reg_31__3_ ( .D(n279), .SIN(rn_reg[2]), .SMC(test_se), .C(
        net12650), .Q(rn_reg[3]) );
  SDFFQX1 rn_reg_reg_31__0_ ( .D(n256), .SIN(rn_reg[15]), .SMC(test_se), .C(
        net12650), .Q(rn_reg[0]) );
  SDFFQX1 rn_reg_reg_15__4_ ( .D(n276), .SIN(rn_reg[131]), .SMC(test_se), .C(
        net12570), .Q(rn_reg[132]) );
  SDFFQX1 rn_reg_reg_4__4_ ( .D(n276), .SIN(rn_reg[219]), .SMC(test_se), .C(
        net12515), .Q(rn_reg[220]) );
  SDFFQX1 rn_reg_reg_20__3_ ( .D(n279), .SIN(rn_reg[90]), .SMC(test_se), .C(
        net12595), .Q(rn_reg[91]) );
  SDFFQX1 rn_reg_reg_20__0_ ( .D(n256), .SIN(rn_reg[103]), .SMC(test_se), .C(
        net12595), .Q(rn_reg[88]) );
  SDFFQX1 rn_reg_reg_28__3_ ( .D(n278), .SIN(rn_reg[26]), .SMC(test_se), .C(
        net12635), .Q(rn_reg[27]) );
  SDFFQX1 rn_reg_reg_28__0_ ( .D(n255), .SIN(rn_reg[39]), .SMC(test_se), .C(
        net12635), .Q(rn_reg[24]) );
  SDFFQX1 rn_reg_reg_12__4_ ( .D(n275), .SIN(rn_reg[155]), .SMC(test_se), .C(
        net12555), .Q(rn_reg[156]) );
  SDFFQX1 rn_reg_reg_5__4_ ( .D(n275), .SIN(rn_reg[211]), .SMC(test_se), .C(
        net12520), .Q(rn_reg[212]) );
  SDFFQX1 rn_reg_reg_21__4_ ( .D(n275), .SIN(rn_reg[83]), .SMC(test_se), .C(
        net12600), .Q(rn_reg[84]) );
  SDFFQX1 rn_reg_reg_21__3_ ( .D(n278), .SIN(rn_reg[82]), .SMC(test_se), .C(
        net12600), .Q(rn_reg[83]) );
  SDFFQX1 rn_reg_reg_21__1_ ( .D(n251), .SIN(rn_reg[80]), .SMC(test_se), .C(
        net12600), .Q(rn_reg[81]) );
  SDFFQX1 rn_reg_reg_21__0_ ( .D(n255), .SIN(rn_reg[95]), .SMC(test_se), .C(
        net12600), .Q(rn_reg[80]) );
  SDFFQX1 rn_reg_reg_29__3_ ( .D(n278), .SIN(rn_reg[18]), .SMC(test_se), .C(
        net12640), .Q(rn_reg[19]) );
  SDFFQX1 rn_reg_reg_29__1_ ( .D(n251), .SIN(rn_reg[16]), .SMC(test_se), .C(
        net12640), .Q(rn_reg[17]) );
  SDFFQX1 rn_reg_reg_29__0_ ( .D(n255), .SIN(rn_reg[31]), .SMC(test_se), .C(
        net12640), .Q(rn_reg[16]) );
  SDFFQX1 rn_reg_reg_13__4_ ( .D(n274), .SIN(rn_reg[147]), .SMC(test_se), .C(
        net12560), .Q(rn_reg[148]) );
  SDFFQX1 dpc_tab_reg_0__5_ ( .D(n2214), .SIN(dpc_tab[4]), .SMC(test_se), .C(
        net12480), .Q(dpc_tab[5]) );
  SDFFQX1 dpc_tab_reg_0__4_ ( .D(n2220), .SIN(dpc_tab[3]), .SMC(test_se), .C(
        net12480), .Q(dpc_tab[4]) );
  SDFFQX1 dpc_tab_reg_4__5_ ( .D(N12692), .SIN(dpc_tab[28]), .SMC(test_se), 
        .C(net12460), .Q(dpc_tab[29]) );
  SDFFQX1 dpc_tab_reg_4__4_ ( .D(n2220), .SIN(dpc_tab[27]), .SMC(test_se), .C(
        net12460), .Q(dpc_tab[28]) );
  SDFFQX1 dpc_tab_reg_1__5_ ( .D(n2214), .SIN(dpc_tab[10]), .SMC(test_se), .C(
        net12475), .Q(dpc_tab[11]) );
  SDFFQX1 dpc_tab_reg_1__4_ ( .D(n2220), .SIN(dpc_tab[9]), .SMC(test_se), .C(
        net12475), .Q(dpc_tab[10]) );
  SDFFQX1 dpc_tab_reg_5__5_ ( .D(N12692), .SIN(dpc_tab[34]), .SMC(test_se), 
        .C(net12455), .Q(dpc_tab[35]) );
  SDFFQX1 dpc_tab_reg_5__4_ ( .D(n2220), .SIN(dpc_tab[33]), .SMC(test_se), .C(
        net12455), .Q(dpc_tab[34]) );
  SDFFQX1 rn_reg_reg_3__7_ ( .D(n2231), .SIN(rn_reg[230]), .SMC(test_se), .C(
        net12510), .Q(rn_reg[231]) );
  SDFFQX1 rn_reg_reg_3__1_ ( .D(n2176), .SIN(rn_reg[224]), .SMC(test_se), .C(
        net12510), .Q(rn_reg[225]) );
  SDFFQX1 rn_reg_reg_3__0_ ( .D(n2177), .SIN(rn_reg[239]), .SMC(test_se), .C(
        net12510), .Q(rn_reg[224]) );
  SDFFQX1 rn_reg_reg_19__7_ ( .D(n2231), .SIN(rn_reg[102]), .SMC(test_se), .C(
        net12590), .Q(rn_reg[103]) );
  SDFFQX1 rn_reg_reg_19__5_ ( .D(n2214), .SIN(rn_reg[100]), .SMC(test_se), .C(
        net12590), .Q(rn_reg[101]) );
  SDFFQX1 rn_reg_reg_19__1_ ( .D(n254), .SIN(rn_reg[96]), .SMC(test_se), .C(
        net12590), .Q(rn_reg[97]) );
  SDFFQX1 rn_reg_reg_27__7_ ( .D(n2231), .SIN(rn_reg[38]), .SMC(test_se), .C(
        net12630), .Q(rn_reg[39]) );
  SDFFQX1 rn_reg_reg_27__5_ ( .D(n273), .SIN(rn_reg[36]), .SMC(test_se), .C(
        net12630), .Q(rn_reg[37]) );
  SDFFQX1 rn_reg_reg_11__7_ ( .D(n2231), .SIN(rn_reg[166]), .SMC(test_se), .C(
        net12550), .Q(rn_reg[167]) );
  SDFFQX1 rn_reg_reg_11__1_ ( .D(n254), .SIN(rn_reg[160]), .SMC(test_se), .C(
        net12550), .Q(rn_reg[161]) );
  SDFFQX1 rn_reg_reg_11__0_ ( .D(n258), .SIN(rn_reg[175]), .SMC(test_se), .C(
        net12550), .Q(rn_reg[160]) );
  SDFFQX1 rn_reg_reg_0__7_ ( .D(n282), .SIN(rn_reg[254]), .SMC(test_se), .C(
        net12495), .Q(rn_reg[255]) );
  SDFFQX1 rn_reg_reg_0__1_ ( .D(n254), .SIN(rn_reg[248]), .SMC(test_se), .C(
        net12495), .Q(rn_reg[249]) );
  SDFFQX1 rn_reg_reg_0__0_ ( .D(n258), .SIN(rmwinstr), .SMC(test_se), .C(
        net12495), .Q(rn_reg[248]) );
  SDFFQX1 rn_reg_reg_16__7_ ( .D(n280), .SIN(rn_reg[126]), .SMC(test_se), .C(
        net12575), .Q(rn_reg[127]) );
  SDFFQX1 rn_reg_reg_16__5_ ( .D(n273), .SIN(rn_reg[124]), .SMC(test_se), .C(
        net12575), .Q(rn_reg[125]) );
  SDFFQX1 dpc_tab_reg_0__0_ ( .D(n258), .SIN(divtempreg[6]), .SMC(test_se), 
        .C(net12480), .Q(dpc_tab[0]) );
  SDFFQX1 dpc_tab_reg_4__0_ ( .D(n258), .SIN(dpc_tab[23]), .SMC(test_se), .C(
        net12460), .Q(dpc_tab[24]) );
  SDFFQX1 rn_reg_reg_24__7_ ( .D(n280), .SIN(rn_reg[62]), .SMC(test_se), .C(
        net12615), .Q(rn_reg[63]) );
  SDFFQX1 rn_reg_reg_24__5_ ( .D(n273), .SIN(rn_reg[60]), .SMC(test_se), .C(
        net12615), .Q(rn_reg[61]) );
  SDFFQX1 rn_reg_reg_8__7_ ( .D(n280), .SIN(rn_reg[190]), .SMC(test_se), .C(
        net12535), .Q(rn_reg[191]) );
  SDFFQX1 rn_reg_reg_8__1_ ( .D(n253), .SIN(rn_reg[184]), .SMC(test_se), .C(
        net12535), .Q(rn_reg[185]) );
  SDFFQX1 rn_reg_reg_8__0_ ( .D(n258), .SIN(rn_reg[199]), .SMC(test_se), .C(
        net12535), .Q(rn_reg[184]) );
  SDFFQX1 rn_reg_reg_1__7_ ( .D(n280), .SIN(rn_reg[246]), .SMC(test_se), .C(
        net12500), .Q(rn_reg[247]) );
  SDFFQX1 rn_reg_reg_1__1_ ( .D(n253), .SIN(rn_reg[240]), .SMC(test_se), .C(
        net12500), .Q(rn_reg[241]) );
  SDFFQX1 rn_reg_reg_1__0_ ( .D(n257), .SIN(rn_reg[255]), .SMC(test_se), .C(
        net12500), .Q(rn_reg[240]) );
  SDFFQX1 rn_reg_reg_17__7_ ( .D(n280), .SIN(rn_reg[118]), .SMC(test_se), .C(
        net12580), .Q(rn_reg[119]) );
  SDFFQX1 rn_reg_reg_17__5_ ( .D(n272), .SIN(rn_reg[116]), .SMC(test_se), .C(
        net12580), .Q(rn_reg[117]) );
  SDFFQX1 dpc_tab_reg_1__0_ ( .D(n257), .SIN(dpc_tab[5]), .SMC(test_se), .C(
        net12475), .Q(dpc_tab[6]) );
  SDFFQX1 rn_reg_reg_26__7_ ( .D(n281), .SIN(rn_reg[46]), .SMC(test_se), .C(
        net12625), .Q(rn_reg[47]) );
  SDFFQX1 rn_reg_reg_26__5_ ( .D(n271), .SIN(rn_reg[44]), .SMC(test_se), .C(
        net12625), .Q(rn_reg[45]) );
  SDFFQX1 rn_reg_reg_10__7_ ( .D(n282), .SIN(rn_reg[174]), .SMC(test_se), .C(
        net12545), .Q(rn_reg[175]) );
  SDFFQX1 rn_reg_reg_10__1_ ( .D(n252), .SIN(rn_reg[168]), .SMC(test_se), .C(
        net12545), .Q(rn_reg[169]) );
  SDFFQX1 rn_reg_reg_10__0_ ( .D(n256), .SIN(rn_reg[183]), .SMC(test_se), .C(
        net12545), .Q(rn_reg[168]) );
  SDFFQX1 rn_reg_reg_3__3_ ( .D(n2221), .SIN(rn_reg[226]), .SMC(test_se), .C(
        net12510), .Q(rn_reg[227]) );
  SDFFQX1 rn_reg_reg_3__4_ ( .D(n2220), .SIN(rn_reg[227]), .SMC(test_se), .C(
        net12510), .Q(rn_reg[228]) );
  SDFFQX1 rn_reg_reg_19__4_ ( .D(n2220), .SIN(rn_reg[99]), .SMC(test_se), .C(
        net12590), .Q(rn_reg[100]) );
  SDFFQX1 rn_reg_reg_19__3_ ( .D(n2221), .SIN(rn_reg[98]), .SMC(test_se), .C(
        net12590), .Q(rn_reg[99]) );
  SDFFQX1 rn_reg_reg_19__0_ ( .D(n256), .SIN(rn_reg[111]), .SMC(test_se), .C(
        net12590), .Q(rn_reg[96]) );
  SDFFQX1 rn_reg_reg_27__4_ ( .D(n276), .SIN(rn_reg[35]), .SMC(test_se), .C(
        net12630), .Q(rn_reg[36]) );
  SDFFQX1 rn_reg_reg_27__3_ ( .D(n279), .SIN(rn_reg[34]), .SMC(test_se), .C(
        net12630), .Q(rn_reg[35]) );
  SDFFQX1 rn_reg_reg_27__1_ ( .D(n252), .SIN(rn_reg[32]), .SMC(test_se), .C(
        net12630), .Q(rn_reg[33]) );
  SDFFQX1 rn_reg_reg_27__0_ ( .D(n256), .SIN(rn_reg[47]), .SMC(test_se), .C(
        net12630), .Q(rn_reg[32]) );
  SDFFQX1 rn_reg_reg_11__4_ ( .D(n276), .SIN(rn_reg[163]), .SMC(test_se), .C(
        net12550), .Q(rn_reg[164]) );
  SDFFQX1 rn_reg_reg_11__3_ ( .D(n279), .SIN(rn_reg[162]), .SMC(test_se), .C(
        net12550), .Q(rn_reg[163]) );
  SDFFQX1 rn_reg_reg_0__3_ ( .D(n279), .SIN(rn_reg[250]), .SMC(test_se), .C(
        net12495), .Q(rn_reg[251]) );
  SDFFQX1 rn_reg_reg_0__4_ ( .D(n276), .SIN(rn_reg[251]), .SMC(test_se), .C(
        net12495), .Q(rn_reg[252]) );
  SDFFQX1 rn_reg_reg_16__4_ ( .D(n276), .SIN(rn_reg[123]), .SMC(test_se), .C(
        net12575), .Q(rn_reg[124]) );
  SDFFQX1 rn_reg_reg_16__3_ ( .D(n279), .SIN(rn_reg[122]), .SMC(test_se), .C(
        net12575), .Q(rn_reg[123]) );
  SDFFQX1 rn_reg_reg_16__1_ ( .D(n252), .SIN(rn_reg[120]), .SMC(test_se), .C(
        net12575), .Q(rn_reg[121]) );
  SDFFQX1 rn_reg_reg_16__0_ ( .D(n256), .SIN(rn_reg[135]), .SMC(test_se), .C(
        net12575), .Q(rn_reg[120]) );
  SDFFQX1 rn_reg_reg_24__4_ ( .D(n276), .SIN(rn_reg[59]), .SMC(test_se), .C(
        net12615), .Q(rn_reg[60]) );
  SDFFQX1 rn_reg_reg_24__3_ ( .D(n279), .SIN(rn_reg[58]), .SMC(test_se), .C(
        net12615), .Q(rn_reg[59]) );
  SDFFQX1 rn_reg_reg_24__1_ ( .D(n252), .SIN(rn_reg[56]), .SMC(test_se), .C(
        net12615), .Q(rn_reg[57]) );
  SDFFQX1 rn_reg_reg_24__0_ ( .D(n256), .SIN(rn_reg[71]), .SMC(test_se), .C(
        net12615), .Q(rn_reg[56]) );
  SDFFQX1 rn_reg_reg_8__4_ ( .D(n275), .SIN(rn_reg[187]), .SMC(test_se), .C(
        net12535), .Q(rn_reg[188]) );
  SDFFQX1 rn_reg_reg_8__3_ ( .D(n278), .SIN(rn_reg[186]), .SMC(test_se), .C(
        net12535), .Q(rn_reg[187]) );
  SDFFQX1 rn_reg_reg_1__3_ ( .D(n278), .SIN(rn_reg[242]), .SMC(test_se), .C(
        net12500), .Q(rn_reg[243]) );
  SDFFQX1 rn_reg_reg_1__4_ ( .D(n275), .SIN(rn_reg[243]), .SMC(test_se), .C(
        net12500), .Q(rn_reg[244]) );
  SDFFQX1 rn_reg_reg_17__4_ ( .D(n275), .SIN(rn_reg[115]), .SMC(test_se), .C(
        net12580), .Q(rn_reg[116]) );
  SDFFQX1 rn_reg_reg_17__3_ ( .D(n278), .SIN(rn_reg[114]), .SMC(test_se), .C(
        net12580), .Q(rn_reg[115]) );
  SDFFQX1 rn_reg_reg_17__1_ ( .D(n251), .SIN(rn_reg[112]), .SMC(test_se), .C(
        net12580), .Q(rn_reg[113]) );
  SDFFQX1 rn_reg_reg_17__0_ ( .D(n255), .SIN(rn_reg[127]), .SMC(test_se), .C(
        net12580), .Q(rn_reg[112]) );
  SDFFQX1 rn_reg_reg_26__4_ ( .D(n274), .SIN(rn_reg[43]), .SMC(test_se), .C(
        net12625), .Q(rn_reg[44]) );
  SDFFQX1 rn_reg_reg_26__3_ ( .D(n277), .SIN(rn_reg[42]), .SMC(test_se), .C(
        net12625), .Q(rn_reg[43]) );
  SDFFQX1 rn_reg_reg_26__1_ ( .D(n251), .SIN(rn_reg[40]), .SMC(test_se), .C(
        net12625), .Q(rn_reg[41]) );
  SDFFQX1 rn_reg_reg_26__0_ ( .D(n255), .SIN(rn_reg[55]), .SMC(test_se), .C(
        net12625), .Q(rn_reg[40]) );
  SDFFQX1 rn_reg_reg_10__4_ ( .D(n274), .SIN(rn_reg[171]), .SMC(test_se), .C(
        net12545), .Q(rn_reg[172]) );
  SDFFQX1 rn_reg_reg_25__7_ ( .D(n281), .SIN(rn_reg[54]), .SMC(test_se), .C(
        net12620), .Q(rn_reg[55]) );
  SDFFQX1 rn_reg_reg_25__5_ ( .D(n272), .SIN(rn_reg[52]), .SMC(test_se), .C(
        net12620), .Q(rn_reg[53]) );
  SDFFQX1 rn_reg_reg_9__7_ ( .D(n281), .SIN(rn_reg[182]), .SMC(test_se), .C(
        net12540), .Q(rn_reg[183]) );
  SDFFQX1 rn_reg_reg_9__1_ ( .D(n253), .SIN(rn_reg[176]), .SMC(test_se), .C(
        net12540), .Q(rn_reg[177]) );
  SDFFQX1 rn_reg_reg_25__4_ ( .D(n275), .SIN(rn_reg[51]), .SMC(test_se), .C(
        net12620), .Q(rn_reg[52]) );
  SDFFQX1 rn_reg_reg_25__3_ ( .D(n278), .SIN(rn_reg[50]), .SMC(test_se), .C(
        net12620), .Q(rn_reg[51]) );
  SDFFQX1 rn_reg_reg_25__1_ ( .D(n251), .SIN(rn_reg[48]), .SMC(test_se), .C(
        net12620), .Q(rn_reg[49]) );
  SDFFQX1 rn_reg_reg_25__0_ ( .D(n255), .SIN(rn_reg[63]), .SMC(test_se), .C(
        net12620), .Q(rn_reg[48]) );
  SDFFQX1 rn_reg_reg_9__4_ ( .D(n275), .SIN(rn_reg[179]), .SMC(test_se), .C(
        net12540), .Q(rn_reg[180]) );
  SDFFQX1 rn_reg_reg_9__3_ ( .D(n278), .SIN(rn_reg[178]), .SMC(test_se), .C(
        net12540), .Q(rn_reg[179]) );
  SDFFQX1 rn_reg_reg_9__0_ ( .D(n255), .SIN(rn_reg[191]), .SMC(test_se), .C(
        net12540), .Q(rn_reg[176]) );
  SDFFQX1 rn_reg_reg_2__7_ ( .D(n281), .SIN(rn_reg[238]), .SMC(test_se), .C(
        net12505), .Q(rn_reg[239]) );
  SDFFQX1 rn_reg_reg_2__1_ ( .D(n253), .SIN(rn_reg[232]), .SMC(test_se), .C(
        net12505), .Q(rn_reg[233]) );
  SDFFQX1 rn_reg_reg_2__0_ ( .D(n257), .SIN(rn_reg[247]), .SMC(test_se), .C(
        net12505), .Q(rn_reg[232]) );
  SDFFQX1 rn_reg_reg_2__6_ ( .D(n269), .SIN(rn_reg[237]), .SMC(test_se), .C(
        net12505), .Q(rn_reg[238]) );
  SDFFQX1 rn_reg_reg_2__5_ ( .D(n271), .SIN(rn_reg[236]), .SMC(test_se), .C(
        net12505), .Q(rn_reg[237]) );
  SDFFQX1 rn_reg_reg_18__7_ ( .D(n281), .SIN(rn_reg[110]), .SMC(test_se), .C(
        net12585), .Q(rn_reg[111]) );
  SDFFQX1 rn_reg_reg_18__5_ ( .D(n271), .SIN(rn_reg[108]), .SMC(test_se), .C(
        net12585), .Q(rn_reg[109]) );
  SDFFQX1 rn_reg_reg_18__2_ ( .D(n264), .SIN(rn_reg[105]), .SMC(test_se), .C(
        net12585), .Q(rn_reg[106]) );
  SDFFQX1 rn_reg_reg_18__0_ ( .D(n255), .SIN(rn_reg[119]), .SMC(test_se), .C(
        net12585), .Q(rn_reg[104]) );
  SDFFQX1 rn_reg_reg_6__7_ ( .D(n281), .SIN(rn_reg[206]), .SMC(test_se), .C(
        net12525), .Q(rn_reg[207]) );
  SDFFQX1 rn_reg_reg_6__1_ ( .D(n253), .SIN(rn_reg[200]), .SMC(test_se), .C(
        net12525), .Q(rn_reg[201]) );
  SDFFQX1 rn_reg_reg_6__0_ ( .D(n257), .SIN(rn_reg[215]), .SMC(test_se), .C(
        net12525), .Q(rn_reg[200]) );
  SDFFQX1 rn_reg_reg_6__5_ ( .D(n271), .SIN(rn_reg[204]), .SMC(test_se), .C(
        net12525), .Q(rn_reg[205]) );
  SDFFQX1 rn_reg_reg_22__7_ ( .D(n281), .SIN(rn_reg[78]), .SMC(test_se), .C(
        net12605), .Q(rn_reg[79]) );
  SDFFQX1 rn_reg_reg_22__5_ ( .D(n271), .SIN(rn_reg[76]), .SMC(test_se), .C(
        net12605), .Q(rn_reg[77]) );
  SDFFQX1 rn_reg_reg_22__2_ ( .D(n264), .SIN(rn_reg[73]), .SMC(test_se), .C(
        net12605), .Q(rn_reg[74]) );
  SDFFQX1 rn_reg_reg_22__1_ ( .D(n253), .SIN(rn_reg[72]), .SMC(test_se), .C(
        net12605), .Q(rn_reg[73]) );
  SDFFQX1 rn_reg_reg_22__0_ ( .D(n257), .SIN(rn_reg[87]), .SMC(test_se), .C(
        net12605), .Q(rn_reg[72]) );
  SDFFQX1 rn_reg_reg_30__7_ ( .D(n281), .SIN(rn_reg[14]), .SMC(test_se), .C(
        net12645), .Q(rn_reg[15]) );
  SDFFQX1 rn_reg_reg_30__5_ ( .D(n271), .SIN(rn_reg[12]), .SMC(test_se), .C(
        net12645), .Q(rn_reg[13]) );
  SDFFQX1 rn_reg_reg_30__1_ ( .D(n252), .SIN(rn_reg[8]), .SMC(test_se), .C(
        net12645), .Q(rn_reg[9]) );
  SDFFQX1 rn_reg_reg_14__7_ ( .D(n282), .SIN(rn_reg[142]), .SMC(test_se), .C(
        net12565), .Q(rn_reg[143]) );
  SDFFQX1 rn_reg_reg_14__1_ ( .D(n252), .SIN(rn_reg[136]), .SMC(test_se), .C(
        net12565), .Q(rn_reg[137]) );
  SDFFQX1 rn_reg_reg_14__0_ ( .D(n256), .SIN(rn_reg[151]), .SMC(test_se), .C(
        net12565), .Q(rn_reg[136]) );
  SDFFQX1 rn_reg_reg_30__4_ ( .D(n274), .SIN(rn_reg[11]), .SMC(test_se), .C(
        net12645), .Q(rn_reg[12]) );
  SDFFQX1 rn_reg_reg_30__0_ ( .D(n255), .SIN(rn_reg[23]), .SMC(test_se), .C(
        net12645), .Q(rn_reg[8]) );
  SDFFQX1 rn_reg_reg_14__4_ ( .D(n274), .SIN(rn_reg[139]), .SMC(test_se), .C(
        net12565), .Q(rn_reg[140]) );
  SDFFQX1 sp_reg_reg_7_ ( .D(N12704), .SIN(sp[6]), .SMC(test_se), .C(net12389), 
        .Q(sp[7]) );
  SDFFQX1 dph_reg_reg_3__2_ ( .D(N12523), .SIN(dph_reg[25]), .SMC(test_se), 
        .C(net12425), .Q(dph_reg[26]) );
  SDFFQX1 dph_reg_reg_7__2_ ( .D(N12559), .SIN(dph_reg[57]), .SMC(test_se), 
        .C(net12405), .Q(dph_reg[58]) );
  SDFFQX1 dph_reg_reg_3__7_ ( .D(N12528), .SIN(dph_reg[30]), .SMC(test_se), 
        .C(net12425), .Q(dph_reg[31]) );
  SDFFQX1 dph_reg_reg_3__5_ ( .D(N12526), .SIN(dph_reg[28]), .SMC(test_se), 
        .C(net12425), .Q(dph_reg[29]) );
  SDFFQX1 dph_reg_reg_3__3_ ( .D(N12524), .SIN(dph_reg[26]), .SMC(test_se), 
        .C(net12425), .Q(dph_reg[27]) );
  SDFFQX1 dph_reg_reg_3__1_ ( .D(N12522), .SIN(dph_reg[24]), .SMC(test_se), 
        .C(net12425), .Q(dph_reg[25]) );
  SDFFQX1 dpl_reg_reg_3__6_ ( .D(N12599), .SIN(dpl_reg[29]), .SMC(test_se), 
        .C(net12425), .Q(dpl_reg[30]) );
  SDFFQX1 dpl_reg_reg_3__5_ ( .D(N12598), .SIN(dpl_reg[28]), .SMC(test_se), 
        .C(net12425), .Q(dpl_reg[29]) );
  SDFFQX1 dpl_reg_reg_3__4_ ( .D(N12597), .SIN(dpl_reg[27]), .SMC(test_se), 
        .C(net12425), .Q(dpl_reg[28]) );
  SDFFQX1 dpl_reg_reg_3__2_ ( .D(N12595), .SIN(dpl_reg[25]), .SMC(test_se), 
        .C(net12425), .Q(dpl_reg[26]) );
  SDFFQX1 dpl_reg_reg_3__1_ ( .D(N12594), .SIN(dpl_reg[24]), .SMC(test_se), 
        .C(net12425), .Q(dpl_reg[25]) );
  SDFFQX1 dpl_reg_reg_3__0_ ( .D(N12593), .SIN(dpl_reg[23]), .SMC(test_se), 
        .C(net12425), .Q(dpl_reg[24]) );
  SDFFQX1 dph_reg_reg_7__6_ ( .D(N12563), .SIN(dph_reg[61]), .SMC(test_se), 
        .C(net12405), .Q(dph_reg[62]) );
  SDFFQX1 dph_reg_reg_7__5_ ( .D(N12562), .SIN(dph_reg[60]), .SMC(test_se), 
        .C(net12405), .Q(dph_reg[61]) );
  SDFFQX1 dph_reg_reg_7__4_ ( .D(N12561), .SIN(dph_reg[59]), .SMC(test_se), 
        .C(net12405), .Q(dph_reg[60]) );
  SDFFQX1 dph_reg_reg_7__3_ ( .D(N12560), .SIN(dph_reg[58]), .SMC(test_se), 
        .C(net12405), .Q(dph_reg[59]) );
  SDFFQX1 dph_reg_reg_7__1_ ( .D(N12558), .SIN(dph_reg[56]), .SMC(test_se), 
        .C(net12405), .Q(dph_reg[57]) );
  SDFFQX1 dpl_reg_reg_7__6_ ( .D(N12635), .SIN(dpl_reg[61]), .SMC(test_se), 
        .C(net12405), .Q(dpl_reg[62]) );
  SDFFQX1 dpl_reg_reg_7__5_ ( .D(N12634), .SIN(dpl_reg[60]), .SMC(test_se), 
        .C(net12405), .Q(dpl_reg[61]) );
  SDFFQX1 dpl_reg_reg_7__4_ ( .D(N12633), .SIN(dpl_reg[59]), .SMC(test_se), 
        .C(net12405), .Q(dpl_reg[60]) );
  SDFFQX1 dpl_reg_reg_7__1_ ( .D(N12630), .SIN(dpl_reg[56]), .SMC(test_se), 
        .C(net12405), .Q(dpl_reg[57]) );
  SDFFQX1 dph_reg_reg_7__0_ ( .D(N12557), .SIN(dph_reg[55]), .SMC(test_se), 
        .C(net12405), .Q(dph_reg[56]) );
  SDFFQX1 dph_reg_reg_3__0_ ( .D(N12521), .SIN(dph_reg[23]), .SMC(test_se), 
        .C(net12425), .Q(dph_reg[24]) );
  SDFFQX1 dpl_reg_reg_7__7_ ( .D(N12636), .SIN(dpl_reg[62]), .SMC(test_se), 
        .C(net12405), .Q(dpl_reg[63]) );
  SDFFQX1 dpl_reg_reg_7__0_ ( .D(N12629), .SIN(dpl_reg[55]), .SMC(test_se), 
        .C(net12405), .Q(dpl_reg[56]) );
  SDFFQX1 dph_reg_reg_1__2_ ( .D(N12505), .SIN(dph_reg[9]), .SMC(test_se), .C(
        net12435), .Q(dph_reg[10]) );
  SDFFQX1 dph_reg_reg_5__2_ ( .D(N12541), .SIN(dph_reg[41]), .SMC(test_se), 
        .C(net12415), .Q(dph_reg[42]) );
  SDFFQX1 dph_reg_reg_6__2_ ( .D(N12550), .SIN(dph_reg[49]), .SMC(test_se), 
        .C(net12410), .Q(dph_reg[50]) );
  SDFFQX1 dph_reg_reg_1__6_ ( .D(N12509), .SIN(dph_reg[13]), .SMC(test_se), 
        .C(net12435), .Q(dph_reg[14]) );
  SDFFQX1 dph_reg_reg_1__5_ ( .D(N12508), .SIN(dph_reg[12]), .SMC(test_se), 
        .C(net12435), .Q(dph_reg[13]) );
  SDFFQX1 dph_reg_reg_1__4_ ( .D(N12507), .SIN(dph_reg[11]), .SMC(test_se), 
        .C(net12435), .Q(dph_reg[12]) );
  SDFFQX1 dph_reg_reg_1__3_ ( .D(N12506), .SIN(dph_reg[10]), .SMC(test_se), 
        .C(net12435), .Q(dph_reg[11]) );
  SDFFQX1 dph_reg_reg_1__1_ ( .D(N12504), .SIN(dph_reg[8]), .SMC(test_se), .C(
        net12435), .Q(dph_reg[9]) );
  SDFFQX1 dpl_reg_reg_1__6_ ( .D(N12581), .SIN(dpl_reg[13]), .SMC(test_se), 
        .C(net12435), .Q(dpl_reg[14]) );
  SDFFQX1 dpl_reg_reg_1__5_ ( .D(N12580), .SIN(dpl_reg[12]), .SMC(test_se), 
        .C(net12435), .Q(dpl_reg[13]) );
  SDFFQX1 dpl_reg_reg_1__4_ ( .D(N12579), .SIN(dpl_reg[11]), .SMC(test_se), 
        .C(net12435), .Q(dpl_reg[12]) );
  SDFFQX1 dpl_reg_reg_1__1_ ( .D(N12576), .SIN(dpl_reg[8]), .SMC(test_se), .C(
        net12435), .Q(dpl_reg[9]) );
  SDFFQX1 dph_reg_reg_5__6_ ( .D(N12545), .SIN(dph_reg[45]), .SMC(test_se), 
        .C(net12415), .Q(dph_reg[46]) );
  SDFFQX1 dph_reg_reg_5__5_ ( .D(N12544), .SIN(dph_reg[44]), .SMC(test_se), 
        .C(net12415), .Q(dph_reg[45]) );
  SDFFQX1 dph_reg_reg_5__4_ ( .D(N12543), .SIN(dph_reg[43]), .SMC(test_se), 
        .C(net12415), .Q(dph_reg[44]) );
  SDFFQX1 dph_reg_reg_5__3_ ( .D(N12542), .SIN(dph_reg[42]), .SMC(test_se), 
        .C(net12415), .Q(dph_reg[43]) );
  SDFFQX1 dph_reg_reg_5__1_ ( .D(N12540), .SIN(dph_reg[40]), .SMC(test_se), 
        .C(net12415), .Q(dph_reg[41]) );
  SDFFQX1 dpl_reg_reg_5__6_ ( .D(N12617), .SIN(dpl_reg[45]), .SMC(test_se), 
        .C(net12415), .Q(dpl_reg[46]) );
  SDFFQX1 dpl_reg_reg_5__5_ ( .D(N12616), .SIN(dpl_reg[44]), .SMC(test_se), 
        .C(net12415), .Q(dpl_reg[45]) );
  SDFFQX1 dpl_reg_reg_5__4_ ( .D(N12615), .SIN(dpl_reg[43]), .SMC(test_se), 
        .C(net12415), .Q(dpl_reg[44]) );
  SDFFQX1 dpl_reg_reg_5__1_ ( .D(N12612), .SIN(dpl_reg[40]), .SMC(test_se), 
        .C(net12415), .Q(dpl_reg[41]) );
  SDFFQX1 dph_reg_reg_1__0_ ( .D(N12503), .SIN(dph_reg[7]), .SMC(test_se), .C(
        net12435), .Q(dph_reg[8]) );
  SDFFQX1 dph_reg_reg_2__7_ ( .D(N12519), .SIN(dph_reg[22]), .SMC(test_se), 
        .C(net12430), .Q(dph_reg[23]) );
  SDFFQX1 dph_reg_reg_2__3_ ( .D(N12515), .SIN(dph_reg[18]), .SMC(test_se), 
        .C(net12430), .Q(dph_reg[19]) );
  SDFFQX1 dph_reg_reg_2__1_ ( .D(N12513), .SIN(dph_reg[16]), .SMC(test_se), 
        .C(net12430), .Q(dph_reg[17]) );
  SDFFQX1 dpl_reg_reg_2__6_ ( .D(N12590), .SIN(dpl_reg[21]), .SMC(test_se), 
        .C(net12430), .Q(dpl_reg[22]) );
  SDFFQX1 dpl_reg_reg_2__5_ ( .D(N12589), .SIN(dpl_reg[20]), .SMC(test_se), 
        .C(net12430), .Q(dpl_reg[21]) );
  SDFFQX1 dpl_reg_reg_2__4_ ( .D(N12588), .SIN(dpl_reg[19]), .SMC(test_se), 
        .C(net12430), .Q(dpl_reg[20]) );
  SDFFQX1 dpl_reg_reg_2__2_ ( .D(N12586), .SIN(dpl_reg[17]), .SMC(test_se), 
        .C(net12430), .Q(dpl_reg[18]) );
  SDFFQX1 dpl_reg_reg_2__1_ ( .D(N12585), .SIN(dpl_reg[16]), .SMC(test_se), 
        .C(net12430), .Q(dpl_reg[17]) );
  SDFFQX1 dpl_reg_reg_2__0_ ( .D(N12584), .SIN(dpl_reg[15]), .SMC(test_se), 
        .C(net12430), .Q(dpl_reg[16]) );
  SDFFQX1 dph_reg_reg_6__6_ ( .D(N12554), .SIN(dph_reg[53]), .SMC(test_se), 
        .C(net12410), .Q(dph_reg[54]) );
  SDFFQX1 dph_reg_reg_6__5_ ( .D(N12553), .SIN(dph_reg[52]), .SMC(test_se), 
        .C(net12410), .Q(dph_reg[53]) );
  SDFFQX1 dph_reg_reg_6__3_ ( .D(N12551), .SIN(dph_reg[50]), .SMC(test_se), 
        .C(net12410), .Q(dph_reg[51]) );
  SDFFQX1 dph_reg_reg_6__1_ ( .D(N12549), .SIN(dph_reg[48]), .SMC(test_se), 
        .C(net12410), .Q(dph_reg[49]) );
  SDFFQX1 dpl_reg_reg_6__6_ ( .D(N12626), .SIN(dpl_reg[53]), .SMC(test_se), 
        .C(net12410), .Q(dpl_reg[54]) );
  SDFFQX1 dpl_reg_reg_6__5_ ( .D(N12625), .SIN(dpl_reg[52]), .SMC(test_se), 
        .C(net12410), .Q(dpl_reg[53]) );
  SDFFQX1 dpl_reg_reg_6__4_ ( .D(N12624), .SIN(dpl_reg[51]), .SMC(test_se), 
        .C(net12410), .Q(dpl_reg[52]) );
  SDFFQX1 dpl_reg_reg_6__2_ ( .D(N12622), .SIN(dpl_reg[49]), .SMC(test_se), 
        .C(net12410), .Q(dpl_reg[50]) );
  SDFFQX1 dpl_reg_reg_6__1_ ( .D(N12621), .SIN(dpl_reg[48]), .SMC(test_se), 
        .C(net12410), .Q(dpl_reg[49]) );
  SDFFQX1 dph_reg_reg_6__0_ ( .D(N12548), .SIN(dph_reg[47]), .SMC(test_se), 
        .C(net12410), .Q(dph_reg[48]) );
  SDFFQX1 dph_reg_reg_2__0_ ( .D(N12512), .SIN(dph_reg[15]), .SMC(test_se), 
        .C(net12430), .Q(dph_reg[16]) );
  SDFFQX1 dpl_reg_reg_1__7_ ( .D(N12582), .SIN(dpl_reg[14]), .SMC(test_se), 
        .C(net12435), .Q(dpl_reg[15]) );
  SDFFQX1 dpl_reg_reg_1__0_ ( .D(N12575), .SIN(dpl_reg[7]), .SMC(test_se), .C(
        net12435), .Q(dpl_reg[8]) );
  SDFFQX1 dpl_reg_reg_5__7_ ( .D(N12618), .SIN(dpl_reg[46]), .SMC(test_se), 
        .C(net12415), .Q(dpl_reg[47]) );
  SDFFQX1 dpl_reg_reg_5__0_ ( .D(N12611), .SIN(dpl_reg[39]), .SMC(test_se), 
        .C(net12415), .Q(dpl_reg[40]) );
  SDFFQX1 dph_reg_reg_6__7_ ( .D(N12555), .SIN(dph_reg[54]), .SMC(test_se), 
        .C(net12410), .Q(dph_reg[55]) );
  SDFFQX1 dpl_reg_reg_6__0_ ( .D(N12620), .SIN(dpl_reg[47]), .SMC(test_se), 
        .C(net12410), .Q(dpl_reg[48]) );
  SDFFQX1 dph_reg_reg_0__2_ ( .D(N12496), .SIN(dph_reg[1]), .SMC(test_se), .C(
        net12440), .Q(dph_reg[2]) );
  SDFFQX1 dph_reg_reg_4__2_ ( .D(N12532), .SIN(dph_reg[33]), .SMC(test_se), 
        .C(net12420), .Q(dph_reg[34]) );
  SDFFQX1 dph_reg_reg_0__6_ ( .D(N12500), .SIN(dph_reg[5]), .SMC(test_se), .C(
        net12440), .Q(dph_reg[6]) );
  SDFFQX1 dph_reg_reg_0__5_ ( .D(N12499), .SIN(dph_reg[4]), .SMC(test_se), .C(
        net12440), .Q(dph_reg[5]) );
  SDFFQX1 dph_reg_reg_0__4_ ( .D(N12498), .SIN(dph_reg[3]), .SMC(test_se), .C(
        net12440), .Q(dph_reg[4]) );
  SDFFQX1 dph_reg_reg_0__3_ ( .D(N12497), .SIN(dph_reg[2]), .SMC(test_se), .C(
        net12440), .Q(dph_reg[3]) );
  SDFFQX1 dph_reg_reg_0__1_ ( .D(N12495), .SIN(dph_reg[0]), .SMC(test_se), .C(
        net12440), .Q(dph_reg[1]) );
  SDFFQX1 dpl_reg_reg_0__6_ ( .D(N12572), .SIN(dpl_reg[5]), .SMC(test_se), .C(
        net12440), .Q(dpl_reg[6]) );
  SDFFQX1 dpl_reg_reg_0__5_ ( .D(N12571), .SIN(dpl_reg[4]), .SMC(test_se), .C(
        net12440), .Q(dpl_reg[5]) );
  SDFFQX1 dpl_reg_reg_0__4_ ( .D(N12570), .SIN(dpl_reg[3]), .SMC(test_se), .C(
        net12440), .Q(dpl_reg[4]) );
  SDFFQX1 dpl_reg_reg_0__1_ ( .D(N12567), .SIN(dpl_reg[0]), .SMC(test_se), .C(
        net12440), .Q(dpl_reg[1]) );
  SDFFQX1 dpl_reg_reg_0__0_ ( .D(N12566), .SIN(dph_reg[63]), .SMC(test_se), 
        .C(net12440), .Q(dpl_reg[0]) );
  SDFFQX1 dph_reg_reg_4__6_ ( .D(N12536), .SIN(dph_reg[37]), .SMC(test_se), 
        .C(net12420), .Q(dph_reg[38]) );
  SDFFQX1 dph_reg_reg_4__5_ ( .D(N12535), .SIN(dph_reg[36]), .SMC(test_se), 
        .C(net12420), .Q(dph_reg[37]) );
  SDFFQX1 dph_reg_reg_4__4_ ( .D(N12534), .SIN(dph_reg[35]), .SMC(test_se), 
        .C(net12420), .Q(dph_reg[36]) );
  SDFFQX1 dph_reg_reg_4__3_ ( .D(N12533), .SIN(dph_reg[34]), .SMC(test_se), 
        .C(net12420), .Q(dph_reg[35]) );
  SDFFQX1 dph_reg_reg_4__1_ ( .D(N12531), .SIN(dph_reg[32]), .SMC(test_se), 
        .C(net12420), .Q(dph_reg[33]) );
  SDFFQX1 dpl_reg_reg_4__6_ ( .D(N12608), .SIN(dpl_reg[37]), .SMC(test_se), 
        .C(net12420), .Q(dpl_reg[38]) );
  SDFFQX1 dpl_reg_reg_4__5_ ( .D(N12607), .SIN(dpl_reg[36]), .SMC(test_se), 
        .C(net12420), .Q(dpl_reg[37]) );
  SDFFQX1 dpl_reg_reg_4__4_ ( .D(N12606), .SIN(dpl_reg[35]), .SMC(test_se), 
        .C(net12420), .Q(dpl_reg[36]) );
  SDFFQX1 dpl_reg_reg_4__1_ ( .D(N12603), .SIN(dpl_reg[32]), .SMC(test_se), 
        .C(net12420), .Q(dpl_reg[33]) );
  SDFFQX1 dph_reg_reg_0__0_ ( .D(N12494), .SIN(dpc_tab[47]), .SMC(test_se), 
        .C(net12440), .Q(dph_reg[0]) );
  SDFFQX1 dpl_reg_reg_0__7_ ( .D(N12573), .SIN(dpl_reg[6]), .SMC(test_se), .C(
        net12440), .Q(dpl_reg[7]) );
  SDFFQX1 dpl_reg_reg_4__7_ ( .D(N12609), .SIN(dpl_reg[38]), .SMC(test_se), 
        .C(net12420), .Q(dpl_reg[39]) );
  SDFFQX1 dpl_reg_reg_4__0_ ( .D(N12602), .SIN(dpl_reg[31]), .SMC(test_se), 
        .C(net12420), .Q(dpl_reg[32]) );
  SDFFQX1 dec_cop_reg_4_ ( .D(N10586), .SIN(dec_cop[3]), .SMC(test_se), .C(
        net12389), .Q(dec_cop[4]) );
  SDFFQX1 dec_cop_reg_7_ ( .D(N10589), .SIN(dec_cop[6]), .SMC(test_se), .C(
        net12389), .Q(dec_cop[7]) );
  SDFFQX1 dec_cop_reg_3_ ( .D(N10585), .SIN(dec_cop[2]), .SMC(test_se), .C(
        net12389), .Q(dec_cop[3]) );
  SDFFQX1 dec_cop_reg_2_ ( .D(N10584), .SIN(dec_cop[1]), .SMC(test_se), .C(
        net12389), .Q(dec_cop[2]) );
  SDFFQX1 dec_cop_reg_1_ ( .D(N10583), .SIN(dec_cop[0]), .SMC(test_se), .C(
        net12389), .Q(dec_cop[1]) );
  SDFFQX1 ckcon_r_reg_7_ ( .D(N12972), .SIN(ckcon[6]), .SMC(test_se), .C(
        net12389), .Q(ckcon[7]) );
  SDFFQX1 ckcon_r_reg_3_ ( .D(N12968), .SIN(ckcon[2]), .SMC(test_se), .C(
        net12389), .Q(ckcon[3]) );
  SDFFQX1 dec_cop_reg_5_ ( .D(N10587), .SIN(dec_cop[4]), .SMC(test_se), .C(
        net12389), .Q(dec_cop[5]) );
  SDFFQX1 rmwinstr_reg ( .D(n2284), .SIN(ramwe), .SMC(test_se), .C(net12389), 
        .Q(rmwinstr) );
  SDFFQX1 dec_cop_reg_6_ ( .D(N10588), .SIN(dec_cop[5]), .SMC(test_se), .C(
        net12389), .Q(dec_cop[6]) );
  SDFFQX1 p2_reg_reg_2_ ( .D(N12487), .SIN(p2[1]), .SMC(test_se), .C(net12389), 
        .Q(p2[2]) );
  SDFFQX1 p2_reg_reg_1_ ( .D(N12486), .SIN(p2[0]), .SMC(test_se), .C(net12389), 
        .Q(p2[1]) );
  SDFFQX1 rn_reg_reg_7__3_ ( .D(n2221), .SIN(rn_reg[194]), .SMC(test_se), .C(
        net12530), .Q(rn_reg[195]) );
  SDFFQX1 rn_reg_reg_23__4_ ( .D(n276), .SIN(rn_reg[67]), .SMC(test_se), .C(
        net12610), .Q(rn_reg[68]) );
  SDFFQX1 rn_reg_reg_15__3_ ( .D(n279), .SIN(rn_reg[130]), .SMC(test_se), .C(
        net12570), .Q(rn_reg[131]) );
  SDFFQX1 rn_reg_reg_4__3_ ( .D(n279), .SIN(rn_reg[218]), .SMC(test_se), .C(
        net12515), .Q(rn_reg[219]) );
  SDFFQX1 rn_reg_reg_20__4_ ( .D(n276), .SIN(rn_reg[91]), .SMC(test_se), .C(
        net12595), .Q(rn_reg[92]) );
  SDFFQX1 rn_reg_reg_28__4_ ( .D(n275), .SIN(rn_reg[27]), .SMC(test_se), .C(
        net12635), .Q(rn_reg[28]) );
  SDFFQX1 rn_reg_reg_12__3_ ( .D(n278), .SIN(rn_reg[154]), .SMC(test_se), .C(
        net12555), .Q(rn_reg[155]) );
  SDFFQX1 rn_reg_reg_5__3_ ( .D(n278), .SIN(rn_reg[210]), .SMC(test_se), .C(
        net12520), .Q(rn_reg[211]) );
  SDFFQX1 rn_reg_reg_29__4_ ( .D(n275), .SIN(rn_reg[19]), .SMC(test_se), .C(
        net12640), .Q(rn_reg[20]) );
  SDFFQX1 rn_reg_reg_13__3_ ( .D(n277), .SIN(rn_reg[146]), .SMC(test_se), .C(
        net12560), .Q(rn_reg[147]) );
  SDFFQX1 rn_reg_reg_10__3_ ( .D(n277), .SIN(rn_reg[170]), .SMC(test_se), .C(
        net12545), .Q(rn_reg[171]) );
  SDFFQX1 rn_reg_reg_18__1_ ( .D(n253), .SIN(rn_reg[104]), .SMC(test_se), .C(
        net12585), .Q(rn_reg[105]) );
  SDFFQX1 rn_reg_reg_2__3_ ( .D(n277), .SIN(rn_reg[234]), .SMC(test_se), .C(
        net12505), .Q(rn_reg[235]) );
  SDFFQX1 rn_reg_reg_2__4_ ( .D(n274), .SIN(rn_reg[235]), .SMC(test_se), .C(
        net12505), .Q(rn_reg[236]) );
  SDFFQX1 rn_reg_reg_18__4_ ( .D(n274), .SIN(rn_reg[107]), .SMC(test_se), .C(
        net12585), .Q(rn_reg[108]) );
  SDFFQX1 rn_reg_reg_18__3_ ( .D(n277), .SIN(rn_reg[106]), .SMC(test_se), .C(
        net12585), .Q(rn_reg[107]) );
  SDFFQX1 rn_reg_reg_6__3_ ( .D(n277), .SIN(rn_reg[202]), .SMC(test_se), .C(
        net12525), .Q(rn_reg[203]) );
  SDFFQX1 rn_reg_reg_6__4_ ( .D(n274), .SIN(rn_reg[203]), .SMC(test_se), .C(
        net12525), .Q(rn_reg[204]) );
  SDFFQX1 rn_reg_reg_22__4_ ( .D(n274), .SIN(rn_reg[75]), .SMC(test_se), .C(
        net12605), .Q(rn_reg[76]) );
  SDFFQX1 rn_reg_reg_22__3_ ( .D(n277), .SIN(rn_reg[74]), .SMC(test_se), .C(
        net12605), .Q(rn_reg[75]) );
  SDFFQX1 rn_reg_reg_30__3_ ( .D(n277), .SIN(rn_reg[10]), .SMC(test_se), .C(
        net12645), .Q(rn_reg[11]) );
  SDFFQX1 rn_reg_reg_14__3_ ( .D(n277), .SIN(rn_reg[138]), .SMC(test_se), .C(
        net12565), .Q(rn_reg[139]) );
  SDFFQX1 dph_reg_reg_3__6_ ( .D(N12527), .SIN(dph_reg[29]), .SMC(test_se), 
        .C(net12425), .Q(dph_reg[30]) );
  SDFFQX1 dph_reg_reg_3__4_ ( .D(N12525), .SIN(dph_reg[27]), .SMC(test_se), 
        .C(net12425), .Q(dph_reg[28]) );
  SDFFQX1 dpl_reg_reg_3__7_ ( .D(N12600), .SIN(dpl_reg[30]), .SMC(test_se), 
        .C(net12425), .Q(dpl_reg[31]) );
  SDFFQX1 dph_reg_reg_2__2_ ( .D(N12514), .SIN(dph_reg[17]), .SMC(test_se), 
        .C(net12430), .Q(dph_reg[18]) );
  SDFFQX1 dph_reg_reg_2__6_ ( .D(N12518), .SIN(dph_reg[21]), .SMC(test_se), 
        .C(net12430), .Q(dph_reg[22]) );
  SDFFQX1 dph_reg_reg_2__5_ ( .D(N12517), .SIN(dph_reg[20]), .SMC(test_se), 
        .C(net12430), .Q(dph_reg[21]) );
  SDFFQX1 dph_reg_reg_2__4_ ( .D(N12516), .SIN(dph_reg[19]), .SMC(test_se), 
        .C(net12430), .Q(dph_reg[20]) );
  SDFFQX1 dph_reg_reg_6__4_ ( .D(N12552), .SIN(dph_reg[51]), .SMC(test_se), 
        .C(net12410), .Q(dph_reg[52]) );
  SDFFQX1 dpl_reg_reg_2__7_ ( .D(N12591), .SIN(dpl_reg[22]), .SMC(test_se), 
        .C(net12430), .Q(dpl_reg[23]) );
  SDFFQX1 dpl_reg_reg_6__7_ ( .D(N12627), .SIN(dpl_reg[54]), .SMC(test_se), 
        .C(net12410), .Q(dpl_reg[55]) );
  SDFFQX1 sp_reg_reg_4_ ( .D(N12701), .SIN(sp[3]), .SMC(test_se), .C(net12389), 
        .Q(sp[4]) );
  SDFFQX1 sp_reg_reg_3_ ( .D(N12700), .SIN(sp[2]), .SMC(test_se), .C(net12389), 
        .Q(sp[3]) );
  SDFFQX1 sp_reg_reg_5_ ( .D(N12702), .SIN(sp[4]), .SMC(test_se), .C(net12389), 
        .Q(sp[5]) );
  SDFFQX1 sp_reg_reg_6_ ( .D(N12703), .SIN(sp[5]), .SMC(test_se), .C(net12389), 
        .Q(sp[6]) );
  SDFFQX1 multempreg_reg_1_ ( .D(N13326), .SIN(multempreg[0]), .SMC(test_se), 
        .C(net12655), .Q(multempreg[1]) );
  SDFFQX1 ramwe_r_reg ( .D(N11487), .SIN(ramsfrwe), .SMC(test_se), .C(net12389), .Q(ramwe) );
  SDFFQX1 pmw_reg_reg ( .D(n2204), .SIN(phase[5]), .SMC(test_se), .C(net12389), 
        .Q(pmw) );
  SDFFQX1 temp2_reg_7_ ( .D(N12730), .SIN(temp2_comb[6]), .SMC(test_se), .C(
        net12389), .Q(temp2_comb[7]) );
  SDFFQX1 bitno_reg_2_ ( .D(n2224), .SIN(N344), .SMC(test_se), .C(net12400), 
        .Q(N345) );
  SDFFQX1 phase_reg_2_ ( .D(N681), .SIN(n263), .SMC(test_se), .C(net12389), 
        .Q(phase[2]) );
  SDFFQX1 ramdatao_r_reg_5_ ( .D(N11503), .SIN(ramdatao[4]), .SMC(test_se), 
        .C(net12389), .Q(ramdatao[5]) );
  SDFFQX1 ramdatao_r_reg_6_ ( .D(N11504), .SIN(ramdatao[5]), .SMC(test_se), 
        .C(net12389), .Q(ramdatao[6]) );
  SDFFQX1 ramdatao_r_reg_7_ ( .D(N11505), .SIN(ramdatao[6]), .SMC(test_se), 
        .C(net12389), .Q(ramdatao[7]) );
  SDFFQX1 sp_reg_reg_2_ ( .D(N12699), .SIN(sp[1]), .SMC(test_se), .C(net12389), 
        .Q(sp[2]) );
  SDFFQX1 sp_reg_reg_1_ ( .D(N12698), .SIN(sp[0]), .SMC(test_se), .C(net12389), 
        .Q(sp[1]) );
  SDFFQX1 sp_reg_reg_0_ ( .D(N12697), .SIN(sfrwe_r), .SMC(test_se), .C(
        net12389), .Q(sp[0]) );
  SDFFQX1 dec_accop_reg_11_ ( .D(N10574), .SIN(dec_accop[10]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[11]) );
  SDFFQX1 multempreg_reg_0_ ( .D(N13325), .SIN(memwr), .SMC(test_se), .C(
        net12655), .Q(multempreg[0]) );
  SDFFQX1 dec_accop_reg_17_ ( .D(n2150), .SIN(dec_accop[16]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[17]) );
  SDFFQX1 sfroe_r_reg ( .D(N11488), .SIN(rs[1]), .SMC(test_se), .C(net12389), 
        .Q(sfroe_r) );
  SDFFQX1 sfrwe_r_reg ( .D(N11489), .SIN(sfroe_r), .SMC(test_se), .C(net12389), 
        .Q(sfrwe_r) );
  SDFFQX1 dps_reg_reg_3_ ( .D(n1884), .SIN(dps[2]), .SMC(test_se), .C(net12389), .Q(dps[3]) );
  SDFFQX1 bitno_reg_1_ ( .D(n2225), .SIN(N343), .SMC(test_se), .C(net12400), 
        .Q(N344) );
  SDFFQX1 temp_reg_0_ ( .D(N12714), .SIN(temp2_comb[7]), .SMC(test_se), .C(
        net12485), .Q(temp[0]) );
  SDFFQX1 temp_reg_1_ ( .D(N12715), .SIN(temp[0]), .SMC(test_se), .C(net12485), 
        .Q(temp[1]) );
  SDFFQX1 temp_reg_5_ ( .D(N12719), .SIN(temp[4]), .SMC(test_se), .C(net12485), 
        .Q(temp[5]) );
  SDFFQX1 temp_reg_6_ ( .D(N12720), .SIN(temp[5]), .SMC(test_se), .C(net12485), 
        .Q(temp[6]) );
  SDFFQX1 temp_reg_2_ ( .D(N12716), .SIN(temp[1]), .SMC(test_se), .C(net12485), 
        .Q(temp[2]) );
  SDFFQX1 dps_reg_reg_0_ ( .D(N12693), .SIN(dpl_reg[63]), .SMC(test_se), .C(
        net12389), .Q(dps[0]) );
  SDFFQX1 dps_reg_reg_1_ ( .D(N12694), .SIN(dps[0]), .SMC(test_se), .C(
        net12389), .Q(dps[1]) );
  SDFFQX1 temp_reg_7_ ( .D(N12721), .SIN(temp[6]), .SMC(test_se), .C(net12485), 
        .Q(temp[7]) );
  SDFFQX1 bitno_reg_0_ ( .D(n2257), .SIN(b[7]), .SMC(test_se), .C(net12400), 
        .Q(N343) );
  SDFFQX1 temp2_reg_6_ ( .D(N12729), .SIN(temp2_comb[5]), .SMC(test_se), .C(
        net12389), .Q(temp2_comb[6]) );
  SDFFQX1 interrupt_reg ( .D(n2275), .SIN(instr[7]), .SMC(test_se), .C(
        net12395), .Q(interrupt) );
  SDFFQX1 ramdatao_r_reg_2_ ( .D(N11500), .SIN(ramdatao[1]), .SMC(test_se), 
        .C(net12389), .Q(ramdatao[2]) );
  SDFFQX1 ramdatao_r_reg_1_ ( .D(N11499), .SIN(ramdatao[0]), .SMC(test_se), 
        .C(net12389), .Q(ramdatao[1]) );
  SDFFQX1 ramdatao_r_reg_0_ ( .D(N11498), .SIN(pmw), .SMC(test_se), .C(
        net12389), .Q(ramdatao[0]) );
  SDFFQX1 dps_reg_reg_2_ ( .D(N12695), .SIN(dps[1]), .SMC(test_se), .C(
        net12389), .Q(n2510) );
  SDFFQX1 dec_accop_reg_14_ ( .D(N10577), .SIN(dec_accop[13]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[14]) );
  SDFFQX1 dec_accop_reg_2_ ( .D(N10565), .SIN(dec_accop[1]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[2]) );
  SDFFQX1 dec_accop_reg_15_ ( .D(N10578), .SIN(dec_accop[14]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[15]) );
  SDFFQX1 dec_accop_reg_13_ ( .D(N10576), .SIN(dec_accop[12]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[13]) );
  SDFFQX1 dec_accop_reg_12_ ( .D(N10575), .SIN(dec_accop[11]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[12]) );
  SDFFQX1 rs_reg_reg_1_ ( .D(N12710), .SIN(rs[0]), .SMC(test_se), .C(net12389), 
        .Q(rs[1]) );
  SDFFQX1 memrd_s_reg ( .D(N584), .SIN(n2499), .SMC(test_se), .C(net12389), 
        .Q(memrd) );
  SDFFQX1 memwr_s_reg ( .D(N585), .SIN(memrd), .SMC(test_se), .C(net12389), 
        .Q(memwr) );
  SDFFQX1 mempsrd_r_reg ( .D(N582), .SIN(israccess), .SMC(test_se), .C(
        net12389), .Q(mempsrd) );
  SDFFQX1 rs_reg_reg_0_ ( .D(N12709), .SIN(rn_reg[7]), .SMC(test_se), .C(
        net12389), .Q(rs[0]) );
  SDFFQX1 temp2_reg_5_ ( .D(N12728), .SIN(temp2_comb[4]), .SMC(test_se), .C(
        net12389), .Q(temp2_comb[5]) );
  SDFFQX1 temp2_reg_4_ ( .D(N12727), .SIN(temp2_comb[3]), .SMC(test_se), .C(
        net12389), .Q(temp2_comb[4]) );
  SDFFQX1 ramdatao_r_reg_4_ ( .D(N11502), .SIN(ramdatao[3]), .SMC(test_se), 
        .C(net12389), .Q(ramdatao[4]) );
  SDFFQX1 ramdatao_r_reg_3_ ( .D(N11501), .SIN(ramdatao[2]), .SMC(test_se), 
        .C(net12389), .Q(n2501) );
  SDFFQX1 mempswr_s_reg ( .D(N583), .SIN(mempsrd), .SMC(test_se), .C(net12389), 
        .Q(n2499) );
  SDFFQX1 phase_reg_0_ ( .D(N679), .SIN(phase0_ff), .SMC(test_se), .C(net12389), .Q(phase[0]) );
  SDFFQX1 dec_accop_reg_0_ ( .D(N10563), .SIN(d_hold), .SMC(test_se), .C(
        net12389), .Q(dec_accop[0]) );
  SDFFQX1 dec_accop_reg_3_ ( .D(N10566), .SIN(dec_accop[2]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[3]) );
  SDFFQX1 ckcon_r_reg_0_ ( .D(N12965), .SIN(n151), .SMC(test_se), .C(net12389), 
        .Q(ckcon[0]) );
  SDFFQX1 dec_accop_reg_4_ ( .D(N10567), .SIN(dec_accop[3]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[4]) );
  SDFFQX1 ckcon_r_reg_4_ ( .D(N12969), .SIN(ckcon[3]), .SMC(test_se), .C(
        net12389), .Q(ckcon[4]) );
  SDFFQX1 dec_accop_reg_1_ ( .D(N10564), .SIN(dec_accop[0]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[1]) );
  SDFFQX1 ckcon_r_reg_1_ ( .D(N12966), .SIN(ckcon[0]), .SMC(test_se), .C(
        net12389), .Q(ckcon[1]) );
  SDFFQX1 ckcon_r_reg_5_ ( .D(N12970), .SIN(ckcon[4]), .SMC(test_se), .C(
        net12389), .Q(ckcon[5]) );
  SDFFQX1 temp2_reg_3_ ( .D(N12726), .SIN(temp2_comb[2]), .SMC(test_se), .C(
        net12389), .Q(temp2_comb[3]) );
  SDFFQX1 waitcnt_reg_2_ ( .D(N12976), .SIN(waitcnt_1_), .SMC(test_se), .C(
        net12490), .Q(test_so) );
  SDFFQX1 ckcon_r_reg_2_ ( .D(N12967), .SIN(ckcon[1]), .SMC(test_se), .C(
        net12389), .Q(ckcon[2]) );
  SDFFQX1 waitcnt_reg_1_ ( .D(N12975), .SIN(waitcnt_0_), .SMC(test_se), .C(
        net12490), .Q(waitcnt_1_) );
  SDFFQX1 waitcnt_reg_0_ ( .D(N12974), .SIN(temp[7]), .SMC(test_se), .C(
        net12490), .Q(waitcnt_0_) );
  SDFFQX1 ckcon_r_reg_6_ ( .D(N12971), .SIN(ckcon[5]), .SMC(test_se), .C(
        net12389), .Q(ckcon[6]) );
  SDFFQX1 acc_reg_reg_5_ ( .D(n2213), .SIN(acc[4]), .SMC(test_se), .C(net12389), .Q(acc[5]) );
  SDFFQX1 acc_reg_reg_4_ ( .D(n2217), .SIN(acc[3]), .SMC(test_se), .C(net12389), .Q(acc[4]) );
  SDFFQX1 accactv_reg ( .D(N10562), .SIN(acc[7]), .SMC(test_se), .C(net12389), 
        .Q(accactv) );
  SDFFQX1 instr_reg_4_ ( .D(N674), .SIN(instr[3]), .SMC(test_se), .C(net12395), 
        .Q(n2506) );
  SDFFQX1 acc_reg_reg_6_ ( .D(n2209), .SIN(acc[5]), .SMC(test_se), .C(net12389), .Q(acc[6]) );
  SDFFQX1 ramsfrwe_reg ( .D(n2254), .SIN(ramsfraddr[7]), .SMC(test_se), .C(
        net12389), .Q(ramsfrwe) );
  SDFFQX1 temp2_reg_2_ ( .D(N12725), .SIN(temp2_comb[1]), .SMC(test_se), .C(
        net12389), .Q(temp2_comb[2]) );
  SDFFQX1 ramsfraddr_s_reg_1_ ( .D(N11479), .SIN(ramsfraddr[0]), .SMC(test_se), 
        .C(net12389), .Q(ramsfraddr[1]) );
  SDFFQX1 ramsfraddr_s_reg_5_ ( .D(N11483), .SIN(ramsfraddr[4]), .SMC(test_se), 
        .C(net12389), .Q(ramsfraddr[5]) );
  SDFFQX1 ramsfraddr_s_reg_4_ ( .D(N11482), .SIN(ramsfraddr[3]), .SMC(test_se), 
        .C(net12389), .Q(ramsfraddr[4]) );
  SDFFQX1 ramsfraddr_s_reg_0_ ( .D(N11478), .SIN(ramoe), .SMC(test_se), .C(
        net12389), .Q(ramsfraddr[0]) );
  SDFFQX1 ramsfraddr_s_reg_6_ ( .D(N11484), .SIN(ramsfraddr[5]), .SMC(test_se), 
        .C(net12389), .Q(ramsfraddr[6]) );
  SDFFQX1 ramsfraddr_s_reg_2_ ( .D(N11480), .SIN(ramsfraddr[1]), .SMC(test_se), 
        .C(net12389), .Q(ramsfraddr[2]) );
  SDFFQX1 ramsfraddr_s_reg_3_ ( .D(N11481), .SIN(ramsfraddr[2]), .SMC(test_se), 
        .C(net12389), .Q(ramsfraddr[3]) );
  SDFFQX1 phase_reg_1_ ( .D(N680), .SIN(n106), .SMC(test_se), .C(net12389), 
        .Q(phase[1]) );
  SDFFQX1 divtempreg_reg_6_ ( .D(N13373), .SIN(divtempreg[5]), .SMC(test_se), 
        .C(net12660), .Q(divtempreg[6]) );
  SDFFQX1 temp2_reg_1_ ( .D(N12724), .SIN(temp2_comb[0]), .SMC(test_se), .C(
        net12389), .Q(temp2_comb[1]) );
  SDFFQX1 ramsfraddr_s_reg_7_ ( .D(N11485), .SIN(ramsfraddr[6]), .SMC(test_se), 
        .C(net12389), .Q(ramsfraddr[7]) );
  SDFFQX1 instr_reg_2_ ( .D(N672), .SIN(n2508), .SMC(test_se), .C(net12395), 
        .Q(instr[2]) );
  SDFFQX1 instr_reg_6_ ( .D(N676), .SIN(instr[5]), .SMC(test_se), .C(net12395), 
        .Q(instr[6]) );
  SDFFQX1 b_reg_reg_7_ ( .D(N12484), .SIN(b[6]), .SMC(test_se), .C(net12389), 
        .Q(b[7]) );
  SDFFQX1 instr_reg_0_ ( .D(N670), .SIN(idle), .SMC(test_se), .C(net12395), 
        .Q(n2509) );
  SDFFQX1 instr_reg_1_ ( .D(N671), .SIN(instr[0]), .SMC(test_se), .C(net12395), 
        .Q(n2508) );
  SDFFQX1 instr_reg_5_ ( .D(N675), .SIN(instr[4]), .SMC(test_se), .C(net12395), 
        .Q(n2505) );
  SDFFQX1 instr_reg_7_ ( .D(N677), .SIN(instr[6]), .SMC(test_se), .C(net12395), 
        .Q(n2504) );
  SDFFQX1 instr_reg_3_ ( .D(N673), .SIN(instr[2]), .SMC(test_se), .C(net12395), 
        .Q(n2507) );
  SDFFQX1 ac_reg_reg ( .D(N12706), .SIN(test_si), .SMC(test_se), .C(net12389), 
        .Q(ac) );
  SDFFQX1 pc_reg_1_ ( .D(N481), .SIN(pc_o[0]), .SMC(test_se), .C(net12389), 
        .Q(memaddr[1]) );
  SDFFQX1 pc_reg_10_ ( .D(N490), .SIN(memaddr[9]), .SMC(test_se), .C(net12389), 
        .Q(memaddr[10]) );
  SDFFQX1 divtempreg_reg_5_ ( .D(N13372), .SIN(divtempreg[4]), .SMC(test_se), 
        .C(net12660), .Q(divtempreg[5]) );
  SDFFQX1 divtempreg_reg_4_ ( .D(N13371), .SIN(divtempreg[3]), .SMC(test_se), 
        .C(net12660), .Q(divtempreg[4]) );
  SDFFQX1 dec_accop_reg_7_ ( .D(N10570), .SIN(dec_accop[6]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[7]) );
  SDFFQX1 dec_accop_reg_18_ ( .D(N10581), .SIN(dec_accop[17]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[18]) );
  SDFFQX1 dec_accop_reg_16_ ( .D(n2175), .SIN(dec_accop[15]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[16]) );
  SDFFQX1 dec_accop_reg_5_ ( .D(N10568), .SIN(dec_accop[4]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[5]) );
  SDFFQX1 dec_accop_reg_6_ ( .D(N10569), .SIN(dec_accop[5]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[6]) );
  SDFFQX1 temp2_reg_0_ ( .D(N12723), .SIN(stop), .SMC(test_se), .C(net12389), 
        .Q(temp2_comb[0]) );
  SDFFQX1 acc_reg_reg_2_ ( .D(n2193), .SIN(acc[1]), .SMC(test_se), .C(net12389), .Q(acc[2]) );
  SDFFQX1 acc_reg_reg_1_ ( .D(N12470), .SIN(acc[0]), .SMC(test_se), .C(
        net12389), .Q(acc[1]) );
  SDFFQX1 acc_reg_reg_0_ ( .D(N12469), .SIN(ac), .SMC(test_se), .C(net12389), 
        .Q(acc[0]) );
  SDFFQX1 acc_reg_reg_3_ ( .D(N12472), .SIN(acc[2]), .SMC(test_se), .C(
        net12389), .Q(acc[3]) );
  SDFFQX1 c_reg_reg ( .D(N12705), .SIN(N345), .SMC(test_se), .C(net12389), .Q(
        c) );
  SDFFQX1 b_reg_reg_6_ ( .D(N12483), .SIN(b[5]), .SMC(test_se), .C(net12389), 
        .Q(b[6]) );
  SDFFQX1 dec_accop_reg_8_ ( .D(N10571), .SIN(dec_accop[7]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[8]) );
  SDFFQX1 divtempreg_reg_3_ ( .D(N13370), .SIN(divtempreg[2]), .SMC(test_se), 
        .C(net12660), .Q(divtempreg[3]) );
  SDFFQX1 dec_accop_reg_9_ ( .D(N10572), .SIN(dec_accop[8]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[9]) );
  SDFFQX1 dec_accop_reg_10_ ( .D(N10573), .SIN(dec_accop[9]), .SMC(test_se), 
        .C(net12389), .Q(dec_accop[10]) );
  SDFFQX1 b_reg_reg_5_ ( .D(N12482), .SIN(b[4]), .SMC(test_se), .C(net12389), 
        .Q(b[5]) );
  SDFFQX1 b_reg_reg_4_ ( .D(N12481), .SIN(b[3]), .SMC(test_se), .C(net12389), 
        .Q(b[4]) );
  SDFFQX1 divtempreg_reg_2_ ( .D(N13369), .SIN(divtempreg[1]), .SMC(test_se), 
        .C(net12660), .Q(divtempreg[2]) );
  SDFFQX1 divtempreg_reg_1_ ( .D(N13368), .SIN(divtempreg[0]), .SMC(test_se), 
        .C(net12660), .Q(divtempreg[1]) );
  SDFFQX1 b_reg_reg_3_ ( .D(N12480), .SIN(b[2]), .SMC(test_se), .C(net12389), 
        .Q(b[3]) );
  SDFFQX1 divtempreg_reg_0_ ( .D(N13367), .SIN(dec_cop[7]), .SMC(test_se), .C(
        net12660), .Q(divtempreg[0]) );
  SDFFQX1 b_reg_reg_1_ ( .D(N12478), .SIN(b[0]), .SMC(test_se), .C(net12389), 
        .Q(b[1]) );
  SDFFQX1 b_reg_reg_2_ ( .D(N12479), .SIN(b[1]), .SMC(test_se), .C(net12389), 
        .Q(b[2]) );
  SDFFQX1 acc_reg_reg_7_ ( .D(n2196), .SIN(acc[6]), .SMC(test_se), .C(net12389), .Q(acc[7]) );
  SDFFQX1 b_reg_reg_0_ ( .D(N12477), .SIN(n123), .SMC(test_se), .C(net12389), 
        .Q(b[0]) );
  MUX4X1 U2264 ( .D0(temp[0]), .D1(temp[1]), .D2(temp[2]), .D3(temp[3]), .S0(
        N343), .S1(N344), .Y(n2032) );
  MUX4X1 U2263 ( .D0(temp[4]), .D1(temp[5]), .D2(temp[6]), .D3(temp[7]), .S0(
        N343), .S1(N344), .Y(n2031) );
  SDFFQX1 pc_reg_4_ ( .D(N484), .SIN(pc_o[3]), .SMC(test_se), .C(net12389), 
        .Q(n2502) );
  SDFFQX1 pc_reg_0_ ( .D(N480), .SIN(p), .SMC(test_se), .C(net12389), .Q(
        memaddr[0]) );
  SDFFQX1 pc_reg_3_ ( .D(N483), .SIN(n2503), .SMC(test_se), .C(net12389), .Q(
        memaddr[3]) );
  MUX2X1 U9 ( .D0(n2503), .D1(n1715), .S(n14), .Y(memaddr_comb[2]) );
  INVX1 U10 ( .A(n2), .Y(n14) );
  INVX4 U11 ( .A(n434), .Y(n1656) );
  MUX2X1 U12 ( .D0(pc_o[1]), .D1(n1714), .S(n15), .Y(memaddr_comb[1]) );
  BUFX1 U13 ( .A(n1443), .Y(n1) );
  INVX3 U14 ( .A(sfrdatai[4]), .Y(n674) );
  OR3X4 U15 ( .A(n174), .B(n175), .C(n176), .Y(n656) );
  NOR2X2 U16 ( .A(n674), .B(n354), .Y(n174) );
  OAI22X1 U17 ( .A(n1504), .B(n354), .C(n353), .D(n904), .Y(n1988) );
  OA222X1 U18 ( .A(n2495), .B(n1934), .C(n787), .D(n1932), .E(n951), .F(n1931), 
        .Y(n184) );
  INVX2 U19 ( .A(n361), .Y(n1858) );
  MUX2IX1 U20 ( .D0(idle), .D1(n1656), .S(n1405), .Y(n454) );
  NOR3XL U21 ( .A(n2366), .B(n2364), .C(n1333), .Y(n1147) );
  NAND21X1 U22 ( .B(n358), .A(n357), .Y(n359) );
  MUX2IX1 U23 ( .D0(n356), .D1(n355), .S(N345), .Y(n357) );
  OR3X1 U24 ( .A(n177), .B(n178), .C(n179), .Y(n695) );
  NOR3XL U25 ( .A(n1332), .B(n2366), .C(n1333), .Y(n1145) );
  NAND21X1 U26 ( .B(n1859), .A(n382), .Y(n416) );
  OA2222XL U27 ( .A(n1531), .B(n487), .C(n1532), .D(n2330), .E(n486), .F(n1859), .G(n1886), .H(n485), .Y(n489) );
  INVX2 U28 ( .A(sfrdatai[7]), .Y(n1504) );
  INVX1 U29 ( .A(sfrdatai[6]), .Y(n975) );
  INVX1 U30 ( .A(sfrdatai[1]), .Y(n775) );
  MUX2IX1 U31 ( .D0(stop), .D1(n1657), .S(n1405), .Y(n496) );
  INVX1 U32 ( .A(sfrdatai[3]), .Y(n639) );
  MUX2X1 U33 ( .D0(n50), .D1(n1718), .S(n15), .Y(memaddr_comb[5]) );
  INVX1 U34 ( .A(n2), .Y(n15) );
  NAND42X1 U35 ( .C(n302), .D(n1637), .A(n301), .B(n300), .Y(n1658) );
  OR2X1 U36 ( .A(n1712), .B(n286), .Y(n2) );
  OA22X1 U37 ( .A(n1435), .B(n180), .C(n1461), .D(n1), .Y(n3) );
  OR3XL U38 ( .A(n2306), .B(dpc[1]), .C(n1170), .Y(n10) );
  AND3X1 U39 ( .A(n599), .B(n600), .C(n601), .Y(n11) );
  INVXL U40 ( .A(n2501), .Y(n12) );
  INVXL U41 ( .A(n12), .Y(ramdatao[3]) );
  INVXL U42 ( .A(n1324), .Y(n16) );
  INVXL U43 ( .A(n16), .Y(n17) );
  INVXL U44 ( .A(n234), .Y(n18) );
  INVXL U45 ( .A(n18), .Y(n19) );
  INVXL U46 ( .A(n233), .Y(n20) );
  INVXL U47 ( .A(n20), .Y(n21) );
  INVXL U48 ( .A(n20), .Y(n22) );
  INVXL U49 ( .A(n231), .Y(n23) );
  INVXL U50 ( .A(n23), .Y(n24) );
  INVXL U51 ( .A(n232), .Y(n25) );
  INVXL U52 ( .A(n25), .Y(n26) );
  INVXL U53 ( .A(n25), .Y(n27) );
  INVXL U54 ( .A(n618), .Y(n28) );
  INVXL U55 ( .A(n618), .Y(n29) );
  INVXL U56 ( .A(n617), .Y(n30) );
  INVXL U57 ( .A(n617), .Y(n31) );
  INVXL U58 ( .A(instr[2]), .Y(n32) );
  INVXL U59 ( .A(instr[2]), .Y(n33) );
  INVXL U60 ( .A(pc_o[15]), .Y(n34) );
  INVXL U61 ( .A(n34), .Y(memaddr[15]) );
  INVXL U62 ( .A(n1132), .Y(n36) );
  INVXL U63 ( .A(n36), .Y(n37) );
  INVXL U64 ( .A(n788), .Y(n38) );
  INVXL U65 ( .A(n38), .Y(n39) );
  INVXL U66 ( .A(memaddr[12]), .Y(n40) );
  INVXL U67 ( .A(n40), .Y(pc_o[12]) );
  INVXL U68 ( .A(n10), .Y(n42) );
  INVXL U69 ( .A(n10), .Y(n43) );
  INVXL U70 ( .A(n2508), .Y(n44) );
  INVXL U71 ( .A(n44), .Y(instr[1]) );
  INVXL U72 ( .A(pc_o[13]), .Y(n46) );
  INVXL U73 ( .A(n46), .Y(memaddr[13]) );
  INVXL U74 ( .A(n37), .Y(n48) );
  INVXL U75 ( .A(memaddr[5]), .Y(n49) );
  INVXL U76 ( .A(n49), .Y(n50) );
  INVXL U77 ( .A(pc_o[9]), .Y(n51) );
  INVXL U78 ( .A(n51), .Y(memaddr[9]) );
  INVXL U79 ( .A(pc_o[8]), .Y(n53) );
  INVXL U80 ( .A(n53), .Y(memaddr[8]) );
  INVXL U81 ( .A(n2502), .Y(n55) );
  INVXL U82 ( .A(n55), .Y(memaddr[4]) );
  INVXL U83 ( .A(pc_o[6]), .Y(n57) );
  INVXL U84 ( .A(n57), .Y(memaddr[6]) );
  INVXL U85 ( .A(n2503), .Y(n59) );
  INVXL U86 ( .A(n59), .Y(memaddr[2]) );
  INVX2 U87 ( .A(n930), .Y(n1712) );
  NAND31X4 U88 ( .C(n417), .A(n416), .B(n415), .Y(n433) );
  INVX1 U89 ( .A(instr[3]), .Y(n61) );
  INVX1 U90 ( .A(instr[0]), .Y(n62) );
  BUFX3 U91 ( .A(n1118), .Y(n63) );
  BUFX3 U92 ( .A(n2448), .Y(n64) );
  BUFX3 U93 ( .A(n2509), .Y(instr[0]) );
  NAND2X1 U94 ( .A(n2011), .B(n2013), .Y(n1798) );
  INVX1 U95 ( .A(n1798), .Y(n66) );
  INVX1 U96 ( .A(n1798), .Y(n67) );
  BUFX3 U97 ( .A(n1105), .Y(n68) );
  BUFX3 U98 ( .A(n2262), .Y(n69) );
  BUFX3 U99 ( .A(n1124), .Y(n70) );
  NAND2X1 U100 ( .A(n2026), .B(n2012), .Y(n1808) );
  INVX1 U101 ( .A(n1808), .Y(n71) );
  INVX1 U102 ( .A(n1808), .Y(n72) );
  NAND2X1 U103 ( .A(n2008), .B(n2013), .Y(n1794) );
  INVX1 U104 ( .A(n1794), .Y(n73) );
  INVX1 U105 ( .A(n1794), .Y(n74) );
  BUFX3 U106 ( .A(n1407), .Y(n75) );
  INVX1 U107 ( .A(n1614), .Y(n76) );
  INVX1 U108 ( .A(n2415), .Y(n77) );
  INVX1 U109 ( .A(n152), .Y(dps[2]) );
  BUFX3 U110 ( .A(n2507), .Y(instr[3]) );
  INVX1 U111 ( .A(n109), .Y(instr[7]) );
  AOI21X1 U112 ( .B(n124), .C(n221), .A(n248), .Y(n1117) );
  INVX1 U113 ( .A(n1117), .Y(n81) );
  INVX1 U114 ( .A(n1117), .Y(n82) );
  AOI21X1 U115 ( .B(n104), .C(n220), .A(n246), .Y(n1123) );
  INVX1 U116 ( .A(n1123), .Y(n83) );
  INVX1 U117 ( .A(n1123), .Y(n84) );
  BUFX3 U118 ( .A(n1116), .Y(n85) );
  INVX1 U119 ( .A(n2304), .Y(n86) );
  NAND2X1 U120 ( .A(n2011), .B(n2012), .Y(n1795) );
  INVX1 U121 ( .A(n1795), .Y(n87) );
  INVX1 U122 ( .A(n1795), .Y(n88) );
  INVX1 U123 ( .A(n596), .Y(n89) );
  AOI211X1 U124 ( .C(n2431), .D(n2436), .A(n170), .B(n902), .Y(n899) );
  INVX1 U125 ( .A(n2489), .Y(n90) );
  AOI21X1 U126 ( .B(n149), .C(n221), .A(n248), .Y(n1113) );
  INVX1 U127 ( .A(n1113), .Y(n91) );
  INVX1 U128 ( .A(n1113), .Y(n92) );
  AOI21X1 U129 ( .B(n148), .C(n220), .A(n247), .Y(n1119) );
  INVX1 U130 ( .A(n1119), .Y(n93) );
  INVX1 U131 ( .A(n1119), .Y(n94) );
  BUFX3 U132 ( .A(n1122), .Y(n95) );
  NAND2X1 U133 ( .A(n2013), .B(n2025), .Y(n1807) );
  INVX1 U134 ( .A(n1807), .Y(n96) );
  INVX1 U135 ( .A(n1807), .Y(n97) );
  NAND2X1 U136 ( .A(n2026), .B(n2010), .Y(n1809) );
  INVX1 U137 ( .A(n1809), .Y(n98) );
  INVX1 U138 ( .A(n1809), .Y(n99) );
  NAND2X1 U139 ( .A(n2008), .B(n2009), .Y(n1793) );
  INVX1 U140 ( .A(n1793), .Y(n100) );
  INVX1 U141 ( .A(n1793), .Y(n101) );
  INVX1 U142 ( .A(n147), .Y(instr[5]) );
  INVX1 U143 ( .A(n2453), .Y(pc_o[11]) );
  NOR3XL U144 ( .A(n1332), .B(n2366), .C(n1333), .Y(n104) );
  NOR3XL U145 ( .A(n1089), .B(n2325), .C(n2364), .Y(n105) );
  NOR3XL U146 ( .A(n1089), .B(n2325), .C(n2364), .Y(n1152) );
  INVX1 U147 ( .A(n168), .Y(n106) );
  INVX1 U148 ( .A(n2403), .Y(n107) );
  BUFX3 U149 ( .A(n2186), .Y(n109) );
  INVX1 U150 ( .A(n153), .Y(n110) );
  AOI21X1 U151 ( .B(n105), .C(n221), .A(n2162), .Y(n1103) );
  INVX1 U152 ( .A(n1103), .Y(n111) );
  INVX1 U153 ( .A(n1103), .Y(n112) );
  AOI21X1 U154 ( .B(n166), .C(n220), .A(n248), .Y(n1111) );
  INVX1 U155 ( .A(n1111), .Y(n113) );
  INVX1 U156 ( .A(n1111), .Y(n114) );
  BUFX3 U157 ( .A(n1114), .Y(n115) );
  NAND2X1 U158 ( .A(n2026), .B(n2013), .Y(n1811) );
  INVX1 U159 ( .A(n1811), .Y(n116) );
  INVX1 U160 ( .A(n1811), .Y(n117) );
  NAND2X1 U161 ( .A(n2009), .B(n2025), .Y(n1804) );
  INVX1 U162 ( .A(n1804), .Y(n118) );
  INVX1 U163 ( .A(n1804), .Y(n119) );
  NAND2X1 U164 ( .A(n2008), .B(n2010), .Y(n1792) );
  INVX1 U165 ( .A(n1792), .Y(n120) );
  INVX1 U166 ( .A(n1792), .Y(n121) );
  INVX1 U167 ( .A(n2464), .Y(pc_o[14]) );
  BUFX3 U168 ( .A(accactv), .Y(n123) );
  NAND2X1 U169 ( .A(n396), .B(pc_o[0]), .Y(n413) );
  NOR3XL U170 ( .A(n2364), .B(n1089), .C(n1333), .Y(n124) );
  NOR3XL U171 ( .A(n2364), .B(n1089), .C(n1333), .Y(n1148) );
  NOR3XL U172 ( .A(n2366), .B(n2325), .C(n1332), .Y(n125) );
  NOR3XL U173 ( .A(n2366), .B(n2325), .C(n1332), .Y(n1149) );
  BUFX3 U174 ( .A(n2506), .Y(n2260) );
  INVX1 U175 ( .A(n2260), .Y(n126) );
  INVX1 U176 ( .A(n2260), .Y(n128) );
  INVX1 U177 ( .A(n458), .Y(n130) );
  BUFX3 U178 ( .A(n2478), .Y(n131) );
  INVX1 U179 ( .A(n2499), .Y(n132) );
  INVX1 U180 ( .A(n132), .Y(mempswr) );
  INVX1 U181 ( .A(n1356), .Y(n134) );
  AOI21X1 U182 ( .B(n125), .C(n220), .A(n2162), .Y(n1115) );
  INVX1 U183 ( .A(n1115), .Y(n135) );
  INVX1 U184 ( .A(n1115), .Y(n136) );
  AOI21X1 U185 ( .B(n165), .C(n221), .A(n248), .Y(n1121) );
  INVX1 U186 ( .A(n1121), .Y(n137) );
  INVX1 U187 ( .A(n1121), .Y(n138) );
  BUFX3 U188 ( .A(n1112), .Y(n139) );
  NAND2X1 U189 ( .A(n2008), .B(n2012), .Y(n1812) );
  INVX1 U190 ( .A(n1812), .Y(n140) );
  INVX1 U191 ( .A(n1812), .Y(n141) );
  NAND2X1 U192 ( .A(n2010), .B(n2025), .Y(n1806) );
  INVX1 U193 ( .A(n1806), .Y(n142) );
  INVX1 U194 ( .A(n1806), .Y(n143) );
  NAND2X1 U195 ( .A(n2011), .B(n2009), .Y(n1797) );
  INVX1 U196 ( .A(n1797), .Y(n144) );
  INVX1 U197 ( .A(n1797), .Y(n145) );
  INVX1 U198 ( .A(n2468), .Y(pc_o[7]) );
  BUFX3 U199 ( .A(n2243), .Y(n147) );
  NOR3XL U200 ( .A(n2366), .B(n2364), .C(n1333), .Y(n148) );
  NOR3XL U201 ( .A(n1089), .B(n2325), .C(n1332), .Y(n149) );
  NOR3XL U202 ( .A(n1089), .B(n2325), .C(n1332), .Y(n1150) );
  INVX1 U203 ( .A(n2473), .Y(n150) );
  INVX1 U204 ( .A(n2484), .Y(n151) );
  BUFX3 U205 ( .A(n2324), .Y(n152) );
  BUFX3 U206 ( .A(n1134), .Y(n153) );
  INVX1 U207 ( .A(acc[1]), .Y(n154) );
  BUFX3 U208 ( .A(n1120), .Y(n155) );
  BUFX3 U209 ( .A(n1829), .Y(n156) );
  NAND2X1 U210 ( .A(n2026), .B(n2009), .Y(n1810) );
  INVX1 U211 ( .A(n1810), .Y(n157) );
  INVX1 U212 ( .A(n1810), .Y(n158) );
  NAND2X1 U213 ( .A(n2025), .B(n2012), .Y(n1805) );
  INVX1 U214 ( .A(n1805), .Y(n159) );
  INVX1 U215 ( .A(n1805), .Y(n160) );
  NAND2X1 U216 ( .A(n2011), .B(n2010), .Y(n1796) );
  INVX1 U217 ( .A(n1796), .Y(n161) );
  INVX1 U218 ( .A(n1796), .Y(n162) );
  INVX1 U219 ( .A(n2465), .Y(pc_o[3]) );
  INVX1 U220 ( .A(n1138), .Y(n222) );
  INVX1 U221 ( .A(n222), .Y(n164) );
  NOR3XL U222 ( .A(n1332), .B(n1089), .C(n1333), .Y(n165) );
  NOR3XL U223 ( .A(n1332), .B(n1089), .C(n1333), .Y(n1146) );
  NOR3XL U224 ( .A(n2364), .B(n2325), .C(n2366), .Y(n166) );
  NOR3XL U225 ( .A(n2364), .B(n2325), .C(n2366), .Y(n1151) );
  BUFX3 U226 ( .A(n2506), .Y(instr[4]) );
  BUFX3 U227 ( .A(phase[0]), .Y(n2183) );
  INVX1 U228 ( .A(n2183), .Y(n168) );
  INVX1 U229 ( .A(n2183), .Y(n169) );
  INVX1 U230 ( .A(n2183), .Y(n170) );
  OR2X2 U231 ( .A(n354), .B(n1462), .Y(n171) );
  OR2X1 U232 ( .A(n2493), .B(n353), .Y(n172) );
  NAND3X1 U233 ( .A(n171), .B(n172), .C(n173), .Y(n1437) );
  AO21X1 U234 ( .B(n336), .C(n337), .A(n2187), .Y(n354) );
  INVX1 U235 ( .A(sfrdatai[2]), .Y(n1462) );
  MUX2XL U236 ( .D0(pc_o[0]), .D1(n1713), .S(n14), .Y(memaddr_comb[0]) );
  OR2X1 U237 ( .A(n938), .B(n352), .Y(n173) );
  NAND2XL U238 ( .A(n354), .B(n352), .Y(n353) );
  INVXL U239 ( .A(n1437), .Y(n1442) );
  NOR2XL U240 ( .A(n353), .B(n654), .Y(n175) );
  NOR2X1 U241 ( .A(n928), .B(n352), .Y(n176) );
  NOR2XL U242 ( .A(n184), .B(n181), .Y(n180) );
  INVX1 U243 ( .A(n394), .Y(n181) );
  AND3X2 U244 ( .A(n1500), .B(n454), .C(n208), .Y(n507) );
  OR3XL U245 ( .A(n1886), .B(n180), .C(n209), .Y(n414) );
  NOR2XL U246 ( .A(n1933), .B(n354), .Y(n177) );
  NOR2XL U247 ( .A(n353), .B(n1954), .Y(n178) );
  NOR2X1 U248 ( .A(n923), .B(n352), .Y(n179) );
  NAND21XL U249 ( .B(n2500), .A(n287), .Y(N370) );
  NAND21XL U250 ( .B(n1712), .A(n237), .Y(n618) );
  NAND21XL U251 ( .B(n247), .A(n1712), .Y(n617) );
  INVXL U252 ( .A(n463), .Y(n474) );
  INVXL U253 ( .A(n2500), .Y(n286) );
  INVXL U254 ( .A(n723), .Y(n727) );
  NAND2X2 U255 ( .A(n619), .B(n616), .Y(n930) );
  NAND21XL U256 ( .B(n394), .A(n184), .Y(n395) );
  AOI31XL U257 ( .A(n1779), .B(n689), .C(n480), .D(n474), .Y(n481) );
  AOI221XL U258 ( .A(n2311), .B(n1778), .C(n1777), .D(memdatai[5]), .E(n1852), 
        .Y(n450) );
  AND2XL U259 ( .A(n241), .B(n1657), .Y(N11499) );
  XNOR3X1 U260 ( .A(n887), .B(n890), .C(n182), .Y(n858) );
  XNOR2XL U261 ( .A(n857), .B(n830), .Y(n182) );
  AND2XL U262 ( .A(n242), .B(n857), .Y(N12470) );
  MUX2IX1 U263 ( .D0(n1409), .D1(n2228), .S(n377), .Y(n372) );
  OAI211XL U264 ( .C(n1738), .D(n787), .A(n430), .B(n429), .Y(n829) );
  OAI222XL U265 ( .A(n440), .B(n1373), .C(n435), .D(n448), .E(n734), .F(n447), 
        .Y(n1693) );
  OAI222XL U266 ( .A(n584), .B(n2245), .C(n170), .D(n187), .E(n1758), .F(n261), 
        .Y(n1653) );
  NAND3XL U267 ( .A(n1624), .B(memack), .C(n1619), .Y(n2155) );
  NAND2X2 U268 ( .A(n507), .B(n496), .Y(n1575) );
  MUX2XL U269 ( .D0(pc_o[6]), .D1(n1719), .S(n14), .Y(memaddr_comb[6]) );
  INVX1 U270 ( .A(n395), .Y(n209) );
  AO2222XL U271 ( .A(pc_o[8]), .B(n411), .C(n2246), .D(temp2_comb[0]), .E(
        n2239), .F(pc_i[0]), .G(n410), .H(n812), .Y(n412) );
  AOI222XL U272 ( .A(n1136), .B(temp[0]), .C(n1137), .D(n2139), .E(dptr_inc[0]), .F(n164), .Y(n736) );
  AOI222XL U273 ( .A(n1136), .B(temp[1]), .C(n1137), .D(n2138), .E(dptr_inc[1]), .F(n164), .Y(n731) );
  AOI222XL U274 ( .A(n1136), .B(temp[2]), .C(n1137), .D(n2137), .E(dptr_inc[2]), .F(n164), .Y(n726) );
  OAI222XL U275 ( .A(n1784), .B(n1783), .C(ramdatao[7]), .D(n1787), .E(n1786), 
        .F(n1785), .Y(n908) );
  AOI222XL U276 ( .A(n1136), .B(temp[5]), .C(n1137), .D(n2135), .E(dptr_inc[5]), .F(n164), .Y(n711) );
  AOI222XL U277 ( .A(n1136), .B(temp[3]), .C(n1137), .D(n2127), .E(dptr_inc[3]), .F(n164), .Y(n721) );
  AOI222XL U278 ( .A(n1136), .B(temp[4]), .C(n1137), .D(n2136), .E(dptr_inc[4]), .F(n164), .Y(n716) );
  OAI222XL U279 ( .A(n1908), .B(n1907), .C(ramdatao[3]), .D(n1787), .E(n1910), 
        .F(n1909), .Y(n933) );
  AOI222XL U280 ( .A(n1136), .B(temp[6]), .C(n1137), .D(n2134), .E(dptr_inc[6]), .F(n164), .Y(n706) );
  OAI222XL U281 ( .A(n1831), .B(n1830), .C(ramdatao[6]), .D(n1787), .E(n1833), 
        .F(n1832), .Y(n918) );
  AOI22AXL U282 ( .A(sp[5]), .B(n156), .D(n1829), .C(ramdatao[5]), .Y(n1855)
         );
  AOI22AXL U283 ( .A(sp[7]), .B(n156), .D(n156), .C(ramdatao[7]), .Y(n1826) );
  AOI222XL U284 ( .A(n1136), .B(temp[7]), .C(n1137), .D(n2144), .E(dptr_inc[7]), .F(n164), .Y(n698) );
  OAI31XL U285 ( .A(n1562), .B(n613), .C(n309), .D(mempsrd), .Y(n588) );
  NOR3XL U286 ( .A(n2442), .B(ramsfraddr[2]), .C(n2443), .Y(n856) );
  INVX1 U287 ( .A(n247), .Y(n237) );
  INVX1 U288 ( .A(n246), .Y(n238) );
  INVX1 U289 ( .A(n246), .Y(n239) );
  INVX1 U290 ( .A(n245), .Y(n243) );
  INVX1 U291 ( .A(n246), .Y(n240) );
  INVX1 U292 ( .A(n245), .Y(n242) );
  INVX1 U293 ( .A(n245), .Y(n241) );
  INVX1 U294 ( .A(n250), .Y(n247) );
  INVX1 U295 ( .A(n250), .Y(n246) );
  INVX1 U296 ( .A(n250), .Y(n245) );
  INVX1 U297 ( .A(n2162), .Y(n244) );
  INVX1 U298 ( .A(n250), .Y(n248) );
  INVX1 U299 ( .A(n2162), .Y(n250) );
  INVX1 U300 ( .A(n2162), .Y(n249) );
  INVX1 U301 ( .A(n2160), .Y(n2233) );
  INVX1 U302 ( .A(n737), .Y(n627) );
  INVX1 U303 ( .A(n2423), .Y(n2255) );
  INVX1 U304 ( .A(n286), .Y(n284) );
  INVX1 U305 ( .A(n957), .Y(n2272) );
  INVX1 U306 ( .A(n2165), .Y(n2193) );
  INVX1 U307 ( .A(n713), .Y(n2213) );
  NAND21X1 U308 ( .B(n292), .A(n283), .Y(n2162) );
  INVX1 U309 ( .A(n286), .Y(waitstaten) );
  INVX1 U310 ( .A(n2067), .Y(n282) );
  INVX1 U311 ( .A(n2279), .Y(n264) );
  INVX1 U312 ( .A(n2280), .Y(n251) );
  INVX1 U313 ( .A(n2283), .Y(n255) );
  INVX1 U314 ( .A(n2278), .Y(n278) );
  INVX1 U315 ( .A(n2277), .Y(n275) );
  INVX1 U316 ( .A(n2278), .Y(n279) );
  INVX1 U317 ( .A(n2277), .Y(n276) );
  INVX1 U318 ( .A(n2280), .Y(n252) );
  INVX1 U319 ( .A(n2283), .Y(n256) );
  INVX1 U320 ( .A(n2067), .Y(n281) );
  INVX1 U321 ( .A(n2283), .Y(n257) );
  INVX1 U322 ( .A(n765), .Y(n269) );
  INVX1 U323 ( .A(n2280), .Y(n253) );
  INVX1 U324 ( .A(n2279), .Y(n265) );
  INVX1 U325 ( .A(n2276), .Y(n272) );
  INVX1 U326 ( .A(n2067), .Y(n280) );
  INVX1 U327 ( .A(n2279), .Y(n266) );
  INVX1 U328 ( .A(n765), .Y(n270) );
  INVX1 U329 ( .A(n2276), .Y(n273) );
  INVX1 U330 ( .A(n2283), .Y(n258) );
  INVX1 U331 ( .A(n2280), .Y(n254) );
  INVX1 U332 ( .A(n2279), .Y(n267) );
  INVX1 U333 ( .A(n1507), .Y(n2254) );
  INVX1 U334 ( .A(n759), .Y(n2211) );
  AND2X1 U335 ( .A(n240), .B(n1694), .Y(N11482) );
  AND2X1 U336 ( .A(n241), .B(n1695), .Y(N11483) );
  AND2X1 U337 ( .A(n241), .B(n1696), .Y(N11484) );
  INVX1 U338 ( .A(n2386), .Y(n2230) );
  INVX1 U339 ( .A(rst), .Y(n287) );
  INVX1 U340 ( .A(rst), .Y(n288) );
  INVX1 U341 ( .A(rst), .Y(n289) );
  INVX1 U342 ( .A(n292), .Y(n290) );
  INVX1 U343 ( .A(n443), .Y(sfrwe_comb_s) );
  INVXL U344 ( .A(n363), .Y(n374) );
  NAND21X1 U345 ( .B(n1994), .A(n375), .Y(n376) );
  NAND21X1 U346 ( .B(n1436), .A(n374), .Y(n375) );
  NAND21X1 U347 ( .B(n1407), .A(n2093), .Y(n2160) );
  NAND21XL U348 ( .B(n1712), .A(n1424), .Y(n929) );
  INVX1 U349 ( .A(n286), .Y(n283) );
  NAND4X1 U350 ( .A(n781), .B(n2233), .C(n1369), .D(n2345), .Y(n737) );
  INVX1 U351 ( .A(n1697), .Y(n1654) );
  INVX1 U352 ( .A(n1777), .Y(n440) );
  NAND21X1 U353 ( .B(n591), .A(n1697), .Y(n443) );
  INVX1 U354 ( .A(n1538), .Y(n1405) );
  NOR21XL U355 ( .B(n2233), .A(n685), .Y(n664) );
  NAND21X1 U356 ( .B(n2433), .A(n2256), .Y(n2423) );
  NAND21X1 U357 ( .B(n2160), .A(n685), .Y(n861) );
  INVX1 U358 ( .A(n1450), .Y(n2328) );
  INVXL U359 ( .A(n1988), .Y(n1995) );
  AO21X1 U360 ( .B(n1534), .C(memdatai[7]), .A(n2275), .Y(N677) );
  AO21X1 U361 ( .B(n1534), .C(memdatai[5]), .A(n2275), .Y(N675) );
  OAI21X1 U362 ( .B(n261), .C(n2387), .A(n444), .Y(n1986) );
  INVX1 U363 ( .A(n1824), .Y(n2339) );
  INVX1 U364 ( .A(n1607), .Y(n2181) );
  NOR2X1 U365 ( .A(n734), .B(n594), .Y(N676) );
  NOR2X1 U366 ( .A(n1373), .B(n594), .Y(N673) );
  NOR2X1 U367 ( .A(n670), .B(n594), .Y(N674) );
  INVX1 U368 ( .A(n2388), .Y(n1702) );
  INVX1 U369 ( .A(n2387), .Y(n1987) );
  NAND21X1 U370 ( .B(n1702), .A(n337), .Y(n398) );
  NAND2X1 U371 ( .A(n2252), .B(n1762), .Y(n798) );
  INVX1 U372 ( .A(n1725), .Y(n446) );
  NAND21X1 U373 ( .B(n2395), .A(n2388), .Y(n366) );
  NAND32X1 U374 ( .B(n367), .C(n366), .A(n694), .Y(n1887) );
  INVX1 U375 ( .A(n364), .Y(n367) );
  INVX1 U376 ( .A(n1532), .Y(n410) );
  INVX1 U377 ( .A(n396), .Y(n432) );
  OR2X1 U378 ( .A(n1625), .B(n1765), .Y(n2046) );
  INVX1 U379 ( .A(n760), .Y(n388) );
  INVX1 U380 ( .A(n1765), .Y(n2393) );
  INVX1 U381 ( .A(n1735), .Y(n386) );
  INVX1 U382 ( .A(n767), .Y(n419) );
  NAND21X1 U383 ( .B(n1661), .A(n237), .Y(n2165) );
  INVX1 U384 ( .A(n1436), .Y(n2228) );
  INVX1 U385 ( .A(n694), .Y(n1994) );
  INVX1 U386 ( .A(n371), .Y(n2226) );
  INVX1 U387 ( .A(n322), .Y(n2244) );
  INVX1 U388 ( .A(n330), .Y(n1746) );
  NAND21X1 U389 ( .B(n366), .A(n336), .Y(n330) );
  INVX1 U390 ( .A(n2395), .Y(n314) );
  NAND3X1 U391 ( .A(n755), .B(n2272), .C(n756), .Y(n754) );
  NAND21X1 U392 ( .B(n1666), .A(n238), .Y(n713) );
  NOR2X1 U393 ( .A(n388), .B(n2434), .Y(n957) );
  INVX1 U394 ( .A(n2166), .Y(n2209) );
  INVX1 U395 ( .A(n2167), .Y(n2217) );
  INVX1 U396 ( .A(n2161), .Y(n2196) );
  NAND21X1 U397 ( .B(n1659), .A(n283), .Y(n1691) );
  INVX1 U398 ( .A(n742), .Y(n2158) );
  INVX1 U399 ( .A(n2121), .Y(n1227) );
  NAND21X1 U400 ( .B(n2093), .A(n237), .Y(n2121) );
  NAND2X1 U401 ( .A(n1227), .B(n166), .Y(n1112) );
  INVX1 U402 ( .A(n765), .Y(n268) );
  INVX1 U403 ( .A(n2277), .Y(n274) );
  INVX1 U404 ( .A(n2278), .Y(n277) );
  INVX1 U405 ( .A(n2276), .Y(n271) );
  NAND21X1 U406 ( .B(n591), .A(n237), .Y(n1507) );
  NAND21X1 U407 ( .B(n2266), .A(n238), .Y(n759) );
  AND2X1 U408 ( .A(n685), .B(n2237), .Y(n183) );
  NAND21X1 U409 ( .B(n1659), .A(n238), .Y(n1490) );
  AO21X1 U410 ( .B(n166), .C(n244), .A(n295), .Y(N12547) );
  OA21X1 U411 ( .B(n957), .C(n2164), .A(n250), .Y(N10572) );
  INVX1 U412 ( .A(n797), .Y(n2164) );
  NOR32XL U413 ( .B(n239), .C(n2180), .A(n2040), .Y(N10576) );
  AND2X1 U414 ( .A(n2254), .B(n1697), .Y(N11489) );
  AND2X1 U415 ( .A(n2168), .B(n2394), .Y(N10568) );
  NOR2X1 U416 ( .A(n2040), .B(n2047), .Y(N10570) );
  AND2X1 U417 ( .A(n241), .B(n1697), .Y(N11485) );
  AND2X1 U418 ( .A(n241), .B(n2357), .Y(N12710) );
  AND2X1 U419 ( .A(n242), .B(n2174), .Y(n2284) );
  NAND32X1 U420 ( .B(n581), .C(n582), .A(n2173), .Y(n2174) );
  NAND31X1 U421 ( .C(n583), .A(n2267), .B(n584), .Y(n582) );
  INVX1 U422 ( .A(n466), .Y(n2224) );
  INVX1 U423 ( .A(n595), .Y(n2225) );
  INVX1 U424 ( .A(n467), .Y(n2257) );
  INVX1 U425 ( .A(n450), .Y(n1695) );
  INVX1 U426 ( .A(n449), .Y(n1696) );
  INVX1 U427 ( .A(n451), .Y(n1694) );
  INVX1 U428 ( .A(n1934), .Y(n2200) );
  INVX1 U429 ( .A(n1932), .Y(n2201) );
  INVX1 U430 ( .A(n1531), .Y(n2240) );
  NAND21X1 U431 ( .B(n2416), .A(n2252), .Y(n2386) );
  OAI21X1 U432 ( .B(n2378), .C(n261), .A(n999), .Y(n977) );
  INVX1 U433 ( .A(n297), .Y(n292) );
  INVX1 U434 ( .A(n939), .Y(n2343) );
  INVX1 U435 ( .A(n906), .Y(n2271) );
  OAI21X1 U436 ( .B(n2434), .C(n2393), .A(n798), .Y(n2064) );
  NOR2X1 U437 ( .A(n2046), .B(n760), .Y(n2045) );
  INVX1 U438 ( .A(n296), .Y(n295) );
  NOR2X1 U439 ( .A(n2266), .B(n291), .Y(n477) );
  INVX1 U440 ( .A(n297), .Y(n293) );
  INVX1 U441 ( .A(n296), .Y(n294) );
  MUX2X1 U442 ( .D0(n2499), .D1(n1703), .S(n283), .Y(mempswr_comb) );
  OAI22X1 U443 ( .A(n975), .B(n354), .C(n2491), .D(n353), .Y(n723) );
  OAI22X1 U444 ( .A(n354), .B(n775), .C(n2494), .D(n353), .Y(n463) );
  OAI222XL U445 ( .A(n775), .B(n1932), .C(n2494), .D(n1934), .E(n944), .F(
        n1931), .Y(n1443) );
  INVX1 U446 ( .A(n1658), .Y(n2500) );
  OAI22X1 U447 ( .A(n354), .B(n639), .C(n2492), .D(n353), .Y(n1743) );
  MUX2X1 U448 ( .D0(n1436), .D1(n2229), .S(n202), .Y(n480) );
  NAND21X1 U449 ( .B(n900), .A(n619), .Y(n1407) );
  INVX1 U450 ( .A(n626), .Y(n1341) );
  NAND32X1 U451 ( .B(n692), .C(n636), .A(n627), .Y(n626) );
  INVX1 U452 ( .A(N13353), .Y(n2273) );
  INVX1 U453 ( .A(n701), .Y(n1371) );
  NOR21XL U454 ( .B(n692), .A(n737), .Y(n701) );
  OAI21X1 U455 ( .B(n1524), .C(n1523), .A(n2202), .Y(n1525) );
  OAI22X1 U456 ( .A(n2285), .B(n440), .C(n1509), .D(n448), .Y(n1697) );
  AOI21X1 U457 ( .B(n2285), .C(n1929), .A(n1778), .Y(n1777) );
  INVX1 U458 ( .A(memdatai[7]), .Y(n2285) );
  OR2X1 U459 ( .A(n1420), .B(n1421), .Y(n1419) );
  NAND5XL U460 ( .A(n450), .B(n449), .C(n453), .D(n451), .E(n452), .Y(n1538)
         );
  INVX1 U461 ( .A(n1693), .Y(n453) );
  AND4X1 U462 ( .A(sfrwe_comb_s), .B(n198), .C(n1692), .D(n197), .Y(n452) );
  INVX1 U463 ( .A(n1705), .Y(n1709) );
  OAI21BBX1 U464 ( .A(n575), .B(n576), .C(n578), .Y(n577) );
  INVX1 U465 ( .A(n1367), .Y(n2481) );
  INVX1 U466 ( .A(n876), .Y(n2311) );
  AOI22AXL U467 ( .A(n1777), .B(memdatai[6]), .D(n880), .C(n1778), .Y(n449) );
  AOI22X1 U468 ( .A(n1777), .B(memdatai[4]), .C(n884), .D(n1778), .Y(n451) );
  INVX1 U469 ( .A(memdatai[3]), .Y(n1373) );
  INVX1 U470 ( .A(memdatai[6]), .Y(n734) );
  INVX1 U471 ( .A(memdatai[0]), .Y(n826) );
  INVX1 U472 ( .A(n1852), .Y(n447) );
  NOR32XL U473 ( .B(n1045), .C(n1358), .A(n1361), .Y(n1450) );
  NAND21X1 U474 ( .B(n259), .A(n2255), .Y(n444) );
  NAND32X1 U475 ( .B(n636), .C(n861), .A(n860), .Y(n1424) );
  INVX1 U476 ( .A(n974), .Y(n2256) );
  INVX1 U477 ( .A(n2050), .Y(n2433) );
  INVX1 U478 ( .A(memdatai[1]), .Y(n791) );
  OR2X1 U479 ( .A(n2232), .B(n2198), .Y(n185) );
  INVX1 U480 ( .A(n1683), .Y(n2350) );
  INVX1 U481 ( .A(n722), .Y(n2053) );
  INVX1 U482 ( .A(n745), .Y(n2432) );
  INVX1 U483 ( .A(n1395), .Y(n2333) );
  OAI21X1 U484 ( .B(n690), .C(n1986), .A(n2341), .Y(n1824) );
  INVX1 U485 ( .A(n1349), .Y(n2334) );
  INVX1 U486 ( .A(n1037), .Y(n2357) );
  OAI222XL U487 ( .A(n1954), .B(n1934), .C(n1933), .D(n1932), .E(n923), .F(
        n1931), .Y(n1955) );
  INVX1 U488 ( .A(n951), .Y(n441) );
  INVX1 U489 ( .A(n1032), .Y(n2351) );
  NOR2X1 U490 ( .A(n2377), .B(n2020), .Y(n2010) );
  NOR2X1 U491 ( .A(n2419), .B(n2377), .Y(n2012) );
  OAI22X1 U492 ( .A(n1686), .B(n1490), .C(n1489), .D(n713), .Y(N11503) );
  INVX1 U493 ( .A(n312), .Y(n316) );
  NAND21X1 U494 ( .B(n259), .A(n311), .Y(n312) );
  INVX1 U495 ( .A(n476), .Y(n2402) );
  INVX1 U496 ( .A(n1850), .Y(n2342) );
  NAND21X1 U497 ( .B(n805), .A(n2252), .Y(n2387) );
  NAND21X1 U498 ( .B(n1573), .A(n237), .Y(n1607) );
  AO21X1 U499 ( .B(n1499), .C(n1705), .A(n292), .Y(n1542) );
  INVX1 U500 ( .A(n2389), .Y(n2252) );
  XNOR2XL U501 ( .A(n1596), .B(n576), .Y(n1595) );
  XOR2X1 U502 ( .A(n575), .B(n578), .Y(n1596) );
  NOR2X1 U503 ( .A(n805), .B(n773), .Y(n1726) );
  NAND2X1 U504 ( .A(n1984), .B(n2388), .Y(n1780) );
  NAND2X1 U505 ( .A(n1702), .B(n1984), .Y(n1781) );
  INVX1 U506 ( .A(n746), .Y(n2434) );
  INVX1 U507 ( .A(n262), .Y(n260) );
  OR2X1 U508 ( .A(n593), .B(n585), .Y(n594) );
  OAI22X1 U509 ( .A(n1665), .B(n1490), .C(n1489), .D(n2167), .Y(N11502) );
  OAI21X1 U510 ( .B(n593), .C(n466), .A(n464), .Y(N672) );
  OAI21X1 U511 ( .B(n593), .C(n467), .A(n464), .Y(N670) );
  INVX1 U512 ( .A(memdatai[5]), .Y(n686) );
  INVX1 U513 ( .A(memdatai[4]), .Y(n670) );
  AND2X1 U514 ( .A(n240), .B(n1664), .Y(N11501) );
  INVX1 U515 ( .A(n464), .Y(n2275) );
  INVX1 U516 ( .A(n772), .Y(n2270) );
  AOI31X1 U517 ( .A(n1546), .B(n1779), .C(n1992), .D(n1767), .Y(n1856) );
  EORX1 U518 ( .A(n2178), .B(n2228), .C(n2178), .D(n2229), .Y(n1546) );
  INVX1 U519 ( .A(n590), .Y(n1534) );
  NAND21X1 U520 ( .B(n593), .A(n237), .Y(n590) );
  INVX1 U521 ( .A(n2020), .Y(n2419) );
  NAND21X1 U522 ( .B(n259), .A(n322), .Y(n2388) );
  NAND21X1 U523 ( .B(n324), .A(n2227), .Y(n1710) );
  AO21X1 U524 ( .B(n1735), .C(n2185), .A(n1987), .Y(n322) );
  NAND43X1 U525 ( .B(n326), .C(n1722), .D(n1690), .A(n358), .Y(n371) );
  INVX1 U526 ( .A(n1710), .Y(n326) );
  NAND21X1 U527 ( .B(n259), .A(n768), .Y(n1744) );
  NAND2X1 U528 ( .A(n2361), .B(n1989), .Y(n1782) );
  NOR2X1 U529 ( .A(n2416), .B(n2396), .Y(n1735) );
  NOR2X1 U530 ( .A(n2436), .B(n772), .Y(n1725) );
  INVX1 U531 ( .A(n338), .Y(n336) );
  INVX1 U532 ( .A(n1014), .Y(n2269) );
  INVX1 U533 ( .A(n813), .Y(n2330) );
  INVX1 U534 ( .A(n262), .Y(n261) );
  NOR2X1 U535 ( .A(n2425), .B(n2427), .Y(n1762) );
  OAI22X1 U536 ( .A(n585), .B(n1570), .C(n586), .D(codefetch_s), .Y(N679) );
  INVX1 U537 ( .A(n1632), .Y(n2385) );
  NOR2X1 U538 ( .A(n1771), .B(n1726), .Y(n1750) );
  INVX1 U539 ( .A(n758), .Y(n2416) );
  NAND2X1 U540 ( .A(n2389), .B(n773), .Y(n1634) );
  INVX1 U541 ( .A(n1486), .Y(n2352) );
  NAND21X1 U542 ( .B(n2389), .A(n2256), .Y(n364) );
  OR4X1 U543 ( .A(n399), .B(n398), .C(n1957), .D(n186), .Y(n1532) );
  AOI21X1 U544 ( .B(n2173), .C(n2267), .A(n261), .Y(n186) );
  NAND21X1 U545 ( .B(n1647), .A(n2242), .Y(n358) );
  OAI211X1 U546 ( .C(n1727), .D(n2434), .A(n313), .B(n446), .Y(n2395) );
  INVX1 U547 ( .A(n1726), .Y(n313) );
  OR2X1 U548 ( .A(n338), .B(n398), .Y(n352) );
  NAND2X1 U549 ( .A(n369), .B(n364), .Y(n327) );
  NAND21X1 U550 ( .B(n259), .A(n2395), .Y(n337) );
  NOR2X1 U551 ( .A(n2100), .B(n2427), .Y(n1765) );
  OR3XL U552 ( .A(n1689), .B(n1414), .C(n319), .Y(n399) );
  INVX1 U553 ( .A(n1489), .Y(n1659) );
  INVX1 U554 ( .A(n324), .Y(n2242) );
  OAI21X1 U555 ( .B(n2437), .C(n2393), .A(n798), .Y(n581) );
  NOR2X1 U556 ( .A(n164), .B(n1136), .Y(n1137) );
  INVX1 U557 ( .A(n325), .Y(n1722) );
  NAND21X1 U558 ( .B(n773), .A(n2256), .Y(n325) );
  NAND2X1 U559 ( .A(n1704), .B(n1698), .Y(n1706) );
  INVX1 U560 ( .A(n1139), .Y(n2401) );
  INVX1 U561 ( .A(n1778), .Y(n448) );
  INVX1 U562 ( .A(n2152), .Y(n1666) );
  INVX1 U563 ( .A(n892), .Y(n1661) );
  AO21X1 U564 ( .B(n1698), .C(n369), .A(n368), .Y(n1436) );
  AO21X1 U565 ( .B(n1704), .C(n365), .A(n368), .Y(n694) );
  NAND32X1 U566 ( .B(n2396), .C(n2429), .A(n2269), .Y(n365) );
  NAND21X1 U567 ( .B(n2250), .A(n384), .Y(n1934) );
  OR2X1 U568 ( .A(n2250), .B(n384), .Y(n1932) );
  NAND21X1 U569 ( .B(n2247), .A(n1533), .Y(n396) );
  AOI21X1 U570 ( .B(n2046), .C(n746), .A(n956), .Y(n797) );
  NOR43XL U571 ( .B(n2244), .C(n776), .D(n743), .A(n777), .Y(n762) );
  NOR2X1 U572 ( .A(n2418), .B(n2392), .Y(n760) );
  INVX1 U573 ( .A(n945), .Y(n2247) );
  AND4X1 U574 ( .A(n761), .B(n762), .C(n763), .D(n764), .Y(n755) );
  AOI211X1 U575 ( .C(n760), .D(n2180), .A(n766), .B(n767), .Y(n764) );
  NOR32XL U576 ( .B(n187), .C(n779), .A(n780), .Y(n761) );
  NOR3XL U577 ( .A(n770), .B(n2395), .C(n580), .Y(n763) );
  OR2X1 U578 ( .A(n1409), .B(n366), .Y(n368) );
  NOR2X1 U579 ( .A(n2393), .B(n2431), .Y(n767) );
  NOR2X1 U580 ( .A(n2437), .B(n772), .Y(n583) );
  INVX1 U581 ( .A(n580), .Y(n2173) );
  INVX1 U582 ( .A(n1647), .Y(n2241) );
  INVX1 U583 ( .A(n900), .Y(n982) );
  INVX1 U584 ( .A(n2431), .Y(n2180) );
  INVX1 U585 ( .A(n1931), .Y(n2250) );
  AOI21X1 U586 ( .B(n2379), .C(n2179), .A(n1706), .Y(n779) );
  INVX1 U587 ( .A(n1550), .Y(n492) );
  INVX1 U588 ( .A(n1372), .Y(n921) );
  NOR2X1 U589 ( .A(n16), .B(n2100), .Y(n1625) );
  AOI21AX1 U590 ( .B(n1765), .C(n2184), .A(n436), .Y(n187) );
  INVX1 U591 ( .A(n2142), .Y(n2093) );
  AND2X1 U592 ( .A(n242), .B(n858), .Y(N12905) );
  XNOR2XL U593 ( .A(n894), .B(n895), .Y(n887) );
  AND2XL U594 ( .A(n242), .B(n1656), .Y(N11498) );
  INVX1 U595 ( .A(n751), .Y(n2392) );
  NOR3XL U596 ( .A(n2428), .B(n972), .C(n2425), .Y(n1626) );
  OR2X1 U597 ( .A(n2114), .B(n2050), .Y(n1635) );
  NAND2X1 U598 ( .A(n1651), .B(n2437), .Y(n1749) );
  INVX1 U599 ( .A(n1644), .Y(n2383) );
  INVX1 U600 ( .A(n601), .Y(n620) );
  INVX1 U601 ( .A(n805), .Y(n2424) );
  NAND21X1 U602 ( .B(n319), .A(n316), .Y(n1531) );
  XOR2X1 U603 ( .A(n2149), .B(n2148), .Y(n894) );
  XOR2X1 U604 ( .A(n2152), .B(n2151), .Y(n895) );
  NAND21X1 U605 ( .B(n1978), .A(n769), .Y(n2104) );
  NAND3X1 U606 ( .A(n2269), .B(n2385), .C(n1623), .Y(n584) );
  INVX1 U607 ( .A(n1496), .Y(n427) );
  INVX1 U608 ( .A(n1414), .Y(n1886) );
  NAND3X1 U609 ( .A(n2424), .B(n2396), .C(n2253), .Y(n1011) );
  INVX1 U610 ( .A(n1690), .Y(n2267) );
  INVX1 U611 ( .A(n829), .Y(n830) );
  NAND4X1 U612 ( .A(n796), .B(n797), .C(n2272), .D(n798), .Y(n807) );
  NAND3X1 U613 ( .A(n2447), .B(n2432), .C(n2436), .Y(n2089) );
  INVX1 U614 ( .A(n1653), .Y(n591) );
  INVX1 U615 ( .A(n1623), .Y(n2426) );
  INVX1 U616 ( .A(n809), .Y(n2381) );
  INVX1 U617 ( .A(n956), .Y(n2382) );
  NAND21X1 U618 ( .B(n2151), .A(n238), .Y(n2167) );
  NAND21X1 U619 ( .B(n2148), .A(n239), .Y(n2161) );
  NAND21X1 U620 ( .B(n2149), .A(n238), .Y(n2166) );
  NAND32X1 U621 ( .B(n621), .C(n2158), .A(n2423), .Y(n1578) );
  INVX1 U622 ( .A(n743), .Y(n621) );
  NAND21X1 U623 ( .B(n768), .A(n769), .Y(n766) );
  NOR2X1 U624 ( .A(n901), .B(n2428), .Y(n794) );
  AND2X1 U625 ( .A(n240), .B(n891), .Y(N12472) );
  NAND2X1 U626 ( .A(n2394), .B(n2185), .Y(n742) );
  NOR31X1 U627 ( .C(n796), .A(n794), .B(n795), .Y(n608) );
  INVX1 U628 ( .A(n2338), .Y(n411) );
  INVX1 U629 ( .A(n1409), .Y(n2229) );
  NOR3XL U630 ( .A(n808), .B(n794), .C(n795), .Y(n756) );
  AND2X1 U631 ( .A(n240), .B(n829), .Y(N12469) );
  INVX1 U632 ( .A(n2039), .Y(n2394) );
  NAND2X1 U633 ( .A(n2039), .B(n772), .Y(n2043) );
  NAND2X1 U634 ( .A(n2433), .B(n2431), .Y(n2112) );
  NAND21X1 U635 ( .B(n1658), .A(n1659), .Y(n1688) );
  NOR2X1 U636 ( .A(n1014), .B(n2428), .Y(n795) );
  INVX1 U637 ( .A(n704), .Y(n2239) );
  INVX1 U638 ( .A(n1533), .Y(n2249) );
  INVX1 U639 ( .A(n2067), .Y(n2231) );
  INVX1 U640 ( .A(n2066), .Y(n1348) );
  NAND21X1 U641 ( .B(n1347), .A(n239), .Y(n2066) );
  NAND2X1 U642 ( .A(n1227), .B(n148), .Y(n1120) );
  NAND2X1 U643 ( .A(n1227), .B(n149), .Y(n1114) );
  NAND2X1 U644 ( .A(n1227), .B(n165), .Y(n1122) );
  NAND2X1 U645 ( .A(n1227), .B(n125), .Y(n1116) );
  NAND2X1 U646 ( .A(n1227), .B(n104), .Y(n1124) );
  NAND2X1 U647 ( .A(n1227), .B(n124), .Y(n1118) );
  NAND2X1 U648 ( .A(n1227), .B(n105), .Y(n1105) );
  NOR2X1 U649 ( .A(n2232), .B(n691), .Y(n781) );
  NOR3XL U650 ( .A(n974), .B(n260), .C(n2437), .Y(n691) );
  INVX1 U651 ( .A(n690), .Y(n2345) );
  OAI22X1 U652 ( .A(n672), .B(n114), .C(n2299), .D(n139), .Y(N12550) );
  OAI22X1 U653 ( .A(n672), .B(n94), .C(n2299), .D(n155), .Y(N12514) );
  OAI22X1 U654 ( .A(n672), .B(n92), .C(n2299), .D(n115), .Y(N12541) );
  OAI22X1 U655 ( .A(n672), .B(n138), .C(n2299), .D(n95), .Y(N12505) );
  OAI22X1 U656 ( .A(n672), .B(n136), .C(n2299), .D(n85), .Y(N12532) );
  OAI22X1 U657 ( .A(n672), .B(n84), .C(n2299), .D(n70), .Y(N12496) );
  OAI22X1 U658 ( .A(n672), .B(n112), .C(n2299), .D(n68), .Y(N12559) );
  OAI22X1 U659 ( .A(n672), .B(n82), .C(n2299), .D(n63), .Y(N12523) );
  INVX1 U660 ( .A(n2276), .Y(n2214) );
  INVX1 U661 ( .A(n2278), .Y(n2221) );
  INVX1 U662 ( .A(n2277), .Y(n2220) );
  INVX1 U663 ( .A(n1236), .Y(n2400) );
  INVX1 U664 ( .A(n2280), .Y(n2176) );
  INVX1 U665 ( .A(n2279), .Y(n2191) );
  INVX1 U666 ( .A(n2147), .Y(n2421) );
  INVX1 U667 ( .A(n765), .Y(n2207) );
  INVX1 U668 ( .A(n2283), .Y(n2177) );
  NAND21X1 U669 ( .B(n2162), .A(memdatai[1]), .Y(n595) );
  NAND21X1 U670 ( .B(n247), .A(memdatai[0]), .Y(n467) );
  NAND21X1 U671 ( .B(n245), .A(memdatai[2]), .Y(n466) );
  NAND21X1 U672 ( .B(n634), .A(n237), .Y(n1339) );
  OR2X1 U673 ( .A(n245), .B(n2052), .Y(n2037) );
  NAND21X1 U674 ( .B(n248), .A(n2050), .Y(n2047) );
  NAND43X1 U675 ( .B(n1563), .C(n1587), .D(n248), .A(n1562), .Y(n586) );
  NOR3XL U676 ( .A(n690), .B(n691), .C(n692), .Y(n685) );
  NAND21X1 U677 ( .B(n246), .A(n2263), .Y(n1079) );
  INVX1 U678 ( .A(n1369), .Y(n2237) );
  AO21X1 U679 ( .B(n244), .C(n2169), .A(n295), .Y(N12698) );
  INVX1 U680 ( .A(n1077), .Y(n2169) );
  AO21X1 U681 ( .B(n244), .C(n2170), .A(n295), .Y(N12697) );
  INVX1 U682 ( .A(n1078), .Y(n2170) );
  AO21X1 U683 ( .B(n244), .C(n2171), .A(n295), .Y(N12699) );
  INVX1 U684 ( .A(n1076), .Y(n2171) );
  AO21X1 U685 ( .B(n104), .C(n249), .A(n294), .Y(N12493) );
  AO21X1 U686 ( .B(n165), .C(n244), .A(n295), .Y(N12502) );
  AO21X1 U687 ( .B(n148), .C(n244), .A(n294), .Y(N12511) );
  AO21X1 U688 ( .B(n124), .C(n249), .A(n294), .Y(N12520) );
  AO21X1 U689 ( .B(n125), .C(n249), .A(n295), .Y(N12529) );
  AO21X1 U690 ( .B(n149), .C(n244), .A(n294), .Y(N12538) );
  AO21X1 U691 ( .B(n105), .C(n249), .A(n295), .Y(N12556) );
  AND3X1 U692 ( .A(n2179), .B(n243), .C(n2172), .Y(N10575) );
  AND3X1 U693 ( .A(n239), .B(n2184), .C(n2394), .Y(N10577) );
  AND3X1 U694 ( .A(n240), .B(n746), .C(n2379), .Y(N10589) );
  INVX1 U695 ( .A(n587), .Y(n1577) );
  OAI21X1 U696 ( .B(n2143), .C(n852), .A(n296), .Y(N13122) );
  OAI21X1 U697 ( .B(n2441), .C(n852), .A(n296), .Y(N13131) );
  OAI21X1 U698 ( .B(n842), .C(n852), .A(n296), .Y(N13149) );
  OAI21X1 U699 ( .B(n2143), .C(n843), .A(n290), .Y(N13266) );
  OAI21X1 U700 ( .B(n2441), .C(n843), .A(n290), .Y(N13275) );
  OAI21X1 U701 ( .B(n842), .C(n843), .A(n298), .Y(N13293) );
  OAI21X1 U702 ( .B(n1099), .C(n1101), .A(n288), .Y(N12637) );
  AND2X1 U703 ( .A(n2204), .B(n11), .Y(N583) );
  AND2X1 U704 ( .A(n2168), .B(n2379), .Y(N10564) );
  AND2X1 U705 ( .A(n1701), .B(n243), .Y(N584) );
  AND2X1 U706 ( .A(n207), .B(n243), .Y(N10578) );
  NOR3XL U707 ( .A(n2034), .B(n2425), .C(n2389), .Y(N10581) );
  NOR3XL U708 ( .A(n2034), .B(n2425), .C(n773), .Y(N10565) );
  NAND2X1 U709 ( .A(n287), .B(n2278), .Y(N12690) );
  NAND2X1 U710 ( .A(n287), .B(n2276), .Y(N12692) );
  NAND2X1 U711 ( .A(n287), .B(n2277), .Y(N12691) );
  INVX1 U712 ( .A(n2163), .Y(n2168) );
  NAND21X1 U713 ( .B(n2437), .A(n237), .Y(n2163) );
  NOR2X1 U714 ( .A(n2389), .B(n2037), .Y(N10582) );
  NOR2X1 U715 ( .A(n773), .B(n2037), .Y(N10583) );
  NAND3X1 U716 ( .A(n585), .B(n288), .C(n586), .Y(N685) );
  NOR21XL U717 ( .B(n250), .A(n2042), .Y(N10574) );
  AOI21X1 U718 ( .B(n2179), .C(n2043), .A(n2044), .Y(n2042) );
  AND2X1 U719 ( .A(n240), .B(n1693), .Y(N11481) );
  AND2X1 U720 ( .A(n241), .B(n198), .Y(N11480) );
  AND2X1 U721 ( .A(n241), .B(n1692), .Y(N11478) );
  AND2X1 U722 ( .A(n242), .B(n197), .Y(N11479) );
  AND2X1 U723 ( .A(n241), .B(n2377), .Y(N12709) );
  NOR21XL U724 ( .B(n242), .A(n1075), .Y(N12700) );
  NOR21XL U725 ( .B(n242), .A(n1074), .Y(N12701) );
  NOR21XL U726 ( .B(n242), .A(n1072), .Y(N12703) );
  NOR21XL U727 ( .B(n242), .A(n1073), .Y(N12702) );
  NOR21XL U728 ( .B(n240), .A(n1004), .Y(N10585) );
  AND2X1 U729 ( .A(n241), .B(n502), .Y(N12704) );
  AND2X1 U730 ( .A(n241), .B(n1655), .Y(N11486) );
  OAI22X1 U731 ( .A(n1531), .B(n2451), .C(n2326), .D(n1532), .Y(n1528) );
  INVX1 U732 ( .A(n1587), .Y(n589) );
  INVX1 U733 ( .A(n728), .Y(n2056) );
  INVX1 U734 ( .A(n1859), .Y(n2055) );
  INVX1 U735 ( .A(n1134), .Y(n2302) );
  AOI21X1 U736 ( .B(n2459), .C(n2302), .A(n1170), .Y(n1157) );
  AOI21X1 U737 ( .B(n1192), .C(n2302), .A(n1170), .Y(n1180) );
  NAND2X1 U738 ( .A(n2291), .B(n2386), .Y(n1374) );
  INVX1 U739 ( .A(n1170), .Y(n2303) );
  AOI221XL U740 ( .A(n2454), .B(n48), .C(n2452), .D(n43), .E(n1170), .Y(n1259)
         );
  MUX2X1 U741 ( .D0(n1436), .D1(n2229), .S(n204), .Y(n1438) );
  INVX1 U742 ( .A(n42), .Y(n2305) );
  INVX1 U743 ( .A(n1739), .Y(n2218) );
  INVX1 U744 ( .A(n2178), .Y(n1766) );
  OAI21X1 U745 ( .B(n1169), .C(n1132), .A(n1157), .Y(n1168) );
  INVX1 U746 ( .A(n1738), .Y(n2219) );
  AOI22AXL U747 ( .A(n659), .B(n2228), .D(n659), .C(n1409), .Y(n1510) );
  AOI22AXL U748 ( .A(n697), .B(n2228), .D(n697), .C(n1409), .Y(n1470) );
  INVX1 U749 ( .A(n2291), .Y(n2206) );
  NOR4XL U750 ( .A(multemp2[9]), .B(multemp2[8]), .C(multemp2[7]), .D(
        multemp2[6]), .Y(n1025) );
  INVX1 U751 ( .A(multemp2[9]), .Y(n2290) );
  OAI21X1 U752 ( .B(n1130), .C(n153), .A(n1300), .Y(n1309) );
  NOR2X1 U753 ( .A(n43), .B(n48), .Y(n1209) );
  INVX1 U754 ( .A(n1255), .Y(n2455) );
  NOR4XL U755 ( .A(multemp2[5]), .B(multemp2[4]), .C(multemp2[3]), .D(
        multemp2[2]), .Y(n1024) );
  INVX1 U756 ( .A(n1177), .Y(n651) );
  INVX1 U757 ( .A(n1257), .Y(n2452) );
  NAND31X1 U758 ( .C(n1010), .A(n584), .B(n1011), .Y(n1009) );
  AND2X1 U759 ( .A(n444), .B(n2349), .Y(n999) );
  INVX1 U760 ( .A(n986), .Y(n2347) );
  INVX1 U761 ( .A(n983), .Y(n2348) );
  NOR2X1 U762 ( .A(n2272), .B(n259), .Y(n906) );
  INVX1 U763 ( .A(n912), .Y(n1384) );
  INVX1 U764 ( .A(n913), .Y(n2344) );
  NAND2X1 U765 ( .A(n952), .B(n2359), .Y(n939) );
  INVX1 U766 ( .A(rst), .Y(n297) );
  NOR2X1 U767 ( .A(n2394), .B(n780), .Y(n2107) );
  INVX1 U768 ( .A(n1001), .Y(n2378) );
  AOI21BBXL U769 ( .B(n1735), .C(n2251), .A(n2447), .Y(n2044) );
  AOI211X1 U770 ( .C(n2111), .D(n1634), .A(n2044), .B(n207), .Y(n2110) );
  OAI21X1 U771 ( .B(n2425), .C(n2428), .A(n2052), .Y(n2111) );
  INVX1 U772 ( .A(n911), .Y(n1385) );
  INVX1 U773 ( .A(n2041), .Y(n2172) );
  NOR21XL U774 ( .B(n2045), .A(n963), .Y(n2041) );
  AOI21X1 U775 ( .B(n1625), .C(n746), .A(n808), .Y(n2119) );
  INVX1 U776 ( .A(n1192), .Y(n2456) );
  NOR2X1 U777 ( .A(n2043), .B(n2048), .Y(n2040) );
  NAND2X1 U778 ( .A(n287), .B(n2399), .Y(n869) );
  INVX1 U779 ( .A(n298), .Y(n291) );
  INVX1 U780 ( .A(rst), .Y(n298) );
  INVX1 U781 ( .A(rst), .Y(n296) );
  INVX1 U782 ( .A(n1015), .Y(n2266) );
  MUX2X1 U783 ( .D0(memwr), .D1(n1700), .S(n284), .Y(memwr_comb) );
  AND2X1 U784 ( .A(n488), .B(n11), .Y(n1703) );
  MUX2X2 U785 ( .D0(n495), .D1(n857), .S(n1659), .Y(n1657) );
  OAI22X1 U786 ( .A(n51), .B(n2338), .C(n2469), .D(n2380), .Y(n490) );
  AO21X1 U787 ( .B(pc_i[1]), .C(n2239), .A(n455), .Y(n491) );
  NAND21X1 U788 ( .B(mempsack), .A(n1621), .Y(n300) );
  INVX1 U789 ( .A(n1624), .Y(n302) );
  NAND21X1 U790 ( .B(memack), .A(n1619), .Y(n301) );
  INVX1 U791 ( .A(pc_i[9]), .Y(n487) );
  NAND21X1 U792 ( .B(n588), .A(n1575), .Y(n615) );
  INVX1 U793 ( .A(sfrdatai[5]), .Y(n1933) );
  NAND21X1 U794 ( .B(n374), .A(n373), .Y(n379) );
  NAND31X1 U795 ( .C(n473), .A(n372), .B(n655), .Y(n373) );
  INVX1 U796 ( .A(sfrdatai[0]), .Y(n787) );
  OA222X1 U797 ( .A(n2495), .B(n492), .C(n921), .D(n826), .E(n951), .F(n1739), 
        .Y(n429) );
  OA22X1 U798 ( .A(n1434), .B(n825), .C(n2291), .D(n2329), .Y(n430) );
  OAI211XL U799 ( .C(n1738), .D(n775), .A(n494), .B(n493), .Y(n857) );
  OA22X1 U800 ( .A(n2469), .B(n1434), .C(n2291), .D(n2330), .Y(n494) );
  OA222X1 U801 ( .A(n2494), .B(n492), .C(n921), .D(n791), .E(n944), .F(n1739), 
        .Y(n493) );
  AOI21BBXL U802 ( .B(cpu_resume), .C(irq), .A(n291), .Y(N13379) );
  MUX2XL U803 ( .D0(n235), .D1(n1728), .S(n15), .Y(memaddr_comb[10]) );
  AO21X1 U804 ( .B(n612), .C(n610), .A(n609), .Y(n619) );
  OA222X1 U805 ( .A(n743), .B(n2245), .C(n260), .D(n608), .E(n2272), .F(n2238), 
        .Y(n609) );
  AOI21X1 U806 ( .B(n803), .C(n807), .A(n607), .Y(n610) );
  AOI21X1 U807 ( .B(n801), .C(n795), .A(n794), .Y(n612) );
  NAND21X1 U808 ( .B(n793), .A(n792), .Y(n1714) );
  OA2222XL U809 ( .A(n781), .B(n791), .C(n2469), .D(n1371), .E(n944), .F(n1369), .G(n2345), .H(n2494), .Y(n792) );
  AO2222XL U810 ( .A(alu_out[1]), .B(n1407), .C(n220), .D(n1187), .E(n1341), 
        .F(pc_o[1]), .G(n1334), .H(pc_i[1]), .Y(n793) );
  AO21X1 U811 ( .B(n130), .C(n2273), .A(n404), .Y(n408) );
  OAI31XL U812 ( .A(n1603), .B(n2489), .C(n1604), .D(n403), .Y(n404) );
  INVX1 U813 ( .A(n628), .Y(n1334) );
  NAND32X1 U814 ( .B(n692), .C(n862), .A(n627), .Y(n628) );
  INVX1 U815 ( .A(N13343), .Y(n2274) );
  NAND2X1 U816 ( .A(n810), .B(n811), .Y(n803) );
  NOR4XL U817 ( .A(n816), .B(n817), .C(n818), .D(n2313), .Y(n810) );
  NOR4XL U818 ( .A(n812), .B(n813), .C(n814), .D(n815), .Y(n811) );
  NOR2XL U819 ( .A(n1712), .B(n1418), .Y(n188) );
  NOR2XL U820 ( .A(n1712), .B(n1412), .Y(n195) );
  MUX2X1 U821 ( .D0(n235), .D1(n1410), .S(n89), .Y(N12851) );
  EORX1 U822 ( .A(n1492), .B(n1491), .C(n1493), .D(n1435), .Y(n196) );
  XNOR2XL U823 ( .A(n1415), .B(n1416), .Y(n1413) );
  XNOR2XL U824 ( .A(n2202), .B(n1417), .Y(n1416) );
  AOI22X1 U825 ( .A(n2202), .B(n1419), .C(n1420), .D(n1421), .Y(n1415) );
  OAI222XL U826 ( .A(n456), .B(n1691), .C(n2148), .D(n1688), .E(n2195), .F(
        waitstaten), .Y(ramdatao_comb[7]) );
  OAI22X1 U827 ( .A(n1956), .B(n1955), .C(n1435), .D(n196), .Y(n1421) );
  AND2X1 U828 ( .A(n196), .B(n1435), .Y(n1956) );
  OAI22X1 U829 ( .A(n1435), .B(n3), .C(n1741), .D(n1740), .Y(n1523) );
  AND2X1 U830 ( .A(n3), .B(n1435), .Y(n1741) );
  OAI221X1 U831 ( .A(n170), .B(n1502), .C(n1501), .D(n1697), .E(n444), .Y(
        n1655) );
  AOI221XL U832 ( .A(n965), .B(n1775), .C(n758), .D(n147), .E(n1776), .Y(n1502) );
  INVX1 U833 ( .A(n1611), .Y(n1501) );
  OAI211X1 U834 ( .C(n2185), .D(n1727), .A(n2423), .B(n2387), .Y(n1776) );
  INVX1 U835 ( .A(n812), .Y(n2329) );
  AND2XL U836 ( .A(n180), .B(n1435), .Y(n1461) );
  AOI22X1 U837 ( .A(N11555), .B(n1456), .C(n1457), .D(n2375), .Y(n1454) );
  NAND2X1 U838 ( .A(n1458), .B(n2404), .Y(n1456) );
  NAND21X1 U839 ( .B(n483), .A(n1495), .Y(n1705) );
  AOI21BBXL U840 ( .B(n1599), .C(n1600), .A(n1601), .Y(n575) );
  AOI21X1 U841 ( .B(n1600), .C(n1599), .A(n1602), .Y(n1601) );
  INVX1 U842 ( .A(n1376), .Y(n2313) );
  XNOR2XL U843 ( .A(n1398), .B(n1401), .Y(n1452) );
  OAI22X1 U844 ( .A(n1398), .B(n1399), .C(n1400), .D(n1401), .Y(n1035) );
  AND2X1 U845 ( .A(n1399), .B(n1398), .Y(n1400) );
  NOR2X1 U846 ( .A(n2483), .B(n1681), .Y(n1367) );
  OAI21X1 U847 ( .B(n1397), .C(n1035), .A(n1070), .Y(n1069) );
  OAI21X1 U848 ( .B(n1367), .C(n2469), .A(n2472), .Y(n578) );
  INVX1 U849 ( .A(n1575), .Y(n1590) );
  NAND2X1 U850 ( .A(n1397), .B(n1035), .Y(n1070) );
  INVX1 U851 ( .A(n1598), .Y(n2483) );
  INVX1 U852 ( .A(n879), .Y(n435) );
  INVX1 U853 ( .A(N11555), .Y(n2439) );
  XNOR2XL U854 ( .A(n1365), .B(n2477), .Y(n576) );
  XNOR2XL U855 ( .A(n1365), .B(n2478), .Y(n1600) );
  XNOR2XL U856 ( .A(n2439), .B(n1458), .Y(n1518) );
  XOR2X1 U857 ( .A(n1479), .B(n1453), .Y(n1478) );
  AOI21X1 U858 ( .B(n2375), .C(n1457), .A(n1484), .Y(n1479) );
  AOI21X1 U859 ( .B(n2404), .C(n1458), .A(n2439), .Y(n1484) );
  AO222X1 U860 ( .A(n1164), .B(n2249), .C(n817), .D(n2056), .E(n1471), .F(
        n1414), .Y(n710) );
  XNOR2XL U861 ( .A(n196), .B(n1488), .Y(n1471) );
  XOR2X1 U862 ( .A(n1955), .B(n2202), .Y(n1488) );
  NOR3XL U863 ( .A(n1742), .B(n2362), .C(memdatai[7]), .Y(n1852) );
  AOI22X1 U864 ( .A(n1429), .B(n1414), .C(n2249), .D(n1153), .Y(n1427) );
  XOR2X1 U865 ( .A(n1421), .B(n1431), .Y(n1429) );
  XNOR2XL U866 ( .A(n1420), .B(n2202), .Y(n1431) );
  OAI222XL U867 ( .A(n1686), .B(n1691), .C(n1666), .D(n1688), .E(n2212), .F(
        waitstaten), .Y(ramdatao_comb[5]) );
  OAI222XL U868 ( .A(n1687), .B(n1691), .C(n2149), .D(n1688), .E(n2208), .F(
        waitstaten), .Y(ramdatao_comb[6]) );
  OAI222XL U869 ( .A(n883), .B(n448), .C(n1373), .D(n447), .E(n1929), .F(n826), 
        .Y(n1692) );
  OAI21X1 U870 ( .B(n1068), .C(n1069), .A(n1070), .Y(n1036) );
  AO222X1 U871 ( .A(memdatai[4]), .B(n1852), .C(n881), .D(n1778), .E(n2362), 
        .F(memdatai[1]), .Y(n197) );
  AO222X1 U872 ( .A(memdatai[5]), .B(n1852), .C(n875), .D(n1778), .E(n2362), 
        .F(memdatai[2]), .Y(n198) );
  INVX1 U873 ( .A(n712), .Y(n1686) );
  NAND41X1 U874 ( .D(n710), .A(n709), .B(n708), .C(n707), .Y(n712) );
  OA222X1 U875 ( .A(n49), .B(n945), .C(n704), .D(n703), .E(n2380), .F(n702), 
        .Y(n708) );
  OA222X1 U876 ( .A(n2386), .B(n1954), .C(n1531), .D(n705), .E(n46), .F(n2338), 
        .Y(n707) );
  INVX1 U877 ( .A(n928), .Y(n2215) );
  NAND21X1 U878 ( .B(n2429), .A(n39), .Y(n974) );
  NOR2X1 U879 ( .A(n2450), .B(n2243), .Y(n2050) );
  OAI211X1 U880 ( .C(n2367), .D(n2335), .A(n1673), .B(n1672), .Y(n1669) );
  NOR3XL U881 ( .A(n1677), .B(n2355), .C(n1603), .Y(n1683) );
  OAI222XL U882 ( .A(n1665), .B(n1691), .C(n2151), .D(n1688), .E(n2216), .F(
        waitstaten), .Y(ramdatao_comb[4]) );
  NOR2X1 U883 ( .A(n1669), .B(n2367), .Y(n1362) );
  AND2X1 U884 ( .A(n1026), .B(n1353), .Y(n1045) );
  INVX1 U885 ( .A(n868), .Y(n2198) );
  NAND32X1 U886 ( .B(n862), .C(n861), .A(n860), .Y(n868) );
  NOR2X1 U887 ( .A(n1392), .B(n2264), .Y(n1044) );
  INVX1 U888 ( .A(n1393), .Y(n2264) );
  INVX1 U889 ( .A(n1737), .Y(n2236) );
  NOR2X1 U890 ( .A(n126), .B(n444), .Y(retiinstr) );
  INVX1 U891 ( .A(n1005), .Y(n2429) );
  INVX1 U892 ( .A(n668), .Y(n1665) );
  NAND41X1 U893 ( .D(n667), .A(n666), .B(n663), .C(n662), .Y(n668) );
  OA222X1 U894 ( .A(n55), .B(n945), .C(n704), .D(n649), .E(n2380), .F(n669), 
        .Y(n666) );
  OA222X1 U895 ( .A(n2386), .B(n654), .C(n728), .D(n652), .E(n1533), .F(n651), 
        .Y(n663) );
  NOR21XL U896 ( .B(n1672), .A(n1673), .Y(n1363) );
  AO222X1 U897 ( .A(n351), .B(n350), .C(n349), .D(n348), .E(n465), .F(n2216), 
        .Y(n928) );
  AND4X1 U898 ( .A(n1894), .B(n1895), .C(n1892), .D(n1893), .Y(n350) );
  AND4X1 U899 ( .A(n1902), .B(n1903), .C(n1900), .D(n1901), .Y(n348) );
  AND4X1 U900 ( .A(n1890), .B(n1891), .C(n1888), .D(n1889), .Y(n351) );
  NAND31X1 U901 ( .C(n1505), .A(n199), .B(irq), .Y(n1587) );
  NAND3X1 U902 ( .A(n873), .B(n1653), .C(n579), .Y(n199) );
  NAND32X1 U903 ( .B(n462), .C(n461), .A(n460), .Y(n813) );
  OAI22X1 U904 ( .A(n1486), .B(n2475), .C(n1393), .D(n2199), .Y(n462) );
  OA2222XL U905 ( .A(n2478), .B(n2351), .C(n1593), .D(n2469), .E(n1595), .F(
        n1450), .G(n2406), .H(n459), .Y(n460) );
  OAI221X1 U906 ( .A(N13343), .B(n458), .C(n2334), .D(n2473), .E(n457), .Y(
        n461) );
  AO222X1 U907 ( .A(n2056), .B(n2313), .C(n2055), .D(n2054), .E(ramdatai[7]), 
        .F(n2230), .Y(n1382) );
  AO21X1 U908 ( .B(n2053), .C(n2038), .A(n2035), .Y(n2054) );
  GEN2XL U909 ( .D(n2228), .E(n1995), .C(n1994), .B(n212), .A(n1993), .Y(n2035) );
  NOR2X1 U910 ( .A(n2418), .B(n33), .Y(n758) );
  MUX2AXL U911 ( .D0(n1526), .D1(n891), .S(n1659), .Y(n1664) );
  NOR4XL U912 ( .A(n1527), .B(n1528), .C(n1529), .D(n1530), .Y(n1526) );
  OAI22X1 U913 ( .A(n2380), .B(n2438), .C(n945), .D(n2465), .Y(n1530) );
  ENOX1 U914 ( .A(n2338), .B(n2453), .C(n2239), .D(pc_i[3]), .Y(n1529) );
  NOR2X1 U915 ( .A(n2243), .B(n2448), .Y(n745) );
  OAI221X1 U916 ( .A(n2405), .B(n1780), .C(n2361), .D(n1037), .E(n1876), .Y(
        n884) );
  OA222X1 U917 ( .A(n2286), .B(n1781), .C(n1074), .D(n2340), .E(n928), .F(
        n1782), .Y(n1876) );
  INVX1 U918 ( .A(n1356), .Y(n2331) );
  OAI222XL U919 ( .A(n1661), .B(n1688), .C(n1660), .D(n1691), .E(n2192), .F(
        waitstaten), .Y(ramdatao_comb[2]) );
  NOR2X1 U920 ( .A(n1033), .B(n1363), .Y(n1395) );
  NOR2X1 U921 ( .A(n874), .B(n875), .Y(n873) );
  AOI33X1 U922 ( .A(n876), .B(n2310), .C(n877), .D(n878), .E(n879), .F(n880), 
        .Y(n874) );
  INVX1 U923 ( .A(n881), .Y(n2310) );
  OAI21X1 U924 ( .B(n876), .C(n881), .A(n882), .Y(n878) );
  NAND3X1 U925 ( .A(n2442), .B(n2444), .C(n2443), .Y(n842) );
  OAI222XL U926 ( .A(n1886), .B(n1885), .C(n1877), .D(n1859), .E(n1533), .F(
        n205), .Y(n1527) );
  GEN2XL U927 ( .D(n1767), .E(n2228), .C(n1994), .B(n1766), .A(n1754), .Y(
        n1857) );
  AOI21X1 U928 ( .B(n1775), .C(n2184), .A(n758), .Y(n2028) );
  INVX1 U929 ( .A(n2430), .Y(n2184) );
  INVX1 U930 ( .A(n263), .Y(n259) );
  INVX1 U931 ( .A(n2182), .Y(n263) );
  NAND2X1 U932 ( .A(n1037), .B(n1787), .Y(n1799) );
  NAND2X1 U933 ( .A(n1787), .B(n2357), .Y(n1817) );
  INVX1 U934 ( .A(n579), .Y(n1509) );
  INVX1 U935 ( .A(n862), .Y(n636) );
  OAI22X1 U936 ( .A(n1199), .B(n1533), .C(n1886), .D(n1463), .Y(n1466) );
  XOR3X1 U937 ( .A(n2202), .B(n3), .C(n1740), .Y(n1463) );
  OAI22X1 U938 ( .A(n456), .B(n1490), .C(n1489), .D(n2161), .Y(N11505) );
  NOR3XL U939 ( .A(n885), .B(n880), .C(n883), .Y(n877) );
  XNOR2XL U940 ( .A(n879), .B(n884), .Y(n885) );
  INVX1 U941 ( .A(n1775), .Y(n2418) );
  NAND3X1 U942 ( .A(n1044), .B(n1353), .C(n1043), .Y(n1031) );
  AOI31X1 U943 ( .A(n1408), .B(n211), .C(n1992), .D(n1995), .Y(n1993) );
  AOI22AXL U944 ( .A(n212), .B(n1409), .D(n212), .C(n2228), .Y(n1408) );
  INVX1 U945 ( .A(n2027), .Y(n2417) );
  INVX1 U946 ( .A(n1458), .Y(n2375) );
  INVX1 U947 ( .A(n908), .Y(n2197) );
  NOR32XL U948 ( .B(n840), .C(n1668), .A(n1669), .Y(n1349) );
  GEN2XL U949 ( .D(n2314), .E(n1828), .C(n1824), .B(n2342), .A(n1826), .Y(
        n1827) );
  INVX1 U950 ( .A(n1825), .Y(n2314) );
  OA2222XL U951 ( .A(n2189), .B(n1780), .C(n2318), .D(n1781), .E(n923), .F(
        n1782), .G(n1073), .H(n2340), .Y(n876) );
  OAI21X1 U952 ( .B(n1603), .C(n1604), .A(n1049), .Y(n1032) );
  AO222X1 U953 ( .A(n335), .B(n334), .C(n333), .D(n332), .E(n465), .F(n2203), 
        .Y(n951) );
  AND4X1 U954 ( .A(n2002), .B(n2003), .C(n2000), .D(n2001), .Y(n334) );
  AND4X1 U955 ( .A(n2023), .B(n2024), .C(n2021), .D(n2022), .Y(n332) );
  AND4X1 U956 ( .A(n1998), .B(n1999), .C(n1996), .D(n1997), .Y(n335) );
  AO222X1 U957 ( .A(n471), .B(n470), .C(n469), .D(n468), .E(n465), .F(n2199), 
        .Y(n944) );
  AND4X1 U958 ( .A(n1964), .B(n1965), .C(n1962), .D(n1963), .Y(n470) );
  AND4X1 U959 ( .A(n1972), .B(n1973), .C(n1970), .D(n1971), .Y(n468) );
  AND4X1 U960 ( .A(n1960), .B(n1961), .C(n1958), .D(n1959), .Y(n471) );
  AO222X1 U961 ( .A(n342), .B(n341), .C(n340), .D(n339), .E(n465), .F(n2192), 
        .Y(n938) );
  AND4X1 U962 ( .A(n1941), .B(n1942), .C(n1939), .D(n1940), .Y(n341) );
  AND4X1 U963 ( .A(n1949), .B(n1950), .C(n1947), .D(n1948), .Y(n339) );
  AND4X1 U964 ( .A(n1937), .B(n1938), .C(n1935), .D(n1936), .Y(n342) );
  MUX2X1 U965 ( .D0(n2216), .D1(n2356), .S(n1015), .Y(n1037) );
  NAND21X1 U966 ( .B(n844), .A(n1222), .Y(n1829) );
  AND2X1 U967 ( .A(n1570), .B(n1587), .Y(n1545) );
  NOR21XL U968 ( .B(n1905), .A(N12773), .Y(n1854) );
  OA2222XL U969 ( .A(n2340), .B(n1072), .C(n918), .D(n1782), .E(n1780), .F(
        n2188), .G(n2319), .H(n1781), .Y(n880) );
  AO222X1 U970 ( .A(n347), .B(n346), .C(n345), .D(n344), .E(n465), .F(n2212), 
        .Y(n923) );
  AND4X1 U971 ( .A(n1866), .B(n1867), .C(n1864), .D(n1865), .Y(n346) );
  AND4X1 U972 ( .A(n1874), .B(n1875), .C(n1872), .D(n1873), .Y(n344) );
  AND4X1 U973 ( .A(n1862), .B(n1863), .C(n1860), .D(n1861), .Y(n347) );
  AO21X1 U974 ( .B(n1621), .C(n2154), .A(n2153), .Y(n1637) );
  INVX1 U975 ( .A(n1544), .Y(n1570) );
  NOR21XL U976 ( .B(n1928), .A(N12772), .Y(n1905) );
  NOR21XL U977 ( .B(n1952), .A(N12771), .Y(n1928) );
  OAI221X1 U978 ( .A(n2442), .B(n1780), .C(n2361), .D(n69), .E(n1953), .Y(n881) );
  OA222X1 U979 ( .A(n2317), .B(n1781), .C(n1077), .D(n2340), .E(n944), .F(
        n1782), .Y(n1953) );
  AND3X1 U980 ( .A(n2189), .B(n2236), .C(n2188), .Y(n1102) );
  AOI222XL U981 ( .A(n2339), .B(n1854), .C(n1904), .D(N12773), .E(N12805), .F(
        n1822), .Y(n1074) );
  OAI21X1 U982 ( .B(n1905), .C(n1824), .A(n2342), .Y(n1904) );
  AOI222XL U983 ( .A(n2339), .B(n1952), .C(n1974), .D(N12770), .E(N12802), .F(
        n1822), .Y(n1077) );
  OAI21X1 U984 ( .B(n1975), .C(n1824), .A(n2342), .Y(n1974) );
  AOI222XL U985 ( .A(n2339), .B(n1905), .C(n1927), .D(N12772), .E(N12804), .F(
        n1822), .Y(n1075) );
  OAI21X1 U986 ( .B(n1928), .C(n1824), .A(n2342), .Y(n1927) );
  AND2X1 U987 ( .A(n1102), .B(n850), .Y(n1222) );
  NAND32X1 U988 ( .B(n397), .C(n316), .A(n2380), .Y(n1689) );
  NOR2X1 U989 ( .A(n32), .B(n1775), .Y(n2020) );
  NAND3X1 U990 ( .A(n1102), .B(n853), .C(n855), .Y(n476) );
  NOR3XL U991 ( .A(n1822), .B(n690), .C(n1986), .Y(n1850) );
  NAND2X1 U992 ( .A(n1752), .B(n2261), .Y(n772) );
  INVX1 U993 ( .A(n1038), .Y(n2377) );
  NAND3X1 U994 ( .A(n1364), .B(n2189), .C(n853), .Y(n1015) );
  AND2X1 U995 ( .A(n970), .B(n774), .Y(n1752) );
  INVX1 U996 ( .A(n1787), .Y(n465) );
  AOI222XL U997 ( .A(n2200), .B(ramdatai[6]), .C(n2201), .D(sfrdatai[6]), .E(
        n2250), .F(n2210), .Y(n1420) );
  INVX1 U998 ( .A(n918), .Y(n2210) );
  NAND2X1 U999 ( .A(n1854), .B(n1855), .Y(n1825) );
  OAI221X1 U1000 ( .A(n2444), .B(n1780), .C(n2361), .D(n33), .E(n1930), .Y(
        n875) );
  OA222X1 U1001 ( .A(n2321), .B(n1781), .C(n1076), .D(n2340), .E(n938), .F(
        n1782), .Y(n1930) );
  NAND3X1 U1002 ( .A(n774), .B(n2261), .C(n1756), .Y(n1757) );
  INVX1 U1003 ( .A(n1975), .Y(n206) );
  INVX1 U1004 ( .A(n1736), .Y(n2437) );
  INVX1 U1005 ( .A(n310), .Y(n311) );
  NAND32X1 U1006 ( .B(n126), .C(n2437), .A(n2256), .Y(n310) );
  NOR3XL U1007 ( .A(n2479), .B(n2367), .C(n2350), .Y(n1361) );
  INVX1 U1008 ( .A(n818), .Y(n2316) );
  INVX1 U1009 ( .A(n1603), .Y(n2354) );
  INVX1 U1010 ( .A(n1457), .Y(n2404) );
  INVX1 U1011 ( .A(n814), .Y(n2327) );
  NOR2X1 U1012 ( .A(n2190), .B(n2417), .Y(n2011) );
  NOR2X1 U1013 ( .A(n2027), .B(n2190), .Y(n2008) );
  NOR2X1 U1014 ( .A(n2419), .B(n1038), .Y(n2009) );
  NOR2X1 U1015 ( .A(n2020), .B(n1038), .Y(n2013) );
  INVX1 U1016 ( .A(n1604), .Y(n2355) );
  OAI22X1 U1017 ( .A(n1687), .B(n1490), .C(n1489), .D(n2166), .Y(N11504) );
  NOR4XL U1018 ( .A(n1824), .B(n1825), .C(n129), .D(n108), .Y(n1823) );
  INVX1 U1019 ( .A(n1332), .Y(n2364) );
  INVX1 U1020 ( .A(n1333), .Y(n2325) );
  NOR2X1 U1021 ( .A(n206), .B(N12770), .Y(n1952) );
  INVX1 U1022 ( .A(n721), .Y(n1368) );
  INVX1 U1023 ( .A(n736), .Y(n1228) );
  INVX1 U1024 ( .A(n731), .Y(n1187) );
  INVX1 U1025 ( .A(n726), .Y(n1126) );
  NAND3X1 U1026 ( .A(n2354), .B(n1604), .C(n1677), .Y(n1049) );
  INVX1 U1027 ( .A(n1359), .Y(n2332) );
  NAND2X1 U1028 ( .A(n1675), .B(n1683), .Y(n1358) );
  NAND4X1 U1029 ( .A(n883), .B(n876), .C(n881), .D(n884), .Y(n882) );
  INVX1 U1030 ( .A(n1663), .Y(n2336) );
  INVX1 U1031 ( .A(n1668), .Y(n2337) );
  INVX1 U1032 ( .A(n1071), .Y(n502) );
  AOI211X1 U1033 ( .C(N12808), .D(n1822), .A(n2308), .B(n1823), .Y(n1071) );
  INVX1 U1034 ( .A(n1827), .Y(n2308) );
  INVX1 U1035 ( .A(n1822), .Y(n2341) );
  NAND32X1 U1036 ( .B(n2434), .C(n1699), .A(n2270), .Y(n945) );
  NAND21X1 U1037 ( .B(n589), .A(n1544), .Y(n593) );
  NAND21X1 U1038 ( .B(n168), .A(n311), .Y(n1533) );
  OR2X1 U1039 ( .A(n126), .B(n1651), .Y(n2389) );
  NAND21X1 U1040 ( .B(n2186), .A(n2106), .Y(n1651) );
  NAND32X1 U1041 ( .B(n248), .C(n1572), .A(n1573), .Y(n1571) );
  AOI21X1 U1042 ( .B(n1393), .C(n1392), .A(n2353), .Y(n1486) );
  GEN2XL U1043 ( .D(n1442), .E(n2228), .C(n1994), .B(n204), .A(n1441), .Y(
        n1467) );
  AND2XL U1044 ( .A(n1858), .B(n1440), .Y(n1441) );
  AOI222XL U1045 ( .A(n1850), .B(n127), .C(N12806), .D(n1822), .E(n2339), .F(
        n1853), .Y(n1073) );
  OAI21X1 U1046 ( .B(n1854), .C(n1855), .A(n1825), .Y(n1853) );
  AOI222XL U1047 ( .A(n2339), .B(n1928), .C(n1951), .D(N12771), .E(N12803), 
        .F(n1822), .Y(n1076) );
  OAI21X1 U1048 ( .B(n1952), .C(n1824), .A(n2342), .Y(n1951) );
  OR2X1 U1049 ( .A(n2162), .B(n200), .Y(n464) );
  AOI21X1 U1050 ( .B(n589), .C(n1544), .A(n588), .Y(n200) );
  AOI222XL U1051 ( .A(n2339), .B(n1975), .C(n1850), .D(n206), .E(N12801), .F(
        n1822), .Y(n1078) );
  GEN2XL U1052 ( .D(n2053), .E(n1440), .C(n730), .B(n2055), .A(n729), .Y(n732)
         );
  OAI22X1 U1053 ( .A(n2491), .B(n2386), .C(n728), .D(n2316), .Y(n729) );
  GEN2XL U1054 ( .D(n727), .E(n2228), .C(n1994), .B(n214), .A(n725), .Y(n730)
         );
  AOI222XL U1055 ( .A(n1850), .B(n129), .C(N12807), .D(n1822), .E(n1851), .F(
        n2339), .Y(n1072) );
  XNOR2XL U1056 ( .A(n129), .B(n1825), .Y(n1851) );
  OA222X1 U1057 ( .A(n700), .B(n699), .C(n697), .D(n696), .E(n2323), .F(n722), 
        .Y(n709) );
  AND3X1 U1058 ( .A(n1470), .B(n211), .C(n689), .Y(n699) );
  INVXL U1059 ( .A(n695), .Y(n700) );
  OA222X1 U1060 ( .A(n661), .B(n660), .C(n659), .D(n658), .E(n2322), .F(n722), 
        .Y(n662) );
  AND3X1 U1061 ( .A(n1510), .B(n211), .C(n655), .Y(n660) );
  NOR2X1 U1062 ( .A(n2243), .B(n2449), .Y(n746) );
  XNOR2XL U1063 ( .A(n1365), .B(n2415), .Y(n1399) );
  XNOR2XL U1064 ( .A(n1365), .B(n2406), .Y(n1455) );
  NOR2X1 U1065 ( .A(n2448), .B(n2186), .Y(n1649) );
  INVX1 U1066 ( .A(n1357), .Y(n459) );
  NOR2X1 U1067 ( .A(n2245), .B(n2423), .Y(n690) );
  NAND2X1 U1068 ( .A(n39), .B(n17), .Y(n805) );
  NAND2X1 U1069 ( .A(n1649), .B(n1723), .Y(n773) );
  NOR3XL U1070 ( .A(n1989), .B(n1982), .C(n1985), .Y(n1984) );
  AND2X1 U1071 ( .A(n510), .B(n287), .Y(N512) );
  INVX1 U1072 ( .A(n1495), .Y(n1573) );
  INVX1 U1073 ( .A(ramdatai[5]), .Y(n1954) );
  INVX1 U1074 ( .A(ramdatai[4]), .Y(n654) );
  OAI32X1 U1075 ( .A(n1608), .B(n483), .C(n1607), .D(n1606), .E(n246), .Y(N582) );
  INVX1 U1076 ( .A(n1708), .Y(n1608) );
  INVX1 U1077 ( .A(n1707), .Y(n1606) );
  INVX1 U1078 ( .A(n815), .Y(n2326) );
  OAI31XL U1079 ( .A(n1573), .B(cs_run), .C(n1572), .D(n1538), .Y(n1535) );
  AND2X1 U1080 ( .A(n1540), .B(n287), .Y(N515) );
  OAI22X1 U1081 ( .A(n1539), .B(n1538), .C(n1537), .D(n1535), .Y(n1540) );
  AND2X1 U1082 ( .A(n1543), .B(n1541), .Y(n1537) );
  INVXL U1083 ( .A(n1657), .Y(n1539) );
  INVX1 U1084 ( .A(ramdatai[6]), .Y(n2491) );
  INVX1 U1085 ( .A(ramdatai[0]), .Y(n2495) );
  OAI22X1 U1086 ( .A(n1571), .B(n1543), .C(n1542), .D(n1541), .Y(n1880) );
  INVX1 U1087 ( .A(ramdatai[1]), .Y(n2494) );
  INVX1 U1088 ( .A(ramdatai[7]), .Y(n904) );
  INVX1 U1089 ( .A(ramdatai[2]), .Y(n2493) );
  INVX1 U1090 ( .A(ramdatai[3]), .Y(n2492) );
  INVX1 U1091 ( .A(n1985), .Y(n2340) );
  INVX1 U1092 ( .A(n1023), .Y(n458) );
  INVX1 U1093 ( .A(n1089), .Y(n2366) );
  INVX1 U1094 ( .A(n716), .Y(n1020) );
  INVX1 U1095 ( .A(n711), .Y(n1012) );
  INVX1 U1096 ( .A(n706), .Y(n997) );
  AOI31X1 U1097 ( .A(n724), .B(n1439), .C(n211), .D(n727), .Y(n725) );
  MUX2X1 U1098 ( .D0(n1436), .D1(n2229), .S(n214), .Y(n724) );
  INVX1 U1099 ( .A(n1034), .Y(n2353) );
  INVX1 U1100 ( .A(n2182), .Y(n262) );
  INVX1 U1101 ( .A(n1855), .Y(n127) );
  AOI222XL U1102 ( .A(memdatai[3]), .B(n1372), .C(n2218), .D(n2194), .E(
        ramdatai[3]), .F(n1550), .Y(n1549) );
  NAND42X1 U1103 ( .C(n1409), .D(n371), .A(n329), .B(n328), .Y(n338) );
  NAND21X1 U1104 ( .B(n259), .A(n327), .Y(n329) );
  NAND21X1 U1105 ( .B(n2245), .A(n1706), .Y(n328) );
  NOR32XL U1106 ( .B(n970), .C(n746), .A(n2262), .Y(n1771) );
  NOR21XL U1107 ( .B(n1222), .A(n848), .Y(n479) );
  AND2X1 U1108 ( .A(n1742), .B(n1929), .Y(n1778) );
  NOR2X1 U1109 ( .A(n2480), .B(n2367), .Y(n840) );
  XNOR2XL U1110 ( .A(n1678), .B(n1602), .Y(n1676) );
  XNOR2XL U1111 ( .A(n1600), .B(n1599), .Y(n1678) );
  NOR3XL U1112 ( .A(n805), .B(n126), .C(n2437), .Y(n1690) );
  NOR2X1 U1113 ( .A(n2243), .B(n126), .Y(n1632) );
  OAI32X1 U1114 ( .A(n1727), .B(n2434), .C(n260), .D(n2028), .E(n168), .Y(
        n1989) );
  NAND2X1 U1115 ( .A(n973), .B(n788), .Y(n1014) );
  NOR2X1 U1116 ( .A(n2478), .B(n2490), .Y(N14336) );
  INVX1 U1117 ( .A(n2205), .Y(n488) );
  NOR2X1 U1118 ( .A(n2030), .B(n2434), .Y(n768) );
  INVX1 U1119 ( .A(n588), .Y(codefetch_s) );
  INVX1 U1120 ( .A(n418), .Y(n2227) );
  OAI22X1 U1121 ( .A(n1660), .B(n1490), .C(n1489), .D(n2165), .Y(N11500) );
  INVX1 U1122 ( .A(n1828), .Y(n129) );
  INVX1 U1123 ( .A(n1982), .Y(n2361) );
  NOR2X1 U1124 ( .A(n2385), .B(n2448), .Y(n2033) );
  NOR3XL U1125 ( .A(n595), .B(n588), .C(n593), .Y(N671) );
  INVX1 U1126 ( .A(n774), .Y(n2427) );
  INVX1 U1127 ( .A(n698), .Y(n995) );
  INVX1 U1128 ( .A(n1826), .Y(n108) );
  INVX1 U1129 ( .A(n2362), .Y(n1929) );
  INVX1 U1130 ( .A(n1063), .Y(n2288) );
  OAI211X1 U1131 ( .C(n2440), .D(n1434), .A(n1558), .B(n1559), .Y(n892) );
  AOI222XL U1132 ( .A(memdatai[2]), .B(n1372), .C(n2218), .D(n2222), .E(
        ramdatai[2]), .F(n1550), .Y(n1559) );
  INVX1 U1133 ( .A(n938), .Y(n2222) );
  NAND21X1 U1134 ( .B(n2432), .A(n2186), .Y(n2431) );
  NAND21X1 U1135 ( .B(n323), .A(n902), .Y(n1409) );
  INVX1 U1136 ( .A(n675), .Y(n2151) );
  OA21X1 U1137 ( .B(n1434), .C(n669), .A(n1494), .Y(n673) );
  OA22X1 U1138 ( .A(n921), .B(n670), .C(n928), .D(n1739), .Y(n671) );
  OR2X1 U1139 ( .A(n169), .B(n201), .Y(n1931) );
  AOI21X1 U1140 ( .B(n2251), .C(n2253), .A(n387), .Y(n201) );
  NAND21X1 U1141 ( .B(n2243), .A(n1006), .Y(n1647) );
  NAND21X1 U1142 ( .B(n603), .A(n2190), .Y(n324) );
  NAND21X1 U1143 ( .B(n1014), .A(n1764), .Y(n369) );
  OAI211X1 U1144 ( .C(n260), .D(n318), .A(n383), .B(n1931), .Y(n1414) );
  OA22X1 U1145 ( .A(n2450), .B(n386), .C(n2437), .D(n388), .Y(n318) );
  INVX1 U1146 ( .A(n317), .Y(n808) );
  NAND21X1 U1147 ( .B(n2261), .A(n2252), .Y(n317) );
  NOR4XL U1148 ( .A(n1759), .B(n1760), .C(n767), .D(n1690), .Y(n1758) );
  AO2222XL U1149 ( .A(n2242), .B(n1006), .C(n1735), .D(n2185), .E(n1763), .F(
        n2270), .G(n1764), .H(n2269), .Y(n1759) );
  ENOX1 U1150 ( .A(n1761), .B(n2435), .C(n1749), .D(n1762), .Y(n1760) );
  NAND5XL U1151 ( .A(n432), .B(n1886), .C(n1859), .D(n2380), .E(n431), .Y(
        n1489) );
  AND4X1 U1152 ( .A(n1531), .B(n2338), .C(n704), .D(n650), .Y(n431) );
  OAI211XL U1153 ( .C(n1738), .D(n1933), .A(n688), .B(n687), .Y(n2152) );
  OA21X1 U1154 ( .B(n1434), .C(n702), .A(n1460), .Y(n688) );
  OA22X1 U1155 ( .A(n921), .B(n686), .C(n923), .D(n1739), .Y(n687) );
  AOI22X1 U1156 ( .A(n817), .B(n1374), .C(ramdatai[5]), .D(n1375), .Y(n1460)
         );
  NOR2X1 U1157 ( .A(n32), .B(n126), .Y(n751) );
  NOR2X1 U1158 ( .A(n2262), .B(n2190), .Y(n1623) );
  INVX1 U1159 ( .A(n926), .Y(n2148) );
  OAI211XL U1160 ( .C(n1738), .D(n1504), .A(n925), .B(n924), .Y(n926) );
  OA22X1 U1161 ( .A(n921), .B(n2285), .C(n908), .D(n1739), .Y(n924) );
  OA21X1 U1162 ( .B(n1434), .C(n920), .A(n1370), .Y(n925) );
  AO21X1 U1163 ( .B(n963), .C(n1736), .A(n808), .Y(n387) );
  INVX1 U1164 ( .A(n2449), .Y(n2185) );
  NAND2X1 U1165 ( .A(n855), .B(n1222), .Y(n1139) );
  NOR2X1 U1166 ( .A(n2243), .B(n2190), .Y(n1335) );
  NOR2X1 U1167 ( .A(n1013), .B(n2245), .Y(n1136) );
  NAND2X1 U1168 ( .A(n1775), .B(n970), .Y(n1727) );
  INVX1 U1169 ( .A(n2450), .Y(n2253) );
  NOR2X1 U1170 ( .A(n2477), .B(n2490), .Y(N14344) );
  INVX1 U1171 ( .A(n789), .Y(n2397) );
  NAND2X1 U1172 ( .A(n2363), .B(n2365), .Y(n1099) );
  NOR2X1 U1173 ( .A(n1099), .B(n2324), .Y(n228) );
  NOR2X1 U1174 ( .A(n1098), .B(n2324), .Y(n224) );
  NOR2X1 U1175 ( .A(n1097), .B(n2324), .Y(n230) );
  NOR2X1 U1176 ( .A(n1095), .B(n2324), .Y(n226) );
  NOR2X1 U1177 ( .A(n1099), .B(n2324), .Y(n227) );
  NOR2X1 U1178 ( .A(n1098), .B(n2324), .Y(n223) );
  NOR2X1 U1179 ( .A(n1099), .B(n152), .Y(n511) );
  NOR2X1 U1180 ( .A(n1098), .B(n152), .Y(n513) );
  NOR2X1 U1181 ( .A(n1097), .B(n2324), .Y(n229) );
  NOR2X1 U1182 ( .A(n1095), .B(n2324), .Y(n225) );
  NOR2X1 U1183 ( .A(n1097), .B(n2324), .Y(n512) );
  NOR2X1 U1184 ( .A(n1095), .B(n152), .Y(n514) );
  INVX1 U1185 ( .A(n1723), .Y(n2396) );
  INVX1 U1186 ( .A(n2091), .Y(n2425) );
  NAND2X1 U1187 ( .A(n751), .B(n2261), .Y(n2100) );
  NOR2X1 U1188 ( .A(n2030), .B(n2449), .Y(n1978) );
  NAND3X1 U1189 ( .A(n2269), .B(n1723), .C(n1623), .Y(n1704) );
  OAI221X1 U1190 ( .A(n2432), .B(n388), .C(n2448), .D(n2383), .E(n1755), .Y(
        n1747) );
  AOI31X1 U1191 ( .A(n1736), .B(n1005), .C(n1756), .D(n2265), .Y(n1755) );
  INVX1 U1192 ( .A(n1757), .Y(n2265) );
  INVX1 U1193 ( .A(n871), .Y(n2399) );
  INVX1 U1194 ( .A(n971), .Y(n2436) );
  INVX1 U1195 ( .A(n739), .Y(n2149) );
  OAI211XL U1196 ( .C(n1738), .D(n975), .A(n738), .B(n735), .Y(n739) );
  OA22X1 U1197 ( .A(n921), .B(n734), .C(n918), .D(n1739), .Y(n735) );
  OA21X1 U1198 ( .B(n1434), .C(n2358), .A(n1423), .Y(n738) );
  INVX1 U1199 ( .A(n1773), .Y(n2420) );
  NAND3X1 U1200 ( .A(n1335), .B(n789), .C(n2269), .Y(n1698) );
  GEN2XL U1201 ( .D(n321), .E(n320), .C(n2182), .B(n370), .A(n399), .Y(n1859)
         );
  AND2X1 U1202 ( .A(n2244), .B(n2267), .Y(n321) );
  AND2X1 U1203 ( .A(n314), .B(n2173), .Y(n320) );
  OR3XL U1204 ( .A(n1372), .B(n2360), .C(n1618), .Y(n1739) );
  NAND32X1 U1205 ( .B(n1497), .C(n427), .A(n424), .Y(n2291) );
  NAND43X1 U1206 ( .B(n323), .C(n304), .D(n327), .A(n2099), .Y(n580) );
  NOR21XL U1207 ( .B(n1710), .A(n1722), .Y(n2099) );
  INVX1 U1208 ( .A(n358), .Y(n304) );
  OR2X1 U1209 ( .A(n2187), .B(n383), .Y(n384) );
  AO21X1 U1210 ( .B(n428), .C(n427), .A(n426), .Y(n1550) );
  INVX1 U1211 ( .A(n1498), .Y(n426) );
  INVX1 U1212 ( .A(n1497), .Y(n428) );
  NAND21X1 U1213 ( .B(n418), .A(n1623), .Y(n2147) );
  OAI221X1 U1214 ( .A(n261), .B(n421), .C(n1620), .D(n170), .E(n420), .Y(n1372) );
  INVX1 U1215 ( .A(n976), .Y(n420) );
  AOI211X1 U1216 ( .C(n2185), .D(n1625), .A(n2384), .B(n1626), .Y(n1620) );
  AND3X1 U1217 ( .A(n2147), .B(n1609), .C(n419), .Y(n421) );
  NAND2X1 U1218 ( .A(n785), .B(n432), .Y(n319) );
  NAND21X1 U1219 ( .B(n2449), .A(n2251), .Y(n436) );
  NAND32X1 U1220 ( .B(n1497), .C(n424), .A(n1496), .Y(n1434) );
  OAI211X1 U1221 ( .C(n1618), .D(n2360), .A(n422), .B(n921), .Y(n1497) );
  NOR42XL U1222 ( .C(n797), .D(n798), .A(n799), .B(n800), .Y(n743) );
  OAI31XL U1223 ( .A(n16), .B(n169), .C(n620), .D(n1090), .Y(n2142) );
  AOI211X1 U1224 ( .C(n128), .D(n745), .A(n1634), .B(n1635), .Y(n1618) );
  NOR2X1 U1225 ( .A(n1773), .B(n2432), .Y(n601) );
  NOR32XL U1226 ( .B(n1006), .C(n1335), .A(n2397), .Y(n1138) );
  NOR2X1 U1227 ( .A(n2383), .B(n2449), .Y(n956) );
  NOR2X1 U1228 ( .A(n2385), .B(n2261), .Y(n1644) );
  INVX1 U1229 ( .A(n370), .Y(n1957) );
  INVX1 U1230 ( .A(n422), .Y(n425) );
  INVX1 U1231 ( .A(n17), .Y(n2428) );
  OAI31XL U1232 ( .A(n901), .B(n2426), .C(n170), .D(n596), .Y(n900) );
  INVX1 U1233 ( .A(n899), .Y(n596) );
  NOR2X1 U1234 ( .A(n2261), .B(n126), .Y(n963) );
  INVX1 U1235 ( .A(n392), .Y(n2251) );
  OAI32X1 U1236 ( .A(n2448), .B(n1632), .C(n33), .D(n2392), .E(n1633), .Y(
        n1631) );
  INVX1 U1237 ( .A(n473), .Y(n1779) );
  OAI211X1 U1238 ( .C(n2431), .D(n2418), .A(n755), .B(n757), .Y(n611) );
  AOI221XL U1239 ( .A(n758), .B(n2253), .C(n760), .D(n147), .E(n2268), .Y(n757) );
  INVX1 U1240 ( .A(n1727), .Y(n2268) );
  AOI32X1 U1241 ( .A(n2185), .B(n128), .C(n1005), .D(n2091), .E(n2105), .Y(
        n2102) );
  OAI21X1 U1242 ( .B(n1335), .C(n2447), .A(n2433), .Y(n2105) );
  INVX1 U1243 ( .A(n1734), .Y(n2179) );
  NAND21X1 U1244 ( .B(n2435), .A(n2186), .Y(n1734) );
  AOI21X1 U1245 ( .B(n2420), .C(n2106), .A(n2241), .Y(n2101) );
  INVX1 U1246 ( .A(n602), .Y(n2315) );
  NOR2X1 U1247 ( .A(n973), .B(n969), .Y(n972) );
  OR2X1 U1248 ( .A(n2179), .B(n971), .Y(n2114) );
  INVX1 U1249 ( .A(n2106), .Y(n2435) );
  INVX1 U1250 ( .A(n1774), .Y(n2398) );
  INVX1 U1251 ( .A(n1627), .Y(n2384) );
  INVX1 U1252 ( .A(n965), .Y(n2391) );
  INVX1 U1253 ( .A(n1054), .Y(n2307) );
  NAND32X1 U1254 ( .B(n2187), .C(n1372), .A(n425), .Y(n1738) );
  NAND32X1 U1255 ( .B(n260), .C(n2416), .A(n1636), .Y(n1496) );
  OAI221X1 U1256 ( .A(n128), .B(n1633), .C(n1632), .D(n64), .E(n2433), .Y(
        n1636) );
  MUX2X1 U1257 ( .D0(n2478), .D1(n2320), .S(n1957), .Y(n377) );
  OAI31XL U1258 ( .A(n16), .B(n169), .C(n620), .D(n1090), .Y(n221) );
  OAI31XL U1259 ( .A(n16), .B(n170), .C(n620), .D(n1090), .Y(n220) );
  NAND21X1 U1260 ( .B(n2226), .A(n2323), .Y(n689) );
  NAND2X1 U1261 ( .A(n2033), .B(n1324), .Y(n809) );
  INVX1 U1262 ( .A(n1435), .Y(n2202) );
  INVX1 U1263 ( .A(n2380), .Y(n2246) );
  AOI221XL U1264 ( .A(n1736), .B(n1765), .C(n973), .D(n1644), .E(n583), .Y(
        n776) );
  OAI211X1 U1265 ( .C(n783), .D(n261), .A(n784), .B(n785), .Y(n692) );
  AOI21X1 U1266 ( .B(n601), .C(n789), .A(n2421), .Y(n783) );
  NAND42X1 U1267 ( .C(n786), .D(n603), .A(n2184), .B(n788), .Y(n784) );
  NAND2X1 U1268 ( .A(n1006), .B(n1723), .Y(n901) );
  OAI211X1 U1269 ( .C(n260), .D(n393), .A(n392), .B(n2202), .Y(n394) );
  AND2X1 U1270 ( .A(n386), .B(n385), .Y(n393) );
  INVX1 U1271 ( .A(n583), .Y(n385) );
  NAND2X1 U1272 ( .A(n788), .B(n774), .Y(n769) );
  MUX2IX1 U1273 ( .D0(n2477), .D1(n2317), .S(n1957), .Y(n202) );
  OAI211X1 U1274 ( .C(n2392), .D(n2072), .A(n798), .B(n2382), .Y(n1010) );
  NAND2X1 U1275 ( .A(n746), .B(n2262), .Y(n2072) );
  NAND3X1 U1276 ( .A(n2115), .B(n1004), .C(n2116), .Y(n780) );
  OAI21X1 U1277 ( .B(n2179), .C(n2112), .A(n2043), .Y(n2115) );
  AOI22X1 U1278 ( .A(n1006), .B(n2117), .C(n2046), .D(n1635), .Y(n2116) );
  OAI22X1 U1279 ( .A(n2396), .B(n2429), .C(n2118), .D(n147), .Y(n2117) );
  OAI22X1 U1280 ( .A(n771), .B(n2425), .C(n772), .D(n2430), .Y(n770) );
  AOI22AXL U1281 ( .A(n2381), .B(n109), .D(n773), .C(n774), .Y(n771) );
  AOI32X1 U1282 ( .A(n1649), .B(n2089), .C(n760), .D(n963), .E(n1763), .Y(
        n2085) );
  INVX1 U1283 ( .A(n2360), .Y(n604) );
  AOI211X1 U1284 ( .C(n109), .D(n147), .A(n2092), .B(n2253), .Y(n2084) );
  AOI211X1 U1285 ( .C(n1623), .D(n32), .A(n2186), .B(n1752), .Y(n2077) );
  INVX1 U1286 ( .A(n973), .Y(n2447) );
  AOI31X1 U1287 ( .A(n742), .B(n2267), .C(n2071), .D(n2238), .Y(n2070) );
  AOI31X1 U1288 ( .A(n788), .B(n2190), .C(n2050), .D(n1010), .Y(n2071) );
  INVX1 U1289 ( .A(n902), .Y(n2379) );
  NAND2X1 U1290 ( .A(n17), .B(n33), .Y(n2078) );
  NOR2X1 U1291 ( .A(n17), .B(n1764), .Y(n2118) );
  NAND21X1 U1292 ( .B(n785), .A(n945), .Y(n2338) );
  NAND21X1 U1293 ( .B(n2246), .A(n397), .Y(n704) );
  NAND32X1 U1294 ( .B(n1014), .C(n147), .A(n2242), .Y(n1004) );
  OAI21X1 U1295 ( .B(n974), .C(n2437), .A(n1013), .Y(n777) );
  NAND21X1 U1296 ( .B(n2226), .A(n2322), .Y(n655) );
  NAND3X1 U1297 ( .A(n970), .B(n61), .C(n17), .Y(n2039) );
  INVX1 U1298 ( .A(n993), .Y(n693) );
  INVX1 U1299 ( .A(n991), .Y(n678) );
  INVX1 U1300 ( .A(n1410), .Y(n672) );
  INVX1 U1301 ( .A(n1699), .Y(intcall) );
  NAND2X1 U1302 ( .A(n1623), .B(n39), .Y(n2052) );
  AOI31X1 U1303 ( .A(n2381), .B(n109), .C(n39), .D(n808), .Y(n796) );
  OAI222XL U1304 ( .A(n2415), .B(n823), .C(n2489), .D(n824), .E(n2406), .F(
        n2323), .Y(n821) );
  OAI221X1 U1305 ( .A(n2473), .B(n824), .C(n823), .D(n2475), .E(n2223), .Y(
        n819) );
  OAI21X1 U1306 ( .B(n62), .C(n2425), .A(n2418), .Y(n753) );
  NOR3XL U1307 ( .A(n2450), .B(n805), .C(n2385), .Y(n800) );
  INVX1 U1308 ( .A(n1610), .Y(n1701) );
  NAND32X1 U1309 ( .B(n169), .C(n1609), .A(n2205), .Y(n1610) );
  NAND2X1 U1310 ( .A(n2482), .B(n2487), .Y(n1067) );
  AOI221XL U1311 ( .A(n984), .B(memdatai[2]), .C(n983), .D(n235), .E(n994), 
        .Y(n1433) );
  OAI22X1 U1312 ( .A(n2327), .B(n986), .C(n2346), .D(n2493), .Y(n994) );
  AOI221XL U1313 ( .A(ramdatai[4]), .B(n980), .C(n2347), .D(n816), .E(n990), 
        .Y(n989) );
  OAI22X1 U1314 ( .A(n2349), .B(n670), .C(n40), .D(n2348), .Y(n990) );
  NAND21X1 U1315 ( .B(n2195), .A(n237), .Y(n2067) );
  MUX2X1 U1316 ( .D0(n2249), .D1(n2247), .S(pc_o[1]), .Y(n455) );
  INVX1 U1317 ( .A(n823), .Y(n1440) );
  INVX1 U1318 ( .A(n2323), .Y(n484) );
  INVX1 U1319 ( .A(n824), .Y(n2038) );
  INVX1 U1320 ( .A(n2322), .Y(n362) );
  OAI22XL U1321 ( .A(n1504), .B(n1503), .C(n979), .D(n294), .Y(N12721) );
  AOI221XL U1322 ( .A(ramdatai[7]), .B(n980), .C(n2347), .D(n2313), .E(n981), 
        .Y(n979) );
  OAI22X1 U1323 ( .A(n2349), .B(n2285), .C(n34), .D(n2348), .Y(n981) );
  OAI22XL U1324 ( .A(n1933), .B(n1503), .C(n987), .D(n294), .Y(N12719) );
  AOI221XL U1325 ( .A(ramdatai[5]), .B(n980), .C(n2347), .D(n817), .E(n988), 
        .Y(n987) );
  OAI22X1 U1326 ( .A(n2349), .B(n686), .C(n46), .D(n2348), .Y(n988) );
  OAI22XL U1327 ( .A(n292), .B(n790), .C(n787), .D(n1503), .Y(N12714) );
  AOI221XL U1328 ( .A(n2347), .B(n812), .C(n980), .D(ramdatai[0]), .E(n998), 
        .Y(n790) );
  ENOX1 U1329 ( .A(n53), .B(n2348), .C(n984), .D(memdatai[0]), .Y(n998) );
  OAI22XL U1330 ( .A(n293), .B(n778), .C(n775), .D(n1503), .Y(N12715) );
  AOI221XL U1331 ( .A(n2347), .B(n813), .C(n980), .D(ramdatai[1]), .E(n996), 
        .Y(n778) );
  ENOX1 U1332 ( .A(n51), .B(n2348), .C(n984), .D(memdatai[1]), .Y(n996) );
  NAND21X1 U1333 ( .B(n2212), .A(n238), .Y(n2276) );
  NAND21X1 U1334 ( .B(n12), .A(n238), .Y(n2278) );
  NAND21X1 U1335 ( .B(n2216), .A(n238), .Y(n2277) );
  NAND21X1 U1336 ( .B(n2199), .A(n238), .Y(n2280) );
  NAND21X1 U1337 ( .B(n2192), .A(n238), .Y(n2279) );
  NAND21X1 U1338 ( .B(n2208), .A(n239), .Y(n765) );
  NAND21X1 U1339 ( .B(n2203), .A(n239), .Y(n2283) );
  AND2X1 U1340 ( .A(n1348), .B(n1350), .Y(n1346) );
  NAND4X1 U1341 ( .A(n1026), .B(n1034), .C(n1351), .D(n1352), .Y(n1350) );
  AOI21X1 U1342 ( .B(n1349), .C(n2258), .A(n1033), .Y(n1351) );
  AOI211X1 U1343 ( .C(n1023), .D(n2259), .A(n1032), .B(n1031), .Y(n1352) );
  NAND2X1 U1344 ( .A(n856), .B(n1222), .Y(n1236) );
  NOR2X1 U1345 ( .A(n2234), .B(n164), .Y(n1235) );
  INVX1 U1346 ( .A(n1572), .Y(n1499) );
  INVX1 U1347 ( .A(n1591), .Y(n1562) );
  OAI22X1 U1348 ( .A(n638), .B(n114), .C(n1223), .D(n139), .Y(N12555) );
  OAI22X1 U1349 ( .A(n638), .B(n92), .C(n1223), .D(n115), .Y(N12546) );
  OAI22X1 U1350 ( .A(n638), .B(n138), .C(n1223), .D(n95), .Y(N12510) );
  OAI22X1 U1351 ( .A(n638), .B(n136), .C(n1223), .D(n85), .Y(N12537) );
  OAI22X1 U1352 ( .A(n638), .B(n84), .C(n1223), .D(n70), .Y(N12501) );
  OAI22X1 U1353 ( .A(n638), .B(n112), .C(n1223), .D(n68), .Y(N12564) );
  OAI22X1 U1354 ( .A(n638), .B(n94), .C(n1223), .D(n155), .Y(N12519) );
  OAI22X1 U1355 ( .A(n638), .B(n82), .C(n1223), .D(n63), .Y(N12528) );
  OAI22X1 U1356 ( .A(n736), .B(n113), .C(n1110), .D(n1112), .Y(N12620) );
  OAI22X1 U1357 ( .A(n698), .B(n113), .C(n1104), .D(n1112), .Y(N12627) );
  OAI22X1 U1358 ( .A(n698), .B(n93), .C(n1104), .D(n1120), .Y(N12591) );
  OAI22X1 U1359 ( .A(n736), .B(n91), .C(n1110), .D(n1114), .Y(N12611) );
  OAI22X1 U1360 ( .A(n698), .B(n91), .C(n1104), .D(n1114), .Y(N12618) );
  OAI22X1 U1361 ( .A(n736), .B(n137), .C(n1110), .D(n1122), .Y(N12575) );
  OAI22X1 U1362 ( .A(n698), .B(n137), .C(n1104), .D(n1122), .Y(N12582) );
  OAI22X1 U1363 ( .A(n736), .B(n135), .C(n1110), .D(n1116), .Y(N12602) );
  OAI22X1 U1364 ( .A(n698), .B(n135), .C(n1104), .D(n1116), .Y(N12609) );
  OAI22X1 U1365 ( .A(n698), .B(n83), .C(n1104), .D(n1124), .Y(N12573) );
  OAI22X1 U1366 ( .A(n736), .B(n111), .C(n1110), .D(n1105), .Y(N12629) );
  OAI22X1 U1367 ( .A(n698), .B(n111), .C(n1104), .D(n1105), .Y(N12636) );
  OAI22X1 U1368 ( .A(n698), .B(n81), .C(n1104), .D(n1118), .Y(N12600) );
  OAI22X1 U1369 ( .A(n693), .B(n94), .C(n2301), .D(n155), .Y(N12512) );
  OAI22X1 U1370 ( .A(n693), .B(n114), .C(n2301), .D(n139), .Y(N12548) );
  OAI22X1 U1371 ( .A(n731), .B(n113), .C(n1109), .D(n1112), .Y(N12621) );
  OAI22X1 U1372 ( .A(n726), .B(n113), .C(n1108), .D(n1112), .Y(N12622) );
  OAI22X1 U1373 ( .A(n716), .B(n113), .C(n1107), .D(n1112), .Y(N12624) );
  OAI22X1 U1374 ( .A(n711), .B(n113), .C(n2293), .D(n1112), .Y(N12625) );
  OAI22X1 U1375 ( .A(n706), .B(n113), .C(n1106), .D(n1112), .Y(N12626) );
  OAI22X1 U1376 ( .A(n678), .B(n114), .C(n1226), .D(n139), .Y(N12549) );
  OAI22X1 U1377 ( .A(n665), .B(n114), .C(n1225), .D(n139), .Y(N12551) );
  OAI22X1 U1378 ( .A(n653), .B(n114), .C(n2297), .D(n139), .Y(N12552) );
  OAI22X1 U1379 ( .A(n648), .B(n114), .C(n2295), .D(n139), .Y(N12553) );
  OAI22X1 U1380 ( .A(n643), .B(n114), .C(n1224), .D(n1112), .Y(N12554) );
  OAI22X1 U1381 ( .A(n736), .B(n93), .C(n1110), .D(n1120), .Y(N12584) );
  OAI22X1 U1382 ( .A(n731), .B(n93), .C(n1109), .D(n1120), .Y(N12585) );
  OAI22X1 U1383 ( .A(n726), .B(n93), .C(n1108), .D(n1120), .Y(N12586) );
  OAI22X1 U1384 ( .A(n716), .B(n93), .C(n1107), .D(n1120), .Y(N12588) );
  OAI22X1 U1385 ( .A(n711), .B(n93), .C(n2293), .D(n1120), .Y(N12589) );
  OAI22X1 U1386 ( .A(n706), .B(n93), .C(n1106), .D(n1120), .Y(N12590) );
  OAI22X1 U1387 ( .A(n678), .B(n94), .C(n1226), .D(n155), .Y(N12513) );
  OAI22X1 U1388 ( .A(n665), .B(n94), .C(n1225), .D(n155), .Y(N12515) );
  OAI22X1 U1389 ( .A(n653), .B(n94), .C(n2297), .D(n155), .Y(N12516) );
  OAI22X1 U1390 ( .A(n648), .B(n94), .C(n2295), .D(n155), .Y(N12517) );
  OAI22X1 U1391 ( .A(n643), .B(n94), .C(n1224), .D(n1120), .Y(N12518) );
  OAI22X1 U1392 ( .A(n693), .B(n138), .C(n2301), .D(n95), .Y(N12503) );
  OAI22X1 U1393 ( .A(n693), .B(n92), .C(n2301), .D(n115), .Y(N12539) );
  OAI22X1 U1394 ( .A(n731), .B(n91), .C(n1109), .D(n1114), .Y(N12612) );
  OAI22X1 U1395 ( .A(n726), .B(n91), .C(n1108), .D(n1114), .Y(N12613) );
  OAI22X1 U1396 ( .A(n716), .B(n91), .C(n1107), .D(n1114), .Y(N12615) );
  OAI22X1 U1397 ( .A(n711), .B(n91), .C(n2293), .D(n1114), .Y(N12616) );
  OAI22X1 U1398 ( .A(n706), .B(n91), .C(n1106), .D(n1114), .Y(N12617) );
  OAI22X1 U1399 ( .A(n678), .B(n92), .C(n1226), .D(n115), .Y(N12540) );
  OAI22X1 U1400 ( .A(n665), .B(n92), .C(n1225), .D(n115), .Y(N12542) );
  OAI22X1 U1401 ( .A(n653), .B(n92), .C(n2297), .D(n115), .Y(N12543) );
  OAI22X1 U1402 ( .A(n648), .B(n92), .C(n2295), .D(n115), .Y(N12544) );
  OAI22X1 U1403 ( .A(n643), .B(n92), .C(n1224), .D(n1114), .Y(N12545) );
  OAI22X1 U1404 ( .A(n731), .B(n137), .C(n1109), .D(n1122), .Y(N12576) );
  OAI22X1 U1405 ( .A(n726), .B(n137), .C(n1108), .D(n1122), .Y(N12577) );
  OAI22X1 U1406 ( .A(n716), .B(n137), .C(n1107), .D(n1122), .Y(N12579) );
  OAI22X1 U1407 ( .A(n711), .B(n137), .C(n2293), .D(n1122), .Y(N12580) );
  OAI22X1 U1408 ( .A(n706), .B(n137), .C(n1106), .D(n1122), .Y(N12581) );
  OAI22X1 U1409 ( .A(n678), .B(n138), .C(n1226), .D(n95), .Y(N12504) );
  OAI22X1 U1410 ( .A(n665), .B(n138), .C(n1225), .D(n95), .Y(N12506) );
  OAI22X1 U1411 ( .A(n653), .B(n138), .C(n2297), .D(n95), .Y(N12507) );
  OAI22X1 U1412 ( .A(n648), .B(n138), .C(n2295), .D(n95), .Y(N12508) );
  OAI22X1 U1413 ( .A(n643), .B(n138), .C(n1224), .D(n1122), .Y(N12509) );
  OAI22X1 U1414 ( .A(n693), .B(n84), .C(n2301), .D(n70), .Y(N12494) );
  OAI22X1 U1415 ( .A(n693), .B(n136), .C(n2301), .D(n85), .Y(N12530) );
  OAI22X1 U1416 ( .A(n731), .B(n135), .C(n1109), .D(n1116), .Y(N12603) );
  OAI22X1 U1417 ( .A(n726), .B(n135), .C(n1108), .D(n1116), .Y(N12604) );
  OAI22X1 U1418 ( .A(n716), .B(n135), .C(n1107), .D(n1116), .Y(N12606) );
  OAI22X1 U1419 ( .A(n711), .B(n135), .C(n2293), .D(n1116), .Y(N12607) );
  OAI22X1 U1420 ( .A(n706), .B(n135), .C(n1106), .D(n1116), .Y(N12608) );
  OAI22X1 U1421 ( .A(n678), .B(n136), .C(n1226), .D(n85), .Y(N12531) );
  OAI22X1 U1422 ( .A(n665), .B(n136), .C(n1225), .D(n85), .Y(N12533) );
  OAI22X1 U1423 ( .A(n653), .B(n136), .C(n2297), .D(n85), .Y(N12534) );
  OAI22X1 U1424 ( .A(n648), .B(n136), .C(n2295), .D(n85), .Y(N12535) );
  OAI22X1 U1425 ( .A(n643), .B(n136), .C(n1224), .D(n1116), .Y(N12536) );
  OAI22X1 U1426 ( .A(n736), .B(n83), .C(n1110), .D(n1124), .Y(N12566) );
  OAI22X1 U1427 ( .A(n731), .B(n83), .C(n1109), .D(n1124), .Y(N12567) );
  OAI22X1 U1428 ( .A(n726), .B(n83), .C(n1108), .D(n1124), .Y(N12568) );
  OAI22X1 U1429 ( .A(n716), .B(n83), .C(n1107), .D(n1124), .Y(N12570) );
  OAI22X1 U1430 ( .A(n711), .B(n83), .C(n2293), .D(n1124), .Y(N12571) );
  OAI22X1 U1431 ( .A(n706), .B(n83), .C(n1106), .D(n1124), .Y(N12572) );
  OAI22X1 U1432 ( .A(n678), .B(n84), .C(n1226), .D(n70), .Y(N12495) );
  OAI22X1 U1433 ( .A(n665), .B(n84), .C(n1225), .D(n70), .Y(N12497) );
  OAI22X1 U1434 ( .A(n653), .B(n84), .C(n2297), .D(n70), .Y(N12498) );
  OAI22X1 U1435 ( .A(n648), .B(n84), .C(n2295), .D(n70), .Y(N12499) );
  OAI22X1 U1436 ( .A(n643), .B(n84), .C(n1224), .D(n1124), .Y(N12500) );
  OAI22X1 U1437 ( .A(n693), .B(n82), .C(n2301), .D(n63), .Y(N12521) );
  OAI22X1 U1438 ( .A(n693), .B(n112), .C(n2301), .D(n68), .Y(N12557) );
  OAI22X1 U1439 ( .A(n731), .B(n111), .C(n1109), .D(n1105), .Y(N12630) );
  OAI22X1 U1440 ( .A(n726), .B(n111), .C(n1108), .D(n1105), .Y(N12631) );
  OAI22X1 U1441 ( .A(n716), .B(n111), .C(n1107), .D(n1105), .Y(N12633) );
  OAI22X1 U1442 ( .A(n711), .B(n111), .C(n2293), .D(n1105), .Y(N12634) );
  OAI22X1 U1443 ( .A(n706), .B(n111), .C(n1106), .D(n1105), .Y(N12635) );
  OAI22X1 U1444 ( .A(n678), .B(n112), .C(n1226), .D(n68), .Y(N12558) );
  OAI22X1 U1445 ( .A(n665), .B(n112), .C(n1225), .D(n68), .Y(N12560) );
  OAI22X1 U1446 ( .A(n653), .B(n112), .C(n2297), .D(n68), .Y(N12561) );
  OAI22X1 U1447 ( .A(n648), .B(n112), .C(n2295), .D(n68), .Y(N12562) );
  OAI22X1 U1448 ( .A(n643), .B(n112), .C(n1224), .D(n1105), .Y(N12563) );
  OAI22X1 U1449 ( .A(n736), .B(n81), .C(n1110), .D(n1118), .Y(N12593) );
  OAI22X1 U1450 ( .A(n731), .B(n81), .C(n1109), .D(n1118), .Y(N12594) );
  OAI22X1 U1451 ( .A(n726), .B(n81), .C(n1108), .D(n1118), .Y(N12595) );
  OAI22X1 U1452 ( .A(n716), .B(n81), .C(n1107), .D(n1118), .Y(N12597) );
  OAI22X1 U1453 ( .A(n711), .B(n81), .C(n2293), .D(n1118), .Y(N12598) );
  OAI22X1 U1454 ( .A(n706), .B(n81), .C(n1106), .D(n1118), .Y(N12599) );
  OAI22X1 U1455 ( .A(n678), .B(n82), .C(n1226), .D(n63), .Y(N12522) );
  OAI22X1 U1456 ( .A(n665), .B(n82), .C(n1225), .D(n63), .Y(N12524) );
  OAI22X1 U1457 ( .A(n653), .B(n82), .C(n2297), .D(n63), .Y(N12525) );
  OAI22X1 U1458 ( .A(n648), .B(n82), .C(n2295), .D(n63), .Y(N12526) );
  OAI22X1 U1459 ( .A(n643), .B(n82), .C(n1224), .D(n1118), .Y(N12527) );
  OAI22X1 U1460 ( .A(n721), .B(n113), .C(n2294), .D(n1112), .Y(N12623) );
  OAI22X1 U1461 ( .A(n721), .B(n93), .C(n2294), .D(n1120), .Y(N12587) );
  OAI22X1 U1462 ( .A(n721), .B(n91), .C(n2294), .D(n1114), .Y(N12614) );
  OAI22X1 U1463 ( .A(n721), .B(n137), .C(n2294), .D(n1122), .Y(N12578) );
  OAI22X1 U1464 ( .A(n721), .B(n135), .C(n2294), .D(n1116), .Y(N12605) );
  OAI22X1 U1465 ( .A(n721), .B(n83), .C(n2294), .D(n1124), .Y(N12569) );
  OAI22X1 U1466 ( .A(n721), .B(n111), .C(n2294), .D(n1105), .Y(N12632) );
  OAI22X1 U1467 ( .A(n721), .B(n81), .C(n2294), .D(n1118), .Y(N12596) );
  OAI21X1 U1468 ( .B(n848), .C(n854), .A(n288), .Y(N13014) );
  OAI21X1 U1469 ( .B(n847), .C(n854), .A(n289), .Y(N13023) );
  OAI21X1 U1470 ( .B(n846), .C(n854), .A(n289), .Y(N13032) );
  OAI21X1 U1471 ( .B(n845), .C(n854), .A(n289), .Y(N13041) );
  OAI21X1 U1472 ( .B(n2143), .C(n854), .A(n289), .Y(N13050) );
  OAI21X1 U1473 ( .B(n2441), .C(n854), .A(n289), .Y(N13059) );
  OAI21X1 U1474 ( .B(n844), .C(n854), .A(n289), .Y(N13068) );
  OAI21X1 U1475 ( .B(n842), .C(n854), .A(n289), .Y(N13077) );
  OAI21X1 U1476 ( .B(n848), .C(n851), .A(n296), .Y(N13158) );
  OAI21X1 U1477 ( .B(n847), .C(n851), .A(n296), .Y(N13167) );
  OAI21X1 U1478 ( .B(n846), .C(n851), .A(n296), .Y(N13176) );
  OAI21X1 U1479 ( .B(n845), .C(n851), .A(n297), .Y(N13185) );
  OAI21X1 U1480 ( .B(n2143), .C(n851), .A(n290), .Y(N13194) );
  OAI21X1 U1481 ( .B(n2441), .C(n851), .A(n290), .Y(N13203) );
  OAI21X1 U1482 ( .B(n844), .C(n851), .A(n290), .Y(N13212) );
  OAI21X1 U1483 ( .B(n842), .C(n851), .A(n290), .Y(N13221) );
  INVX1 U1484 ( .A(n1344), .Y(n2281) );
  INVX1 U1485 ( .A(n1343), .Y(n2282) );
  NAND32X1 U1486 ( .B(n170), .C(n69), .A(n601), .Y(n1369) );
  NAND32X1 U1487 ( .B(n1562), .C(n248), .A(n588), .Y(n587) );
  NOR21XL U1488 ( .B(multemp2[2]), .A(n839), .Y(N13325) );
  NOR21XL U1489 ( .B(multemp2[3]), .A(n839), .Y(N13326) );
  NOR21XL U1490 ( .B(multemp2[4]), .A(n839), .Y(N13327) );
  NOR21XL U1491 ( .B(multemp2[5]), .A(n839), .Y(N13328) );
  NOR21XL U1492 ( .B(multemp2[6]), .A(n839), .Y(N13329) );
  NOR21XL U1493 ( .B(multemp2[7]), .A(n839), .Y(N13330) );
  NOR21XL U1494 ( .B(multemp2[8]), .A(n839), .Y(N13331) );
  NAND21X1 U1495 ( .B(n245), .A(n17), .Y(n2034) );
  NAND21X1 U1496 ( .B(n588), .A(n237), .Y(n585) );
  NAND21X1 U1497 ( .B(n247), .A(n1090), .Y(n1080) );
  AO21X1 U1498 ( .B(n244), .C(n1645), .A(n294), .Y(N12722) );
  NAND43X1 U1499 ( .B(n977), .C(n976), .D(n2359), .A(n945), .Y(n1645) );
  AO21X1 U1500 ( .B(n244), .C(n1646), .A(n295), .Y(N11491) );
  INVX1 U1501 ( .A(n1742), .Y(n1646) );
  INVX1 U1502 ( .A(n859), .Y(n2232) );
  AND3X1 U1503 ( .A(n240), .B(n971), .C(n2172), .Y(N10573) );
  AND3X1 U1504 ( .A(n240), .B(n2205), .C(n11), .Y(N585) );
  AND3X1 U1505 ( .A(n1764), .B(n2241), .C(n243), .Y(N10584) );
  NOR32XL U1506 ( .B(n239), .C(n1005), .A(n901), .Y(N10586) );
  INVX1 U1507 ( .A(n2146), .Y(n1100) );
  NAND43X1 U1508 ( .B(n2162), .C(n2145), .D(n2143), .A(n853), .Y(n2146) );
  INVX1 U1509 ( .A(n856), .Y(n2143) );
  INVX1 U1510 ( .A(n1102), .Y(n2145) );
  AND2X1 U1511 ( .A(n1511), .B(n1582), .Y(N12912) );
  OAI32X1 U1512 ( .A(n1509), .B(n1508), .C(n1507), .D(n1506), .E(n245), .Y(
        n1511) );
  INVX1 U1513 ( .A(n1505), .Y(n1506) );
  INVX1 U1514 ( .A(n873), .Y(n1508) );
  OAI32X1 U1515 ( .A(n2383), .B(n2450), .C(n246), .D(n2045), .E(n2047), .Y(
        N10571) );
  NAND2X1 U1516 ( .A(n849), .B(n850), .Y(n843) );
  NAND2X1 U1517 ( .A(n849), .B(n853), .Y(n852) );
  OAI221X1 U1518 ( .A(n1339), .B(n1411), .C(n2279), .D(n684), .E(n298), .Y(
        N12487) );
  OAI22AX1 U1519 ( .D(dpc[3]), .C(n1079), .A(n1089), .B(n1080), .Y(N12693) );
  OAI22AX1 U1520 ( .D(dpc[4]), .C(n1079), .A(n2364), .B(n1080), .Y(N12694) );
  OAI22AX1 U1521 ( .D(dpc[5]), .C(n1079), .A(n2325), .B(n1080), .Y(N12695) );
  OAI22AX1 U1522 ( .D(n1652), .C(n2162), .A(n1697), .B(n1507), .Y(N11487) );
  OAI22X1 U1523 ( .A(n759), .B(n2287), .C(n1015), .D(n2067), .Y(N12705) );
  OAI22X1 U1524 ( .A(n947), .B(n246), .C(n910), .D(n467), .Y(N12723) );
  NOR3XL U1525 ( .A(n948), .B(n949), .C(n950), .Y(n947) );
  OAI211X1 U1526 ( .C(n2460), .D(n939), .A(n945), .B(n955), .Y(n948) );
  OAI22X1 U1527 ( .A(n2495), .B(n2271), .C(n951), .D(n909), .Y(n950) );
  OAI22X1 U1528 ( .A(n940), .B(n247), .C(n910), .D(n595), .Y(N12724) );
  NOR3XL U1529 ( .A(n941), .B(n942), .C(n943), .Y(n940) );
  OAI211X1 U1530 ( .C(n2466), .D(n939), .A(n945), .B(n946), .Y(n941) );
  OAI22X1 U1531 ( .A(n2494), .B(n2271), .C(n944), .D(n909), .Y(n943) );
  OAI22X1 U1532 ( .A(n292), .B(n475), .C(n476), .D(n2278), .Y(n1884) );
  AND2X1 U1533 ( .A(n2150), .B(n613), .Y(N372) );
  AND2X1 U1534 ( .A(n2175), .B(n613), .Y(N371) );
  OAI21X1 U1535 ( .B(n848), .C(n852), .A(n289), .Y(N13086) );
  OAI21X1 U1536 ( .B(n847), .C(n852), .A(n289), .Y(N13095) );
  OAI21X1 U1537 ( .B(n846), .C(n852), .A(n289), .Y(N13104) );
  OAI21X1 U1538 ( .B(n845), .C(n852), .A(n297), .Y(N13113) );
  OAI21X1 U1539 ( .B(n844), .C(n852), .A(n297), .Y(N13140) );
  OAI21X1 U1540 ( .B(n848), .C(n843), .A(n290), .Y(N13230) );
  OAI21X1 U1541 ( .B(n847), .C(n843), .A(n290), .Y(N13239) );
  OAI21X1 U1542 ( .B(n843), .C(n846), .A(n290), .Y(N13248) );
  OAI21X1 U1543 ( .B(n843), .C(n845), .A(n290), .Y(N13257) );
  OAI21X1 U1544 ( .B(n844), .C(n843), .A(n296), .Y(N13284) );
  OAI21X1 U1545 ( .B(n1098), .C(n1101), .A(n288), .Y(N12644) );
  OAI21X1 U1546 ( .B(n1097), .C(n1101), .A(n288), .Y(N12651) );
  OAI21X1 U1547 ( .B(n1095), .C(n1101), .A(n288), .Y(N12658) );
  OAI21X1 U1548 ( .B(n1099), .C(n1096), .A(n288), .Y(N12665) );
  OAI21X1 U1549 ( .B(n1098), .C(n1096), .A(n297), .Y(N12672) );
  OAI21X1 U1550 ( .B(n1097), .C(n1096), .A(n288), .Y(N12679) );
  OAI21X1 U1551 ( .B(n1095), .C(n1096), .A(n288), .Y(N12686) );
  AND2X1 U1552 ( .A(sfroe_comb_s), .B(n243), .Y(N11488) );
  INVX1 U1553 ( .A(n1612), .Y(sfroe_comb_s) );
  NAND21X1 U1554 ( .B(n1654), .A(n1611), .Y(n1612) );
  INVX1 U1555 ( .A(n2159), .Y(n2175) );
  NAND32X1 U1556 ( .B(n147), .C(n245), .A(n2158), .Y(n2159) );
  NOR3XL U1557 ( .A(n2034), .B(n2385), .C(n2422), .Y(N10588) );
  INVX1 U1558 ( .A(n1006), .Y(n2422) );
  NOR3XL U1559 ( .A(n2037), .B(n2396), .C(n2450), .Y(N10563) );
  NAND2X1 U1560 ( .A(n1100), .B(n152), .Y(n1101) );
  INVX1 U1561 ( .A(n782), .Y(n2204) );
  NAND21X1 U1562 ( .B(n2205), .A(n239), .Y(n782) );
  NOR2X1 U1563 ( .A(n839), .B(n2290), .Y(N13332) );
  NOR2X1 U1564 ( .A(n838), .B(n832), .Y(N13367) );
  NOR2X1 U1565 ( .A(n837), .B(n832), .Y(N13368) );
  NOR2X1 U1566 ( .A(n835), .B(n832), .Y(N13370) );
  NOR2X1 U1567 ( .A(n836), .B(n832), .Y(N13369) );
  NOR2X1 U1568 ( .A(n834), .B(n832), .Y(N13371) );
  NOR2X1 U1569 ( .A(n833), .B(n832), .Y(N13372) );
  NOR2X1 U1570 ( .A(n831), .B(n832), .Y(N13373) );
  NOR2X1 U1571 ( .A(n2245), .B(n587), .Y(N682) );
  NOR2X1 U1572 ( .A(n902), .B(n2047), .Y(N10567) );
  NOR21XL U1573 ( .B(n249), .A(n2049), .Y(N10569) );
  AOI211X1 U1574 ( .C(n1736), .D(n1625), .A(n808), .B(n2390), .Y(n2049) );
  INVX1 U1575 ( .A(n798), .Y(n2390) );
  NAND2X1 U1576 ( .A(n287), .B(n866), .Y(n864) );
  AO21X1 U1577 ( .B(n2155), .C(n2154), .A(n2153), .Y(n866) );
  OR2X1 U1578 ( .A(n292), .B(n203), .Y(N13366) );
  AOI21X1 U1579 ( .B(n2157), .C(n2259), .A(n248), .Y(n203) );
  AOI22X1 U1580 ( .A(n1374), .B(n2313), .C(ramdatai[7]), .D(n1375), .Y(n1370)
         );
  INVX1 U1581 ( .A(n933), .Y(n2194) );
  NOR2X1 U1582 ( .A(n865), .B(n864), .Y(N12975) );
  XNOR2XL U1583 ( .A(n2369), .B(n2368), .Y(n865) );
  AOI22X1 U1584 ( .A(n818), .B(n1374), .C(ramdatai[6]), .D(n1375), .Y(n1423)
         );
  NAND43X1 U1585 ( .B(n1643), .C(n1642), .D(n293), .A(n1638), .Y(N12977) );
  INVX1 U1586 ( .A(n1637), .Y(n1638) );
  AND3X1 U1587 ( .A(mempsack), .B(n1624), .C(n1621), .Y(n1642) );
  INVX1 U1588 ( .A(n2155), .Y(n1643) );
  AND2X1 U1589 ( .A(n588), .B(n1582), .Y(n1583) );
  OAI22X1 U1590 ( .A(n2329), .B(n934), .C(n2320), .D(n2344), .Y(n949) );
  INVX1 U1591 ( .A(n613), .Y(n1582) );
  AOI22X1 U1592 ( .A(n816), .B(n1374), .C(ramdatai[4]), .D(n1375), .Y(n1494)
         );
  INVX1 U1593 ( .A(n816), .Y(n652) );
  AOI22X1 U1594 ( .A(n2120), .B(N13353), .C(N13346), .D(n2273), .Y(n837) );
  AOI22X1 U1595 ( .A(n191), .B(N13353), .C(N13349), .D(n2273), .Y(n834) );
  AOI22X1 U1596 ( .A(n192), .B(N13353), .C(N13350), .D(n2273), .Y(n833) );
  AOI22X1 U1597 ( .A(n193), .B(N13353), .C(N13351), .D(n2273), .Y(n831) );
  INVX1 U1598 ( .A(n635), .Y(n860) );
  NAND21X1 U1599 ( .B(n2237), .A(n859), .Y(n635) );
  AOI22X1 U1600 ( .A(n189), .B(N13353), .C(N13347), .D(n2273), .Y(n836) );
  AOI22X1 U1601 ( .A(n190), .B(N13353), .C(N13348), .D(n2273), .Y(n835) );
  INVX1 U1602 ( .A(n2141), .Y(n638) );
  INVX1 U1603 ( .A(n2125), .Y(n643) );
  INVX1 U1604 ( .A(n684), .Y(n634) );
  OAI22X1 U1605 ( .A(n933), .B(n909), .C(n1373), .D(n910), .Y(n932) );
  OAI22X1 U1606 ( .A(n923), .B(n909), .C(n686), .D(n910), .Y(n922) );
  OAI22X1 U1607 ( .A(n908), .B(n909), .C(n2285), .D(n910), .Y(n907) );
  OR2X1 U1608 ( .A(n2230), .B(n650), .Y(n728) );
  NAND21X1 U1609 ( .B(n2226), .A(n824), .Y(n1992) );
  INVX1 U1610 ( .A(n2122), .Y(n665) );
  INVX1 U1611 ( .A(n2123), .Y(n653) );
  INVX1 U1612 ( .A(n2124), .Y(n648) );
  INVX1 U1613 ( .A(n1579), .Y(n1581) );
  MUX2X1 U1614 ( .D0(n2473), .D1(n2289), .S(n1957), .Y(n2178) );
  INVX1 U1615 ( .A(n235), .Y(n2467) );
  NAND3X1 U1616 ( .A(dpc[1]), .B(n2306), .C(n2303), .Y(n1134) );
  NAND3X1 U1617 ( .A(dpc[1]), .B(dpc[2]), .C(n2303), .Y(n1132) );
  NAND2X1 U1618 ( .A(n2263), .B(dpc[0]), .Y(n1170) );
  INVX1 U1619 ( .A(pc_i[11]), .Y(n2451) );
  INVX1 U1620 ( .A(pc_i[13]), .Y(n705) );
  OAI31XL U1621 ( .A(n1496), .B(n2230), .C(n1497), .D(n1498), .Y(n1375) );
  AOI221XL U1622 ( .A(n1135), .B(n48), .C(n1290), .D(n42), .E(n1170), .Y(n1300) );
  AOI221XL U1623 ( .A(n2462), .B(n48), .C(n1269), .D(n43), .E(n1170), .Y(n1278) );
  OAI211X1 U1624 ( .C(n235), .D(n2305), .A(n1278), .B(n1279), .Y(n1276) );
  AOI22X1 U1625 ( .A(n2302), .B(n1280), .C(n48), .D(n235), .Y(n1279) );
  INVX1 U1626 ( .A(n1090), .Y(n2263) );
  NOR2X1 U1627 ( .A(n154), .B(n2445), .Y(N14351) );
  NOR2X1 U1628 ( .A(n2477), .B(n2486), .Y(N14346) );
  NOR2X1 U1629 ( .A(n2477), .B(n2485), .Y(N14347) );
  NOR2X1 U1630 ( .A(n154), .B(n2474), .Y(N14348) );
  NOR2X1 U1631 ( .A(n154), .B(n2471), .Y(N14349) );
  NOR2X1 U1632 ( .A(n154), .B(n2470), .Y(N14350) );
  NOR2X1 U1633 ( .A(n2477), .B(n2488), .Y(N14345) );
  MUX2X1 U1634 ( .D0(n2403), .D1(n2286), .S(n1957), .Y(n659) );
  MUX2X1 U1635 ( .D0(n2406), .D1(n2318), .S(n1957), .Y(n697) );
  NAND21X1 U1636 ( .B(n2226), .A(n823), .Y(n1439) );
  OAI21X1 U1637 ( .B(n2460), .C(n1134), .A(n2303), .Y(n1200) );
  OAI211X1 U1638 ( .C(n1231), .D(n2305), .A(n2303), .B(n1243), .Y(n1233) );
  AOI21X1 U1639 ( .B(n48), .C(n1244), .A(n1245), .Y(n1243) );
  AOI21X1 U1640 ( .B(n2455), .C(n46), .A(n1134), .Y(n1245) );
  OAI21X1 U1641 ( .B(n1191), .C(n37), .A(n1180), .Y(n1190) );
  AOI211X1 U1642 ( .C(n43), .D(n40), .A(n1258), .B(n2296), .Y(n1252) );
  OAI22X1 U1643 ( .A(n40), .B(n1132), .C(n2455), .D(n153), .Y(n1258) );
  INVX1 U1644 ( .A(n1259), .Y(n2296) );
  AOI21X1 U1645 ( .B(n1192), .C(n1202), .A(n1134), .Y(n1201) );
  NOR3XL U1646 ( .A(dpc[1]), .B(dpc[2]), .C(n1170), .Y(n1127) );
  OA21X1 U1647 ( .B(n1215), .C(n2460), .A(n1216), .Y(n1110) );
  OAI21X1 U1648 ( .B(n110), .C(n86), .A(n2460), .Y(n1216) );
  NOR21XL U1649 ( .B(n1209), .A(n1170), .Y(n1215) );
  AND2X1 U1650 ( .A(n1133), .B(n2468), .Y(n1130) );
  INVX1 U1651 ( .A(n1286), .Y(n2299) );
  AO2222XL U1652 ( .A(n86), .B(pc_i[10]), .C(n2458), .D(n110), .E(memaddr[10]), 
        .F(n1287), .G(n1288), .H(n2467), .Y(n1286) );
  INVX1 U1653 ( .A(n1280), .Y(n2458) );
  OAI22X1 U1654 ( .A(n2305), .B(n1269), .C(n37), .D(n2462), .Y(n1288) );
  AOI211X1 U1655 ( .C(n2063), .D(n613), .A(n906), .B(n1614), .Y(n1615) );
  INVX1 U1656 ( .A(n909), .Y(n1614) );
  NAND4X1 U1657 ( .A(n2107), .B(n2108), .C(n2109), .D(n2110), .Y(n2063) );
  AOI221XL U1658 ( .A(n2048), .B(n2112), .C(n2379), .D(n746), .E(n2113), .Y(
        n2109) );
  NAND2X1 U1659 ( .A(n1191), .B(n2460), .Y(n1192) );
  NAND2X1 U1660 ( .A(n1130), .B(n53), .Y(n1302) );
  NAND2X1 U1661 ( .A(n1289), .B(n2467), .Y(n1280) );
  NAND2X1 U1662 ( .A(n1268), .B(n40), .Y(n1255) );
  MUX2IX1 U1663 ( .D0(n2475), .D1(n2321), .S(n1957), .Y(n204) );
  NOR2X1 U1664 ( .A(n2465), .B(n1202), .Y(n1430) );
  OAI22X1 U1665 ( .A(n2330), .B(n934), .C(n2317), .D(n2344), .Y(n942) );
  OAI21X1 U1666 ( .B(n1289), .C(n153), .A(n1278), .Y(n1287) );
  AOI21X1 U1667 ( .B(n1132), .C(n153), .A(n2464), .Y(n1234) );
  XNOR2XL U1668 ( .A(n2468), .B(n1422), .Y(n1125) );
  NOR2X1 U1669 ( .A(n1311), .B(n57), .Y(n1422) );
  INVX1 U1670 ( .A(n1167), .Y(n2459) );
  XNOR2XL U1671 ( .A(n55), .B(n1430), .Y(n1177) );
  NOR3XL U1672 ( .A(n2467), .B(n2453), .C(n1269), .Y(n1257) );
  INVX1 U1673 ( .A(pc_i[4]), .Y(n649) );
  INVX1 U1674 ( .A(pc_i[5]), .Y(n703) );
  AND2X1 U1675 ( .A(n1156), .B(n57), .Y(n1131) );
  NAND2X1 U1676 ( .A(n1131), .B(n2468), .Y(n1135) );
  AND2X1 U1677 ( .A(n1179), .B(n55), .Y(n1169) );
  AND2X1 U1678 ( .A(n1191), .B(n2465), .Y(n1179) );
  AND2X1 U1679 ( .A(n1169), .B(n49), .Y(n1156) );
  NOR3XL U1680 ( .A(n40), .B(n46), .C(n2452), .Y(n1231) );
  INVX1 U1681 ( .A(pc_i[15]), .Y(n2373) );
  XNOR2XL U1682 ( .A(n2465), .B(n1202), .Y(n205) );
  NAND3X1 U1683 ( .A(n40), .B(n46), .C(n1256), .Y(n1244) );
  NAND3X1 U1684 ( .A(n1043), .B(n1044), .C(n2351), .Y(n1042) );
  INVX1 U1685 ( .A(n1291), .Y(n2462) );
  INVX1 U1686 ( .A(pc_o[1]), .Y(n2466) );
  NOR2X1 U1687 ( .A(n977), .B(n953), .Y(n983) );
  NAND3X1 U1688 ( .A(n953), .B(n976), .C(n999), .Y(n986) );
  INVX1 U1689 ( .A(n1588), .Y(n1563) );
  INVX1 U1690 ( .A(n984), .Y(n2349) );
  NAND4X1 U1691 ( .A(n1023), .B(n2490), .C(n2488), .D(n2486), .Y(n1021) );
  INVX1 U1692 ( .A(n980), .Y(n2346) );
  INVX1 U1693 ( .A(n1256), .Y(n2454) );
  INVX1 U1694 ( .A(dpc[2]), .Y(n2306) );
  NOR32XL U1695 ( .B(n952), .C(n953), .A(n954), .Y(n913) );
  NOR43XL U1696 ( .B(n952), .C(n954), .D(n953), .A(n911), .Y(n912) );
  OAI211X1 U1697 ( .C(n2428), .D(n1647), .A(n1003), .B(n1004), .Y(n1001) );
  NAND3X1 U1698 ( .A(n1005), .B(n128), .C(n1006), .Y(n1003) );
  NAND32X1 U1699 ( .B(n2187), .C(n631), .A(n1002), .Y(n1503) );
  NOR3XL U1700 ( .A(n259), .B(n292), .C(n2378), .Y(n1002) );
  INVX1 U1701 ( .A(n999), .Y(n631) );
  AND4X1 U1702 ( .A(n934), .B(n909), .C(n958), .D(n945), .Y(n952) );
  AND2X1 U1703 ( .A(n910), .B(n2271), .Y(n958) );
  NAND2X1 U1704 ( .A(n691), .B(n128), .Y(n910) );
  AOI22X1 U1705 ( .A(n969), .B(n970), .C(n971), .D(n751), .Y(n968) );
  AOI22X1 U1706 ( .A(n969), .B(n2428), .C(n973), .D(n147), .Y(n966) );
  AOI21X1 U1707 ( .B(n774), .C(n751), .A(n963), .Y(n962) );
  INVX1 U1708 ( .A(n953), .Y(n2359) );
  OAI21X1 U1709 ( .B(n128), .C(n2428), .A(n603), .Y(n599) );
  OAI22X1 U1710 ( .A(n2315), .B(n261), .C(n170), .D(n602), .Y(n600) );
  NOR21XL U1711 ( .B(n2232), .A(n128), .Y(n911) );
  AOI222XL U1712 ( .A(n760), .B(n1635), .C(n1736), .D(n1625), .E(n963), .F(
        n2114), .Y(n2108) );
  INVX1 U1713 ( .A(n934), .Y(n1402) );
  AOI21X1 U1714 ( .B(n2383), .C(n2052), .A(n2450), .Y(n2113) );
  NOR32XL U1715 ( .B(n853), .C(n1364), .A(n2189), .Y(n1347) );
  NAND2X1 U1716 ( .A(n1727), .B(n2030), .Y(n2048) );
  NOR3XL U1717 ( .A(n2425), .B(n109), .C(n809), .Y(n207) );
  NAND2X1 U1718 ( .A(n871), .B(n287), .Y(n870) );
  OAI22X1 U1719 ( .A(n2192), .B(n870), .C(n2372), .D(n869), .Y(N12967) );
  OAI22X1 U1720 ( .A(n2208), .B(n870), .C(n2371), .D(n869), .Y(N12971) );
  NAND3X1 U1721 ( .A(n2470), .B(n2445), .C(n2471), .Y(n1022) );
  INVX1 U1722 ( .A(n855), .Y(n2441) );
  INVX1 U1723 ( .A(n483), .Y(cs_run) );
  AND2X1 U1724 ( .A(n2205), .B(n11), .Y(n1700) );
  MUX2XL U1725 ( .D0(pc_o[3]), .D1(n1716), .S(n15), .Y(memaddr_comb[3]) );
  OAI21AX1 U1726 ( .B(sfroe_r), .C(sfrwe_r), .A(sfrack), .Y(n1624) );
  MUX2XL U1727 ( .D0(n2502), .D1(n1717), .S(n14), .Y(memaddr_comb[4]) );
  NAND4X1 U1728 ( .A(n531), .B(n532), .C(n533), .D(n534), .Y(dpl[2]) );
  AOI22X1 U1729 ( .A(n224), .B(dpl_reg[42]), .C(n226), .D(dpl_reg[58]), .Y(
        n531) );
  NAND2X1 U1730 ( .A(cpu_hold), .B(n613), .Y(n208) );
  NAND4X1 U1731 ( .A(n523), .B(n524), .C(n525), .D(n526), .Y(dpl[4]) );
  NAND4X1 U1732 ( .A(n555), .B(n556), .C(n557), .D(n558), .Y(dph[4]) );
  AOI22X1 U1733 ( .A(n223), .B(dpl_reg[44]), .C(n225), .D(dpl_reg[60]), .Y(
        n523) );
  NAND4X1 U1734 ( .A(n519), .B(n520), .C(n521), .D(n522), .Y(dpl[5]) );
  NAND4X1 U1735 ( .A(n551), .B(n552), .C(n553), .D(n554), .Y(dph[5]) );
  AOI22X1 U1736 ( .A(n224), .B(dpl_reg[45]), .C(n226), .D(dpl_reg[61]), .Y(
        n519) );
  NAND4X1 U1737 ( .A(n563), .B(n564), .C(n565), .D(n566), .Y(dph[2]) );
  AOI22X1 U1738 ( .A(n513), .B(dph_reg[42]), .C(n514), .D(dph_reg[58]), .Y(
        n563) );
  AOI22X1 U1739 ( .A(n231), .B(dph_reg[10]), .C(n27), .D(dph_reg[26]), .Y(n565) );
  NOR32XL U1740 ( .B(n1746), .C(acc[1]), .A(n944), .Y(n472) );
  NOR21XL U1741 ( .B(n151), .A(n1710), .Y(n360) );
  NOR32XL U1742 ( .B(acc[0]), .C(n1746), .A(n951), .Y(n381) );
  NAND21X1 U1743 ( .B(n377), .A(n376), .Y(n378) );
  NAND4X1 U1744 ( .A(n515), .B(n516), .C(n517), .D(n518), .Y(dpl[6]) );
  NAND4X1 U1745 ( .A(n547), .B(n548), .C(n549), .D(n550), .Y(dph[6]) );
  NAND4X1 U1746 ( .A(n543), .B(n544), .C(n545), .D(n546), .Y(dph[7]) );
  AOI22X1 U1747 ( .A(n224), .B(dph_reg[47]), .C(n226), .D(dph_reg[63]), .Y(
        n543) );
  NAND4X1 U1748 ( .A(n535), .B(n536), .C(n537), .D(n538), .Y(dpl[1]) );
  AOI22X1 U1749 ( .A(n223), .B(dpl_reg[41]), .C(n225), .D(dpl_reg[57]), .Y(
        n535) );
  NAND4X1 U1750 ( .A(n527), .B(n528), .C(n529), .D(n530), .Y(dpl[3]) );
  AOI22X1 U1751 ( .A(n513), .B(dpl_reg[43]), .C(n514), .D(dpl_reg[59]), .Y(
        n527) );
  AND2X1 U1752 ( .A(sfrwe_r), .B(n2500), .Y(sfrwe) );
  NAND4X1 U1753 ( .A(n567), .B(n568), .C(n569), .D(n570), .Y(dph[1]) );
  AOI22X1 U1754 ( .A(n224), .B(dph_reg[41]), .C(n226), .D(dph_reg[57]), .Y(
        n567) );
  AOI22X1 U1755 ( .A(n24), .B(dph_reg[9]), .C(n27), .D(dph_reg[25]), .Y(n569)
         );
  NAND4X1 U1756 ( .A(n559), .B(n560), .C(n561), .D(n562), .Y(dph[3]) );
  AOI22X1 U1757 ( .A(n223), .B(dph_reg[43]), .C(n225), .D(dph_reg[59]), .Y(
        n559) );
  AOI22X1 U1758 ( .A(n509), .B(dph_reg[11]), .C(n26), .D(dph_reg[27]), .Y(n561) );
  NAND4X1 U1759 ( .A(n571), .B(n572), .C(n573), .D(n574), .Y(dph[0]) );
  NAND4X1 U1760 ( .A(n539), .B(n540), .C(n541), .D(n542), .Y(dpl[0]) );
  AOI22X1 U1761 ( .A(n223), .B(dph_reg[40]), .C(n225), .D(dph_reg[56]), .Y(
        n571) );
  MUX2XL U1762 ( .D0(pc_o[7]), .D1(n1720), .S(n15), .Y(memaddr_comb[7]) );
  MUX2X1 U1763 ( .D0(pc_o[11]), .D1(n1729), .S(n283), .Y(memaddr_comb[11]) );
  MUX2XL U1764 ( .D0(pc_o[8]), .D1(n1721), .S(n15), .Y(memaddr_comb[8]) );
  MUX2X1 U1765 ( .D0(pc_o[12]), .D1(n1730), .S(n283), .Y(memaddr_comb[12]) );
  MUX2XL U1766 ( .D0(pc_o[9]), .D1(n1724), .S(n15), .Y(memaddr_comb[9]) );
  AO2222XL U1767 ( .A(alu_out[12]), .B(n75), .C(n2123), .D(n221), .E(pc_i[12]), 
        .F(n185), .G(n664), .H(temp[4]), .Y(n647) );
  AO2222XL U1768 ( .A(alu_out[11]), .B(n75), .C(n2122), .D(n220), .E(pc_i[11]), 
        .F(n185), .G(n664), .H(temp[3]), .Y(n637) );
  NAND43X1 U1769 ( .B(n409), .C(n408), .D(n407), .A(n406), .Y(n812) );
  OAI22X1 U1770 ( .A(n1486), .B(n2477), .C(n1393), .D(n2203), .Y(n409) );
  OA222X1 U1771 ( .A(n2475), .B(n2334), .C(n1676), .D(n1450), .E(n1049), .F(
        n2484), .Y(n406) );
  AO21X1 U1772 ( .B(n1357), .C(acc[4]), .A(n405), .Y(n407) );
  MUX2BXL U1773 ( .D0(ramwe), .D1(n210), .S(waitstaten), .Y(ramwe_comb) );
  AOI21X1 U1774 ( .B(n1654), .C(n1653), .A(n1652), .Y(n210) );
  MUX2X1 U1775 ( .D0(memrd), .D1(n1701), .S(n283), .Y(memrd_comb) );
  MUX2XL U1776 ( .D0(ramoe), .D1(n1655), .S(waitstaten), .Y(ramoe_comb) );
  NAND21X1 U1777 ( .B(n903), .A(n898), .Y(n1715) );
  OA2222XL U1778 ( .A(n781), .B(n897), .C(n2440), .D(n1371), .E(n938), .F(
        n1369), .G(n2345), .H(n2493), .Y(n898) );
  AO2222XL U1779 ( .A(alu_out[2]), .B(n1407), .C(n2142), .D(n1126), .E(n1341), 
        .F(n2503), .G(pc_i[2]), .H(n1334), .Y(n903) );
  INVX1 U1780 ( .A(memdatai[2]), .Y(n897) );
  NAND21X1 U1781 ( .B(n677), .A(n676), .Y(n1718) );
  OA2222XL U1782 ( .A(n781), .B(n686), .C(n702), .D(n1371), .E(n923), .F(n1369), .G(n2345), .H(n1954), .Y(n676) );
  AO2222XL U1783 ( .A(alu_out[5]), .B(n1407), .C(n220), .D(n1012), .E(n1341), 
        .F(n50), .G(pc_i[5]), .H(n1334), .Y(n677) );
  NAND21X1 U1784 ( .B(n1381), .A(n1380), .Y(n1716) );
  OA2222XL U1785 ( .A(n781), .B(n1373), .C(n2438), .D(n1371), .E(n933), .F(
        n1369), .G(n2345), .H(n2492), .Y(n1380) );
  AO2222XL U1786 ( .A(alu_out[3]), .B(n1407), .C(n221), .D(n1368), .E(n1341), 
        .F(pc_o[3]), .G(pc_i[3]), .H(n1334), .Y(n1381) );
  NAND21X1 U1787 ( .B(n630), .A(n629), .Y(n1717) );
  OA2222XL U1788 ( .A(n781), .B(n670), .C(n669), .D(n1371), .E(n928), .F(n1369), .G(n2345), .H(n654), .Y(n629) );
  AO2222XL U1789 ( .A(alu_out[4]), .B(n1407), .C(n221), .D(n1020), .E(n1341), 
        .F(n2502), .G(pc_i[4]), .H(n1334), .Y(n630) );
  ENOX1 U1790 ( .A(n2489), .B(n2274), .C(N13336), .D(n2274), .Y(n2120) );
  OAI21X1 U1791 ( .B(n2287), .C(n2396), .A(n802), .Y(n801) );
  AOI33X1 U1792 ( .A(instr[5]), .B(n128), .C(n2312), .D(instr[4]), .E(n147), 
        .F(n2287), .Y(n802) );
  INVX1 U1793 ( .A(n804), .Y(n2287) );
  INVX1 U1794 ( .A(n803), .Y(n2312) );
  MUX2X1 U1795 ( .D0(pc_o[13]), .D1(n1731), .S(n283), .Y(memaddr_comb[13]) );
  MUX2X1 U1796 ( .D0(pc_o[14]), .D1(n1732), .S(n283), .Y(memaddr_comb[14]) );
  AO2222XL U1797 ( .A(alu_out[13]), .B(n75), .C(n2124), .D(n220), .E(pc_i[13]), 
        .F(n185), .G(n664), .H(temp[5]), .Y(n683) );
  AO2222XL U1798 ( .A(alu_out[14]), .B(n75), .C(n2125), .D(n220), .E(pc_i[14]), 
        .F(n185), .G(n664), .H(temp[6]), .Y(n931) );
  MUX2X1 U1799 ( .D0(n815), .D1(temp[3]), .S(n982), .Y(N12827) );
  MUX2X1 U1800 ( .D0(pc_o[3]), .D1(n1368), .S(n899), .Y(N12844) );
  MUX2X1 U1801 ( .D0(memaddr[4]), .D1(n1020), .S(n899), .Y(N12845) );
  MUX2X1 U1802 ( .D0(n816), .D1(temp[4]), .S(n982), .Y(N12828) );
  MUX2X1 U1803 ( .D0(pc_o[5]), .D1(n1012), .S(n899), .Y(N12846) );
  MUX2X1 U1804 ( .D0(n817), .D1(temp[5]), .S(n982), .Y(N12829) );
  MUX2X1 U1805 ( .D0(memaddr[11]), .D1(n2122), .S(n89), .Y(N12852) );
  MUX2X1 U1806 ( .D0(n814), .D1(temp[2]), .S(n982), .Y(N12826) );
  MUX2X1 U1807 ( .D0(memaddr[2]), .D1(n1126), .S(n899), .Y(N12843) );
  MUX2X1 U1808 ( .D0(pc_o[12]), .D1(n2123), .S(n89), .Y(N12853) );
  MUX2X1 U1809 ( .D0(pc_o[13]), .D1(n2124), .S(n89), .Y(N12854) );
  MUX2X1 U1810 ( .D0(pc_o[7]), .D1(n995), .S(n899), .Y(N12848) );
  AO21X1 U1811 ( .B(n2313), .C(n900), .A(n2235), .Y(N12831) );
  MUX2X1 U1812 ( .D0(memaddr[8]), .D1(n993), .S(n899), .Y(N12849) );
  MUX2X1 U1813 ( .D0(memaddr[9]), .D1(n991), .S(n89), .Y(N12850) );
  MUX2X1 U1814 ( .D0(n813), .D1(temp[1]), .S(n982), .Y(N12825) );
  MUX2X1 U1815 ( .D0(pc_o[1]), .D1(n1187), .S(n899), .Y(N12842) );
  MUX2X1 U1816 ( .D0(memaddr[6]), .D1(n997), .S(n899), .Y(N12847) );
  MUX2X1 U1817 ( .D0(n818), .D1(temp[6]), .S(n982), .Y(N12830) );
  MUX2X1 U1818 ( .D0(memaddr[14]), .D1(n2125), .S(n89), .Y(N12855) );
  MUX2X1 U1819 ( .D0(n812), .D1(temp[0]), .S(n982), .Y(N12824) );
  AO22X1 U1820 ( .A(divtempreg[0]), .B(N13343), .C(N13337), .D(n2274), .Y(n189) );
  NAND21X1 U1821 ( .B(n828), .A(n827), .Y(n1713) );
  OA2222XL U1822 ( .A(n781), .B(n826), .C(n825), .D(n1371), .E(n951), .F(n1369), .G(n2345), .H(n2495), .Y(n827) );
  AO2222XL U1823 ( .A(alu_out[0]), .B(n1407), .C(n221), .D(n1228), .E(n1341), 
        .F(pc_o[0]), .G(n1334), .H(pc_i[0]), .Y(n828) );
  NAND21X1 U1824 ( .B(n715), .A(n714), .Y(n1719) );
  OA2222XL U1825 ( .A(n781), .B(n734), .C(n2358), .D(n1371), .E(n918), .F(
        n1369), .G(n2345), .H(n2491), .Y(n714) );
  AO2222XL U1826 ( .A(alu_out[6]), .B(n1407), .C(n221), .D(n997), .E(n1341), 
        .F(pc_o[6]), .G(pc_i[6]), .H(n1334), .Y(n715) );
  AO2222XL U1827 ( .A(alu_out[15]), .B(n75), .C(n2141), .D(n221), .E(pc_i[15]), 
        .F(n185), .G(n664), .H(temp[7]), .Y(n741) );
  MUX2X1 U1828 ( .D0(pc_o[15]), .D1(n2141), .S(n89), .Y(N12856) );
  MUX2X1 U1829 ( .D0(mempsrd), .D1(n1711), .S(n283), .Y(mempsrd_comb) );
  AO21X1 U1830 ( .B(n1709), .C(n1708), .A(n1707), .Y(n1711) );
  MUX2X1 U1831 ( .D0(pc_o[15]), .D1(n1733), .S(n284), .Y(memaddr_comb[15]) );
  AO22X1 U1832 ( .A(divtempreg[1]), .B(N13343), .C(N13338), .D(n2274), .Y(n190) );
  AO22X1 U1833 ( .A(divtempreg[2]), .B(N13343), .C(N13339), .D(n2274), .Y(n191) );
  NAND21X1 U1834 ( .B(n1432), .A(n1426), .Y(n1728) );
  OA2222XL U1835 ( .A(n2467), .B(n1424), .C(n2093), .D(n672), .E(n2192), .F(
        n1418), .G(n1412), .H(n1411), .Y(n1426) );
  AO2222XL U1836 ( .A(n2232), .B(instr[7]), .C(alu_out[10]), .D(n75), .E(n664), 
        .F(temp[2]), .G(pc_i[10]), .H(n2198), .Y(n1432) );
  AND3X1 U1837 ( .A(n1377), .B(n1378), .C(n1379), .Y(n456) );
  AOI222XL U1838 ( .A(pc_i[15]), .B(n2240), .C(pc_o[7]), .D(n2247), .E(n2246), 
        .F(temp2_comb[7]), .Y(n1378) );
  AOI221XL U1839 ( .A(pc_o[15]), .B(n411), .C(pc_i[7]), .D(n2239), .E(n1382), 
        .Y(n1379) );
  AOI22X1 U1840 ( .A(n2249), .B(n1125), .C(n1413), .D(n1414), .Y(n1377) );
  XNOR2XL U1841 ( .A(acc[3]), .B(n1365), .Y(N11544) );
  AO21X1 U1842 ( .B(n2481), .C(temp2_comb[3]), .A(n1366), .Y(N11525) );
  NOR43XL U1843 ( .B(n1386), .C(n1387), .D(n1388), .A(n1389), .Y(n1376) );
  AOI22X1 U1844 ( .A(n1023), .B(acc[5]), .C(n2264), .D(ramdatao[7]), .Y(n1387)
         );
  AOI222XL U1845 ( .A(c), .B(n2353), .C(n2332), .D(n2489), .E(multemp2[1]), 
        .F(n1349), .Y(n1388) );
  OAI21BX1 U1846 ( .C(temp2_comb[7]), .B(n1390), .A(n1391), .Y(n1389) );
  NAND21X1 U1847 ( .B(n501), .A(n500), .Y(n1495) );
  MUX2X1 U1848 ( .D0(cs_run), .D1(n1562), .S(codefetch_s), .Y(n501) );
  MUX2X1 U1849 ( .D0(n499), .D1(n498), .S(n1499), .Y(n500) );
  INVX1 U1850 ( .A(state[0]), .Y(n499) );
  MUX2X1 U1851 ( .D0(ramsfraddr[2]), .D1(n198), .S(n284), .Y(
        ramsfraddr_comb[2]) );
  NOR32XL U1852 ( .B(n1598), .C(dec_accop[18]), .A(dec_accop[5]), .Y(n1481) );
  NAND3X1 U1853 ( .A(n1444), .B(n1445), .C(n1446), .Y(n818) );
  AOI22X1 U1854 ( .A(n1023), .B(acc[4]), .C(n2264), .D(ramdatao[6]), .Y(n1444)
         );
  AOI222XL U1855 ( .A(acc[7]), .B(n2352), .C(n2332), .D(n2415), .E(multemp1_0_), .F(n1349), .Y(n1445) );
  AOI221XL U1856 ( .A(acc[5]), .B(n1032), .C(acc[2]), .D(n1357), .E(n1447), 
        .Y(n1446) );
  AO22X1 U1857 ( .A(divtempreg[3]), .B(N13343), .C(N13340), .D(n2274), .Y(n192) );
  MUX2X1 U1858 ( .D0(ramsfraddr[1]), .D1(n197), .S(n284), .Y(
        ramsfraddr_comb[1]) );
  MUX2X1 U1859 ( .D0(ramsfraddr[0]), .D1(n1692), .S(n284), .Y(
        ramsfraddr_comb[0]) );
  NOR2X1 U1860 ( .A(n1680), .B(dec_accop[9]), .Y(n1598) );
  NAND21X1 U1861 ( .B(n888), .A(n886), .Y(n1724) );
  OA2222XL U1862 ( .A(n51), .B(n1424), .C(n2093), .D(n678), .E(n2199), .F(
        n1418), .G(n1412), .H(n872), .Y(n886) );
  AO2222XL U1863 ( .A(instr[6]), .B(n2232), .C(alu_out[9]), .D(n75), .E(n664), 
        .F(temp[1]), .G(n2198), .H(pc_i[9]), .Y(n888) );
  INVX1 U1864 ( .A(p2[1]), .Y(n872) );
  NAND21X1 U1865 ( .B(n896), .A(n893), .Y(n1721) );
  OA2222XL U1866 ( .A(n53), .B(n1424), .C(n2093), .D(n693), .E(n2203), .F(
        n1418), .G(n1412), .H(n889), .Y(n893) );
  AO2222XL U1867 ( .A(n2232), .B(instr[5]), .C(alu_out[8]), .D(n75), .E(n664), 
        .F(temp[0]), .G(n2198), .H(pc_i[8]), .Y(n896) );
  INVX1 U1868 ( .A(p2[0]), .Y(n889) );
  INVX1 U1869 ( .A(n1597), .Y(n2472) );
  GEN2XL U1870 ( .D(n150), .E(n2476), .C(ac), .B(n1481), .A(n1366), .Y(n1597)
         );
  INVX1 U1871 ( .A(n1482), .Y(n2476) );
  AOI221XL U1872 ( .A(n2481), .B(temp2_comb[0]), .C(dec_accop[5]), .D(n1598), 
        .E(n1366), .Y(n1599) );
  NOR3XL U1873 ( .A(n2479), .B(dec_accop[5]), .C(n2483), .Y(n1366) );
  XNOR2XL U1874 ( .A(acc[2]), .B(n1365), .Y(N11543) );
  OAI21X1 U1875 ( .B(n1367), .C(n2440), .A(n2472), .Y(N11524) );
  OAI21X1 U1876 ( .B(n575), .C(n576), .A(n577), .Y(
        add_1_root_add_5140_2_carry[2]) );
  OAI222XL U1877 ( .A(n1448), .B(n2358), .C(n1449), .D(n2415), .E(n1450), .F(
        n1451), .Y(n1447) );
  AOI221XL U1878 ( .A(n2331), .B(n2415), .C(acc[6]), .D(n1360), .E(n1363), .Y(
        n1448) );
  AOI21X1 U1879 ( .B(n2331), .C(n2358), .A(n2333), .Y(n1449) );
  XNOR2XL U1880 ( .A(n1452), .B(n1399), .Y(n1451) );
  AOI222XL U1881 ( .A(n1357), .B(acc[3]), .C(n1396), .D(n2328), .E(acc[6]), 
        .F(n1032), .Y(n1386) );
  XOR2X1 U1882 ( .A(n1069), .B(n1068), .Y(n1396) );
  OAI32X1 U1883 ( .A(n1605), .B(n169), .C(n483), .D(n1592), .E(n1591), .Y(
        n1707) );
  OA21X1 U1884 ( .B(n2205), .C(n1609), .A(n2147), .Y(n1605) );
  AOI32X1 U1885 ( .A(n1590), .B(n2248), .C(n1589), .D(n1588), .E(n1587), .Y(
        n1592) );
  INVX1 U1886 ( .A(pdmode), .Y(n1589) );
  OR2X1 U1887 ( .A(dec_accop[8]), .B(dec_accop[10]), .Y(n1680) );
  OAI211X1 U1888 ( .C(n1045), .D(n1046), .A(n1047), .B(n1048), .Y(n804) );
  AOI22AXL U1889 ( .A(n2353), .B(acc[0]), .D(n1049), .C(acc[7]), .Y(n1048) );
  AOI22AXL U1890 ( .A(n1033), .B(n1050), .D(n1051), .C(c), .Y(n1047) );
  XNOR2XL U1891 ( .A(n1067), .B(n1036), .Y(n1046) );
  AO22X1 U1892 ( .A(divtempreg[4]), .B(N13343), .C(N13341), .D(n2274), .Y(n193) );
  AO22X1 U1893 ( .A(divtempreg[5]), .B(N13343), .C(N13342), .D(n2274), .Y(n194) );
  INVX1 U1894 ( .A(acc[0]), .Y(n2478) );
  NAND4X1 U1895 ( .A(n1681), .B(n2480), .C(n1682), .D(n2479), .Y(n1365) );
  NOR2X1 U1896 ( .A(dec_accop[8]), .B(dec_accop[7]), .Y(n1682) );
  NAND21X1 U1897 ( .B(n914), .A(n905), .Y(n1720) );
  OA2222XL U1898 ( .A(n781), .B(n2285), .C(n920), .D(n1371), .E(n908), .F(
        n1369), .G(n2345), .H(n904), .Y(n905) );
  AO2222XL U1899 ( .A(alu_out[7]), .B(n1407), .C(n220), .D(n995), .E(n1341), 
        .F(pc_o[7]), .G(pc_i[7]), .H(n1334), .Y(n914) );
  NAND2X1 U1900 ( .A(n1512), .B(n1513), .Y(n816) );
  AOI221XL U1901 ( .A(acc[2]), .B(n1023), .C(n2264), .D(ramdatao[4]), .E(n1519), .Y(n1512) );
  AOI221XL U1902 ( .A(acc[3]), .B(n1032), .C(n1357), .D(acc[0]), .E(n1514), 
        .Y(n1513) );
  OAI222XL U1903 ( .A(n2415), .B(n2334), .C(acc[4]), .D(n1359), .E(n1486), .F(
        n2406), .Y(n1519) );
  NOR2X1 U1904 ( .A(acc[2]), .B(acc[1]), .Y(n1482) );
  OAI222XL U1905 ( .A(n1515), .B(n669), .C(n1516), .D(n2403), .E(n1450), .F(
        n1517), .Y(n1514) );
  AOI221XL U1906 ( .A(n2331), .B(n2403), .C(acc[4]), .D(n1360), .E(n1363), .Y(
        n1515) );
  AOI21X1 U1907 ( .B(n134), .C(n669), .A(n2333), .Y(n1516) );
  XNOR2XL U1908 ( .A(n1518), .B(n2404), .Y(n1517) );
  OAI222XL U1909 ( .A(n1475), .B(n702), .C(n1476), .D(n2406), .E(n1450), .F(
        n1477), .Y(n1474) );
  AOI221XL U1910 ( .A(n2331), .B(n2406), .C(acc[5]), .D(n1360), .E(n1363), .Y(
        n1475) );
  AOI21X1 U1911 ( .B(n2331), .C(n702), .A(n2333), .Y(n1476) );
  XOR2X1 U1912 ( .A(n1455), .B(n1478), .Y(n1477) );
  NAND2X1 U1913 ( .A(n1472), .B(n1473), .Y(n817) );
  AOI221XL U1914 ( .A(n1023), .B(acc[3]), .C(n2264), .D(ramdatao[5]), .E(n1485), .Y(n1472) );
  AOI221XL U1915 ( .A(acc[4]), .B(n1032), .C(acc[1]), .D(n1357), .E(n1474), 
        .Y(n1473) );
  OAI222XL U1916 ( .A(n2489), .B(n2334), .C(acc[5]), .D(n1359), .E(n1486), .F(
        n2415), .Y(n1485) );
  NOR2X1 U1917 ( .A(dec_accop[5]), .B(dec_accop[18]), .Y(n1681) );
  INVX1 U1918 ( .A(dec_accop[6]), .Y(n2479) );
  INVX1 U1919 ( .A(dec_accop[16]), .Y(n2480) );
  XNOR2XL U1920 ( .A(n1679), .B(n1365), .Y(n1602) );
  NAND2X1 U1921 ( .A(c), .B(n1680), .Y(n1679) );
  INVX1 U1922 ( .A(n733), .Y(n1687) );
  NAND41X1 U1923 ( .D(n732), .A(n1428), .B(n1425), .C(n1427), .Y(n733) );
  AOI22X1 U1924 ( .A(pc_o[14]), .B(n411), .C(pc_i[6]), .D(n2239), .Y(n1425) );
  AOI222XL U1925 ( .A(pc_i[14]), .B(n2240), .C(pc_o[6]), .D(n2247), .E(n2246), 
        .F(temp2_comb[6]), .Y(n1428) );
  NAND21X1 U1926 ( .B(instr[6]), .A(n2186), .Y(n2450) );
  NOR32XL U1927 ( .B(n2236), .C(ramsfraddr[6]), .A(n842), .Y(n1364) );
  NAND21X1 U1928 ( .B(n2187), .A(ramsfrwe), .Y(n1737) );
  NOR2X1 U1929 ( .A(n2507), .B(instr[2]), .Y(n788) );
  AO222X1 U1930 ( .A(n411), .B(pc_o[12]), .C(pc_i[12]), .D(n2240), .E(n1521), 
        .F(n1414), .Y(n667) );
  OAI21BBX1 U1931 ( .A(accactv), .B(dec_accop[1]), .C(n1044), .Y(n1603) );
  INVX1 U1932 ( .A(n2505), .Y(n2243) );
  INVX1 U1933 ( .A(n2504), .Y(n2186) );
  INVX1 U1934 ( .A(instr[1]), .Y(n2262) );
  INVX1 U1935 ( .A(acc[1]), .Y(n2477) );
  NOR2X1 U1936 ( .A(n2262), .B(n2509), .Y(n1005) );
  NAND3X1 U1937 ( .A(n850), .B(n1364), .C(ramsfraddr[5]), .Y(n1393) );
  AOI211X1 U1938 ( .C(accactv), .D(dec_accop[6]), .A(n1675), .B(n2350), .Y(
        n1672) );
  INVX1 U1939 ( .A(ramsfraddr[7]), .Y(n2187) );
  INVX1 U1940 ( .A(temp2_comb[1]), .Y(n2469) );
  NAND3X1 U1941 ( .A(n2336), .B(dec_accop[18]), .C(n1362), .Y(n1353) );
  NAND43X1 U1942 ( .B(ramsfraddr[7]), .C(ramsfraddr[5]), .D(ramsfraddr[6]), 
        .A(n331), .Y(n1787) );
  AND4X1 U1943 ( .A(n2016), .B(ramwe), .C(n2014), .D(n2015), .Y(n331) );
  XNOR2XL U1944 ( .A(n2357), .B(ramsfraddr[4]), .Y(n2015) );
  XNOR2XL U1945 ( .A(n2377), .B(ramsfraddr[3]), .Y(n2014) );
  AO2222XL U1946 ( .A(ramsfraddr[7]), .B(n439), .C(temp[7]), .D(n438), .E(
        n2197), .F(n437), .G(n1985), .H(n502), .Y(n579) );
  INVX1 U1947 ( .A(n1782), .Y(n437) );
  INVX1 U1948 ( .A(n1780), .Y(n439) );
  INVX1 U1949 ( .A(n1781), .Y(n438) );
  NAND21X1 U1950 ( .B(n2432), .A(n2504), .Y(n2430) );
  NOR43XL U1951 ( .B(n1354), .C(n1355), .D(n1356), .A(n1357), .Y(n1043) );
  AOI21X1 U1952 ( .B(dec_accop[14]), .C(n1362), .A(n1363), .Y(n1354) );
  NOR42XL U1953 ( .C(n1358), .D(n1359), .A(n1360), .B(n1361), .Y(n1355) );
  AOI21X1 U1954 ( .B(n2481), .C(temp2_comb[4]), .A(n1366), .Y(n1458) );
  NAND4X1 U1955 ( .A(n1923), .B(n1924), .C(n1925), .D(n1926), .Y(n1907) );
  NAND4X1 U1956 ( .A(n1915), .B(n1916), .C(n1917), .D(n1918), .Y(n1909) );
  NAND4X1 U1957 ( .A(n1919), .B(n1920), .C(n1921), .D(n1922), .Y(n1908) );
  NAND4X1 U1958 ( .A(n1818), .B(n1819), .C(n1820), .D(n1821), .Y(n1783) );
  NAND4X1 U1959 ( .A(n1800), .B(n1801), .C(n1802), .D(n1803), .Y(n1785) );
  NAND4X1 U1960 ( .A(n1813), .B(n1814), .C(n1815), .D(n1816), .Y(n1784) );
  OAI221X1 U1961 ( .A(n2407), .B(n1780), .C(n2361), .D(n1038), .E(n1906), .Y(
        n879) );
  INVX1 U1962 ( .A(ramsfraddr[3]), .Y(n2407) );
  OA222X1 U1963 ( .A(n2289), .B(n1781), .C(n1075), .D(n2340), .E(n933), .F(
        n1782), .Y(n1906) );
  MUX2XL U1964 ( .D0(n2501), .D1(n1664), .S(n2500), .Y(ramdatao_comb[3]) );
  NOR2X1 U1965 ( .A(n2262), .B(n2507), .Y(n1775) );
  MUX2X1 U1966 ( .D0(n1359), .D1(n1594), .S(acc[1]), .Y(n457) );
  AOI21X1 U1967 ( .B(n134), .C(n2469), .A(n2333), .Y(n1594) );
  MUX2X1 U1968 ( .D0(n2332), .D1(n1670), .S(acc[0]), .Y(n405) );
  OAI21X1 U1969 ( .B(temp2_comb[0]), .C(n1356), .A(n1395), .Y(n1670) );
  AO21X1 U1970 ( .B(n402), .C(n401), .A(n825), .Y(n403) );
  INVX1 U1971 ( .A(n1363), .Y(n401) );
  MUX2X1 U1972 ( .D0(n1356), .D1(n400), .S(acc[0]), .Y(n402) );
  INVX1 U1973 ( .A(n1360), .Y(n400) );
  NOR2X1 U1974 ( .A(ramsfraddr[4]), .B(ramsfraddr[3]), .Y(n850) );
  NAND41X1 U1975 ( .D(dec_accop[15]), .A(n1362), .B(n1685), .C(n1667), .Y(
        n1026) );
  NAND21X1 U1976 ( .B(dec_accop[7]), .A(n1598), .Y(n1685) );
  INVX1 U1977 ( .A(instr[6]), .Y(n2448) );
  AOI211X1 U1978 ( .C(accactv), .D(dec_accop[17]), .A(n840), .B(n1671), .Y(
        n1033) );
  OR2X1 U1979 ( .A(n1669), .B(n2337), .Y(n1671) );
  NAND3X1 U1980 ( .A(n1362), .B(n1667), .C(dec_accop[15]), .Y(n1359) );
  AND4X1 U1981 ( .A(n1898), .B(n1899), .C(n1896), .D(n1897), .Y(n349) );
  AOI22X1 U1982 ( .A(rn_reg[36]), .B(n73), .C(rn_reg[84]), .D(n87), .Y(n1898)
         );
  AOI22X1 U1983 ( .A(rn_reg[100]), .B(n120), .C(rn_reg[4]), .D(n100), .Y(n1899) );
  AOI22X1 U1984 ( .A(rn_reg[116]), .B(n161), .C(rn_reg[20]), .D(n144), .Y(
        n1897) );
  NAND3X1 U1985 ( .A(n1552), .B(n1553), .C(n1554), .Y(n815) );
  AOI22X1 U1986 ( .A(acc[1]), .B(n1023), .C(n2264), .D(n2501), .Y(n1552) );
  AOI222XL U1987 ( .A(acc[4]), .B(n2352), .C(n1349), .D(acc[5]), .E(
        adder_out[3]), .F(n2328), .Y(n1553) );
  AOI221XL U1988 ( .A(n1357), .B(acc[7]), .C(n2332), .D(n2473), .E(n1555), .Y(
        n1554) );
  NAND3X1 U1989 ( .A(n1564), .B(n1565), .C(n1566), .Y(n814) );
  AOI22X1 U1990 ( .A(n1023), .B(acc[0]), .C(n2264), .D(ramdatao[2]), .Y(n1564)
         );
  AOI222XL U1991 ( .A(acc[3]), .B(n2352), .C(n1349), .D(acc[4]), .E(
        adder_out[2]), .F(n2328), .Y(n1565) );
  AOI221XL U1992 ( .A(n1357), .B(acc[6]), .C(n2332), .D(n2475), .E(n1567), .Y(
        n1566) );
  NAND2X1 U1993 ( .A(n2028), .B(n2508), .Y(n2027) );
  NAND2X1 U1994 ( .A(dec_accop[13]), .B(n1362), .Y(n1356) );
  INVX1 U1995 ( .A(acc[7]), .Y(n2489) );
  INVX1 U1996 ( .A(phase[1]), .Y(n2182) );
  OAI222XL U1997 ( .A(n1556), .B(n2438), .C(n1557), .D(n2473), .E(n2351), .F(
        n2475), .Y(n1555) );
  AOI221XL U1998 ( .A(n2331), .B(n2473), .C(acc[3]), .D(n1360), .E(n1363), .Y(
        n1556) );
  AOI21X1 U1999 ( .B(n2331), .C(n2438), .A(n2333), .Y(n1557) );
  OAI222XL U2000 ( .A(n1568), .B(n2440), .C(n1569), .D(n2475), .E(n2351), .F(
        n2477), .Y(n1567) );
  AOI221XL U2001 ( .A(n2331), .B(n2475), .C(acc[2]), .D(n1360), .E(n1363), .Y(
        n1568) );
  AOI21X1 U2002 ( .B(n2331), .C(n2440), .A(n2333), .Y(n1569) );
  INVX1 U2003 ( .A(ramsfraddr[1]), .Y(n2442) );
  AOI21X1 U2004 ( .B(rn_reg[179]), .C(n66), .A(n1799), .Y(n1911) );
  AOI21X1 U2005 ( .B(rn_reg[51]), .C(n66), .A(n1817), .Y(n1919) );
  AOI21X1 U2006 ( .B(rn_reg[183]), .C(n66), .A(n1799), .Y(n1788) );
  INVX1 U2007 ( .A(n1469), .Y(n1660) );
  NAND43X1 U2008 ( .B(n1468), .C(n1467), .D(n1466), .A(n1465), .Y(n1469) );
  AOI221XL U2009 ( .A(n410), .B(n814), .C(n2246), .D(temp2_comb[2]), .E(n1464), 
        .Y(n1465) );
  AOI31X1 U2010 ( .A(n1779), .B(n1439), .C(n1438), .D(n1442), .Y(n1468) );
  INVX1 U2011 ( .A(ramsfraddr[2]), .Y(n2444) );
  AOI221XL U2012 ( .A(n1052), .B(n1053), .C(n2355), .D(n2354), .E(n1031), .Y(
        n1051) );
  NOR43XL U2013 ( .B(n1054), .C(n1055), .D(n1056), .A(n840), .Y(n1053) );
  AOI221XL U2014 ( .A(dec_cop[7]), .B(n123), .C(n123), .D(n1057), .E(n2337), 
        .Y(n1052) );
  OR4X1 U2015 ( .A(dec_accop[17]), .B(dec_cop[6]), .C(dec_accop[1]), .D(
        dec_accop[4]), .Y(n1057) );
  AOI32X1 U2016 ( .A(n1392), .B(n1393), .C(acc[0]), .D(acc[7]), .E(n1394), .Y(
        n1391) );
  OAI21X1 U2017 ( .B(temp2_comb[7]), .C(n1356), .A(n1395), .Y(n1394) );
  INVX1 U2018 ( .A(ramsfraddr[0]), .Y(n2443) );
  MUX2BXL U2019 ( .D0(n625), .D1(n624), .S(codefetch_s), .Y(n862) );
  NAND21X1 U2020 ( .B(n623), .A(n622), .Y(n625) );
  AND2X1 U2021 ( .A(n1587), .B(n1543), .Y(n624) );
  AO2222XL U2022 ( .A(n1578), .B(phase[3]), .C(n614), .D(phase[2]), .E(n754), 
        .F(n106), .G(n611), .H(n262), .Y(n622) );
  AOI21X1 U2023 ( .B(rn_reg[52]), .C(n66), .A(n1817), .Y(n1896) );
  AOI21X1 U2024 ( .B(rn_reg[180]), .C(n66), .A(n1799), .Y(n1888) );
  NOR3XL U2025 ( .A(n2017), .B(n2018), .C(n2019), .Y(n2016) );
  XNOR2XL U2026 ( .A(n2190), .B(ramsfraddr[0]), .Y(n2017) );
  XNOR2XL U2027 ( .A(n2444), .B(n2020), .Y(n2018) );
  XNOR2XL U2028 ( .A(n2442), .B(n2417), .Y(n2019) );
  INVX1 U2029 ( .A(temp2_comb[2]), .Y(n2440) );
  NAND4X1 U2030 ( .A(n1911), .B(n1912), .C(n1913), .D(n1914), .Y(n1910) );
  AOI22X1 U2031 ( .A(rn_reg[243]), .B(n161), .C(rn_reg[147]), .D(n144), .Y(
        n1912) );
  AOI22X1 U2032 ( .A(rn_reg[227]), .B(n120), .C(rn_reg[131]), .D(n100), .Y(
        n1914) );
  AOI22X1 U2033 ( .A(rn_reg[163]), .B(n73), .C(rn_reg[211]), .D(n87), .Y(n1913) );
  NAND4X1 U2034 ( .A(n1788), .B(n1789), .C(n1790), .D(n1791), .Y(n1786) );
  AOI22X1 U2035 ( .A(rn_reg[247]), .B(n161), .C(rn_reg[151]), .D(n144), .Y(
        n1789) );
  AOI22X1 U2036 ( .A(rn_reg[167]), .B(n73), .C(rn_reg[215]), .D(n87), .Y(n1790) );
  AOI22X1 U2037 ( .A(rn_reg[231]), .B(n120), .C(rn_reg[135]), .D(n100), .Y(
        n1791) );
  NOR32XL U2038 ( .B(n1362), .C(dec_accop[2]), .A(dec_accop[13]), .Y(n1357) );
  NOR43XL U2039 ( .B(n1674), .C(n2479), .D(n123), .A(n1675), .Y(n1360) );
  NOR2X1 U2040 ( .A(n2350), .B(n2335), .Y(n1674) );
  NAND21X1 U2041 ( .B(n1757), .A(phase[1]), .Y(n2380) );
  MUX2BXL U2042 ( .D0(n12), .D1(rs[0]), .S(n1015), .Y(n1038) );
  NAND43X1 U2043 ( .B(n772), .C(n2434), .D(n260), .A(interrupt), .Y(n785) );
  AND3X1 U2044 ( .A(n1362), .B(dec_accop[17]), .C(n1662), .Y(n1023) );
  NOR3XL U2045 ( .A(n1663), .B(dec_accop[18]), .C(n840), .Y(n1662) );
  MUX2X1 U2046 ( .D0(pc_o[0]), .D1(n1228), .S(n899), .Y(N12841) );
  NOR21XL U2047 ( .B(dec_accop[0]), .A(n2367), .Y(n1392) );
  NAND4X1 U2048 ( .A(n1846), .B(n1847), .C(n1848), .D(n1849), .Y(n1830) );
  NAND4X1 U2049 ( .A(n1838), .B(n1839), .C(n1840), .D(n1841), .Y(n1832) );
  NAND4X1 U2050 ( .A(n1842), .B(n1843), .C(n1844), .D(n1845), .Y(n1831) );
  XNOR2XL U2051 ( .A(n1365), .B(n107), .Y(n1457) );
  OAI221X1 U2052 ( .A(n1037), .B(n475), .C(n2356), .D(n1336), .E(n1337), .Y(
        n1333) );
  AOI33X1 U2053 ( .A(n2402), .B(n1336), .C(ramdatao[2]), .D(n476), .E(n2374), 
        .F(n2510), .Y(n1337) );
  OAI221X1 U2054 ( .A(n1038), .B(n475), .C(n2376), .D(n1336), .E(n1338), .Y(
        n1332) );
  INVX1 U2055 ( .A(rs[0]), .Y(n2376) );
  AOI33X1 U2056 ( .A(n2402), .B(n1336), .C(ramdatao[1]), .D(n476), .E(n2374), 
        .F(dps[1]), .Y(n1338) );
  GEN2XL U2057 ( .D(acc[7]), .E(n1480), .C(c), .B(n1481), .A(n1366), .Y(n1459)
         );
  OAI31XL U2058 ( .A(n2403), .B(n1482), .C(n2473), .D(n1483), .Y(n1480) );
  NOR2X1 U2059 ( .A(acc[6]), .B(acc[5]), .Y(n1483) );
  INVX1 U2060 ( .A(n445), .Y(n883) );
  NAND21X1 U2061 ( .B(n1983), .A(n442), .Y(n445) );
  OAI222XL U2062 ( .A(n1780), .B(n2443), .C(n1078), .D(n2340), .E(n2320), .F(
        n1781), .Y(n1983) );
  AOI22X1 U2063 ( .A(n1982), .B(instr[0]), .C(n437), .D(n441), .Y(n442) );
  NOR21XL U2064 ( .B(dec_accop[4]), .A(n2367), .Y(n1677) );
  OAI22X1 U2065 ( .A(n2401), .B(n1217), .C(n2203), .D(n1139), .Y(n2139) );
  AND4X1 U2066 ( .A(n1218), .B(n1219), .C(n1220), .D(n1221), .Y(n1217) );
  AOI22X1 U2067 ( .A(n1151), .B(dpl_reg[48]), .C(n1152), .D(dpl_reg[56]), .Y(
        n1218) );
  AOI22X1 U2068 ( .A(n1149), .B(dpl_reg[32]), .C(n1150), .D(dpl_reg[40]), .Y(
        n1219) );
  OAI21X1 U2069 ( .B(n1684), .C(n2367), .A(n1667), .Y(n1663) );
  NOR3XL U2070 ( .A(n2483), .B(dec_accop[7]), .C(dec_accop[15]), .Y(n1684) );
  MUX2XL U2071 ( .D0(ramdatao[1]), .D1(n1657), .S(waitstaten), .Y(
        ramdatao_comb[1]) );
  AOI22AXL U2072 ( .A(sp[0]), .B(n1829), .D(n1829), .C(ramdatao[0]), .Y(n1975)
         );
  NOR2X1 U2073 ( .A(n2190), .B(n2508), .Y(n774) );
  AOI21X1 U2074 ( .B(accactv), .C(dec_accop[18]), .A(n1663), .Y(n1668) );
  INVX1 U2075 ( .A(n2509), .Y(n2190) );
  INVX1 U2076 ( .A(n299), .Y(n2153) );
  OAI211X1 U2077 ( .C(ckcon[2]), .D(n2370), .A(n2057), .B(n1619), .Y(n299) );
  OAI22X1 U2078 ( .A(n2058), .B(n2059), .C(test_so), .D(n2372), .Y(n2057) );
  NOR2X1 U2079 ( .A(ckcon[1]), .B(n2369), .Y(n2058) );
  INVX1 U2080 ( .A(accactv), .Y(n2367) );
  NOR2X1 U2081 ( .A(n2450), .B(n2505), .Y(n1736) );
  MUX2X1 U2082 ( .D0(n1561), .D1(pdmode), .S(n1560), .Y(n2036) );
  AOI211X1 U2083 ( .C(n1551), .D(n588), .A(n291), .B(n1570), .Y(n1560) );
  AND2X1 U2084 ( .A(n1547), .B(n287), .Y(n1561) );
  OAI22X1 U2085 ( .A(idle_r), .B(stop_r), .C(n1563), .D(n1591), .Y(n1551) );
  NAND4X1 U2086 ( .A(n785), .B(n1533), .C(n945), .D(n1991), .Y(n1822) );
  AOI21X1 U2087 ( .B(n1726), .C(phase[1]), .A(n1689), .Y(n1991) );
  NOR3XL U2088 ( .A(ramsfraddr[0]), .B(ramsfraddr[2]), .C(n2442), .Y(n855) );
  ENOX1 U2089 ( .A(n1829), .B(n2199), .C(sp[1]), .D(n1829), .Y(N12770) );
  INVX1 U2090 ( .A(n867), .Y(n2154) );
  GEN2XL U2091 ( .D(n2060), .E(n2371), .C(test_so), .B(n2061), .A(n2062), .Y(
        n867) );
  NAND21X1 U2092 ( .B(n2060), .A(ckcon[6]), .Y(n2061) );
  AOI222XL U2093 ( .A(ckcon[6]), .B(n2370), .C(ckcon[4]), .D(n2368), .E(
        ckcon[5]), .F(n2369), .Y(n2062) );
  AO22X1 U2094 ( .A(n249), .B(n1733), .C(pc_ini[15]), .D(n291), .Y(N495) );
  AND4X1 U2095 ( .A(n1870), .B(n1871), .C(n1868), .D(n1869), .Y(n345) );
  AOI22X1 U2096 ( .A(rn_reg[37]), .B(n74), .C(rn_reg[85]), .D(n88), .Y(n1870)
         );
  AOI22X1 U2097 ( .A(rn_reg[101]), .B(n121), .C(rn_reg[5]), .D(n101), .Y(n1871) );
  AOI22X1 U2098 ( .A(rn_reg[117]), .B(n162), .C(rn_reg[21]), .D(n145), .Y(
        n1869) );
  AND4X1 U2099 ( .A(n2006), .B(n2007), .C(n2004), .D(n2005), .Y(n333) );
  AOI22X1 U2100 ( .A(rn_reg[32]), .B(n74), .C(rn_reg[80]), .D(n88), .Y(n2006)
         );
  AOI22X1 U2101 ( .A(rn_reg[96]), .B(n121), .C(rn_reg[0]), .D(n101), .Y(n2007)
         );
  AOI22X1 U2102 ( .A(rn_reg[112]), .B(n162), .C(rn_reg[16]), .D(n145), .Y(
        n2005) );
  AND4X1 U2103 ( .A(n1968), .B(n1969), .C(n1966), .D(n1967), .Y(n469) );
  AOI22X1 U2104 ( .A(rn_reg[97]), .B(n121), .C(rn_reg[1]), .D(n101), .Y(n1969)
         );
  AOI22X1 U2105 ( .A(rn_reg[113]), .B(n162), .C(rn_reg[17]), .D(n145), .Y(
        n1967) );
  AOI22X1 U2106 ( .A(rn_reg[33]), .B(n74), .C(rn_reg[81]), .D(n88), .Y(n1968)
         );
  AND4X1 U2107 ( .A(n1945), .B(n1946), .C(n1943), .D(n1944), .Y(n340) );
  AOI22X1 U2108 ( .A(rn_reg[34]), .B(n74), .C(rn_reg[82]), .D(n88), .Y(n1945)
         );
  AOI22X1 U2109 ( .A(rn_reg[98]), .B(n121), .C(rn_reg[2]), .D(n101), .Y(n1946)
         );
  AOI22X1 U2110 ( .A(rn_reg[114]), .B(n162), .C(rn_reg[18]), .D(n145), .Y(
        n1944) );
  NOR2X1 U2111 ( .A(n2405), .B(ramsfraddr[3]), .Y(n853) );
  AOI21X1 U2112 ( .B(n2481), .C(temp2_comb[6]), .A(n1459), .Y(n1398) );
  OAI22X1 U2113 ( .A(n2199), .B(n1139), .C(n2401), .D(n1210), .Y(n2138) );
  AND4X1 U2114 ( .A(n1211), .B(n1212), .C(n1213), .D(n1214), .Y(n1210) );
  AOI22X1 U2115 ( .A(n1151), .B(dpl_reg[49]), .C(n1152), .D(dpl_reg[57]), .Y(
        n1211) );
  AOI22X1 U2116 ( .A(n1149), .B(dpl_reg[33]), .C(n1150), .D(dpl_reg[41]), .Y(
        n1212) );
  OAI22X1 U2117 ( .A(n2192), .B(n1139), .C(n2401), .D(n1203), .Y(n2137) );
  AND4X1 U2118 ( .A(n1204), .B(n1205), .C(n1206), .D(n1207), .Y(n1203) );
  AOI22X1 U2119 ( .A(n1151), .B(dpl_reg[50]), .C(n1152), .D(dpl_reg[58]), .Y(
        n1204) );
  AOI22X1 U2120 ( .A(n1149), .B(dpl_reg[34]), .C(n1150), .D(dpl_reg[42]), .Y(
        n1205) );
  OAI31XL U2121 ( .A(dec_accop[13]), .B(dec_accop[2]), .C(dec_accop[14]), .D(
        accactv), .Y(n1667) );
  AOI222XL U2122 ( .A(rn_reg[139]), .B(n118), .C(rn_reg[203]), .D(n159), .E(
        rn_reg[235]), .F(n142), .Y(n1918) );
  AOI222XL U2123 ( .A(rn_reg[11]), .B(n118), .C(rn_reg[75]), .D(n159), .E(
        rn_reg[107]), .F(n142), .Y(n1926) );
  NAND2X1 U2124 ( .A(dec_accop[3]), .B(accactv), .Y(n1604) );
  AOI22X1 U2125 ( .A(rn_reg[99]), .B(n120), .C(rn_reg[3]), .D(n100), .Y(n1922)
         );
  AOI22X1 U2126 ( .A(rn_reg[35]), .B(n73), .C(rn_reg[83]), .D(n87), .Y(n1921)
         );
  AOI22X1 U2127 ( .A(rn_reg[171]), .B(n96), .C(rn_reg[219]), .D(n71), .Y(n1917) );
  AOI22X1 U2128 ( .A(rn_reg[43]), .B(n96), .C(rn_reg[91]), .D(n71), .Y(n1925)
         );
  AOI22X1 U2129 ( .A(rn_reg[115]), .B(n161), .C(rn_reg[19]), .D(n144), .Y(
        n1920) );
  AOI22X1 U2130 ( .A(rn_reg[251]), .B(n98), .C(rn_reg[155]), .D(n157), .Y(
        n1916) );
  AOI22X1 U2131 ( .A(rn_reg[123]), .B(n98), .C(rn_reg[27]), .D(n157), .Y(n1924) );
  INVX1 U2132 ( .A(n315), .Y(n397) );
  NAND21X1 U2133 ( .B(n1757), .A(phase[0]), .Y(n315) );
  AOI21X1 U2134 ( .B(n2481), .C(temp2_comb[5]), .A(n1459), .Y(n1453) );
  AOI22X1 U2135 ( .A(rn_reg[187]), .B(n116), .C(rn_reg[195]), .D(n140), .Y(
        n1915) );
  AOI22X1 U2136 ( .A(rn_reg[59]), .B(n116), .C(rn_reg[67]), .D(n140), .Y(n1923) );
  INVX1 U2137 ( .A(ramsfraddr[5]), .Y(n2189) );
  AOI21X1 U2138 ( .B(rn_reg[55]), .C(n66), .A(n1817), .Y(n1813) );
  AOI21X1 U2139 ( .B(rn_reg[182]), .C(n67), .A(n1799), .Y(n1834) );
  NOR2X1 U2140 ( .A(n126), .B(instr[2]), .Y(n1756) );
  AOI222XL U2141 ( .A(rn_reg[12]), .B(n118), .C(rn_reg[76]), .D(n159), .E(
        rn_reg[108]), .F(n142), .Y(n1903) );
  AOI222XL U2142 ( .A(rn_reg[140]), .B(n118), .C(rn_reg[204]), .D(n159), .E(
        rn_reg[236]), .F(n142), .Y(n1895) );
  AOI222XL U2143 ( .A(rn_reg[9]), .B(n119), .C(rn_reg[73]), .D(n160), .E(
        rn_reg[105]), .F(n143), .Y(n1973) );
  AOI222XL U2144 ( .A(rn_reg[137]), .B(n119), .C(rn_reg[201]), .D(n160), .E(
        rn_reg[233]), .F(n143), .Y(n1965) );
  INVX1 U2145 ( .A(acc[3]), .Y(n2473) );
  NOR2X1 U2146 ( .A(n2417), .B(n2509), .Y(n2026) );
  NOR2X1 U2147 ( .A(n2027), .B(n2509), .Y(n2025) );
  AOI221XL U2148 ( .A(n134), .B(n2477), .C(acc[1]), .D(n1360), .E(n1363), .Y(
        n1593) );
  NAND3X1 U2149 ( .A(n2442), .B(n2444), .C(ramsfraddr[0]), .Y(n844) );
  AOI221XL U2150 ( .A(n134), .B(n2489), .C(n1360), .D(acc[7]), .E(n1363), .Y(
        n1390) );
  INVX1 U2151 ( .A(waitcnt_1_), .Y(n2369) );
  INVX1 U2152 ( .A(acc[4]), .Y(n2403) );
  AOI22X1 U2153 ( .A(rn_reg[124]), .B(n98), .C(rn_reg[28]), .D(n157), .Y(n1901) );
  AOI22X1 U2154 ( .A(n1145), .B(dpl_reg[0]), .C(n1146), .D(dpl_reg[8]), .Y(
        n1221) );
  AOI22X1 U2155 ( .A(n1145), .B(dpl_reg[1]), .C(n1146), .D(dpl_reg[9]), .Y(
        n1214) );
  AOI22X1 U2156 ( .A(n1145), .B(dpl_reg[2]), .C(n1146), .D(dpl_reg[10]), .Y(
        n1207) );
  AOI22X1 U2157 ( .A(rn_reg[60]), .B(n116), .C(rn_reg[68]), .D(n140), .Y(n1900) );
  AOI22X1 U2158 ( .A(rn_reg[188]), .B(n116), .C(rn_reg[196]), .D(n140), .Y(
        n1892) );
  AOI22X1 U2159 ( .A(n1147), .B(dpl_reg[16]), .C(n1148), .D(dpl_reg[24]), .Y(
        n1220) );
  AOI22X1 U2160 ( .A(n1147), .B(dpl_reg[17]), .C(n1148), .D(dpl_reg[25]), .Y(
        n1213) );
  AOI22X1 U2161 ( .A(rn_reg[44]), .B(n96), .C(rn_reg[92]), .D(n71), .Y(n1902)
         );
  AOI22X1 U2162 ( .A(rn_reg[172]), .B(n96), .C(rn_reg[220]), .D(n71), .Y(n1894) );
  AOI21X1 U2163 ( .B(rn_reg[53]), .C(n67), .A(n1817), .Y(n1868) );
  AOI21X1 U2164 ( .B(rn_reg[181]), .C(n67), .A(n1799), .Y(n1860) );
  AOI21X1 U2165 ( .B(rn_reg[48]), .C(n67), .A(n1817), .Y(n2004) );
  AOI21X1 U2166 ( .B(rn_reg[176]), .C(n67), .A(n1799), .Y(n1996) );
  AOI21X1 U2167 ( .B(rn_reg[49]), .C(n67), .A(n1817), .Y(n1966) );
  AOI21X1 U2168 ( .B(rn_reg[177]), .C(n67), .A(n1799), .Y(n1958) );
  AOI21X1 U2169 ( .B(rn_reg[50]), .C(n67), .A(n1817), .Y(n1943) );
  AOI21X1 U2170 ( .B(rn_reg[178]), .C(n67), .A(n1799), .Y(n1935) );
  AOI22X1 U2171 ( .A(ckcon[0]), .B(n2368), .C(ckcon[1]), .D(n2369), .Y(n2059)
         );
  NAND2X1 U2172 ( .A(n2501), .B(n2402), .Y(n1336) );
  INVX1 U2173 ( .A(ramsfraddr[4]), .Y(n2405) );
  INVX1 U2174 ( .A(ramsfraddr[6]), .Y(n2188) );
  NAND2X1 U2175 ( .A(dps[3]), .B(n476), .Y(n475) );
  INVX1 U2176 ( .A(waitcnt_0_), .Y(n2368) );
  NAND4X1 U2177 ( .A(n1834), .B(n1835), .C(n1836), .D(n1837), .Y(n1833) );
  AOI22X1 U2178 ( .A(rn_reg[246]), .B(n162), .C(rn_reg[150]), .D(n145), .Y(
        n1835) );
  AOI22X1 U2179 ( .A(rn_reg[230]), .B(n121), .C(rn_reg[134]), .D(n101), .Y(
        n1837) );
  AOI22X1 U2180 ( .A(rn_reg[166]), .B(n74), .C(rn_reg[214]), .D(n88), .Y(n1836) );
  NOR2X1 U2181 ( .A(n2369), .B(ckcon[5]), .Y(n2060) );
  INVX1 U2182 ( .A(ckcon[6]), .Y(n2371) );
  INVX1 U2183 ( .A(test_so), .Y(n2370) );
  INVX1 U2184 ( .A(ckcon[2]), .Y(n2372) );
  NAND21X1 U2185 ( .B(instr[6]), .A(n2504), .Y(n2449) );
  NOR2X1 U2186 ( .A(instr[1]), .B(n2509), .Y(n1324) );
  NAND21X1 U2187 ( .B(n168), .A(interrupt), .Y(n1699) );
  AOI22X1 U2188 ( .A(n476), .B(dps[0]), .C(n2402), .D(ramdatao[0]), .Y(n1089)
         );
  OR2X1 U2189 ( .A(memwr), .B(memrd), .Y(n1619) );
  AO222X1 U2190 ( .A(n30), .B(n235), .C(n28), .D(n1728), .E(pc_ini[10]), .F(
        n291), .Y(N490) );
  BUFX3 U2191 ( .A(memaddr[10]), .Y(n235) );
  AO222X1 U2192 ( .A(n31), .B(pc_o[1]), .C(n29), .D(n1714), .E(pc_ini[1]), .F(
        n293), .Y(N481) );
  BUFX3 U2193 ( .A(memaddr[1]), .Y(pc_o[1]) );
  AO222X1 U2194 ( .A(n30), .B(pc_o[9]), .C(n28), .D(n1724), .E(pc_ini[9]), .F(
        n293), .Y(N489) );
  AO222X1 U2195 ( .A(n31), .B(pc_o[8]), .C(n29), .D(n1721), .E(pc_ini[8]), .F(
        n293), .Y(N488) );
  AO222X1 U2196 ( .A(n30), .B(pc_o[7]), .C(n28), .D(n1720), .E(pc_ini[7]), .F(
        n293), .Y(N487) );
  AO222X1 U2197 ( .A(n31), .B(pc_o[6]), .C(n29), .D(n1719), .E(pc_ini[6]), .F(
        n291), .Y(N486) );
  AO222X1 U2198 ( .A(n30), .B(pc_o[5]), .C(n28), .D(n1718), .E(pc_ini[5]), .F(
        n291), .Y(N485) );
  AO222X1 U2199 ( .A(n31), .B(memaddr[4]), .C(n29), .D(n1717), .E(pc_ini[4]), 
        .F(n291), .Y(N484) );
  AO222X1 U2200 ( .A(n30), .B(pc_o[3]), .C(n28), .D(n1716), .E(pc_ini[3]), .F(
        n293), .Y(N483) );
  AO222X1 U2201 ( .A(n31), .B(memaddr[2]), .C(n29), .D(n1715), .E(pc_ini[2]), 
        .F(n293), .Y(N482) );
  AO222X1 U2202 ( .A(n30), .B(pc_o[0]), .C(n28), .D(n1713), .E(pc_ini[0]), .F(
        n293), .Y(N480) );
  NAND21X1 U2203 ( .B(n2499), .A(n623), .Y(n1621) );
  AOI22AXL U2204 ( .A(sp[6]), .B(n156), .D(n156), .C(ramdatao[6]), .Y(n1828)
         );
  INVX1 U2205 ( .A(n2507), .Y(n2261) );
  INVX1 U2206 ( .A(n1571), .Y(n1576) );
  GEN2XL U2207 ( .D(n1573), .E(n1590), .C(n1572), .B(newinstrlock), .A(n295), 
        .Y(n1574) );
  NOR2X1 U2208 ( .A(n2506), .B(n2505), .Y(n1723) );
  ENOX1 U2209 ( .A(n156), .B(n2216), .C(sp[4]), .D(n156), .Y(N12773) );
  ENOX1 U2210 ( .A(n1829), .B(n12), .C(sp[3]), .D(n1829), .Y(N12772) );
  ENOX1 U2211 ( .A(n1829), .B(n2192), .C(sp[2]), .D(n1829), .Y(N12771) );
  AND2X1 U2212 ( .A(dec_accop[5]), .B(accactv), .Y(n1675) );
  NOR2X1 U2213 ( .A(n2448), .B(n2505), .Y(n2106) );
  NAND3X1 U2214 ( .A(dec_accop[1]), .B(n123), .C(n1044), .Y(n1034) );
  AO21X1 U2215 ( .B(waitstaten), .C(n1406), .A(n294), .Y(N520) );
  MUX2X1 U2216 ( .D0(p2sel), .D1(n1664), .S(n1405), .Y(n1406) );
  AO22X1 U2217 ( .A(n243), .B(n1732), .C(pc_ini[14]), .D(n294), .Y(N494) );
  AO22X1 U2218 ( .A(n249), .B(n1731), .C(pc_ini[13]), .D(n291), .Y(N493) );
  AO22X1 U2219 ( .A(n243), .B(n1730), .C(pc_ini[12]), .D(n293), .Y(N492) );
  AO22X1 U2220 ( .A(n249), .B(n1729), .C(pc_ini[11]), .D(n295), .Y(N491) );
  INVX1 U2221 ( .A(acc[6]), .Y(n2415) );
  NOR2X1 U2222 ( .A(n32), .B(n2506), .Y(n970) );
  OAI22X1 U2223 ( .A(n12), .B(n1139), .C(n2401), .D(n1193), .Y(n2127) );
  AND4X1 U2224 ( .A(n1194), .B(n1195), .C(n1196), .D(n1197), .Y(n1193) );
  AOI22X1 U2225 ( .A(n1151), .B(dpl_reg[51]), .C(n1152), .D(dpl_reg[59]), .Y(
        n1194) );
  AOI22X1 U2226 ( .A(n1149), .B(dpl_reg[35]), .C(n1150), .D(dpl_reg[43]), .Y(
        n1195) );
  NAND3X1 U2227 ( .A(n1990), .B(n444), .C(n2341), .Y(n1985) );
  OAI21X1 U2228 ( .B(n1987), .C(n2255), .A(phase[0]), .Y(n1990) );
  AOI222XL U2229 ( .A(rn_reg[143]), .B(n118), .C(rn_reg[207]), .D(n159), .E(
        rn_reg[239]), .F(n142), .Y(n1803) );
  AOI222XL U2230 ( .A(rn_reg[15]), .B(n118), .C(rn_reg[79]), .D(n159), .E(
        rn_reg[111]), .F(n142), .Y(n1821) );
  AOI222XL U2231 ( .A(rn_reg[142]), .B(n119), .C(rn_reg[206]), .D(n160), .E(
        rn_reg[238]), .F(n143), .Y(n1841) );
  AOI222XL U2232 ( .A(rn_reg[14]), .B(n119), .C(rn_reg[78]), .D(n160), .E(
        rn_reg[110]), .F(n143), .Y(n1849) );
  INVX1 U2233 ( .A(ramdatao[4]), .Y(n2216) );
  AOI22X1 U2234 ( .A(rn_reg[103]), .B(n120), .C(rn_reg[7]), .D(n100), .Y(n1816) );
  AOI22X1 U2235 ( .A(rn_reg[39]), .B(n73), .C(rn_reg[87]), .D(n87), .Y(n1815)
         );
  AOI22X1 U2236 ( .A(rn_reg[175]), .B(n96), .C(rn_reg[223]), .D(n71), .Y(n1802) );
  AOI22X1 U2237 ( .A(rn_reg[47]), .B(n96), .C(rn_reg[95]), .D(n71), .Y(n1820)
         );
  AOI22X1 U2238 ( .A(rn_reg[119]), .B(n161), .C(rn_reg[23]), .D(n144), .Y(
        n1814) );
  AOI22X1 U2239 ( .A(rn_reg[255]), .B(n98), .C(rn_reg[159]), .D(n157), .Y(
        n1801) );
  AOI22X1 U2240 ( .A(rn_reg[127]), .B(n98), .C(rn_reg[31]), .D(n157), .Y(n1819) );
  AOI22X1 U2241 ( .A(rn_reg[191]), .B(n116), .C(rn_reg[199]), .D(n140), .Y(
        n1800) );
  AOI22X1 U2242 ( .A(rn_reg[63]), .B(n116), .C(rn_reg[71]), .D(n140), .Y(n1818) );
  AOI21X1 U2243 ( .B(rn_reg[54]), .C(n67), .A(n1817), .Y(n1842) );
  AOI222XL U2244 ( .A(rn_reg[13]), .B(n119), .C(rn_reg[77]), .D(n160), .E(
        rn_reg[109]), .F(n143), .Y(n1875) );
  AOI222XL U2245 ( .A(rn_reg[141]), .B(n119), .C(rn_reg[205]), .D(n160), .E(
        rn_reg[237]), .F(n143), .Y(n1867) );
  AOI222XL U2246 ( .A(rn_reg[8]), .B(n119), .C(rn_reg[72]), .D(n160), .E(
        rn_reg[104]), .F(n143), .Y(n2024) );
  AOI222XL U2247 ( .A(rn_reg[136]), .B(n119), .C(rn_reg[200]), .D(n160), .E(
        rn_reg[232]), .F(n143), .Y(n2003) );
  AOI222XL U2248 ( .A(rn_reg[10]), .B(n119), .C(rn_reg[74]), .D(n160), .E(
        rn_reg[106]), .F(n143), .Y(n1950) );
  AOI222XL U2249 ( .A(rn_reg[138]), .B(n119), .C(rn_reg[202]), .D(n160), .E(
        rn_reg[234]), .F(n143), .Y(n1942) );
  INVX1 U2250 ( .A(acc[5]), .Y(n2406) );
  OAI22AX1 U2251 ( .D(idle), .C(n1542), .A(n1571), .B(n1500), .Y(n1879) );
  AOI22X1 U2252 ( .A(rn_reg[245]), .B(n162), .C(rn_reg[149]), .D(n145), .Y(
        n1861) );
  AOI22X1 U2253 ( .A(rn_reg[125]), .B(n99), .C(rn_reg[29]), .D(n158), .Y(n1873) );
  AOI22X1 U2254 ( .A(rn_reg[253]), .B(n99), .C(rn_reg[157]), .D(n158), .Y(
        n1865) );
  AOI22X1 U2255 ( .A(rn_reg[244]), .B(n161), .C(rn_reg[148]), .D(n144), .Y(
        n1889) );
  AOI22X1 U2256 ( .A(rn_reg[252]), .B(n98), .C(rn_reg[156]), .D(n157), .Y(
        n1893) );
  AOI22X1 U2257 ( .A(rn_reg[240]), .B(n162), .C(rn_reg[144]), .D(n145), .Y(
        n1997) );
  AOI22X1 U2258 ( .A(rn_reg[120]), .B(n99), .C(rn_reg[24]), .D(n158), .Y(n2022) );
  AOI22X1 U2259 ( .A(rn_reg[248]), .B(n99), .C(rn_reg[152]), .D(n158), .Y(
        n2001) );
  AOI22X1 U2260 ( .A(rn_reg[241]), .B(n162), .C(rn_reg[145]), .D(n145), .Y(
        n1959) );
  AOI22X1 U2261 ( .A(rn_reg[121]), .B(n99), .C(rn_reg[25]), .D(n158), .Y(n1971) );
  AOI22X1 U2262 ( .A(rn_reg[249]), .B(n99), .C(rn_reg[153]), .D(n158), .Y(
        n1963) );
  AOI22X1 U2265 ( .A(rn_reg[122]), .B(n99), .C(rn_reg[26]), .D(n158), .Y(n1948) );
  AOI22X1 U2266 ( .A(n1145), .B(dpl_reg[3]), .C(n1146), .D(dpl_reg[11]), .Y(
        n1197) );
  AOI22X1 U2267 ( .A(rn_reg[61]), .B(n117), .C(rn_reg[69]), .D(n141), .Y(n1872) );
  AOI22X1 U2268 ( .A(rn_reg[189]), .B(n117), .C(rn_reg[197]), .D(n141), .Y(
        n1864) );
  AOI22X1 U2269 ( .A(rn_reg[56]), .B(n117), .C(rn_reg[64]), .D(n141), .Y(n2021) );
  AOI22X1 U2270 ( .A(rn_reg[184]), .B(n117), .C(rn_reg[192]), .D(n141), .Y(
        n2000) );
  AOI22X1 U2271 ( .A(rn_reg[57]), .B(n117), .C(rn_reg[65]), .D(n141), .Y(n1970) );
  AOI22X1 U2272 ( .A(rn_reg[185]), .B(n117), .C(rn_reg[193]), .D(n141), .Y(
        n1962) );
  AOI22X1 U2273 ( .A(rn_reg[58]), .B(n117), .C(rn_reg[66]), .D(n141), .Y(n1947) );
  AOI22X1 U2274 ( .A(n1147), .B(dpl_reg[18]), .C(n1148), .D(dpl_reg[26]), .Y(
        n1206) );
  AOI22X1 U2275 ( .A(n1147), .B(dpl_reg[19]), .C(n1148), .D(dpl_reg[27]), .Y(
        n1196) );
  AOI22X1 U2276 ( .A(rn_reg[165]), .B(n74), .C(rn_reg[213]), .D(n88), .Y(n1862) );
  AOI22X1 U2277 ( .A(rn_reg[45]), .B(n97), .C(rn_reg[93]), .D(n72), .Y(n1874)
         );
  AOI22X1 U2278 ( .A(rn_reg[173]), .B(n97), .C(rn_reg[221]), .D(n72), .Y(n1866) );
  AOI22X1 U2279 ( .A(rn_reg[164]), .B(n73), .C(rn_reg[212]), .D(n87), .Y(n1890) );
  AOI22X1 U2280 ( .A(rn_reg[160]), .B(n74), .C(rn_reg[208]), .D(n88), .Y(n1998) );
  AOI22X1 U2281 ( .A(rn_reg[40]), .B(n97), .C(rn_reg[88]), .D(n72), .Y(n2023)
         );
  AOI22X1 U2282 ( .A(rn_reg[168]), .B(n97), .C(rn_reg[216]), .D(n72), .Y(n2002) );
  AOI22X1 U2283 ( .A(rn_reg[161]), .B(n74), .C(rn_reg[209]), .D(n88), .Y(n1960) );
  AOI22X1 U2284 ( .A(rn_reg[41]), .B(n97), .C(rn_reg[89]), .D(n72), .Y(n1972)
         );
  AOI22X1 U2285 ( .A(rn_reg[169]), .B(n97), .C(rn_reg[217]), .D(n72), .Y(n1964) );
  AOI22X1 U2286 ( .A(rn_reg[42]), .B(n97), .C(rn_reg[90]), .D(n72), .Y(n1949)
         );
  AOI22X1 U2287 ( .A(rn_reg[229]), .B(n121), .C(rn_reg[133]), .D(n101), .Y(
        n1863) );
  AOI22X1 U2288 ( .A(rn_reg[228]), .B(n120), .C(rn_reg[132]), .D(n100), .Y(
        n1891) );
  AOI22X1 U2289 ( .A(rn_reg[224]), .B(n121), .C(rn_reg[128]), .D(n101), .Y(
        n1999) );
  AOI22X1 U2290 ( .A(rn_reg[225]), .B(n121), .C(rn_reg[129]), .D(n101), .Y(
        n1961) );
  NAND2X1 U2291 ( .A(dec_accop[11]), .B(accactv), .Y(n1673) );
  INVX1 U2292 ( .A(mempsrd), .Y(n623) );
  INVX1 U2293 ( .A(dec_accop[12]), .Y(n2335) );
  INVX1 U2294 ( .A(rs[1]), .Y(n2356) );
  MUX2AXL U2295 ( .D0(pmw), .D1(n2216), .S(n479), .Y(n2205) );
  NOR6XL U2296 ( .A(phase[5]), .B(phase[3]), .C(phase[1]), .D(phase[0]), .E(
        phase[4]), .F(phase[2]), .Y(n309) );
  AO222X1 U2297 ( .A(n2234), .B(temp[0]), .C(dptr_inc[8]), .D(n1138), .E(n2140), .F(n1235), .Y(n993) );
  NOR2X1 U2298 ( .A(n2478), .B(n2488), .Y(N14337) );
  OAI22X1 U2299 ( .A(n871), .B(n2095), .C(n2096), .D(n2399), .Y(n602) );
  AOI22X1 U2300 ( .A(ckcon[7]), .B(n488), .C(ckcon[3]), .D(n2205), .Y(n2095)
         );
  AOI22X1 U2301 ( .A(n488), .B(ramdatao[7]), .C(n2501), .D(n2205), .Y(n2096)
         );
  NAND21X1 U2302 ( .B(n2505), .A(n1006), .Y(n418) );
  GEN3XL U2303 ( .F(dec_cop[4]), .G(c), .E(n2307), .D(n2288), .C(n1058), .B(
        n1056), .A(n1059), .Y(n1050) );
  NOR4XL U2304 ( .A(n1064), .B(n2367), .C(dec_cop[5]), .D(n1065), .Y(n1058) );
  AOI21BBXL U2305 ( .B(n1060), .C(dec_cop[0]), .A(n2367), .Y(n1059) );
  OAI211X1 U2306 ( .C(c), .D(n1066), .A(n1055), .B(n1054), .Y(n1064) );
  OAI22X1 U2307 ( .A(n1976), .B(n170), .C(n261), .D(n446), .Y(n2362) );
  NOR4XL U2308 ( .A(n1977), .B(n1725), .C(n1765), .D(n1978), .Y(n1976) );
  NAND2X1 U2309 ( .A(n1979), .B(n1750), .Y(n1977) );
  AOI32X1 U2310 ( .A(n2508), .B(n2385), .C(n2269), .D(n1762), .E(n2449), .Y(
        n1979) );
  OAI21X1 U2311 ( .B(n169), .C(n2029), .A(n1744), .Y(n1982) );
  OAI31XL U2312 ( .A(n1634), .B(n1736), .C(n2033), .D(n2507), .Y(n2029) );
  NOR2X1 U2313 ( .A(n1773), .B(instr[6]), .Y(n1006) );
  OAI22X1 U2314 ( .A(n2031), .B(n2223), .C(n2032), .D(N345), .Y(n1063) );
  OAI221X1 U2315 ( .A(n2504), .B(n2078), .C(n2392), .D(n2427), .E(n2081), .Y(
        n750) );
  GEN2XL U2316 ( .D(n2506), .E(n602), .C(n2186), .B(n2397), .A(instr[2]), .Y(
        n2081) );
  XNOR2XL U2317 ( .A(n1365), .B(acc[7]), .Y(n1397) );
  NOR2X1 U2318 ( .A(n2448), .B(n2504), .Y(n973) );
  NAND21X1 U2319 ( .B(n308), .A(n307), .Y(n613) );
  AOI222XL U2320 ( .A(n2068), .B(phase[0]), .C(n306), .D(phase[1]), .E(n1579), 
        .F(phase[4]), .Y(n307) );
  AO21X1 U2321 ( .B(n2069), .C(phase[2]), .A(n2070), .Y(n308) );
  OAI211X1 U2322 ( .C(n2084), .D(n61), .A(n2085), .B(n2086), .Y(n2068) );
  NAND2X1 U2323 ( .A(n39), .B(n2504), .Y(n1773) );
  NOR2X1 U2324 ( .A(n1097), .B(n2510), .Y(n234) );
  NOR2X1 U2325 ( .A(n1097), .B(n2510), .Y(n508) );
  OAI22X1 U2326 ( .A(n2216), .B(n1139), .C(n2401), .D(n1181), .Y(n2136) );
  AND4X1 U2327 ( .A(n1182), .B(n1183), .C(n1184), .D(n1185), .Y(n1181) );
  AOI22X1 U2328 ( .A(n1151), .B(dpl_reg[52]), .C(n1152), .D(dpl_reg[60]), .Y(
        n1182) );
  AOI22X1 U2329 ( .A(n1149), .B(dpl_reg[36]), .C(n1150), .D(dpl_reg[44]), .Y(
        n1183) );
  OAI22X1 U2330 ( .A(n2212), .B(n1139), .C(n2401), .D(n1171), .Y(n2135) );
  AND4X1 U2331 ( .A(n1172), .B(n1173), .C(n1174), .D(n1175), .Y(n1171) );
  AOI22X1 U2332 ( .A(n1151), .B(dpl_reg[53]), .C(n1152), .D(dpl_reg[61]), .Y(
        n1172) );
  AOI22X1 U2333 ( .A(n1149), .B(dpl_reg[37]), .C(n1150), .D(dpl_reg[45]), .Y(
        n1173) );
  INVX1 U2334 ( .A(b[0]), .Y(n2490) );
  NAND2X1 U2335 ( .A(dps[1]), .B(n2365), .Y(n1097) );
  INVX1 U2336 ( .A(b[1]), .Y(n2488) );
  INVX1 U2337 ( .A(ramdatao[1]), .Y(n2199) );
  INVX1 U2338 ( .A(ramdatao[2]), .Y(n2192) );
  AOI22X1 U2339 ( .A(rn_reg[102]), .B(n121), .C(rn_reg[6]), .D(n101), .Y(n1845) );
  AOI22X1 U2340 ( .A(n21), .B(dph_reg[4]), .C(n508), .D(dph_reg[20]), .Y(n558)
         );
  AOI22X1 U2341 ( .A(n22), .B(dph_reg[6]), .C(n234), .D(dph_reg[22]), .Y(n550)
         );
  AOI22X1 U2342 ( .A(n233), .B(dpl_reg[7]), .C(n508), .D(dpl_reg[23]), .Y(n506) );
  AOI22X1 U2343 ( .A(rn_reg[38]), .B(n74), .C(rn_reg[86]), .D(n88), .Y(n1844)
         );
  AOI22X1 U2344 ( .A(rn_reg[174]), .B(n97), .C(rn_reg[222]), .D(n72), .Y(n1840) );
  AOI22X1 U2345 ( .A(rn_reg[46]), .B(n97), .C(rn_reg[94]), .D(n72), .Y(n1848)
         );
  AOI21X1 U2346 ( .B(n2481), .C(temp2_comb[7]), .A(n1366), .Y(n1068) );
  AOI22X1 U2347 ( .A(rn_reg[118]), .B(n162), .C(rn_reg[22]), .D(n145), .Y(
        n1843) );
  AOI22X1 U2348 ( .A(rn_reg[254]), .B(n99), .C(rn_reg[158]), .D(n158), .Y(
        n1839) );
  AOI22X1 U2349 ( .A(rn_reg[126]), .B(n99), .C(rn_reg[30]), .D(n158), .Y(n1847) );
  AOI22X1 U2350 ( .A(rn_reg[190]), .B(n117), .C(rn_reg[198]), .D(n141), .Y(
        n1838) );
  AOI22X1 U2351 ( .A(rn_reg[62]), .B(n117), .C(rn_reg[70]), .D(n141), .Y(n1846) );
  AOI21X1 U2352 ( .B(dec_cop[6]), .C(n1063), .A(n2484), .Y(n1065) );
  OAI21AX1 U2353 ( .B(n2073), .C(n2074), .A(n748), .Y(n2069) );
  AOI22X1 U2354 ( .A(n744), .B(n745), .C(n1639), .D(n774), .Y(n2073) );
  AOI32X1 U2355 ( .A(n970), .B(n64), .C(interrupt), .D(instr[6]), .E(n750), 
        .Y(n2074) );
  AOI211X1 U2356 ( .C(n1061), .D(n1062), .A(n2307), .B(n2309), .Y(n1060) );
  INVX1 U2357 ( .A(n1056), .Y(n2309) );
  OAI211X1 U2358 ( .C(c), .D(n1063), .A(n1055), .B(dec_cop[5]), .Y(n1062) );
  OAI21X1 U2359 ( .B(n2288), .C(c), .A(dec_cop[3]), .Y(n1061) );
  AOI22X1 U2360 ( .A(rn_reg[242]), .B(n162), .C(rn_reg[146]), .D(n145), .Y(
        n1936) );
  AOI22X1 U2361 ( .A(rn_reg[250]), .B(n99), .C(rn_reg[154]), .D(n158), .Y(
        n1940) );
  AOI22X1 U2362 ( .A(n1145), .B(dpl_reg[4]), .C(n1146), .D(dpl_reg[12]), .Y(
        n1185) );
  AOI22X1 U2363 ( .A(n1145), .B(dpl_reg[5]), .C(n1146), .D(dpl_reg[13]), .Y(
        n1175) );
  AOI22X1 U2364 ( .A(rn_reg[186]), .B(n117), .C(rn_reg[194]), .D(n141), .Y(
        n1939) );
  AOI22X1 U2365 ( .A(n1147), .B(dpl_reg[20]), .C(n1148), .D(dpl_reg[28]), .Y(
        n1184) );
  AOI22X1 U2366 ( .A(rn_reg[162]), .B(n74), .C(rn_reg[210]), .D(n88), .Y(n1937) );
  AOI22X1 U2367 ( .A(rn_reg[170]), .B(n97), .C(rn_reg[218]), .D(n72), .Y(n1941) );
  AOI22X1 U2368 ( .A(rn_reg[226]), .B(n121), .C(rn_reg[130]), .D(n101), .Y(
        n1938) );
  INVX1 U2369 ( .A(dps[0]), .Y(n2365) );
  NAND4X1 U2370 ( .A(n503), .B(n504), .C(n505), .D(n506), .Y(dpl[7]) );
  AOI22X1 U2371 ( .A(n223), .B(dpl_reg[47]), .C(n225), .D(dpl_reg[63]), .Y(
        n503) );
  AOI22X1 U2372 ( .A(n509), .B(dpl_reg[15]), .C(n232), .D(dpl_reg[31]), .Y(
        n505) );
  AOI22X1 U2373 ( .A(n227), .B(dpl_reg[39]), .C(n229), .D(dpl_reg[55]), .Y(
        n504) );
  INVX1 U2374 ( .A(dps[3]), .Y(n2374) );
  AO222X1 U2375 ( .A(n2234), .B(temp[3]), .C(dptr_inc[11]), .D(n1138), .E(
        n1235), .F(n2132), .Y(n2122) );
  AO222X1 U2376 ( .A(n2234), .B(temp[2]), .C(dptr_inc[10]), .D(n1138), .E(
        n2126), .F(n1235), .Y(n1410) );
  AO222X1 U2377 ( .A(n2234), .B(temp[1]), .C(dptr_inc[9]), .D(n1138), .E(n2133), .F(n1235), .Y(n991) );
  NAND43X1 U2378 ( .B(n2509), .C(n38), .D(n169), .A(n1980), .Y(n1742) );
  OAI221X1 U2379 ( .A(instr[1]), .B(n1774), .C(n603), .D(n2431), .E(n1981), 
        .Y(n1980) );
  OAI21BBX1 U2380 ( .A(n1633), .B(n2449), .C(n2508), .Y(n1981) );
  NAND21X1 U2381 ( .B(n1532), .A(n1520), .Y(n650) );
  OAI21X1 U2382 ( .B(n773), .C(n2360), .A(n1648), .Y(n1520) );
  AOI32X1 U2383 ( .A(phase[0]), .B(n1649), .C(n1644), .D(phase[1]), .E(n1650), 
        .Y(n1648) );
  OAI32X1 U2384 ( .A(n773), .B(n62), .C(n2425), .D(n1651), .E(n2416), .Y(n1650) );
  INVX1 U2385 ( .A(n303), .Y(n323) );
  NAND32X1 U2386 ( .B(n2505), .C(n1014), .A(n2242), .Y(n303) );
  NOR42XL U2387 ( .C(ramsfraddr[3]), .D(n1102), .A(ramsfraddr[4]), .B(n847), 
        .Y(n871) );
  NAND43X1 U2388 ( .B(n2246), .C(n606), .D(n605), .A(n1745), .Y(n1652) );
  NAND3X1 U2389 ( .A(intcall), .B(n1752), .C(n1639), .Y(n1745) );
  INVX1 U2390 ( .A(n1744), .Y(n606) );
  AO222X1 U2391 ( .A(n1747), .B(phase[0]), .C(n1749), .D(n604), .E(n1748), .F(
        phase[1]), .Y(n605) );
  INVX1 U2392 ( .A(n2510), .Y(n2324) );
  OAI31XL U2393 ( .A(n581), .B(n768), .C(n583), .D(phase[1]), .Y(n383) );
  OAI31XL U2394 ( .A(n305), .B(n2418), .C(n147), .D(n2094), .Y(n1579) );
  NAND4X1 U2395 ( .A(n601), .B(n1324), .C(instr[4]), .D(n602), .Y(n2094) );
  AOI32X1 U2396 ( .A(n1649), .B(n602), .C(n1756), .D(n965), .E(n2504), .Y(n305) );
  NAND3X1 U2397 ( .A(n1775), .B(n2509), .C(n1756), .Y(n902) );
  AOI22X1 U2398 ( .A(n2448), .B(n2505), .C(n2506), .D(n2253), .Y(n1774) );
  NOR2X1 U2399 ( .A(n2262), .B(n2506), .Y(n789) );
  NOR2X1 U2400 ( .A(n2449), .B(n2505), .Y(n971) );
  NOR2X1 U2401 ( .A(n33), .B(n2507), .Y(n2091) );
  NOR2X1 U2402 ( .A(n1099), .B(n2510), .Y(n233) );
  NOR2X1 U2403 ( .A(n1098), .B(n2510), .Y(n231) );
  NOR2X1 U2404 ( .A(n1098), .B(n2510), .Y(n509) );
  NAND4X1 U2405 ( .A(n1316), .B(n1317), .C(n1318), .D(n1319), .Y(dpc[2]) );
  AOI22X1 U2406 ( .A(dpc_tab[32]), .B(n224), .C(dpc_tab[44]), .D(n226), .Y(
        n1316) );
  AOI22X1 U2407 ( .A(dpc_tab[8]), .B(n24), .C(dpc_tab[20]), .D(n232), .Y(n1318) );
  AOI22X1 U2408 ( .A(dpc_tab[26]), .B(n228), .C(dpc_tab[38]), .D(n230), .Y(
        n1317) );
  NOR2X1 U2409 ( .A(n1095), .B(n2510), .Y(n232) );
  OAI22X1 U2410 ( .A(n2208), .B(n1139), .C(n2401), .D(n1158), .Y(n2134) );
  AND4X1 U2411 ( .A(n1159), .B(n1160), .C(n1161), .D(n1162), .Y(n1158) );
  AOI22X1 U2412 ( .A(n1151), .B(dpl_reg[54]), .C(n1152), .D(dpl_reg[62]), .Y(
        n1159) );
  AOI22X1 U2413 ( .A(n1149), .B(dpl_reg[38]), .C(n1150), .D(dpl_reg[46]), .Y(
        n1160) );
  OAI21X1 U2414 ( .B(dec_cop[3]), .C(dec_cop[4]), .A(n123), .Y(n1055) );
  NAND2X1 U2415 ( .A(dps[1]), .B(dps[0]), .Y(n1095) );
  NAND2X1 U2416 ( .A(dps[0]), .B(n2363), .Y(n1098) );
  NOR2X1 U2417 ( .A(n2397), .B(n2509), .Y(n1764) );
  INVX1 U2418 ( .A(phase[2]), .Y(n2245) );
  NAND3X1 U2419 ( .A(ramsfraddr[1]), .B(ramsfraddr[2]), .C(ramsfraddr[0]), .Y(
        n848) );
  AOI22X1 U2420 ( .A(dpc_tab[0]), .B(n22), .C(dpc_tab[12]), .D(n234), .Y(n1315) );
  AOI22X1 U2421 ( .A(dpc_tab[4]), .B(n22), .C(dpc_tab[16]), .D(n234), .Y(n1088) );
  AOI22X1 U2422 ( .A(dpc_tab[5]), .B(n22), .C(dpc_tab[17]), .D(n19), .Y(n1084)
         );
  AOI22X1 U2423 ( .A(dpc_tab[2]), .B(n233), .C(dpc_tab[14]), .D(n19), .Y(n1319) );
  AOI22X1 U2424 ( .A(n22), .B(dph_reg[1]), .C(n19), .D(dph_reg[17]), .Y(n570)
         );
  AOI22X1 U2425 ( .A(n233), .B(dph_reg[3]), .C(n508), .D(dph_reg[19]), .Y(n562) );
  AOI22X1 U2426 ( .A(n21), .B(dpl_reg[0]), .C(n508), .D(dpl_reg[16]), .Y(n542)
         );
  AOI22X1 U2427 ( .A(n22), .B(dph_reg[0]), .C(n234), .D(dph_reg[16]), .Y(n574)
         );
  AOI22X1 U2428 ( .A(n21), .B(dpl_reg[4]), .C(n508), .D(dpl_reg[20]), .Y(n526)
         );
  AOI22X1 U2429 ( .A(n22), .B(dph_reg[5]), .C(n19), .D(dph_reg[21]), .Y(n554)
         );
  AOI22X1 U2430 ( .A(n233), .B(dpl_reg[5]), .C(n508), .D(dpl_reg[21]), .Y(n522) );
  AOI22X1 U2431 ( .A(n21), .B(dpl_reg[6]), .C(n234), .D(dpl_reg[22]), .Y(n518)
         );
  AOI22X1 U2432 ( .A(n22), .B(dph_reg[2]), .C(n508), .D(dph_reg[18]), .Y(n566)
         );
  AOI22X1 U2433 ( .A(n21), .B(dpl_reg[2]), .C(n508), .D(dpl_reg[18]), .Y(n534)
         );
  AOI22X1 U2434 ( .A(n509), .B(dpl_reg[8]), .C(n26), .D(dpl_reg[24]), .Y(n541)
         );
  AOI22X1 U2435 ( .A(n509), .B(dph_reg[12]), .C(n26), .D(dph_reg[28]), .Y(n557) );
  AOI22X1 U2436 ( .A(n509), .B(dpl_reg[12]), .C(n26), .D(dpl_reg[28]), .Y(n525) );
  AOI22X1 U2437 ( .A(n24), .B(dph_reg[13]), .C(n27), .D(dph_reg[29]), .Y(n553)
         );
  AOI22X1 U2438 ( .A(n509), .B(dpl_reg[13]), .C(n26), .D(dpl_reg[29]), .Y(n521) );
  AOI22X1 U2439 ( .A(n231), .B(dph_reg[14]), .C(n27), .D(dph_reg[30]), .Y(n549) );
  AOI22X1 U2440 ( .A(n509), .B(dpl_reg[14]), .C(n26), .D(dpl_reg[30]), .Y(n517) );
  AOI22X1 U2441 ( .A(n228), .B(dph_reg[33]), .C(n230), .D(dph_reg[49]), .Y(
        n568) );
  AOI22X1 U2442 ( .A(n227), .B(dph_reg[35]), .C(n229), .D(dph_reg[51]), .Y(
        n560) );
  AOI22X1 U2443 ( .A(n511), .B(dpl_reg[32]), .C(n512), .D(dpl_reg[48]), .Y(
        n540) );
  AOI22X1 U2444 ( .A(n227), .B(dph_reg[32]), .C(n229), .D(dph_reg[48]), .Y(
        n572) );
  AOI22X1 U2445 ( .A(n228), .B(dph_reg[36]), .C(n230), .D(dph_reg[52]), .Y(
        n556) );
  AOI22X1 U2446 ( .A(n227), .B(dpl_reg[36]), .C(n229), .D(dpl_reg[52]), .Y(
        n524) );
  AOI22X1 U2447 ( .A(n511), .B(dph_reg[37]), .C(n512), .D(dph_reg[53]), .Y(
        n552) );
  AOI22X1 U2448 ( .A(n228), .B(dpl_reg[37]), .C(n230), .D(dpl_reg[53]), .Y(
        n520) );
  AOI22X1 U2449 ( .A(n227), .B(dph_reg[38]), .C(n229), .D(dph_reg[54]), .Y(
        n548) );
  AOI22X1 U2450 ( .A(n511), .B(dpl_reg[38]), .C(n512), .D(dpl_reg[54]), .Y(
        n516) );
  AOI22X1 U2451 ( .A(n511), .B(dph_reg[34]), .C(n512), .D(dph_reg[50]), .Y(
        n564) );
  AOI22X1 U2452 ( .A(n228), .B(dpl_reg[34]), .C(n230), .D(dpl_reg[50]), .Y(
        n532) );
  AOI22X1 U2453 ( .A(n513), .B(dpl_reg[40]), .C(n514), .D(dpl_reg[56]), .Y(
        n539) );
  AOI22X1 U2454 ( .A(n224), .B(dph_reg[44]), .C(n226), .D(dph_reg[60]), .Y(
        n555) );
  AOI22X1 U2455 ( .A(n513), .B(dph_reg[45]), .C(n514), .D(dph_reg[61]), .Y(
        n551) );
  AOI22X1 U2456 ( .A(n223), .B(dph_reg[46]), .C(n225), .D(dph_reg[62]), .Y(
        n547) );
  AOI22X1 U2457 ( .A(n513), .B(dpl_reg[46]), .C(n514), .D(dpl_reg[62]), .Y(
        n515) );
  INVX1 U2458 ( .A(acc[2]), .Y(n2475) );
  NAND2X1 U2459 ( .A(n2507), .B(n126), .Y(n2030) );
  NOR2X1 U2460 ( .A(n2434), .B(n2507), .Y(n1639) );
  NAND3X1 U2461 ( .A(ramsfraddr[2]), .B(n2443), .C(ramsfraddr[1]), .Y(n847) );
  NAND2X1 U2462 ( .A(instr[1]), .B(n2506), .Y(n603) );
  AOI22X1 U2463 ( .A(n1145), .B(dpl_reg[6]), .C(n1146), .D(dpl_reg[14]), .Y(
        n1162) );
  AOI22X1 U2464 ( .A(n1147), .B(dpl_reg[21]), .C(n1148), .D(dpl_reg[29]), .Y(
        n1174) );
  AOI22X1 U2465 ( .A(n1147), .B(dpl_reg[22]), .C(n1148), .D(dpl_reg[30]), .Y(
        n1161) );
  NAND4X1 U2466 ( .A(n1312), .B(n1313), .C(n1314), .D(n1315), .Y(dpc[0]) );
  AOI22X1 U2467 ( .A(dpc_tab[30]), .B(n513), .C(dpc_tab[42]), .D(n514), .Y(
        n1312) );
  AOI22X1 U2468 ( .A(dpc_tab[6]), .B(n231), .C(dpc_tab[18]), .D(n27), .Y(n1314) );
  AOI22X1 U2469 ( .A(dpc_tab[24]), .B(n511), .C(dpc_tab[36]), .D(n512), .Y(
        n1313) );
  NAND3X1 U2470 ( .A(n17), .B(n2506), .C(n2227), .Y(n1013) );
  INVX1 U2471 ( .A(dps[1]), .Y(n2363) );
  OAI211X1 U2472 ( .C(n1651), .D(n2416), .A(n1750), .B(n1751), .Y(n1748) );
  AOI32X1 U2473 ( .A(interrupt), .B(n1752), .C(n1639), .D(n1736), .E(n1753), 
        .Y(n1751) );
  ENOX1 U2474 ( .A(n2425), .B(n2262), .C(n2261), .D(n2242), .Y(n1753) );
  GEN2XL U2475 ( .D(n744), .E(n745), .C(n746), .B(n747), .A(n748), .Y(n614) );
  EORX1 U2476 ( .A(n749), .B(n64), .C(n750), .D(n64), .Y(n747) );
  OAI211X1 U2477 ( .C(n751), .D(n69), .A(n752), .B(n753), .Y(n749) );
  OAI21X1 U2478 ( .B(instr[4]), .C(n2248), .A(n69), .Y(n752) );
  AOI31X1 U2479 ( .A(instr[4]), .B(n2190), .C(n2420), .D(n2256), .Y(n1761) );
  NAND4X1 U2480 ( .A(n1085), .B(n1086), .C(n1087), .D(n1088), .Y(dpc[4]) );
  AOI22X1 U2481 ( .A(dpc_tab[34]), .B(n224), .C(dpc_tab[46]), .D(n226), .Y(
        n1085) );
  AOI22X1 U2482 ( .A(dpc_tab[10]), .B(n231), .C(dpc_tab[22]), .D(n27), .Y(
        n1087) );
  AOI22X1 U2483 ( .A(dpc_tab[28]), .B(n228), .C(dpc_tab[40]), .D(n230), .Y(
        n1086) );
  NAND4X1 U2484 ( .A(n1081), .B(n1082), .C(n1083), .D(n1084), .Y(dpc[5]) );
  AOI22X1 U2485 ( .A(dpc_tab[35]), .B(n513), .C(dpc_tab[47]), .D(n514), .Y(
        n1081) );
  AOI22X1 U2486 ( .A(dpc_tab[11]), .B(n24), .C(dpc_tab[23]), .D(n27), .Y(n1083) );
  AOI22X1 U2487 ( .A(dpc_tab[29]), .B(n511), .C(dpc_tab[41]), .D(n512), .Y(
        n1082) );
  INVX1 U2488 ( .A(temp2_comb[3]), .Y(n2438) );
  INVX1 U2489 ( .A(temp2_comb[6]), .Y(n2358) );
  INVX1 U2490 ( .A(N345), .Y(n2223) );
  GEN2XL U2491 ( .D(n1627), .E(n436), .C(n261), .B(n423), .A(n2264), .Y(n424)
         );
  AOI32X1 U2492 ( .A(n1639), .B(phase[3]), .C(n751), .D(n1640), .E(phase[2]), 
        .Y(n423) );
  NAND41X1 U2493 ( .D(n767), .A(n2382), .B(n1011), .C(n1641), .Y(n1640) );
  AOI31X1 U2494 ( .A(n774), .B(instr[2]), .C(n2252), .D(n808), .Y(n1641) );
  AO222X1 U2495 ( .A(n2234), .B(temp[4]), .C(dptr_inc[12]), .D(n1138), .E(
        n1235), .F(n2131), .Y(n2123) );
  AO222X1 U2496 ( .A(n2234), .B(temp[5]), .C(dptr_inc[13]), .D(n1138), .E(
        n1235), .F(n2130), .Y(n2124) );
  AO222X1 U2497 ( .A(n2234), .B(temp[6]), .C(dptr_inc[14]), .D(n1138), .E(
        n1235), .F(n2129), .Y(n2125) );
  AO21X1 U2498 ( .B(n371), .C(N345), .A(n1887), .Y(n473) );
  NAND21X1 U2499 ( .B(n2396), .A(n2507), .Y(n392) );
  NAND32X1 U2500 ( .B(ramsfraddr[7]), .C(n1372), .A(n425), .Y(n1498) );
  NAND21X1 U2501 ( .B(n779), .A(phase[2]), .Y(n370) );
  AOI32X1 U2502 ( .A(n2180), .B(n751), .C(n2508), .D(n973), .E(n1644), .Y(
        n1627) );
  NOR21XL U2503 ( .B(dec_cop[7]), .A(dec_cop[6]), .Y(n1066) );
  OR3XL U2504 ( .A(n2506), .B(n620), .C(n774), .Y(n1609) );
  NAND43X1 U2505 ( .B(n2098), .C(n2097), .D(n580), .A(n776), .Y(n306) );
  OAI222XL U2506 ( .A(n1632), .B(n2416), .C(n2100), .D(n2436), .E(n603), .F(
        n2431), .Y(n2098) );
  OAI211X1 U2507 ( .C(instr[1]), .D(n2101), .A(n2102), .B(n2103), .Y(n2097) );
  AOI31X1 U2508 ( .A(n2092), .B(n2261), .C(n774), .D(n2104), .Y(n2103) );
  NAND2X1 U2509 ( .A(n956), .B(phase[0]), .Y(n909) );
  NOR2X1 U2510 ( .A(n2392), .B(instr[6]), .Y(n965) );
  NAND2X1 U2511 ( .A(n2420), .B(n1325), .Y(n1090) );
  OAI21X1 U2512 ( .B(n786), .C(n809), .A(n1326), .Y(n1325) );
  NAND4X1 U2513 ( .A(n745), .B(phase[1]), .C(n1324), .D(n128), .Y(n1326) );
  OAI22X1 U2514 ( .A(n2195), .B(n1139), .C(n2401), .D(n1140), .Y(n2144) );
  AND4X1 U2515 ( .A(n1141), .B(n1142), .C(n1143), .D(n1144), .Y(n1140) );
  AOI22X1 U2516 ( .A(n1151), .B(dpl_reg[55]), .C(n1152), .D(dpl_reg[63]), .Y(
        n1141) );
  AOI22X1 U2517 ( .A(n1149), .B(dpl_reg[39]), .C(n1150), .D(dpl_reg[47]), .Y(
        n1142) );
  NAND2X1 U2518 ( .A(dec_cop[2]), .B(n123), .Y(n1054) );
  NAND2X1 U2519 ( .A(n76), .B(n1622), .Y(n976) );
  NAND4X1 U2520 ( .A(phase[0]), .B(n2508), .C(n751), .D(n746), .Y(n1622) );
  NAND2X1 U2521 ( .A(dec_cop[1]), .B(n123), .Y(n1056) );
  AND2XL U2522 ( .A(sfroe_r), .B(n283), .Y(sfroe) );
  AOI22X1 U2523 ( .A(dpc_tab[1]), .B(n21), .C(dpc_tab[13]), .D(n508), .Y(n1323) );
  AOI22X1 U2524 ( .A(dpc_tab[3]), .B(n233), .C(dpc_tab[15]), .D(n234), .Y(
        n1094) );
  AOI22X1 U2525 ( .A(n21), .B(dpl_reg[1]), .C(n19), .D(dpl_reg[17]), .Y(n538)
         );
  AOI22X1 U2526 ( .A(n233), .B(dpl_reg[3]), .C(n234), .D(dpl_reg[19]), .Y(n530) );
  AOI22X1 U2527 ( .A(n233), .B(dph_reg[7]), .C(n508), .D(dph_reg[23]), .Y(n546) );
  AOI22X1 U2528 ( .A(n231), .B(dph_reg[8]), .C(n27), .D(dph_reg[24]), .Y(n573)
         );
  AOI22X1 U2529 ( .A(n24), .B(dpl_reg[9]), .C(n232), .D(dpl_reg[25]), .Y(n537)
         );
  AOI22X1 U2530 ( .A(n231), .B(dpl_reg[11]), .C(n232), .D(dpl_reg[27]), .Y(
        n529) );
  AOI22X1 U2531 ( .A(n509), .B(dph_reg[15]), .C(n232), .D(dph_reg[31]), .Y(
        n545) );
  AOI22X1 U2532 ( .A(n509), .B(dpl_reg[10]), .C(n26), .D(dpl_reg[26]), .Y(n533) );
  AOI22X1 U2533 ( .A(n227), .B(dpl_reg[33]), .C(n229), .D(dpl_reg[49]), .Y(
        n536) );
  AOI22X1 U2534 ( .A(n511), .B(dpl_reg[35]), .C(n512), .D(dpl_reg[51]), .Y(
        n528) );
  AOI22X1 U2535 ( .A(n228), .B(dph_reg[39]), .C(n230), .D(dph_reg[55]), .Y(
        n544) );
  AOI22X1 U2536 ( .A(n602), .B(phase[3]), .C(phase[1]), .D(n2315), .Y(n786) );
  NAND4X1 U2537 ( .A(n1320), .B(n1321), .C(n1322), .D(n1323), .Y(dpc[1]) );
  AOI22X1 U2538 ( .A(dpc_tab[31]), .B(n224), .C(dpc_tab[43]), .D(n226), .Y(
        n1320) );
  AOI22X1 U2539 ( .A(dpc_tab[25]), .B(n228), .C(dpc_tab[37]), .D(n230), .Y(
        n1321) );
  AOI22X1 U2540 ( .A(dpc_tab[7]), .B(n509), .C(dpc_tab[19]), .D(n26), .Y(n1322) );
  NOR2X1 U2541 ( .A(n2243), .B(n2504), .Y(n969) );
  AOI32X1 U2542 ( .A(instr[6]), .B(n2190), .C(n1723), .D(n1005), .E(n2432), 
        .Y(n1772) );
  NAND43X1 U2543 ( .B(instr[1]), .C(instr[3]), .D(n260), .A(n1628), .Y(n422)
         );
  OAI21X1 U2544 ( .B(n1629), .C(n62), .A(n1630), .Y(n1628) );
  NAND4X1 U2545 ( .A(n2253), .B(n2396), .C(n62), .D(n32), .Y(n1630) );
  AOI221XL U2546 ( .A(n969), .B(n970), .C(n965), .D(instr[5]), .E(n1631), .Y(
        n1629) );
  AOI22X1 U2547 ( .A(n1145), .B(dpl_reg[7]), .C(n1146), .D(dpl_reg[15]), .Y(
        n1144) );
  AOI22X1 U2548 ( .A(n1147), .B(dpl_reg[23]), .C(n1148), .D(dpl_reg[31]), .Y(
        n1143) );
  OAI22X1 U2549 ( .A(n1768), .B(n169), .C(n584), .D(n261), .Y(n1611) );
  NOR4XL U2550 ( .A(n1769), .B(n1770), .C(n768), .D(n1771), .Y(n1768) );
  AO2222XL U2551 ( .A(n2270), .B(n2449), .C(n1005), .D(n2269), .E(n2424), .F(
        n2398), .G(n1762), .H(n2243), .Y(n1769) );
  OAI32X1 U2552 ( .A(n2391), .B(instr[3]), .C(n2427), .D(n1772), .E(n1773), 
        .Y(n1770) );
  NAND4X1 U2553 ( .A(n1091), .B(n1092), .C(n1093), .D(n1094), .Y(dpc[3]) );
  AOI22X1 U2554 ( .A(dpc_tab[33]), .B(n223), .C(dpc_tab[45]), .D(n225), .Y(
        n1091) );
  AOI22X1 U2555 ( .A(dpc_tab[9]), .B(n231), .C(dpc_tab[21]), .D(n232), .Y(
        n1093) );
  AOI22X1 U2556 ( .A(dpc_tab[27]), .B(n227), .C(dpc_tab[39]), .D(n229), .Y(
        n1092) );
  INVX1 U2557 ( .A(c), .Y(n2484) );
  NAND2X1 U2558 ( .A(n2504), .B(n2243), .Y(n1633) );
  INVX1 U2559 ( .A(temp2_comb[0]), .Y(n825) );
  NAND21X1 U2560 ( .B(n391), .A(n390), .Y(n1435) );
  AND2X1 U2561 ( .A(n387), .B(phase[0]), .Y(n391) );
  NAND21X1 U2562 ( .B(n259), .A(n389), .Y(n390) );
  NAND21X1 U2563 ( .B(n581), .A(n388), .Y(n389) );
  NAND21X1 U2564 ( .B(n169), .A(n2507), .Y(n2360) );
  INVX1 U2565 ( .A(temp[4]), .Y(n2286) );
  INVX1 U2566 ( .A(temp[3]), .Y(n2289) );
  OAI22X1 U2567 ( .A(n2400), .B(n1327), .C(n2203), .D(n1236), .Y(n2140) );
  AND4X1 U2568 ( .A(n1328), .B(n1329), .C(n1330), .D(n1331), .Y(n1327) );
  AOI22X1 U2569 ( .A(n1151), .B(dph_reg[48]), .C(n1152), .D(dph_reg[56]), .Y(
        n1328) );
  AOI22X1 U2570 ( .A(n1149), .B(dph_reg[32]), .C(n1150), .D(dph_reg[40]), .Y(
        n1329) );
  OAI22X1 U2571 ( .A(n2199), .B(n1236), .C(n2400), .D(n1303), .Y(n2133) );
  AND4X1 U2572 ( .A(n1304), .B(n1305), .C(n1306), .D(n1307), .Y(n1303) );
  AOI22X1 U2573 ( .A(n166), .B(dph_reg[49]), .C(n105), .D(dph_reg[57]), .Y(
        n1304) );
  AOI22X1 U2574 ( .A(n125), .B(dph_reg[33]), .C(n149), .D(dph_reg[41]), .Y(
        n1305) );
  OAI21X1 U2575 ( .B(instr[4]), .C(n2448), .A(n2430), .Y(n2092) );
  OAI31XL U2576 ( .A(n2433), .B(instr[4]), .C(n805), .D(n2267), .Y(n799) );
  INVX1 U2577 ( .A(ramdatao[0]), .Y(n2203) );
  INVX1 U2578 ( .A(ramdatao[5]), .Y(n2212) );
  OAI21X1 U2579 ( .B(n2435), .C(n2075), .A(n2076), .Y(n748) );
  GEN2XL U2580 ( .D(n2426), .E(n2428), .C(instr[7]), .B(n2261), .A(n2080), .Y(
        n2075) );
  GEN2XL U2581 ( .D(instr[0]), .E(n109), .C(n2077), .B(n2078), .A(n2079), .Y(
        n2076) );
  AOI21X1 U2582 ( .B(instr[7]), .C(instr[4]), .A(n788), .Y(n2080) );
  EORX1 U2583 ( .A(n2087), .B(n2088), .C(n2052), .D(n2089), .Y(n2086) );
  OAI222XL U2584 ( .A(interrupt), .B(n2449), .C(n1756), .D(n2504), .E(instr[0]), .F(n2446), .Y(n2088) );
  OAI21X1 U2585 ( .B(n2428), .C(n2437), .A(n2090), .Y(n2087) );
  INVX1 U2586 ( .A(n1649), .Y(n2446) );
  AOI33X1 U2587 ( .A(n2091), .B(n2262), .C(n1649), .D(n2270), .E(instr[7]), 
        .F(n2505), .Y(n2090) );
  AOI22X1 U2588 ( .A(n1145), .B(dph_reg[0]), .C(n1146), .D(dph_reg[8]), .Y(
        n1331) );
  AOI22X1 U2589 ( .A(n104), .B(dph_reg[1]), .C(n165), .D(dph_reg[9]), .Y(n1307) );
  AOI32X1 U2590 ( .A(instr[1]), .B(n39), .C(n1763), .D(n971), .E(n2261), .Y(
        n2079) );
  AOI22X1 U2591 ( .A(n1147), .B(dph_reg[16]), .C(n1148), .D(dph_reg[24]), .Y(
        n1330) );
  AOI22X1 U2592 ( .A(n148), .B(dph_reg[17]), .C(n124), .D(dph_reg[25]), .Y(
        n1306) );
  NOR2X1 U2593 ( .A(instr[6]), .B(n2505), .Y(n1763) );
  AO222X1 U2594 ( .A(n2234), .B(temp[7]), .C(n1138), .D(dptr_inc[15]), .E(
        n1235), .F(n2128), .Y(n2141) );
  OAI22X1 U2595 ( .A(n1236), .B(n2195), .C(n1237), .D(n2400), .Y(n2128) );
  AND4X1 U2596 ( .A(n1238), .B(n1239), .C(n1240), .D(n1241), .Y(n1237) );
  NAND21X1 U2597 ( .B(N344), .A(N343), .Y(n2323) );
  NAND21X1 U2598 ( .B(N343), .A(N344), .Y(n823) );
  NAND21X1 U2599 ( .B(n343), .A(N344), .Y(n824) );
  AOI21BBXL U2600 ( .B(n2082), .C(n2083), .A(instr[3]), .Y(n744) );
  XNOR2XL U2601 ( .A(n2262), .B(n2186), .Y(n2082) );
  XNOR2XL U2602 ( .A(n2186), .B(n2509), .Y(n2083) );
  MUX2X1 U2603 ( .D0(n799), .D1(n800), .S(n806), .Y(n607) );
  OAI22X1 U2604 ( .A(n819), .B(n820), .C(n821), .D(n822), .Y(n806) );
  OAI22X1 U2605 ( .A(n2478), .B(n2322), .C(n2323), .D(n2477), .Y(n820) );
  OAI21X1 U2606 ( .B(n2403), .C(n2322), .A(N345), .Y(n822) );
  OAI22X1 U2607 ( .A(n2192), .B(n1236), .C(n2400), .D(n1292), .Y(n2126) );
  AND4X1 U2608 ( .A(n1293), .B(n1294), .C(n1295), .D(n1296), .Y(n1292) );
  AOI22X1 U2609 ( .A(n166), .B(dph_reg[50]), .C(n105), .D(dph_reg[58]), .Y(
        n1293) );
  AOI22X1 U2610 ( .A(n125), .B(dph_reg[34]), .C(n149), .D(dph_reg[42]), .Y(
        n1294) );
  INVX1 U2611 ( .A(N343), .Y(n343) );
  AOI22X1 U2612 ( .A(n104), .B(dph_reg[2]), .C(n165), .D(dph_reg[10]), .Y(
        n1296) );
  AOI22X1 U2613 ( .A(n148), .B(dph_reg[18]), .C(n124), .D(dph_reg[26]), .Y(
        n1295) );
  INVX1 U2614 ( .A(dec_accop[9]), .Y(n2482) );
  INVX1 U2615 ( .A(dec_accop[10]), .Y(n2487) );
  INVX1 U2616 ( .A(temp[1]), .Y(n2317) );
  INVX1 U2617 ( .A(temp[0]), .Y(n2320) );
  INVX1 U2618 ( .A(temp[5]), .Y(n2318) );
  AOI221XL U2619 ( .A(n984), .B(memdatai[3]), .C(n983), .D(pc_o[11]), .E(n992), 
        .Y(n640) );
  OAI22X1 U2620 ( .A(n2326), .B(n986), .C(n2346), .D(n2492), .Y(n992) );
  NAND21X1 U2621 ( .B(N344), .A(n343), .Y(n2322) );
  MUX2X1 U2622 ( .D0(ramsfraddr[4]), .D1(n1694), .S(n284), .Y(
        ramsfraddr_comb[4]) );
  AO21X1 U2623 ( .B(n2255), .C(instr[4]), .A(israccess), .Y(n1505) );
  OAI22X1 U2624 ( .A(n1236), .B(n12), .C(n1281), .D(n2400), .Y(n2132) );
  AND4X1 U2625 ( .A(n1282), .B(n1283), .C(n1284), .D(n1285), .Y(n1281) );
  AOI22X1 U2626 ( .A(n166), .B(dph_reg[51]), .C(n105), .D(dph_reg[59]), .Y(
        n1282) );
  AOI22X1 U2628 ( .A(n125), .B(dph_reg[35]), .C(n149), .D(dph_reg[43]), .Y(
        n1283) );
  OAI22X1 U2629 ( .A(n1236), .B(n2216), .C(n1270), .D(n2400), .Y(n2131) );
  AND4X1 U2630 ( .A(n1271), .B(n1272), .C(n1273), .D(n1274), .Y(n1270) );
  AOI22X1 U2631 ( .A(n166), .B(dph_reg[52]), .C(n105), .D(dph_reg[60]), .Y(
        n1271) );
  AOI22X1 U2632 ( .A(n125), .B(dph_reg[36]), .C(n149), .D(dph_reg[44]), .Y(
        n1272) );
  OAI22XL U2633 ( .A(n292), .B(n978), .C(n975), .D(n1503), .Y(N12720) );
  AOI221XL U2634 ( .A(n984), .B(memdatai[6]), .C(n983), .D(pc_o[14]), .E(n985), 
        .Y(n978) );
  OAI22X1 U2635 ( .A(n2316), .B(n986), .C(n2346), .D(n2491), .Y(n985) );
  AOI22X1 U2636 ( .A(n104), .B(dph_reg[3]), .C(n165), .D(dph_reg[11]), .Y(
        n1285) );
  AOI22X1 U2637 ( .A(n104), .B(dph_reg[4]), .C(n165), .D(dph_reg[12]), .Y(
        n1274) );
  AOI22X1 U2638 ( .A(n148), .B(dph_reg[19]), .C(n124), .D(dph_reg[27]), .Y(
        n1284) );
  OAI221X1 U2639 ( .A(n1342), .B(n1343), .C(n2290), .D(n1344), .E(n1345), .Y(
        N12484) );
  AOI22X1 U2640 ( .A(N13353), .B(n194), .C(N13352), .D(n2273), .Y(n1342) );
  AOI22X1 U2641 ( .A(n1346), .B(b[7]), .C(n1347), .D(n282), .Y(n1345) );
  INVX1 U2642 ( .A(interrupt), .Y(n2248) );
  INVX1 U2643 ( .A(temp[6]), .Y(n2319) );
  INVX1 U2644 ( .A(temp[2]), .Y(n2321) );
  MUX2X1 U2645 ( .D0(ramsfraddr[6]), .D1(n1696), .S(n284), .Y(
        ramsfraddr_comb[6]) );
  MUX2X1 U2646 ( .D0(ramsfraddr[5]), .D1(n1695), .S(n284), .Y(
        ramsfraddr_comb[5]) );
  OR2X1 U2647 ( .A(state[1]), .B(state[2]), .Y(n1572) );
  MUX2X1 U2648 ( .D0(ramsfraddr[7]), .D1(n1697), .S(n284), .Y(
        ramsfraddr_comb[7]) );
  MUX2X1 U2649 ( .D0(ramsfraddr[3]), .D1(n1693), .S(n284), .Y(
        ramsfraddr_comb[3]) );
  NAND21X1 U2650 ( .B(state[0]), .A(n1499), .Y(n1591) );
  INVX1 U2651 ( .A(n2156), .Y(n849) );
  NAND5XL U2652 ( .A(ramwe), .B(n2187), .C(n2189), .D(n243), .E(n2188), .Y(
        n2156) );
  INVX1 U2653 ( .A(n597), .Y(n2235) );
  NAND21X1 U2654 ( .B(n900), .A(temp[7]), .Y(n597) );
  AO2222XL U2655 ( .A(n1346), .B(b[2]), .C(n2281), .D(multemp2[4]), .E(n2282), 
        .F(n2412), .G(n1347), .H(n264), .Y(N12479) );
  INVX1 U2656 ( .A(n836), .Y(n2412) );
  AO2222XL U2657 ( .A(n1346), .B(b[3]), .C(n2281), .D(multemp2[5]), .E(n2282), 
        .F(n2411), .G(n1347), .H(n277), .Y(N12480) );
  INVX1 U2658 ( .A(n835), .Y(n2411) );
  AO2222XL U2659 ( .A(n1347), .B(n255), .C(n1346), .D(b[0]), .E(n2281), .F(
        multemp2[2]), .G(n2282), .H(n2414), .Y(N12477) );
  INVX1 U2660 ( .A(n838), .Y(n2414) );
  AO2222XL U2661 ( .A(n1347), .B(n251), .C(n1346), .D(b[1]), .E(n2281), .F(
        multemp2[3]), .G(n2282), .H(n2413), .Y(N12478) );
  INVX1 U2662 ( .A(n837), .Y(n2413) );
  AO2222XL U2663 ( .A(n1347), .B(n274), .C(n1346), .D(b[4]), .E(n2281), .F(
        multemp2[6]), .G(n2282), .H(n2410), .Y(N12481) );
  INVX1 U2664 ( .A(n834), .Y(n2410) );
  AO2222XL U2665 ( .A(n1346), .B(b[5]), .C(n2281), .D(multemp2[7]), .E(n1347), 
        .F(n271), .G(n2282), .H(n2409), .Y(N12482) );
  INVX1 U2666 ( .A(n833), .Y(n2409) );
  AO2222XL U2667 ( .A(n1347), .B(n268), .C(n1346), .D(b[6]), .E(n2281), .F(
        multemp2[8]), .G(n2282), .H(n2408), .Y(N12483) );
  INVX1 U2668 ( .A(n831), .Y(n2408) );
  INVX1 U2669 ( .A(n633), .Y(n2234) );
  NAND21X1 U2670 ( .B(n1013), .A(n262), .Y(n633) );
  MUX2X1 U2671 ( .D0(n264), .D1(gf0), .S(n478), .Y(n1881) );
  NOR2X1 U2672 ( .A(n291), .B(n479), .Y(n478) );
  AO22X1 U2673 ( .A(n1039), .B(n2211), .C(n268), .D(n2266), .Y(N12706) );
  OAI22AX1 U2674 ( .D(ac), .C(n1040), .A(n1041), .B(n1026), .Y(n1039) );
  AOI32X1 U2675 ( .A(n2487), .B(n2482), .C(N11555), .D(dec_accop[10]), .E(
        n2439), .Y(n1041) );
  NOR4XL U2676 ( .A(n1042), .B(n2336), .C(n1027), .D(n2353), .Y(n1040) );
  OAI22X1 U2677 ( .A(n1236), .B(n2212), .C(n1260), .D(n2400), .Y(n2130) );
  AND4X1 U2678 ( .A(n1261), .B(n1262), .C(n1263), .D(n1264), .Y(n1260) );
  AOI22X1 U2679 ( .A(n166), .B(dph_reg[53]), .C(n105), .D(dph_reg[61]), .Y(
        n1261) );
  AOI22X1 U2680 ( .A(n125), .B(dph_reg[37]), .C(n149), .D(dph_reg[45]), .Y(
        n1262) );
  NAND3X1 U2681 ( .A(finishdiv), .B(n1023), .C(n1348), .Y(n1343) );
  NAND3X1 U2682 ( .A(n1348), .B(n1349), .C(finishmul), .Y(n1344) );
  NAND3X1 U2683 ( .A(ramsfraddr[3]), .B(ramsfraddr[4]), .C(n849), .Y(n854) );
  NAND3X1 U2684 ( .A(ramsfraddr[3]), .B(n2405), .C(n849), .Y(n851) );
  INVX1 U2685 ( .A(ramdatao[6]), .Y(n2208) );
  AOI22X1 U2686 ( .A(n104), .B(dph_reg[5]), .C(n165), .D(dph_reg[13]), .Y(
        n1264) );
  AOI22X1 U2687 ( .A(n148), .B(dph_reg[20]), .C(n124), .D(dph_reg[28]), .Y(
        n1273) );
  AOI22X1 U2688 ( .A(n148), .B(dph_reg[21]), .C(n124), .D(dph_reg[29]), .Y(
        n1263) );
  INVX1 U2689 ( .A(phase[3]), .Y(n2238) );
  NAND31X1 U2690 ( .C(finishmul), .A(n840), .B(n239), .Y(n839) );
  OR3XL U2691 ( .A(finishdiv), .B(n248), .C(n2157), .Y(n832) );
  NAND21X1 U2692 ( .B(n769), .A(n106), .Y(n859) );
  NAND32X1 U2693 ( .B(p2sel), .C(n634), .A(n183), .Y(n1412) );
  AND2XL U2694 ( .A(phase0_ff), .B(n2500), .Y(newinstr) );
  NAND32X1 U2695 ( .B(p2sel), .C(n684), .A(n183), .Y(n1418) );
  INVX1 U2696 ( .A(n1613), .Y(n2150) );
  NAND32X1 U2697 ( .B(instr[5]), .C(n245), .A(n2158), .Y(n1613) );
  NOR32XL U2698 ( .B(n239), .C(n789), .A(n2051), .Y(N10566) );
  NAND3X1 U2699 ( .A(n39), .B(instr[0]), .C(n2050), .Y(n2051) );
  OA21X1 U2700 ( .B(n1404), .C(n1403), .A(n250), .Y(N12726) );
  AO2222XL U2701 ( .A(n2343), .B(pc_o[3]), .C(intvect[0]), .D(n2247), .E(n815), 
        .F(n1402), .G(ramdatai[3]), .H(n906), .Y(n1403) );
  OAI221X1 U2702 ( .A(n2451), .B(n1385), .C(n2438), .D(n1384), .E(n1383), .Y(
        n1404) );
  AOI21X1 U2703 ( .B(n913), .C(temp[3]), .A(n932), .Y(n1383) );
  OA21X1 U2704 ( .B(n645), .C(n644), .A(n250), .Y(N12727) );
  AO2222XL U2705 ( .A(n2343), .B(n2502), .C(intvect[1]), .D(n2247), .E(n816), 
        .F(n1402), .G(ramdatai[4]), .H(n906), .Y(n644) );
  OAI221X1 U2706 ( .A(n642), .B(n1385), .C(n669), .D(n1384), .E(n641), .Y(n645) );
  INVX1 U2707 ( .A(pc_i[12]), .Y(n642) );
  OA21X1 U2708 ( .B(n681), .C(n680), .A(n250), .Y(N12728) );
  AO2222XL U2709 ( .A(n2343), .B(n50), .C(intvect[2]), .D(n2247), .E(n817), 
        .F(n1402), .G(ramdatai[5]), .H(n906), .Y(n680) );
  OAI221X1 U2710 ( .A(n705), .B(n1385), .C(n702), .D(n1384), .E(n679), .Y(n681) );
  AOI21X1 U2711 ( .B(n913), .C(temp[5]), .A(n922), .Y(n679) );
  OA21X1 U2712 ( .B(n720), .C(n719), .A(n244), .Y(N12729) );
  AO2222XL U2713 ( .A(n2343), .B(memaddr[6]), .C(intvect[3]), .D(n2247), .E(
        n818), .F(n1402), .G(ramdatai[6]), .H(n906), .Y(n719) );
  OAI221X1 U2714 ( .A(n718), .B(n1385), .C(n2358), .D(n1384), .E(n717), .Y(
        n720) );
  INVX1 U2715 ( .A(pc_i[14]), .Y(n718) );
  OA21X1 U2716 ( .B(n919), .C(n916), .A(n250), .Y(N12730) );
  AO2222XL U2717 ( .A(n2313), .B(n1402), .C(intvect[4]), .D(n2247), .E(
        ramdatai[7]), .F(n906), .G(n2343), .H(pc_o[7]), .Y(n916) );
  OAI221X1 U2718 ( .A(n2373), .B(n1385), .C(n920), .D(n1384), .E(n915), .Y(
        n919) );
  AOI21X1 U2719 ( .B(n913), .C(temp[7]), .A(n907), .Y(n915) );
  OAI22X1 U2720 ( .A(n1236), .B(n2208), .C(n1246), .D(n2400), .Y(n2129) );
  AND4X1 U2721 ( .A(n1247), .B(n1248), .C(n1249), .D(n1250), .Y(n1246) );
  AOI22X1 U2722 ( .A(n166), .B(dph_reg[54]), .C(n105), .D(dph_reg[62]), .Y(
        n1247) );
  AOI22X1 U2723 ( .A(n125), .B(dph_reg[38]), .C(n149), .D(dph_reg[46]), .Y(
        n1248) );
  NOR32XL U2724 ( .B(n240), .C(n106), .A(newinstrlock), .Y(N689) );
  INVX1 U2725 ( .A(ramdatao[7]), .Y(n2195) );
  OAI221X1 U2726 ( .A(n1339), .B(n740), .C(n684), .D(n765), .E(n298), .Y(
        N12491) );
  INVX1 U2727 ( .A(p2[6]), .Y(n740) );
  OAI221X1 U2728 ( .A(n889), .B(n1339), .C(n684), .D(n2283), .E(n298), .Y(
        N12485) );
  OAI221X1 U2729 ( .A(n1339), .B(n598), .C(n684), .D(n2067), .E(n298), .Y(
        N12492) );
  INVX1 U2730 ( .A(p2[7]), .Y(n598) );
  OAI221X1 U2731 ( .A(n872), .B(n1339), .C(n2280), .D(n684), .E(n298), .Y(
        N12486) );
  OAI221X1 U2732 ( .A(n1339), .B(n646), .C(n2277), .D(n684), .E(n298), .Y(
        N12489) );
  INVX1 U2733 ( .A(p2[4]), .Y(n646) );
  OAI221X1 U2734 ( .A(n1339), .B(n632), .C(n2278), .D(n684), .E(n298), .Y(
        N12488) );
  INVX1 U2735 ( .A(p2[3]), .Y(n632) );
  OAI221X1 U2736 ( .A(n1339), .B(n682), .C(n2276), .D(n684), .E(n298), .Y(
        N12490) );
  INVX1 U2737 ( .A(p2[5]), .Y(n682) );
  AND2X1 U2738 ( .A(n1577), .B(n106), .Y(N680) );
  OAI22X1 U2739 ( .A(n935), .B(n2162), .C(n910), .D(n466), .Y(N12725) );
  AOI211X1 U2740 ( .C(n906), .D(ramdatai[2]), .A(n936), .B(n937), .Y(n935) );
  AO2222XL U2741 ( .A(n913), .B(temp[2]), .C(n911), .D(pc_i[10]), .E(n912), 
        .F(temp2_comb[2]), .G(n2343), .H(n2503), .Y(n936) );
  OAI22X1 U2742 ( .A(n938), .B(n909), .C(n2327), .D(n934), .Y(n937) );
  AND2X1 U2743 ( .A(n1577), .B(n262), .Y(N681) );
  OAI21X1 U2744 ( .B(n1015), .C(n2279), .A(n1016), .Y(N12711) );
  OAI31XL U2745 ( .A(n1017), .B(n1018), .C(n1019), .D(n2211), .Y(n1016) );
  NOR4XL U2746 ( .A(n1021), .B(n1022), .C(b[4]), .D(b[3]), .Y(n1019) );
  AOI21X1 U2747 ( .B(n1024), .C(n1025), .A(n2334), .Y(n1018) );
  AND2X1 U2748 ( .A(n1577), .B(phase[3]), .Y(N683) );
  AND2X1 U2749 ( .A(state[2]), .B(n243), .Y(N590) );
  AOI22X1 U2750 ( .A(n104), .B(dph_reg[6]), .C(n165), .D(dph_reg[14]), .Y(
        n1250) );
  AND2X1 U2751 ( .A(state[1]), .B(n243), .Y(N589) );
  AOI22X1 U2752 ( .A(n148), .B(dph_reg[22]), .C(n124), .D(dph_reg[30]), .Y(
        n1249) );
  NOR3XL U2753 ( .A(n2034), .B(instr[4]), .C(n1647), .Y(N10587) );
  ENOX1 U2754 ( .A(n477), .B(n2280), .C(f1), .D(n477), .Y(n1883) );
  ENOX1 U2755 ( .A(n477), .B(n2276), .C(f0), .D(n477), .Y(n1882) );
  NAND2X1 U2756 ( .A(n1100), .B(dps[2]), .Y(n1096) );
  NOR21XL U2757 ( .B(phase[4]), .A(n587), .Y(N684) );
  OAI21X1 U2758 ( .B(n841), .C(n245), .A(n296), .Y(N13324) );
  NOR2X1 U2759 ( .A(n840), .B(finishmul), .Y(n841) );
  AOI22X1 U2760 ( .A(n104), .B(dph_reg[7]), .C(n165), .D(dph_reg[15]), .Y(
        n1241) );
  AND2X1 U2761 ( .A(n242), .B(n1617), .Y(N10562) );
  NAND32X1 U2762 ( .B(n2065), .C(n1616), .A(n1615), .Y(n1617) );
  AOI31X1 U2763 ( .A(n259), .B(n2245), .C(n169), .D(n742), .Y(n2065) );
  AO22AXL U2764 ( .A(n2064), .B(n262), .C(n106), .D(n2119), .Y(n1616) );
  AOI22X1 U2765 ( .A(n148), .B(dph_reg[23]), .C(n124), .D(dph_reg[31]), .Y(
        n1240) );
  AOI22X1 U2766 ( .A(n166), .B(dph_reg[55]), .C(n105), .D(dph_reg[63]), .Y(
        n1238) );
  AOI22X1 U2767 ( .A(n125), .B(dph_reg[39]), .C(n149), .D(dph_reg[47]), .Y(
        n1239) );
  AOI21X1 U2768 ( .B(n2370), .C(n863), .A(n864), .Y(N12976) );
  NAND2X1 U2769 ( .A(waitcnt_0_), .B(waitcnt_1_), .Y(n863) );
  INVX1 U2770 ( .A(stop_r), .Y(n1543) );
  NOR2X1 U2771 ( .A(waitcnt_0_), .B(n864), .Y(N12974) );
  INVX1 U2772 ( .A(idle_r), .Y(n1500) );
  INVX1 U2773 ( .A(temp2_comb[5]), .Y(n702) );
  NAND42X1 U2774 ( .C(n1586), .D(n1585), .A(n1584), .B(n1583), .Y(n1708) );
  AND2X1 U2775 ( .A(n1578), .B(phase[2]), .Y(n1585) );
  AOI21BBXL U2776 ( .B(n1581), .C(n2238), .A(n1580), .Y(n1584) );
  AND2X1 U2777 ( .A(n262), .B(n614), .Y(n1586) );
  INVX1 U2778 ( .A(temp2_comb[4]), .Y(n669) );
  AOI22X1 U2779 ( .A(acc[6]), .B(N13353), .C(N13345), .D(n2273), .Y(n838) );
  NAND43X1 U2780 ( .B(n1737), .C(n592), .D(n2189), .A(n1340), .Y(n684) );
  NOR2X1 U2781 ( .A(ramsfraddr[6]), .B(n842), .Y(n1340) );
  INVX1 U2782 ( .A(n850), .Y(n592) );
  AO21X1 U2783 ( .B(d_hold), .C(n497), .A(cpu_resume_fff), .Y(n1588) );
  INVX1 U2784 ( .A(cpu_hold), .Y(n497) );
  AOI21BBXL U2785 ( .B(N345), .C(n2226), .A(n1887), .Y(n211) );
  AND3X1 U2786 ( .A(n1746), .B(acc[3]), .C(n2194), .Y(n1754) );
  MUX2AXL U2787 ( .D0(n2489), .D1(temp[7]), .S(n1957), .Y(n212) );
  AOI21X1 U2788 ( .B(n913), .C(temp[4]), .A(n927), .Y(n641) );
  OAI22X1 U2789 ( .A(n928), .B(n909), .C(n670), .D(n910), .Y(n927) );
  AOI21X1 U2790 ( .B(n913), .C(temp[6]), .A(n917), .Y(n717) );
  OAI22X1 U2791 ( .A(n918), .B(n909), .C(n734), .D(n910), .Y(n917) );
  OAI21BBX1 U2792 ( .A(n2247), .B(n2503), .C(n213), .Y(n1464) );
  AOI222XL U2793 ( .A(n411), .B(n235), .C(n2240), .D(pc_i[10]), .E(n2239), .F(
        pc_i[2]), .Y(n213) );
  AND2X1 U2794 ( .A(n106), .B(n611), .Y(n1580) );
  INVX1 U2795 ( .A(temp2_comb[7]), .Y(n920) );
  AOI221X1 U2796 ( .A(n1167), .B(n110), .C(pc_i[4]), .D(n1127), .E(n1176), .Y(
        n1107) );
  AO222X1 U2797 ( .A(n42), .B(n1177), .C(n2502), .D(n1178), .E(n36), .F(n1169), 
        .Y(n1176) );
  OAI221X1 U2798 ( .A(n2465), .B(n1134), .C(n1179), .D(n1132), .E(n1180), .Y(
        n1178) );
  AOI221X1 U2799 ( .A(n1153), .B(n42), .C(pc_i[6]), .D(n1127), .E(n1154), .Y(
        n1106) );
  AO222X1 U2800 ( .A(n1133), .B(n2302), .C(pc_o[6]), .D(n1155), .E(n1131), .F(
        n36), .Y(n1154) );
  OAI221X1 U2801 ( .A(n49), .B(n1134), .C(n1156), .D(n37), .E(n1157), .Y(n1155) );
  AOI221X1 U2802 ( .A(n48), .B(n1291), .C(pc_i[9]), .D(n1127), .E(n2300), .Y(
        n1226) );
  INVX1 U2803 ( .A(n1297), .Y(n2300) );
  AOI221XL U2804 ( .A(n1289), .B(n2302), .C(memaddr[9]), .D(n1298), .E(n1299), 
        .Y(n1297) );
  NOR4XL U2805 ( .A(pc_o[9]), .B(n53), .C(n2305), .D(n1290), .Y(n1299) );
  AOI221X1 U2806 ( .A(n36), .B(n1256), .C(pc_i[11]), .D(n1127), .E(n2298), .Y(
        n1225) );
  INVX1 U2807 ( .A(n1275), .Y(n2298) );
  AOI221XL U2808 ( .A(n1268), .B(n2302), .C(pc_o[11]), .D(n1276), .E(n1277), 
        .Y(n1275) );
  NOR4XL U2809 ( .A(pc_o[11]), .B(n2467), .C(n2305), .D(n1269), .Y(n1277) );
  OAI31XL U2810 ( .A(n1026), .B(n1027), .C(n1028), .D(n1029), .Y(n1017) );
  OAI31XL U2811 ( .A(n1030), .B(n1031), .C(n1032), .D(ov), .Y(n1029) );
  XNOR2XL U2812 ( .A(n1035), .B(n1036), .Y(n1028) );
  NAND32X1 U2813 ( .B(n1033), .C(n1027), .A(n1034), .Y(n1030) );
  OAI211X1 U2814 ( .C(pc_o[8]), .D(n2305), .A(n1300), .B(n1301), .Y(n1298) );
  AOI22X1 U2815 ( .A(n2302), .B(n1302), .C(n48), .D(pc_o[8]), .Y(n1301) );
  INVX1 U2816 ( .A(p2[2]), .Y(n1411) );
  NOR2X1 U2817 ( .A(n131), .B(n2471), .Y(N14341) );
  NOR2X1 U2818 ( .A(n131), .B(n2470), .Y(N14342) );
  NOR2X1 U2819 ( .A(n2478), .B(n2486), .Y(N14338) );
  NOR2X1 U2820 ( .A(n2478), .B(n2485), .Y(N14339) );
  NOR2X1 U2821 ( .A(n2478), .B(n2474), .Y(N14340) );
  NOR2X1 U2822 ( .A(n131), .B(n2445), .Y(N14343) );
  OA222X1 U2823 ( .A(n1229), .B(n34), .C(pc_o[15]), .D(n1230), .E(n2373), .F(
        n2304), .Y(n1223) );
  INVX1 U2824 ( .A(n1127), .Y(n2304) );
  AOI32X1 U2825 ( .A(n43), .B(pc_o[14]), .C(n1231), .D(n1232), .E(n2464), .Y(
        n1230) );
  AOI211X1 U2826 ( .C(n42), .D(n2464), .A(n1233), .B(n1234), .Y(n1229) );
  AOI221X1 U2827 ( .A(n1125), .B(n43), .C(pc_i[7]), .D(n1127), .E(n1128), .Y(
        n1104) );
  AO222X1 U2828 ( .A(n2461), .B(n48), .C(pc_o[7]), .D(n1129), .E(n1130), .F(
        n2302), .Y(n1128) );
  INVX1 U2829 ( .A(n1135), .Y(n2461) );
  OAI221X1 U2830 ( .A(n1131), .B(n37), .C(n1133), .D(n1134), .E(n2303), .Y(
        n1129) );
  AOI222XL U2831 ( .A(n1233), .B(pc_o[14]), .C(n2464), .D(n1242), .E(pc_i[14]), 
        .F(n1127), .Y(n1224) );
  AO21X1 U2832 ( .B(n1231), .C(n42), .A(n1232), .Y(n1242) );
  INVX1 U2833 ( .A(n1186), .Y(n2294) );
  OAI211X1 U2834 ( .C(n205), .D(n2305), .A(n1188), .B(n1189), .Y(n1186) );
  AOI22X1 U2835 ( .A(n48), .B(n1179), .C(n86), .D(pc_i[3]), .Y(n1189) );
  AOI32X1 U2836 ( .A(n2456), .B(n2465), .C(n2302), .D(pc_o[3]), .E(n1190), .Y(
        n1188) );
  INVX1 U2837 ( .A(n1251), .Y(n2295) );
  OAI211X1 U2838 ( .C(n1252), .D(n46), .A(n1253), .B(n1254), .Y(n1251) );
  NAND4X1 U2839 ( .A(n1257), .B(n43), .C(pc_o[12]), .D(n46), .Y(n1253) );
  AOI21X1 U2840 ( .B(n86), .C(pc_i[13]), .A(n1232), .Y(n1254) );
  OAI32X1 U2841 ( .A(n1255), .B(pc_o[13]), .C(n1134), .D(n1132), .E(n1244), 
        .Y(n1232) );
  MUX2BXL U2842 ( .D0(acc[6]), .D1(n2319), .S(n1957), .Y(n214) );
  INVX1 U2843 ( .A(n1265), .Y(n2297) );
  AO2222XL U2844 ( .A(n86), .B(pc_i[12]), .C(n2455), .D(n110), .E(pc_o[12]), 
        .F(n1266), .G(n1267), .H(n40), .Y(n1265) );
  OAI22X1 U2845 ( .A(n2305), .B(n2452), .C(n37), .D(n2454), .Y(n1267) );
  OAI21X1 U2846 ( .B(n1268), .C(n153), .A(n1259), .Y(n1266) );
  INVX1 U2847 ( .A(n1163), .Y(n2293) );
  OAI2B11X1 U2848 ( .D(n1164), .C(n2305), .A(n1165), .B(n1166), .Y(n1163) );
  AOI22X1 U2849 ( .A(n36), .B(n1156), .C(n1127), .D(pc_i[5]), .Y(n1166) );
  AOI32X1 U2850 ( .A(n1167), .B(n49), .C(n2302), .D(n50), .E(n1168), .Y(n1165)
         );
  AOI221X1 U2851 ( .A(n2463), .B(n42), .C(pc_i[2]), .D(n1127), .E(n2292), .Y(
        n1108) );
  INVX1 U2852 ( .A(n1199), .Y(n2463) );
  INVX1 U2853 ( .A(n1198), .Y(n2292) );
  AOI221XL U2854 ( .A(n1199), .B(n36), .C(n2503), .D(n1200), .E(n1201), .Y(
        n1198) );
  NAND21X1 U2855 ( .B(n1572), .A(state[0]), .Y(n483) );
  AOI222XL U2856 ( .A(n1200), .B(memaddr[1]), .C(n2466), .D(n1208), .E(pc_i[1]), .F(n1127), .Y(n1109) );
  OAI21X1 U2857 ( .B(n1134), .C(pc_o[0]), .A(n1209), .Y(n1208) );
  NOR3XL U2858 ( .A(n2502), .B(pc_o[3]), .C(n1192), .Y(n1167) );
  INVX1 U2859 ( .A(n1308), .Y(n2301) );
  AO2222XL U2860 ( .A(n86), .B(pc_i[8]), .C(n2457), .D(n110), .E(memaddr[8]), 
        .F(n1309), .G(n1310), .H(n53), .Y(n1308) );
  INVX1 U2861 ( .A(n1302), .Y(n2457) );
  OAI22X1 U2862 ( .A(n2305), .B(n1290), .C(n1132), .D(n1135), .Y(n1310) );
  INVX1 U2863 ( .A(b[2]), .Y(n2486) );
  INVX1 U2864 ( .A(b[3]), .Y(n2485) );
  NOR3XL U2865 ( .A(n50), .B(pc_o[6]), .C(n2459), .Y(n1133) );
  NOR2X1 U2866 ( .A(pc_o[1]), .B(memaddr[2]), .Y(n1191) );
  NOR2X1 U2867 ( .A(n1302), .B(pc_o[9]), .Y(n1289) );
  NOR2X1 U2868 ( .A(n1280), .B(pc_o[11]), .Y(n1268) );
  NAND3X1 U2869 ( .A(n50), .B(n1430), .C(n2502), .Y(n1311) );
  NAND2X1 U2870 ( .A(pc_o[1]), .B(n2503), .Y(n1202) );
  NAND32X1 U2871 ( .B(n1290), .C(n53), .A(memaddr[9]), .Y(n1269) );
  NAND32X1 U2872 ( .B(n1311), .C(n2468), .A(pc_o[6]), .Y(n1290) );
  INVX1 U2873 ( .A(memaddr[3]), .Y(n2465) );
  INVX1 U2874 ( .A(memaddr[0]), .Y(n2460) );
  XNOR2XL U2875 ( .A(n1311), .B(memaddr[6]), .Y(n1153) );
  NOR3XL U2876 ( .A(n235), .B(pc_o[11]), .C(n2462), .Y(n1256) );
  NOR3XL U2877 ( .A(memaddr[8]), .B(pc_o[9]), .C(n1135), .Y(n1291) );
  INVX1 U2878 ( .A(b[4]), .Y(n2474) );
  XNOR2XL U2879 ( .A(n1487), .B(pc_o[5]), .Y(n1164) );
  NAND2X1 U2880 ( .A(memaddr[4]), .B(n1430), .Y(n1487) );
  INVX1 U2881 ( .A(memaddr[7]), .Y(n2468) );
  XOR2X1 U2882 ( .A(n2466), .B(memaddr[2]), .Y(n1199) );
  OAI211X1 U2883 ( .C(n1007), .D(n170), .A(n633), .B(n1008), .Y(n984) );
  AOI22X1 U2884 ( .A(n262), .B(n1009), .C(n957), .D(phase[2]), .Y(n1008) );
  NOR32XL U2885 ( .B(n756), .C(n2244), .A(n777), .Y(n1007) );
  NAND2X1 U2886 ( .A(n444), .B(n1000), .Y(n980) );
  NAND4X1 U2887 ( .A(n2349), .B(n262), .C(n1001), .D(n2187), .Y(n1000) );
  INVX1 U2888 ( .A(b[5]), .Y(n2471) );
  INVX1 U2889 ( .A(b[6]), .Y(n2470) );
  AOI22X1 U2890 ( .A(n912), .B(temp2_comb[1]), .C(n911), .D(pc_i[9]), .Y(n946)
         );
  AOI22X1 U2891 ( .A(n912), .B(temp2_comb[0]), .C(n911), .D(pc_i[8]), .Y(n955)
         );
  AOI21X1 U2892 ( .B(n106), .C(n2421), .A(n2237), .Y(n953) );
  INVX1 U2893 ( .A(memaddr[11]), .Y(n2453) );
  OAI31XL U2894 ( .A(n959), .B(n960), .C(n961), .D(n106), .Y(n934) );
  OAI22X1 U2895 ( .A(n2428), .B(n2433), .C(n962), .D(n2435), .Y(n961) );
  OAI211X1 U2896 ( .C(n966), .D(n32), .A(n967), .B(n968), .Y(n959) );
  OAI31XL U2897 ( .A(n2450), .B(n128), .C(n805), .D(n964), .Y(n960) );
  AOI22X1 U2898 ( .A(n262), .B(n956), .C(phase[2]), .D(n957), .Y(n954) );
  INVX1 U2899 ( .A(b[7]), .Y(n2445) );
  OAI21BBX1 U2900 ( .A(n2436), .B(n972), .C(instr[3]), .Y(n967) );
  NAND4X1 U2901 ( .A(n965), .B(instr[5]), .C(n61), .D(n69), .Y(n964) );
  INVX1 U2902 ( .A(memaddr[14]), .Y(n2464) );
  NOR2X1 U2903 ( .A(n2482), .B(dec_accop[10]), .Y(n1027) );
  OAI22AX1 U2904 ( .D(ckcon[1]), .C(n869), .A(n2199), .B(n870), .Y(N12966) );
  OAI22AX1 U2905 ( .D(ckcon[5]), .C(n869), .A(n2212), .B(n870), .Y(N12970) );
  OAI22AX1 U2906 ( .D(ckcon[4]), .C(n869), .A(n2216), .B(n870), .Y(N12969) );
  OAI22AX1 U2907 ( .D(ckcon[0]), .C(n869), .A(n2203), .B(n870), .Y(N12965) );
  OAI22AX1 U2908 ( .D(ckcon[7]), .C(n869), .A(n2195), .B(n870), .Y(N12972) );
  OAI22AX1 U2909 ( .D(ckcon[3]), .C(n869), .A(n12), .B(n870), .Y(N12968) );
  AND2X1 U2910 ( .A(cpu_resume_ff1), .B(n288), .Y(N13380) );
  INVX1 U2911 ( .A(finishdiv), .Y(n2259) );
  INVX1 U2912 ( .A(finishmul), .Y(n2258) );
  NAND21X1 U2913 ( .B(n2367), .A(dec_accop[17]), .Y(n2157) );
  INVX1 U2914 ( .A(stop), .Y(n1541) );
  NAND3X1 U2915 ( .A(n2443), .B(n2442), .C(ramsfraddr[2]), .Y(n845) );
  NAND3X1 U2916 ( .A(ramsfraddr[2]), .B(n2442), .C(ramsfraddr[0]), .Y(n846) );
  BUFX3 U2917 ( .A(memaddr[10]), .Y(pc_o[10]) );
  BUFX3 U2918 ( .A(n50), .Y(pc_o[5]) );
  BUFX3 U2919 ( .A(n2502), .Y(pc_o[4]) );
  BUFX3 U2920 ( .A(n2503), .Y(pc_o[2]) );
  BUFX3 U2921 ( .A(memaddr[0]), .Y(pc_o[0]) );
  AO2222XL U2922 ( .A(n188), .B(ramdatao[6]), .C(n931), .D(n930), .E(p2[6]), 
        .F(n195), .G(n929), .H(pc_o[14]), .Y(n1732) );
  AO2222XL U2923 ( .A(n188), .B(ramdatao[7]), .C(n741), .D(n930), .E(p2[7]), 
        .F(n195), .G(n929), .H(pc_o[15]), .Y(n1733) );
  AO2222XL U2924 ( .A(n188), .B(ramdatao[5]), .C(n683), .D(n930), .E(p2[5]), 
        .F(n195), .G(n929), .H(pc_o[13]), .Y(n1731) );
  AO2222XL U2925 ( .A(n188), .B(ramdatao[4]), .C(n647), .D(n930), .E(p2[4]), 
        .F(n195), .G(n929), .H(pc_o[12]), .Y(n1730) );
  AO2222XL U2926 ( .A(n188), .B(ramdatao[3]), .C(n637), .D(n930), .E(p2[3]), 
        .F(n195), .G(n929), .H(pc_o[11]), .Y(n1729) );
  OAI22XL U2927 ( .A(n434), .B(n1538), .C(n507), .D(n1535), .Y(n510) );
  NAND32XL U2928 ( .B(n260), .C(n2223), .A(n657), .Y(n722) );
  NAND32X2 U2929 ( .B(N345), .C(n260), .A(n657), .Y(n361) );
  NAND32X2 U2930 ( .B(n360), .C(n367), .A(n359), .Y(n657) );
  AOI22XL U2931 ( .A(n2206), .B(n814), .C(sfrdatai[2]), .D(n2219), .Y(n1558)
         );
  INVX1 U2932 ( .A(n1743), .Y(n1767) );
  NOR2X1 U2933 ( .A(n1492), .B(n1491), .Y(n1493) );
  XNOR2XL U2934 ( .A(n1492), .B(n2202), .Y(n1522) );
  OAI22XL U2935 ( .A(n674), .B(n1503), .C(n989), .D(n294), .Y(N12718) );
  OAI21BBX1 U2936 ( .A(n1523), .B(n1524), .C(n1525), .Y(n1491) );
  XNOR2XL U2937 ( .A(n1524), .B(n1435), .Y(n1536) );
  OAI211XL U2938 ( .C(n2438), .D(n1434), .A(n1548), .B(n1549), .Y(n891) );
  OAI22XL U2939 ( .A(n292), .B(n640), .C(n639), .D(n1503), .Y(N12717) );
  XOR2XL U2940 ( .A(n1491), .B(n1522), .Y(n1521) );
  XOR2XL U2941 ( .A(n1523), .B(n1536), .Y(n1885) );
  XNOR2XL U2942 ( .A(n891), .B(n892), .Y(n890) );
  OAI22X1 U2943 ( .A(n354), .B(n787), .C(n2495), .D(n353), .Y(n363) );
  XOR3X1 U2944 ( .A(n2202), .B(n180), .C(n1), .Y(n485) );
  INVXL U2945 ( .A(n656), .Y(n661) );
  AOI222XL U2946 ( .A(n2200), .B(ramdatai[3]), .C(n2201), .D(sfrdatai[3]), .E(
        n2250), .F(n2194), .Y(n1524) );
  AOI22XL U2947 ( .A(n2206), .B(n815), .C(sfrdatai[3]), .D(n2219), .Y(n1548)
         );
  OAI211XL U2948 ( .C(n1738), .D(n674), .A(n673), .B(n671), .Y(n675) );
  AOI222XL U2949 ( .A(n2201), .B(sfrdatai[7]), .C(ramdatai[7]), .D(n2200), .E(
        n2197), .F(n2250), .Y(n1417) );
  OAI22XL U2950 ( .A(n292), .B(n1433), .C(n1462), .D(n1503), .Y(N12716) );
  OAI222XL U2951 ( .A(n1462), .B(n1932), .C(n2493), .D(n1934), .E(n938), .F(
        n1931), .Y(n1740) );
  AOI211XL U2952 ( .C(n1858), .D(n2038), .A(n1857), .B(n1856), .Y(n1877) );
  NAND32X1 U2953 ( .B(n491), .C(n490), .A(n489), .Y(n495) );
  AOI211X1 U2954 ( .C(n1858), .D(n484), .A(n482), .B(n481), .Y(n486) );
  OA21XL U2955 ( .B(n1436), .C(n695), .A(n694), .Y(n696) );
  AOI222XL U2956 ( .A(n2200), .B(ramdatai[4]), .C(n2201), .D(sfrdatai[4]), .E(
        n2250), .F(n2215), .Y(n1492) );
  MUX2XL U2957 ( .D0(ramdatao[0]), .D1(n1656), .S(waitstaten), .Y(
        ramdatao_comb[0]) );
  OA21XL U2958 ( .B(n1436), .C(n656), .A(n694), .Y(n658) );
  AO21XL U2959 ( .B(n1576), .C(n1575), .A(n1574), .Y(n1878) );
  GEN2XL U2960 ( .D(n1563), .E(n1575), .C(n1545), .B(n1562), .A(codefetch_s), 
        .Y(n1547) );
  NAND21XL U2961 ( .B(pdmode), .A(n1575), .Y(n1544) );
  AOI32XL U2962 ( .A(n1590), .B(codefetch_s), .C(n1543), .D(n1588), .E(n615), 
        .Y(n498) );
  INVX2 U2963 ( .A(n615), .Y(n616) );
  NAND42X1 U2964 ( .C(n381), .D(n380), .A(n379), .B(n378), .Y(n382) );
  AND2X1 U2965 ( .A(n1858), .B(n362), .Y(n380) );
  AO2222X1 U2966 ( .A(n1743), .B(n2038), .C(n463), .D(n484), .E(n1437), .F(
        n1440), .G(n363), .H(n362), .Y(n356) );
  AO2222X1 U2967 ( .A(n695), .B(n484), .C(n656), .D(n362), .E(n723), .F(n1440), 
        .G(n1988), .H(n2038), .Y(n355) );
  NOR21X4 U2968 ( .B(pc_i[8]), .A(n1531), .Y(n417) );
  NOR32X4 U2969 ( .B(n414), .C(n413), .A(n412), .Y(n415) );
  MUX2IX4 U2970 ( .D0(n433), .D1(n829), .S(n1659), .Y(n434) );
  GEN2X1 U2971 ( .D(n474), .E(n2228), .C(n1994), .B(n202), .A(n472), .Y(n482)
         );
endmodule


module mcu51_cpu_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  NOR21XL U2 ( .B(A[0]), .A(n2), .Y(carry[1]) );
  INVX1 U3 ( .A(B[0]), .Y(n2) );
endmodule


module mcu51_cpu_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  NOR21XL U1 ( .B(A[0]), .A(n2), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
endmodule


module mcu51_cpu_a0_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
endmodule


module mcu51_cpu_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n13), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n15), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  INVX1 U1 ( .A(B[2]), .Y(n14) );
  INVX1 U2 ( .A(B[3]), .Y(n13) );
  INVX1 U3 ( .A(B[4]), .Y(n12) );
  INVX1 U4 ( .A(B[5]), .Y(n11) );
  INVX1 U5 ( .A(B[1]), .Y(n15) );
  NAND21X1 U6 ( .B(n17), .A(n16), .Y(carry[1]) );
  INVX1 U7 ( .A(A[0]), .Y(n16) );
  INVX1 U8 ( .A(B[6]), .Y(n10) );
  AOI21X1 U9 ( .B(carry[7]), .C(A[7]), .A(n9), .Y(DIFF[8]) );
  AOI21BBXL U10 ( .B(A[7]), .C(carry[7]), .A(B[7]), .Y(n9) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U12 ( .A(B[0]), .Y(n17) );
endmodule


module mcu51_cpu_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [8:1] carry;

  FAD1X1 U2_7 ( .A(A[7]), .B(n11), .CI(carry[7]), .CO(carry[8]), .SO(DIFF[7])
         );
  FAD1X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n13), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n14), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n16), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n17), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  INVX1 U1 ( .A(carry[8]), .Y(DIFF[8]) );
  INVX1 U2 ( .A(B[7]), .Y(n11) );
  INVX1 U3 ( .A(B[2]), .Y(n16) );
  INVX1 U4 ( .A(B[3]), .Y(n15) );
  INVX1 U5 ( .A(B[4]), .Y(n14) );
  INVX1 U6 ( .A(B[5]), .Y(n13) );
  INVX1 U7 ( .A(B[6]), .Y(n12) );
  INVX1 U8 ( .A(B[1]), .Y(n17) );
  NAND21X1 U9 ( .B(n18), .A(n10), .Y(carry[1]) );
  INVX1 U10 ( .A(A[0]), .Y(n10) );
  INVX1 U11 ( .A(B[0]), .Y(n18) );
  XOR2X1 U12 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module mcu51_cpu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [15:1] carry;

  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  INVX1 U1 ( .A(B[0]), .Y(n2) );
  NOR21XL U2 ( .B(A[0]), .A(n2), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mpb_a0 ( i_rd, i_wr, wdat0, wdat1, addr0, addr1, r_i2c_attr, esfrm_oe, 
        esfrm_we, sfrack, esfrm_wdat, esfrm_adr, mcu_esfr_rdat, delay_rdat, 
        delay_rrdy, esfrm_rrdy, esfrm_rdat, channel_sel, r_pg0_sel, dma_w, 
        dma_r, dma_addr, dma_wdat, dma_ack, memaddr, memaddr_c, memwr, memrd, 
        memrd_c, cpurst, memdatao, memack, hit_xd, hit_xr, hit_ps, hit_ps_c, 
        idat_r, idat_w, idat_adr, idat_wdat, iram_ce, xram_ce, regx_re, 
        iram_we, xram_we, regx_we, iram_a, xram_a, iram_d, xram_d, iram_rdat, 
        xram_rdat, regx_rdat, bist_en, bist_wr, bist_adr, bist_wdat, bist_xram, 
        mclk, srstz, test_si, test_so, test_se );
  input [1:0] i_rd;
  input [1:0] i_wr;
  input [7:0] wdat0;
  input [7:0] wdat1;
  input [7:0] addr0;
  input [7:0] addr1;
  output [7:0] esfrm_wdat;
  output [6:0] esfrm_adr;
  input [7:0] mcu_esfr_rdat;
  input [7:0] delay_rdat;
  output [7:0] esfrm_rdat;
  input [3:0] r_pg0_sel;
  input [10:0] dma_addr;
  input [7:0] dma_wdat;
  input [15:0] memaddr;
  input [15:0] memaddr_c;
  input [7:0] memdatao;
  input [7:0] idat_adr;
  input [7:0] idat_wdat;
  output [10:0] iram_a;
  output [10:0] xram_a;
  output [7:0] iram_d;
  output [7:0] xram_d;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  input [7:0] regx_rdat;
  input [10:0] bist_adr;
  input [7:0] bist_wdat;
  input r_i2c_attr, delay_rrdy, channel_sel, dma_w, dma_r, memwr, memrd,
         memrd_c, cpurst, idat_r, idat_w, bist_en, bist_wr, bist_xram, mclk,
         srstz, test_si, test_se;
  output esfrm_oe, esfrm_we, sfrack, esfrm_rrdy, dma_ack, memack, hit_xd,
         hit_xr, hit_ps, hit_ps_c, iram_ce, xram_ce, regx_re, iram_we, xram_we,
         regx_we, test_so;
  wire   n238, pg0_rdwait, pg0_wrwait, N44, N45, r_pg0_rdrdy, N46,
         xram_rdsel_0_, n55, n91, n110, n112, n114, n128, n129, n130, n132,
         n133, n134, n136, n137, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n30, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n111, n113, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n131, n135, n138, n139, n140, n141, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237;

  SDFFRQX1 r_pg0_rdrdy_reg ( .D(N46), .SIN(pg0_wrwait), .SMC(test_se), .C(mclk), .XR(srstz), .Q(r_pg0_rdrdy) );
  SDFFRQX1 xram_rdsel_reg_1_ ( .D(n229), .SIN(xram_rdsel_0_), .SMC(test_se), 
        .C(mclk), .XR(srstz), .Q(test_so) );
  SDFFRQX1 xram_rdsel_reg_0_ ( .D(n230), .SIN(n5), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(xram_rdsel_0_) );
  SDFFRQX1 pg0_rdwait_reg ( .D(N45), .SIN(test_si), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(pg0_rdwait) );
  SDFFRQX1 pg0_wrwait_reg ( .D(N44), .SIN(pg0_rdwait), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(pg0_wrwait) );
  BUFX1 U3 ( .A(n53), .Y(n1) );
  AND2XL U4 ( .A(n228), .B(n227), .Y(sfrack) );
  NAND21X1 U5 ( .B(i_wr[1]), .A(n39), .Y(n38) );
  BUFX3 U6 ( .A(n238), .Y(xram_a[0]) );
  INVX1 U7 ( .A(n222), .Y(n223) );
  MUX2IX2 U8 ( .D0(addr0[7]), .D1(addr1[7]), .S(n38), .Y(n222) );
  NOR2X1 U9 ( .A(n33), .B(cpurst), .Y(memack) );
  OAI31XL U10 ( .A(r_i2c_attr), .B(n42), .C(n223), .D(n41), .Y(n53) );
  NAND21X1 U11 ( .B(n156), .A(dma_addr[6]), .Y(n111) );
  AND3X1 U12 ( .A(n13), .B(n14), .C(n15), .Y(n102) );
  AND3X1 U13 ( .A(n22), .B(n23), .C(n24), .Y(n100) );
  OAI2B11X1 U14 ( .D(dma_addr[3]), .C(n156), .A(n163), .B(n104), .Y(xram_a[3])
         );
  AND3X1 U15 ( .A(n19), .B(n20), .C(n21), .Y(n104) );
  AND3X1 U16 ( .A(n25), .B(n26), .C(n27), .Y(n105) );
  OA33X1 U17 ( .A(n194), .B(n192), .C(n185), .D(bist_en), .E(n184), .F(n183), 
        .Y(n3) );
  INVX1 U18 ( .A(n192), .Y(n4) );
  BUFX3 U19 ( .A(r_pg0_rdrdy), .Y(n5) );
  INVX1 U20 ( .A(n181), .Y(n6) );
  INVX1 U21 ( .A(n193), .Y(n7) );
  BUFX3 U22 ( .A(bist_en), .Y(n8) );
  NAND2X1 U23 ( .A(r_pg0_sel[2]), .B(n40), .Y(n35) );
  INVX1 U24 ( .A(n35), .Y(n9) );
  INVX1 U25 ( .A(n35), .Y(n10) );
  BUFX3 U26 ( .A(bist_en), .Y(n196) );
  INVX1 U27 ( .A(n196), .Y(n11) );
  INVX1 U28 ( .A(n196), .Y(n12) );
  NAND21XL U29 ( .B(n222), .A(n221), .Y(n227) );
  NAND2X1 U30 ( .A(memaddr_c[5]), .B(n127), .Y(n18) );
  NAND2X2 U31 ( .A(memaddr_c[1]), .B(n127), .Y(n15) );
  NAND2X1 U32 ( .A(memaddr[1]), .B(n120), .Y(n13) );
  NAND2X1 U33 ( .A(n131), .B(esfrm_adr[1]), .Y(n14) );
  OAI2B11X1 U34 ( .D(dma_addr[1]), .C(n156), .A(n159), .B(n102), .Y(xram_a[1])
         );
  INVX1 U35 ( .A(n141), .Y(n127) );
  NAND2X1 U36 ( .A(memaddr[5]), .B(n120), .Y(n16) );
  NAND2X1 U37 ( .A(n131), .B(esfrm_adr[5]), .Y(n17) );
  AND3X1 U38 ( .A(n16), .B(n17), .C(n18), .Y(n106) );
  NAND2X1 U39 ( .A(memaddr[3]), .B(n120), .Y(n19) );
  NAND2X1 U40 ( .A(n131), .B(esfrm_adr[3]), .Y(n20) );
  NAND2X1 U41 ( .A(memaddr_c[3]), .B(n127), .Y(n21) );
  NAND2X1 U42 ( .A(dma_addr[0]), .B(n121), .Y(n22) );
  NAND2X1 U43 ( .A(memaddr_c[0]), .B(n127), .Y(n23) );
  NAND2X1 U44 ( .A(memaddr[0]), .B(n120), .Y(n24) );
  OAI211X1 U45 ( .C(n101), .D(n152), .A(n157), .B(n100), .Y(n238) );
  NAND2X1 U46 ( .A(memaddr[4]), .B(n120), .Y(n25) );
  NAND2XL U47 ( .A(n131), .B(esfrm_adr[4]), .Y(n26) );
  NAND2X1 U48 ( .A(memaddr_c[4]), .B(n127), .Y(n27) );
  INVXL U49 ( .A(n168), .Y(esfrm_adr[4]) );
  OAI2B11X1 U50 ( .D(dma_addr[4]), .C(n156), .A(n166), .B(n105), .Y(xram_a[4])
         );
  MUX2IX2 U51 ( .D0(addr1[6]), .D1(addr0[6]), .S(n107), .Y(n174) );
  INVXL U52 ( .A(n38), .Y(n107) );
  INVXL U53 ( .A(i_rd[1]), .Y(n39) );
  INVXL U54 ( .A(n171), .Y(esfrm_adr[5]) );
  INVXL U55 ( .A(n101), .Y(esfrm_adr[0]) );
  OR2X2 U56 ( .A(n1), .B(n202), .Y(n182) );
  OAI21BXL U57 ( .C(n218), .B(n110), .A(n200), .Y(regx_we) );
  INVX1 U58 ( .A(addr0[2]), .Y(n30) );
  AO21XL U59 ( .B(n222), .C(n221), .A(pg0_rdwait), .Y(n202) );
  AO22XL U60 ( .A(idat_adr[2]), .B(n198), .C(n179), .D(esfrm_adr[2]), .Y(n162)
         );
  INVX1 U61 ( .A(n189), .Y(n97) );
  INVX1 U62 ( .A(n152), .Y(n131) );
  INVX1 U63 ( .A(n192), .Y(n179) );
  INVX1 U64 ( .A(n181), .Y(n198) );
  INVX1 U65 ( .A(n156), .Y(n121) );
  INVX1 U66 ( .A(n227), .Y(esfrm_oe) );
  INVX1 U67 ( .A(n154), .Y(n120) );
  INVX1 U68 ( .A(n96), .Y(n99) );
  INVX1 U69 ( .A(n57), .Y(n72) );
  NAND32X1 U70 ( .B(bist_en), .C(n99), .A(n56), .Y(n57) );
  NOR2X1 U71 ( .A(memaddr_c[10]), .B(n204), .Y(n28) );
  AND3X1 U72 ( .A(n215), .B(n214), .C(n213), .Y(n207) );
  NAND21X1 U73 ( .B(bist_en), .A(n189), .Y(n98) );
  NAND21X1 U74 ( .B(bist_en), .A(n97), .Y(n152) );
  OR2X1 U75 ( .A(bist_en), .B(n56), .Y(n75) );
  NAND21X1 U76 ( .B(bist_en), .A(n78), .Y(n192) );
  INVX1 U77 ( .A(n77), .Y(n78) );
  INVX1 U78 ( .A(n193), .Y(n231) );
  NAND21X1 U79 ( .B(bist_en), .A(n77), .Y(n181) );
  NAND21X1 U80 ( .B(n11), .A(bist_wdat[0]), .Y(n79) );
  NAND21X1 U81 ( .B(n11), .A(bist_wdat[1]), .Y(n81) );
  NAND21X1 U82 ( .B(n11), .A(bist_wdat[4]), .Y(n87) );
  NAND21X1 U83 ( .B(n12), .A(bist_wdat[2]), .Y(n83) );
  NAND21X1 U84 ( .B(n12), .A(bist_wdat[3]), .Y(n85) );
  NAND21X1 U85 ( .B(n12), .A(bist_wdat[6]), .Y(n92) );
  NAND21X1 U86 ( .B(n232), .A(n193), .Y(n43) );
  NAND32X1 U87 ( .B(n97), .C(n96), .A(n12), .Y(n156) );
  INVX1 U88 ( .A(n54), .Y(n73) );
  NAND32X1 U89 ( .B(n8), .C(n96), .A(n56), .Y(n54) );
  NAND31X1 U90 ( .C(n8), .A(n203), .B(n219), .Y(n211) );
  INVX1 U91 ( .A(n236), .Y(n117) );
  INVX1 U92 ( .A(n165), .Y(esfrm_adr[3]) );
  AOI21BBXL U93 ( .B(n174), .C(n152), .A(n108), .Y(n109) );
  AND2X1 U94 ( .A(memaddr_c[6]), .B(n127), .Y(n108) );
  INVX1 U95 ( .A(n184), .Y(n218) );
  INVX1 U96 ( .A(n228), .Y(esfrm_we) );
  OR2X1 U97 ( .A(idat_r), .B(idat_w), .Y(n77) );
  OR3XL U98 ( .A(n99), .B(n37), .C(n98), .Y(n154) );
  AO21X1 U99 ( .B(n205), .C(n190), .A(n230), .Y(n96) );
  NAND32X1 U100 ( .B(n99), .C(n98), .A(n37), .Y(n141) );
  NAND21X1 U101 ( .B(memaddr_c[9]), .A(n124), .Y(n204) );
  OAI221XL U102 ( .A(n168), .B(n192), .C(n181), .D(n167), .E(n166), .Y(
        iram_a[4]) );
  INVX1 U103 ( .A(idat_adr[4]), .Y(n167) );
  INVX1 U104 ( .A(memaddr_c[8]), .Y(n124) );
  INVX1 U105 ( .A(memaddr_c[13]), .Y(n213) );
  INVX1 U106 ( .A(memaddr_c[11]), .Y(n215) );
  INVX1 U107 ( .A(memaddr_c[12]), .Y(n214) );
  NAND5XL U108 ( .A(n28), .B(n216), .C(n215), .D(n214), .E(n213), .Y(n217) );
  INVX1 U109 ( .A(memaddr_c[7]), .Y(n216) );
  AOI211X1 U110 ( .C(memaddr_c[10]), .D(n204), .A(memaddr_c[14]), .B(
        memaddr_c[15]), .Y(n206) );
  INVX1 U111 ( .A(idat_adr[6]), .Y(n173) );
  OAI221XL U112 ( .A(n165), .B(n192), .C(n181), .D(n164), .E(n163), .Y(
        iram_a[3]) );
  INVX1 U113 ( .A(idat_adr[3]), .Y(n164) );
  OAI221XL U114 ( .A(n171), .B(n192), .C(n181), .D(n170), .E(n169), .Y(
        iram_a[5]) );
  INVX1 U115 ( .A(idat_adr[5]), .Y(n170) );
  OA222X1 U116 ( .A(n154), .B(n236), .C(n153), .D(n152), .E(n151), .F(n141), 
        .Y(n155) );
  INVX1 U117 ( .A(memaddr_c[10]), .Y(n151) );
  INVX1 U118 ( .A(memaddr[10]), .Y(n236) );
  NAND4X1 U119 ( .A(memaddr_c[14]), .B(memaddr_c[13]), .C(memaddr_c[15]), .D(
        n114), .Y(n112) );
  AND3X1 U120 ( .A(memaddr_c[12]), .B(memaddr_c[11]), .C(memaddr_c[7]), .Y(
        n114) );
  NOR43XL U121 ( .B(n230), .C(n200), .D(n199), .A(n112), .Y(n201) );
  AND4X1 U122 ( .A(memaddr_c[9]), .B(memaddr_c[10]), .C(memaddr_c[8]), .D(n229), .Y(n199) );
  NAND21X1 U123 ( .B(n194), .A(n9), .Y(n200) );
  INVX1 U124 ( .A(n110), .Y(hit_xr) );
  INVX1 U125 ( .A(hit_xd), .Y(n183) );
  INVX1 U126 ( .A(n205), .Y(n229) );
  NAND21X1 U127 ( .B(n9), .A(n185), .Y(n193) );
  OAI211X1 U128 ( .C(n55), .D(n237), .A(n3), .B(n211), .Y(xram_we) );
  NAND2X1 U129 ( .A(bist_wr), .B(n8), .Y(n55) );
  NAND21XL U130 ( .B(esfrm_oe), .A(n36), .Y(esfrm_rrdy) );
  INVX1 U131 ( .A(n153), .Y(n40) );
  AO21X1 U132 ( .B(idat_w), .C(n198), .A(n197), .Y(iram_we) );
  OAI33XL U133 ( .A(bist_xram), .B(n12), .C(n195), .D(n194), .E(n193), .F(n192), .Y(n197) );
  INVX1 U134 ( .A(bist_wr), .Y(n195) );
  INVX1 U135 ( .A(idat_adr[7]), .Y(n176) );
  NAND21X1 U136 ( .B(n12), .A(bist_wdat[5]), .Y(n89) );
  INVX1 U137 ( .A(iram_a[9]), .Y(n135) );
  INVX1 U138 ( .A(n185), .Y(n232) );
  INVX1 U139 ( .A(n191), .Y(n219) );
  NAND32X1 U140 ( .B(n212), .C(n190), .A(n189), .Y(n191) );
  OA21X1 U141 ( .B(idat_adr[4]), .C(idat_adr[3]), .A(idat_adr[5]), .Y(n129) );
  AO21X1 U142 ( .B(test_so), .C(n220), .A(n219), .Y(dma_ack) );
  AOI31X1 U143 ( .A(idat_adr[4]), .B(idat_adr[6]), .C(idat_adr[5]), .D(
        idat_adr[7]), .Y(n130) );
  INVX1 U144 ( .A(n91), .Y(n116) );
  AO21X1 U145 ( .B(n188), .C(n187), .A(n186), .Y(n203) );
  MUX2BXL U146 ( .D0(addr1[2]), .D1(n30), .S(n107), .Y(esfrm_adr[2]) );
  MUX2XL U147 ( .D0(addr1[1]), .D1(addr0[1]), .S(n107), .Y(esfrm_adr[1]) );
  NAND4X1 U148 ( .A(n32), .B(n172), .C(n111), .D(n109), .Y(xram_a[6]) );
  NAND2X1 U149 ( .A(memaddr[6]), .B(n120), .Y(n32) );
  INVX1 U150 ( .A(pg0_wrwait), .Y(n41) );
  INVXL U151 ( .A(n224), .Y(n42) );
  NAND43X1 U152 ( .B(dma_r), .C(dma_w), .D(n182), .A(memwr), .Y(n184) );
  OAI2B11X1 U153 ( .D(dma_addr[5]), .C(n156), .A(n169), .B(n106), .Y(xram_a[5]) );
  OAI211X1 U154 ( .C(n226), .D(n225), .A(n224), .B(n223), .Y(n228) );
  INVX1 U155 ( .A(r_i2c_attr), .Y(n225) );
  INVX1 U156 ( .A(n174), .Y(esfrm_adr[6]) );
  AOI21X1 U157 ( .B(xram_rdsel_0_), .C(test_so), .A(n218), .Y(n33) );
  GEN3XL U158 ( .F(xram_rdsel_0_), .G(n52), .E(n51), .D(n50), .C(n97), .B(n49), 
        .A(n212), .Y(n205) );
  INVX1 U159 ( .A(dma_r), .Y(n51) );
  OAI211X1 U160 ( .C(dma_r), .D(memrd_c), .A(xram_rdsel_0_), .B(n48), .Y(n49)
         );
  AND2X1 U161 ( .A(n190), .B(n52), .Y(n48) );
  INVX1 U162 ( .A(n47), .Y(n230) );
  MUX3X1 U163 ( .D0(n44), .D1(n34), .D2(n194), .S0(xram_rdsel_0_), .S1(test_so), .Y(n45) );
  INVX1 U164 ( .A(n212), .Y(n46) );
  NAND21X1 U165 ( .B(dma_w), .A(memrd_c), .Y(n50) );
  NOR2X1 U166 ( .A(dma_r), .B(n50), .Y(n34) );
  INVX1 U167 ( .A(esfrm_wdat[0]), .Y(n59) );
  AOI22X1 U168 ( .A(dma_wdat[0]), .B(n73), .C(memdatao[0]), .D(n72), .Y(n58)
         );
  OAI211X1 U169 ( .C(n229), .D(n3), .A(n211), .B(n210), .Y(xram_ce) );
  MUX3IX1 U170 ( .D0(n209), .D1(n208), .D2(bist_xram), .S0(n230), .S1(bist_en), 
        .Y(n210) );
  AND2X1 U171 ( .A(n229), .B(n203), .Y(n209) );
  AO21X1 U172 ( .B(n207), .C(n206), .A(n205), .Y(n208) );
  AOI211X1 U173 ( .C(memaddr_c[14]), .D(n217), .A(memaddr_c[15]), .B(cpurst), 
        .Y(hit_ps_c) );
  NAND21X1 U174 ( .B(n162), .A(n161), .Y(iram_a[2]) );
  NAND21X1 U175 ( .B(n160), .A(n159), .Y(iram_a[1]) );
  AO22XL U176 ( .A(idat_adr[1]), .B(n198), .C(n179), .D(esfrm_adr[1]), .Y(n160) );
  NAND21X1 U177 ( .B(n158), .A(n157), .Y(iram_a[0]) );
  AO22XL U178 ( .A(idat_adr[0]), .B(n198), .C(n179), .D(esfrm_adr[0]), .Y(n158) );
  OAI211X1 U179 ( .C(n154), .D(n140), .A(n139), .B(n138), .Y(xram_a[9]) );
  INVX1 U180 ( .A(memaddr[9]), .Y(n140) );
  OA21X1 U181 ( .B(n156), .C(n187), .A(n135), .Y(n138) );
  NAND32X1 U182 ( .B(n4), .C(n6), .A(n178), .Y(iram_a[8]) );
  OAI221X1 U183 ( .A(n126), .B(n152), .C(n12), .D(n178), .E(n125), .Y(
        xram_a[8]) );
  INVX1 U184 ( .A(bist_adr[8]), .Y(n178) );
  OAI221X1 U185 ( .A(n192), .B(n177), .C(n181), .D(n176), .E(n175), .Y(
        iram_a[7]) );
  OAI211X1 U186 ( .C(n177), .D(n152), .A(n175), .B(n122), .Y(xram_a[7]) );
  INVX1 U187 ( .A(r_pg0_sel[0]), .Y(n177) );
  OAI2B11X1 U188 ( .D(n128), .C(n181), .A(n192), .B(n180), .Y(iram_a[10]) );
  OAI211X1 U189 ( .C(n186), .D(n156), .A(n180), .B(n155), .Y(xram_a[10]) );
  OAI211X1 U190 ( .C(n129), .D(idat_adr[6]), .A(n130), .B(channel_sel), .Y(
        n128) );
  AOI222XL U191 ( .A(dma_addr[7]), .B(n121), .C(n120), .D(n119), .E(n127), .F(
        n118), .Y(n122) );
  OAI31XL U192 ( .A(n117), .B(n116), .C(n115), .D(n113), .Y(n119) );
  AO21X1 U193 ( .B(channel_sel), .C(n28), .A(memaddr_c[7]), .Y(n118) );
  INVX1 U194 ( .A(channel_sel), .Y(n115) );
  INVX1 U195 ( .A(esfrm_wdat[1]), .Y(n61) );
  AOI22X1 U196 ( .A(dma_wdat[1]), .B(n73), .C(memdatao[1]), .D(n72), .Y(n60)
         );
  OA222X1 U197 ( .A(n156), .B(n188), .C(n124), .D(n141), .E(n154), .F(n123), 
        .Y(n125) );
  INVX1 U198 ( .A(memaddr[8]), .Y(n123) );
  AOI32X1 U199 ( .A(n131), .B(r_pg0_sel[2]), .C(n226), .D(n127), .E(
        memaddr_c[9]), .Y(n139) );
  INVX1 U200 ( .A(esfrm_wdat[2]), .Y(n63) );
  AOI22X1 U201 ( .A(dma_wdat[2]), .B(n73), .C(memdatao[2]), .D(n72), .Y(n62)
         );
  OAI211X1 U202 ( .C(n67), .D(n75), .A(n87), .B(n66), .Y(xram_d[4]) );
  INVX1 U203 ( .A(esfrm_wdat[4]), .Y(n67) );
  AOI22X1 U204 ( .A(dma_wdat[4]), .B(n73), .C(memdatao[4]), .D(n72), .Y(n66)
         );
  OAI211X1 U205 ( .C(n65), .D(n75), .A(n85), .B(n64), .Y(xram_d[3]) );
  INVX1 U206 ( .A(esfrm_wdat[3]), .Y(n65) );
  AOI22X1 U207 ( .A(dma_wdat[3]), .B(n73), .C(memdatao[3]), .D(n72), .Y(n64)
         );
  INVX1 U208 ( .A(memaddr[11]), .Y(n234) );
  OAI211X1 U209 ( .C(r_pg0_sel[1]), .D(r_pg0_sel[0]), .A(r_pg0_sel[2]), .B(
        r_pg0_sel[3]), .Y(n226) );
  AOI211X1 U210 ( .C(memaddr[14]), .D(n136), .A(memaddr[15]), .B(cpurst), .Y(
        hit_ps) );
  NAND4X1 U211 ( .A(n234), .B(n236), .C(n91), .D(n137), .Y(n136) );
  NOR3XL U212 ( .A(memaddr[12]), .B(memaddr[7]), .C(memaddr[13]), .Y(n137) );
  NOR2X1 U213 ( .A(memaddr[8]), .B(memaddr[9]), .Y(n91) );
  OAI211X1 U214 ( .C(n76), .D(n75), .A(n94), .B(n74), .Y(xram_d[7]) );
  INVX1 U215 ( .A(esfrm_wdat[7]), .Y(n76) );
  AOI22X1 U216 ( .A(dma_wdat[7]), .B(n73), .C(memdatao[7]), .D(n72), .Y(n74)
         );
  OAI211X1 U217 ( .C(n69), .D(n75), .A(n89), .B(n68), .Y(xram_d[5]) );
  INVX1 U218 ( .A(esfrm_wdat[5]), .Y(n69) );
  AOI22X1 U219 ( .A(dma_wdat[5]), .B(n73), .C(memdatao[5]), .D(n72), .Y(n68)
         );
  OAI211X1 U220 ( .C(n71), .D(n75), .A(n92), .B(n70), .Y(xram_d[6]) );
  INVX1 U221 ( .A(esfrm_wdat[6]), .Y(n71) );
  AOI22X1 U222 ( .A(dma_wdat[6]), .B(n73), .C(memdatao[6]), .D(n72), .Y(n70)
         );
  NOR4XL U223 ( .A(memaddr[14]), .B(memaddr[15]), .C(memaddr[13]), .D(n134), 
        .Y(hit_xd) );
  OAI211X1 U224 ( .C(n236), .D(n91), .A(n235), .B(n234), .Y(n134) );
  INVX1 U225 ( .A(memaddr[12]), .Y(n235) );
  NAND4X1 U226 ( .A(memaddr[11]), .B(memaddr[7]), .C(n132), .D(n133), .Y(n110)
         );
  NOR43XL U227 ( .B(memaddr[15]), .C(memaddr[13]), .D(memaddr[14]), .A(n235), 
        .Y(n133) );
  AND3X1 U228 ( .A(memaddr[8]), .B(memaddr[9]), .C(memaddr[10]), .Y(n132) );
  AO222X1 U229 ( .A(xram_rdat[7]), .B(n232), .C(iram_rdat[7]), .D(n231), .E(
        regx_rdat[7]), .F(n10), .Y(n142) );
  NOR21XL U230 ( .B(delay_rrdy), .A(r_pg0_rdrdy), .Y(n143) );
  AO21X1 U231 ( .B(r_pg0_sel[1]), .C(n40), .A(n9), .Y(n185) );
  NAND2X1 U232 ( .A(n226), .B(r_pg0_sel[3]), .Y(n153) );
  NOR2X1 U233 ( .A(r_pg0_rdrdy), .B(delay_rrdy), .Y(n36) );
  AO222X1 U234 ( .A(xram_rdat[2]), .B(n232), .C(iram_rdat[2]), .D(n231), .E(
        regx_rdat[2]), .F(n10), .Y(n148) );
  MUX2BXL U235 ( .D0(n212), .D1(bist_xram), .S(n8), .Y(iram_ce) );
  AO222X1 U236 ( .A(xram_rdat[5]), .B(n232), .C(iram_rdat[5]), .D(n231), .E(
        regx_rdat[5]), .F(n10), .Y(n145) );
  AO222X1 U237 ( .A(xram_rdat[3]), .B(n232), .C(iram_rdat[3]), .D(n231), .E(
        regx_rdat[3]), .F(n10), .Y(n147) );
  AO222X1 U238 ( .A(xram_rdat[4]), .B(n232), .C(iram_rdat[4]), .D(n231), .E(
        regx_rdat[4]), .F(n10), .Y(n146) );
  AO222XL U239 ( .A(mcu_esfr_rdat[6]), .B(n36), .C(r_pg0_rdrdy), .D(n144), .E(
        delay_rdat[6]), .F(n143), .Y(esfrm_rdat[6]) );
  AO222X1 U240 ( .A(xram_rdat[6]), .B(n232), .C(iram_rdat[6]), .D(n231), .E(
        regx_rdat[6]), .F(n10), .Y(n144) );
  AO222XL U241 ( .A(mcu_esfr_rdat[1]), .B(n36), .C(r_pg0_rdrdy), .D(n149), .E(
        delay_rdat[1]), .F(n143), .Y(esfrm_rdat[1]) );
  AO222X1 U242 ( .A(xram_rdat[1]), .B(n232), .C(iram_rdat[1]), .D(n231), .E(
        regx_rdat[1]), .F(n10), .Y(n149) );
  AO222XL U243 ( .A(mcu_esfr_rdat[0]), .B(n36), .C(n5), .D(n150), .E(
        delay_rdat[0]), .F(n143), .Y(esfrm_rdat[0]) );
  AO222X1 U244 ( .A(xram_rdat[0]), .B(n232), .C(iram_rdat[0]), .D(n231), .E(
        regx_rdat[0]), .F(n10), .Y(n150) );
  NAND21X1 U245 ( .B(n11), .A(bist_adr[6]), .Y(n172) );
  NAND21X1 U246 ( .B(n11), .A(bist_adr[1]), .Y(n159) );
  NAND21X1 U247 ( .B(n11), .A(bist_adr[2]), .Y(n161) );
  NAND21X1 U248 ( .B(n11), .A(bist_adr[0]), .Y(n157) );
  NAND21X1 U249 ( .B(n11), .A(bist_adr[5]), .Y(n169) );
  NAND21X1 U250 ( .B(n11), .A(bist_adr[3]), .Y(n163) );
  NAND21X1 U251 ( .B(n11), .A(bist_adr[4]), .Y(n166) );
  INVX1 U252 ( .A(test_so), .Y(n52) );
  NOR2X1 U253 ( .A(memrd), .B(memwr), .Y(n37) );
  NAND21X1 U254 ( .B(n12), .A(bist_wdat[7]), .Y(n94) );
  AND2X1 U255 ( .A(bist_adr[9]), .B(n8), .Y(iram_a[9]) );
  NAND21X1 U256 ( .B(n12), .A(bist_adr[10]), .Y(n180) );
  NAND21X1 U257 ( .B(n12), .A(bist_adr[7]), .Y(n175) );
  INVX1 U258 ( .A(memaddr[7]), .Y(n113) );
  INVX1 U259 ( .A(r_pg0_sel[1]), .Y(n126) );
  INVX1 U260 ( .A(xram_rdsel_0_), .Y(n220) );
  INVX1 U261 ( .A(bist_xram), .Y(n237) );
  INVX1 U262 ( .A(dma_w), .Y(n190) );
  INVX1 U263 ( .A(dma_addr[10]), .Y(n186) );
  INVX1 U264 ( .A(dma_addr[8]), .Y(n188) );
  INVX1 U265 ( .A(dma_addr[9]), .Y(n187) );
  OA21XL U266 ( .B(n10), .C(n78), .A(n202), .Y(N46) );
  AND3XL U267 ( .A(n77), .B(n202), .C(n43), .Y(N45) );
  AO21XL U268 ( .B(n10), .C(n202), .A(n201), .Y(regx_re) );
  OAI211XL U269 ( .C(n34), .D(n202), .A(n46), .B(n45), .Y(n47) );
  NAND21XL U270 ( .B(n202), .A(n97), .Y(n44) );
  NAND21XL U271 ( .B(n7), .A(n182), .Y(n189) );
  AO21XL U272 ( .B(n231), .C(n182), .A(n77), .Y(n212) );
  AND3XL U273 ( .A(n77), .B(n1), .C(n43), .Y(N44) );
  NAND21XL U274 ( .B(n231), .A(n1), .Y(n56) );
  INVXL U275 ( .A(n1), .Y(n194) );
  AO222XL U276 ( .A(mcu_esfr_rdat[2]), .B(n36), .C(r_pg0_rdrdy), .D(n148), .E(
        delay_rdat[2]), .F(n143), .Y(esfrm_rdat[2]) );
  OAI221XL U277 ( .A(n174), .B(n192), .C(n181), .D(n173), .E(n172), .Y(
        iram_a[6]) );
  AO222XL U278 ( .A(mcu_esfr_rdat[3]), .B(n36), .C(r_pg0_rdrdy), .D(n147), .E(
        delay_rdat[3]), .F(n143), .Y(esfrm_rdat[3]) );
  AO222XL U279 ( .A(mcu_esfr_rdat[7]), .B(n36), .C(r_pg0_rdrdy), .D(n142), .E(
        delay_rdat[7]), .F(n143), .Y(esfrm_rdat[7]) );
  AO222XL U280 ( .A(mcu_esfr_rdat[5]), .B(n36), .C(r_pg0_rdrdy), .D(n145), .E(
        delay_rdat[5]), .F(n143), .Y(esfrm_rdat[5]) );
  INVX1 U281 ( .A(i_wr[1]), .Y(n233) );
  NAND21XL U282 ( .B(i_wr[0]), .A(n233), .Y(n224) );
  AO22XL U283 ( .A(idat_wdat[1]), .B(n198), .C(esfrm_wdat[1]), .D(n179), .Y(
        n82) );
  AO22XL U284 ( .A(idat_wdat[2]), .B(n198), .C(esfrm_wdat[2]), .D(n179), .Y(
        n84) );
  AO22XL U285 ( .A(idat_wdat[4]), .B(n6), .C(esfrm_wdat[4]), .D(n179), .Y(n88)
         );
  AO22XL U286 ( .A(idat_wdat[5]), .B(n6), .C(esfrm_wdat[5]), .D(n4), .Y(n90)
         );
  AO22XL U287 ( .A(idat_wdat[6]), .B(n198), .C(esfrm_wdat[6]), .D(n179), .Y(
        n93) );
  AO22XL U288 ( .A(idat_wdat[7]), .B(n198), .C(esfrm_wdat[7]), .D(n179), .Y(
        n95) );
  AO22XL U289 ( .A(idat_wdat[0]), .B(n198), .C(esfrm_wdat[0]), .D(n179), .Y(
        n80) );
  AO22XL U290 ( .A(idat_wdat[3]), .B(n198), .C(esfrm_wdat[3]), .D(n179), .Y(
        n86) );
  NAND21X1 U291 ( .B(n82), .A(n81), .Y(iram_d[1]) );
  OAI211XL U292 ( .C(n61), .D(n75), .A(n81), .B(n60), .Y(xram_d[1]) );
  NAND21X1 U293 ( .B(n84), .A(n83), .Y(iram_d[2]) );
  OAI211XL U294 ( .C(n63), .D(n75), .A(n83), .B(n62), .Y(xram_d[2]) );
  NAND21X1 U295 ( .B(n88), .A(n87), .Y(iram_d[4]) );
  NAND21X1 U296 ( .B(n90), .A(n89), .Y(iram_d[5]) );
  NAND21X1 U297 ( .B(n93), .A(n92), .Y(iram_d[6]) );
  NAND21X1 U298 ( .B(n95), .A(n94), .Y(iram_d[7]) );
  NAND21X1 U299 ( .B(n80), .A(n79), .Y(iram_d[0]) );
  OAI211XL U300 ( .C(n59), .D(n75), .A(n79), .B(n58), .Y(xram_d[0]) );
  NAND21X1 U301 ( .B(n86), .A(n85), .Y(iram_d[3]) );
  NAND21XL U302 ( .B(i_rd[0]), .A(n39), .Y(n221) );
  AO222XL U303 ( .A(mcu_esfr_rdat[4]), .B(n36), .C(r_pg0_rdrdy), .D(n146), .E(
        delay_rdat[4]), .F(n143), .Y(esfrm_rdat[4]) );
  AOI222XL U304 ( .A(memaddr[2]), .B(n120), .C(n131), .D(esfrm_adr[2]), .E(
        memaddr_c[2]), .F(n127), .Y(n103) );
  AO22XL U305 ( .A(wdat1[1]), .B(i_wr[1]), .C(wdat0[1]), .D(n233), .Y(
        esfrm_wdat[1]) );
  AO22XL U306 ( .A(wdat1[2]), .B(i_wr[1]), .C(wdat0[2]), .D(n233), .Y(
        esfrm_wdat[2]) );
  AO22XL U307 ( .A(wdat1[4]), .B(i_wr[1]), .C(wdat0[4]), .D(n233), .Y(
        esfrm_wdat[4]) );
  AO22XL U308 ( .A(wdat1[5]), .B(i_wr[1]), .C(wdat0[5]), .D(n233), .Y(
        esfrm_wdat[5]) );
  AO22XL U309 ( .A(wdat1[6]), .B(i_wr[1]), .C(wdat0[6]), .D(n233), .Y(
        esfrm_wdat[6]) );
  AO22XL U310 ( .A(wdat1[7]), .B(i_wr[1]), .C(wdat0[7]), .D(n233), .Y(
        esfrm_wdat[7]) );
  OA22XL U311 ( .A(wdat1[0]), .B(n233), .C(wdat0[0]), .D(i_wr[1]), .Y(
        esfrm_wdat[0]) );
  AO22XL U312 ( .A(wdat1[3]), .B(i_wr[1]), .C(wdat0[3]), .D(n233), .Y(
        esfrm_wdat[3]) );
  MUX2IXL U313 ( .D0(addr1[5]), .D1(addr0[5]), .S(n107), .Y(n171) );
  MUX2IXL U314 ( .D0(addr1[4]), .D1(addr0[4]), .S(n107), .Y(n168) );
  MUX2IXL U315 ( .D0(addr1[3]), .D1(addr0[3]), .S(n107), .Y(n165) );
  MUX2IXL U316 ( .D0(addr1[0]), .D1(addr0[0]), .S(n107), .Y(n101) );
  OAI2B11X4 U317 ( .D(dma_addr[2]), .C(n156), .A(n161), .B(n103), .Y(xram_a[2]) );
endmodule


module ATO0008KX8MX180LBX4DA ( A, CSB, CLK, PGM, RE, TWLB, VSS, VDD, VDDP, SAP, 
        Q );
  input [15:0] A;
  input [1:0] TWLB;
  input [1:0] SAP;
  output [7:0] Q;
  input CSB, CLK, PGM, RE, VSS, VDD, VDDP;


endmodule


module MSL18B_1536X8_RW10TM4_16_20221107 ( DO, CK, CSB, OEB, WEB, A, DI );
  output [7:0] DO;
  input [10:0] A;
  input [7:0] DI;
  input CK, CSB, OEB, WEB;


endmodule


module IOBMURUDA_A1 ( PAD, IE, DI, OE, DO, PU, PD, ANA_R, RSTB_5, VB, ANA_P );
  input IE, OE, DO, PU, PD, RSTB_5, VB, ANA_P;
  output DI, ANA_R;
  inout PAD;


endmodule


module IOBMURUDA_A0 ( PAD, IE, DI, OE, DO, PU, PD, ANA_R, RSTB_5, VB );
  input IE, OE, DO, PU, PD, RSTB_5, VB;
  output DI, ANA_R;
  inout PAD;


endmodule


module IODMURUDA_A0 ( PAD, IE, DI, OE, DO, PU, PD, ANA_R, RSTB_5, VB );
  input IE, OE, DO, PU, PD, RSTB_5, VB;
  output DI, ANA_R;
  inout PAD;


endmodule


module anatop_1127a0 ( CC1, CC2, DP, DN, VFB, CSP, CSN, COM, SW, BST, VDRV, LG, 
        HG, GATE, BST_SET, DCM_SEL, HGOFF, HGON, LGOFF, LGON, EN_DRV, FSW, 
        EN_OSC, MAXDS, EN_GM, EN_ODLDO, EN_IBUK, CP_EN, EXT_CP, INT_CP, 
        ANTI_INRUSH, PWREN_HOLD, RP_SEL, RP1_EN, RP2_EN, VCONN1_EN, VCONN2_EN, 
        SGP, S20U, S100U, TX_EN, TX_DAT, CC_SEL, TRA, TFA, LSR, RX_DAT, RX_SQL, 
        SEL_RX_TH, DAC1_EN, DPDN_SHORT, DP_2V7_EN, DN_2V7_EN, DP_0P6V_EN, 
        DN_0P6V_EN, DP_DWN_EN, DN_DWN_EN, PWR_I, DAC3, DAC1, CV2, LFOSC_ENB, 
        VO_DISCHG, DISCHG_SEL, CMP_SEL_VO10, CMP_SEL_VO20, CMP_SEL_GP1, 
        CMP_SEL_GP2, CMP_SEL_GP3, CMP_SEL_GP4, CMP_SEL_GP5, CMP_SEL_VIN20, 
        CMP_SEL_TS, CMP_SEL_IS, CMP_SEL_CC2, CMP_SEL_CC1, CMP_SEL_CC2_4, 
        CMP_SEL_CC1_4, CMP_SEL_DP, CMP_SEL_DP_3, CMP_SEL_DN, CMP_SEL_DN_3, 
        OCP_EN, CS_EN, COMP_O, CCI2C_EN, UVP_SEL, TM, V5OCP, RSTB, DAC0, SLEEP, 
        OSC_LOW, OSC_STOP, PWRDN, VPP_ZERO, OSC_O, RD_DET, IMP_OSC, DRP_OSC, 
        STB_RP, RD_ENB, OCP, SCP, UVP, LDO3P9V, VPP_SEL, CC1_DOB, CC2_DOB, 
        CC1_DI, CC2_DI, OTPI, OVP_SEL, OVP, DN_COMP, DP_COMP, DPDN_VTH, DPDEN, 
        DPDO, DPIE, DNDEN, DNDO, DNIE, DUMMY_IN, CP_CLKX2, SEL_CONST_OVP, 
        LP_EN, DNCHK_EN, IRP_EN, CCBFEN, REGTRM, AD_RST, AD_HOLD, DN_FAULT, 
        SEL_CCGAIN, VFB_SW, CPVSEL, CLAMPV_EN, HVNG_CPEN, OCP_SEL, OCP_80M, 
        OCP_160M, OPTO1, OPTO2, VPP_OTP, RSTB_5, V1P1, TS_ANA_R, GP5_ANA_R, 
        GP4_ANA_R, GP3_ANA_R, GP2_ANA_R, GP1_ANA_R, TS_ANA_P, GP5_ANA_P, 
        GP4_ANA_P, GP3_ANA_P, GP2_ANA_P, GP1_ANA_P );
  input [1:0] FSW;
  input [1:0] RP_SEL;
  input [5:1] SGP;
  input [7:0] PWR_I;
  input [5:0] DAC3;
  input [9:0] DAC1;
  input [3:0] TM;
  input [10:0] DAC0;
  input [1:0] OVP_SEL;
  input [7:0] DUMMY_IN;
  input [55:0] REGTRM;
  input BST_SET, DCM_SEL, HGOFF, HGON, LGOFF, LGON, EN_DRV, EN_OSC, MAXDS,
         EN_GM, EN_ODLDO, EN_IBUK, CP_EN, EXT_CP, INT_CP, ANTI_INRUSH,
         PWREN_HOLD, RP1_EN, RP2_EN, VCONN1_EN, VCONN2_EN, S20U, S100U, TX_EN,
         TX_DAT, CC_SEL, TRA, TFA, LSR, SEL_RX_TH, DAC1_EN, DPDN_SHORT,
         DP_2V7_EN, DN_2V7_EN, DP_0P6V_EN, DN_0P6V_EN, DP_DWN_EN, DN_DWN_EN,
         CV2, LFOSC_ENB, VO_DISCHG, DISCHG_SEL, CMP_SEL_VO10, CMP_SEL_VO20,
         CMP_SEL_GP1, CMP_SEL_GP2, CMP_SEL_GP3, CMP_SEL_GP4, CMP_SEL_GP5,
         CMP_SEL_VIN20, CMP_SEL_TS, CMP_SEL_IS, CMP_SEL_CC2, CMP_SEL_CC1,
         CMP_SEL_CC2_4, CMP_SEL_CC1_4, CMP_SEL_DP, CMP_SEL_DP_3, CMP_SEL_DN,
         CMP_SEL_DN_3, OCP_EN, CS_EN, CCI2C_EN, UVP_SEL, SLEEP, OSC_LOW,
         OSC_STOP, PWRDN, VPP_ZERO, STB_RP, RD_ENB, LDO3P9V, VPP_SEL, CC1_DOB,
         CC2_DOB, DPDN_VTH, DPDEN, DPDO, DPIE, DNDEN, DNDO, DNIE, CP_CLKX2,
         SEL_CONST_OVP, LP_EN, DNCHK_EN, IRP_EN, CCBFEN, AD_RST, AD_HOLD,
         SEL_CCGAIN, VFB_SW, CPVSEL, CLAMPV_EN, HVNG_CPEN, OCP_SEL, TS_ANA_R,
         GP5_ANA_R, GP4_ANA_R, GP3_ANA_R, GP2_ANA_R, GP1_ANA_R;
  output LG, HG, GATE, RX_DAT, RX_SQL, COMP_O, V5OCP, RSTB, OSC_O, RD_DET,
         IMP_OSC, DRP_OSC, OCP, SCP, UVP, CC1_DI, CC2_DI, OTPI, OVP, DN_COMP,
         DP_COMP, DN_FAULT, OCP_80M, OCP_160M, OPTO1, OPTO2, VPP_OTP, RSTB_5,
         V1P1, TS_ANA_P, GP5_ANA_P, GP4_ANA_P, GP3_ANA_P, GP2_ANA_P, GP1_ANA_P;
  inout CC1,  CC2,  DP,  DN,  VFB,  CSP,  CSN,  COM,  SW,  BST,  VDRV;


endmodule

