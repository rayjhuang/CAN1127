
module chiptop_1127a0 ( CSP, CSN, VFB, COM, LG, SW, HG, BST, GATE, VDRV, DP, 
        DN, CC1, CC2, TST, GPIO_TS, SCL, SDA, GPIO1, GPIO2, GPIO3, GPIO4, 
        GPIO5 );
  input TST;
  inout CSP,  CSN,  VFB,  COM,  LG,  SW,  HG,  BST,  GATE,  VDRV,  DP,  DN, 
     CC1,  CC2,  GPIO_TS,  SCL,  SDA,  GPIO1,  GPIO2,  GPIO3,  GPIO4,  GPIO5;
  wire   SRAM_WEB, SRAM_CEB, SRAM_OEB, RD_ENB, STB_RP, DRP_OSC, IMP_OSC, TX_EN,
         TX_DAT, RX_DAT, RX_SQL, DAC1_EN, AD_RST, AD_HOLD, COMP_O, CCI2C_EN,
         RSTB, SLEEP, OSC_LOW, OSC_STOP, PWRDN, VPP_0V, VPP_SEL, LDO3P9V,
         OSC_O, RD_DET, OCP_SEL, CC1_DOB, CC2_DOB, CC1_DI, CC2_DI, DP_COMP,
         DN_COMP, DN_FAULT, PWREN_HOLD, LFOSC_ENB, VPP_OTP, IO_RSTB5, V1P1,
         ANAP_TS, TS_ANA_R, ANAP_GP1, GP1_ANA_R, ANAP_GP2, GP2_ANA_R, ANAP_GP3,
         GP3_ANA_R, ANAP_GP4, GP4_ANA_R, ANAP_GP5, GP5_ANA_R, DI_TST, DI_TS,
         SRAM_CLK, PMEM_RE, PMEM_PGM, PMEM_CSB, do_ccctl_0_, do_srcctl_0,
         tm_atpg, n1, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, net1, net2, net3, net4;
  wire   [10:0] SRAM_A;
  wire   [7:0] SRAM_D;
  wire   [7:0] xdat_o;
  wire   [7:0] ANAOPT;
  wire   [1:0] FSW;
  wire   [1:0] RP_EN;
  wire   [1:0] VCONN_EN;
  wire   [17:0] SAMPL_SEL;
  wire   [7:0] DUMMY_IN;
  wire   [55:0] REGTRM;
  wire   [7:0] PWR_I;
  wire   [1:0] OVP_SEL;
  wire   [5:0] DAC3_V;
  wire   [10:0] DAC0;
  wire   [3:0] ANA_TM;
  wire   [9:0] DAC1;
  wire   [1:0] RP_SEL;
  wire   [1:0] IE_GPIO;
  wire   [6:0] DI_GPIO;
  wire   [6:0] OE_GPIO;
  wire   [6:0] DO_GPIO;
  wire   [6:0] PU_GPIO;
  wire   [6:0] PD_GPIO;
  wire   [3:0] DO_TS;
  wire   [1:0] PMEM_CLK;
  wire   [7:0] PMEM_Q1;
  wire   [7:0] PMEM_Q0;
  wire   [1:0] PMEM_SAP;
  wire   [1:0] PMEM_TWLB;
  wire   [15:0] PMEM_A;
  wire   [6:0] bck_regx0;
  wire   [7:2] do_xana1;
  wire   [7:0] do_xana0;
  wire   [3:0] do_regx_xtm;
  wire   [5:2] do_cvctl;
  wire   [3:0] do_vooc;
  wire   [5:0] do_dpdm;
  wire   [5:4] do_srcctl;
  wire   [7:0] do_cctrx;
  wire   [3:0] di_xanav;
  wire   [5:0] srci;
  tri   VFB;
  tri   COM;
  tri   LG;
  tri   SW;
  tri   HG;
  tri   BST;
  tri   GATE;
  tri   VDRV;
  tri   DP;
  tri   DN;
  tri   CC1;
  tri   CC2;
  tri   TST;
  tri   GPIO_TS;
  tri   SCL;
  tri   SDA;
  tri   GPIO1;
  tri   GPIO2;
  tri   GPIO3;
  tri   GPIO4;
  tri   GPIO5;

  anatop_1127a0 U0_ANALOG_TOP ( .CC1(CC1), .CC2(CC2), .DP(DP), .DN(DN), .VFB(
        VFB), .CSP(), .CSN(), .COM(COM), .LG(LG), .SW(SW), .HG(HG), .BST(BST), 
        .GATE(GATE), .VDRV(VDRV), .BST_SET(bck_regx0[0]), .DCM_SEL(
        bck_regx0[1]), .HGOFF(bck_regx0[2]), .HGLGOFF(bck_regx0[3]), .HGON(
        bck_regx0[4]), .LGON(bck_regx0[5]), .ENDRV(bck_regx0[6]), .FSW(FSW), 
        .EN_OSC(bck_regx0[2]), .MAXDS(bck_regx0[3]), .EN_GM(bck_regx0[4]), 
        .EN_ODLDO(bck_regx0[5]), .EN_IBUK(bck_regx0[6]), .RP_SEL(RP_SEL), 
        .RP1_EN(RP_EN[0]), .RP2_EN(RP_EN[1]), .VCONN1_EN(VCONN_EN[0]), 
        .VCONN2_EN(VCONN_EN[1]), .SGP({do_cctrx[0], do_regx_xtm}), .S20U(
        do_cctrx[1]), .S100U(do_cctrx[2]), .TX_EN(TX_EN), .TX_DAT(TX_DAT), 
        .CC_SEL(do_ccctl_0_), .TRA(do_cctrx[4]), .TFA(do_cctrx[5]), .LSR(
        do_cctrx[6]), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .SEL_RX_TH(do_cctrx[7]), .DAC1_EN(DAC1_EN), .DPDN_SHORT(do_dpdm[0]), .DP_2V7_EN(do_dpdm[4]), 
        .DN_2V7_EN(do_dpdm[3]), .DP_0P6V_EN(do_xana1[3]), .DN_0P6V_EN(
        do_xana1[2]), .DP_DWN_EN(do_dpdm[2]), .DN_DWN_EN(do_dpdm[1]), .PWR_I(
        PWR_I), .DAC3(DAC3_V), .DAC1(DAC1), .CV2(do_xana0[0]), .LFOSC_ENB(
        LFOSC_ENB), .VO_DISCHG(do_srcctl[4]), .DISCHG_SEL(do_srcctl[5]), 
        .CMP_SEL_VO10(SAMPL_SEL[0]), .CMP_SEL_VO20(SAMPL_SEL[10]), 
        .CMP_SEL_GP1(SAMPL_SEL[17]), .CMP_SEL_GP2(SAMPL_SEL[16]), 
        .CMP_SEL_GP3(SAMPL_SEL[15]), .CMP_SEL_GP4(SAMPL_SEL[14]), 
        .CMP_SEL_GP5(SAMPL_SEL[13]), .CMP_SEL_VIN20(SAMPL_SEL[1]), 
        .CMP_SEL_TS(SAMPL_SEL[3]), .CMP_SEL_IS(SAMPL_SEL[2]), .CMP_SEL_CC2(
        SAMPL_SEL[7]), .CMP_SEL_CC1(SAMPL_SEL[6]), .CMP_SEL_CC2_4(
        SAMPL_SEL[12]), .CMP_SEL_CC1_4(SAMPL_SEL[11]), .CMP_SEL_DP(
        SAMPL_SEL[4]), .CMP_SEL_DP_3(SAMPL_SEL[8]), .CMP_SEL_DN(SAMPL_SEL[5]), 
        .CMP_SEL_DN_3(SAMPL_SEL[9]), .OCP_EN(do_cvctl[2]), .CS_EN(do_cctrx[3]), 
        .COMP_O(COMP_O), .CCI2C_EN(CCI2C_EN), .UVP_SEL(do_xana0[7]), .TM(
        ANA_TM), .V5OCP(srci[4]), .RSTB(RSTB), .DAC0(DAC0), .SLEEP(SLEEP), 
        .OSC_LOW(OSC_LOW), .OSC_STOP(OSC_STOP), .PWRDN(PWRDN), .VPP_ZERO(
        VPP_0V), .OSC_O(OSC_O), .RD_DET(RD_DET), .IMP_OSC(IMP_OSC), .DRP_OSC(
        DRP_OSC), .STB_RP(STB_RP), .RD_ENB(RD_ENB), .PWREN(do_srcctl_0), .OCP(
        srci[1]), .SCP(srci[3]), .UVP(srci[0]), .LDO3P9V(LDO3P9V), .VPP_SEL(
        VPP_SEL), .CC1_DOB(CC1_DOB), .CC2_DOB(CC2_DOB), .CC1_DI(CC1_DI), 
        .CC2_DI(CC2_DI), .ANTI_INRUSH(do_cvctl[5]), .OTPI(srci[5]), .OVP_SEL(
        OVP_SEL), .OVP(srci[2]), .DN_COMP(DN_COMP), .DP_COMP(DP_COMP), 
        .DPDN_VTH(do_xana0[5]), .DPDEN(do_vooc[3]), .DPDO(do_vooc[2]), .DPIE(
        do_dpdm[5]), .DNDEN(do_vooc[1]), .DNDO(do_vooc[0]), .DNIE(do_dpdm[5]), 
        .DUMMY_IN(DUMMY_IN), .CP_CLKX2(ANAOPT[7]), .SEL_CONST_OVP(ANAOPT[6]), 
        .LP_EN(ANAOPT[5]), .DNCHK_EN(ANAOPT[3]), .IRP_EN(ANAOPT[2]), .CCBFEN(
        ANAOPT[0]), .REGTRM(REGTRM), .AD_RST(AD_RST), .AD_HOLD(AD_HOLD), 
        .DN_FAULT(DN_FAULT), .SEL_CCGAIN(do_xana0[3]), .VFB_SW(do_xana0[1]), 
        .CPV_SEL(do_xana1[6]), .CLAMPV_EN(do_xana1[5]), .HVNG_CPEN(do_xana1[7]), .PWREN_HOLD(PWREN_HOLD), .OCP_SEL(OCP_SEL), .OCP_80M(di_xanav[1]), 
        .OCP_160M(di_xanav[0]), .OPTO1(di_xanav[2]), .OPTO2(di_xanav[3]), 
        .VPP_OTP(VPP_OTP), .VDD_OTP(), .RSTB_5(IO_RSTB5), .V1P1(V1P1), 
        .TS_ANA_R(TS_ANA_R), .GP5_ANA_R(GP5_ANA_R), .GP4_ANA_R(GP4_ANA_R), 
        .GP3_ANA_R(GP3_ANA_R), .GP2_ANA_R(GP2_ANA_R), .GP1_ANA_R(GP1_ANA_R), 
        .TS_ANA_P(ANAP_TS), .GP5_ANA_P(ANAP_GP5), .GP4_ANA_P(ANAP_GP4), 
        .GP3_ANA_P(ANAP_GP3), .GP2_ANA_P(ANAP_GP2), .GP1_ANA_P(ANAP_GP1) );
  IODMURUDA_A0 PAD_SCL ( .PAD(SCL), .IE(IE_GPIO[1]), .DI(DI_GPIO[0]), .OE(
        OE_GPIO[0]), .DO(DO_GPIO[0]), .PU(PU_GPIO[0]), .PD(PD_GPIO[0]), 
        .ANA_R(), .RSTB_5(IO_RSTB5), .VB(V1P1) );
  IODMURUDA_A0 PAD_SDA ( .PAD(SDA), .IE(IE_GPIO[1]), .DI(DI_GPIO[1]), .OE(
        OE_GPIO[1]), .DO(DO_GPIO[1]), .PU(PU_GPIO[1]), .PD(PD_GPIO[1]), 
        .ANA_R(), .RSTB_5(IO_RSTB5), .VB(V1P1) );
  IOBMURUDA_A0 PAD_TST ( .PAD(TST), .IE(1'b1), .DI(DI_TST), .OE(1'b0), .DO(
        1'b0), .PU(1'b0), .PD(1'b1), .ANA_R(), .RSTB_5(IO_RSTB5), .VB(V1P1) );
  IOBMURUDA_A1 PAD_GPIO1 ( .PAD(GPIO1), .IE(IE_GPIO[0]), .DI(DI_GPIO[2]), .OE(
        OE_GPIO[2]), .DO(DO_GPIO[2]), .PU(PU_GPIO[2]), .PD(PD_GPIO[2]), 
        .ANA_R(GP1_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP1) );
  IOBMURUDA_A1 PAD_GPIO2 ( .PAD(GPIO2), .IE(IE_GPIO[0]), .DI(DI_GPIO[3]), .OE(
        OE_GPIO[3]), .DO(DO_GPIO[3]), .PU(PU_GPIO[3]), .PD(PD_GPIO[3]), 
        .ANA_R(GP2_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP2) );
  IOBMURUDA_A1 PAD_GPIO3 ( .PAD(GPIO3), .IE(IE_GPIO[0]), .DI(DI_GPIO[4]), .OE(
        OE_GPIO[4]), .DO(DO_GPIO[4]), .PU(PU_GPIO[4]), .PD(PD_GPIO[4]), 
        .ANA_R(GP3_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP3) );
  IOBMURUDA_A1 PAD_GPIO4 ( .PAD(GPIO4), .IE(IE_GPIO[0]), .DI(DI_GPIO[5]), .OE(
        OE_GPIO[5]), .DO(DO_GPIO[5]), .PU(PU_GPIO[5]), .PD(PD_GPIO[5]), 
        .ANA_R(GP4_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP4) );
  IOBMURUDA_A1 PAD_GPIO5 ( .PAD(GPIO5), .IE(IE_GPIO[0]), .DI(DI_GPIO[6]), .OE(
        OE_GPIO[6]), .DO(DO_GPIO[6]), .PU(PU_GPIO[6]), .PD(PD_GPIO[6]), 
        .ANA_R(GP5_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_GP5) );
  IOBMURUDA_A1 PAD_GPIO_TS ( .PAD(GPIO_TS), .IE(IE_GPIO[0]), .DI(DI_TS), .OE(
        DO_TS[2]), .DO(DO_TS[3]), .PU(DO_TS[1]), .PD(DO_TS[0]), .ANA_R(
        TS_ANA_R), .RSTB_5(IO_RSTB5), .VB(V1P1), .ANA_P(ANAP_TS) );
  MSL18B_1536X8_RW10TM4_16 U0_SRAM ( .DO(xdat_o), .CK(SRAM_CLK), .CSB(SRAM_CEB), .OEB(SRAM_OEB), .WEB(SRAM_WEB), .A(SRAM_A), .DI(SRAM_D) );
  ATO0008KX8MX180LBX4DA U0_CODE_0_ ( .A(PMEM_A), .CSB(PMEM_CSB), .CLK(
        PMEM_CLK[0]), .PGM(n1), .RE(PMEM_RE), .TWLB(PMEM_TWLB), .VSS(net3), 
        .VDD(net4), .VDDP(VPP_OTP), .SAP(PMEM_SAP), .Q(PMEM_Q0) );
  ATO0008KX8MX180LBX4DA U0_CODE_1_ ( .A(PMEM_A), .CSB(PMEM_CSB), .CLK(
        PMEM_CLK[1]), .PGM(PMEM_PGM), .RE(PMEM_RE), .TWLB(PMEM_TWLB), .VSS(
        net1), .VDD(net2), .VDDP(VPP_OTP), .SAP(PMEM_SAP), .Q(PMEM_Q1) );
  core_a0 U0_CORE ( .SRCI(srci), .XANAV({1'b0, di_xanav}), .BCK_REGX({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        FSW, SYNOPSYS_UNCONNECTED_7, bck_regx0}), .ANA_REGX({do_xana1[7:5], 
        SYNOPSYS_UNCONNECTED_8, do_xana1[3:2], SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, do_xana0[7], SYNOPSYS_UNCONNECTED_11, 
        do_xana0[5], SYNOPSYS_UNCONNECTED_12, do_xana0[3], 
        SYNOPSYS_UNCONNECTED_13, do_xana0[1:0]}), .LFOSC_ENB(LFOSC_ENB), 
        .STB_RP(STB_RP), .RD_ENB(RD_ENB), .OCP_SEL(OCP_SEL), .PWREN_HOLD(
        PWREN_HOLD), .CC1_DI(CC1_DI), .CC2_DI(CC2_DI), .DRP_OSC(DRP_OSC), 
        .IMP_OSC(IMP_OSC), .CC1_DOB(CC1_DOB), .CC2_DOB(CC2_DOB), .DAC1_EN(
        DAC1_EN), .SH_RST(AD_RST), .SH_HOLD(AD_HOLD), .LDO3P9V(LDO3P9V), .XTM(
        do_regx_xtm), .DO_CVCTL({OVP_SEL, do_cvctl[5], SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, do_cvctl[2], SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17}), .DO_CCTRX(do_cctrx), .DO_SRCCTL({
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, do_srcctl, VCONN_EN, 
        SYNOPSYS_UNCONNECTED_20, do_srcctl_0}), .DO_CCCTL({RP_EN, RP_SEL, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, do_ccctl_0_}), .DO_DAC0(DAC0), .DO_DPDN(
        do_dpdm), .DO_VOOC(do_vooc), .DO_PWR_I(PWR_I), .PMEM_A(PMEM_A), 
        .PMEM_Q0(PMEM_Q0), .PMEM_Q1(PMEM_Q1), .PMEM_TWLB(PMEM_TWLB), 
        .PMEM_SAP(PMEM_SAP), .PMEM_CLK(PMEM_CLK), .PMEM_CSB(PMEM_CSB), 
        .PMEM_RE(PMEM_RE), .PMEM_PGM(PMEM_PGM), .VPP_SEL(VPP_SEL), .VPP_0V(
        VPP_0V), .SRAM_WEB(SRAM_WEB), .SRAM_CEB(SRAM_CEB), .SRAM_OEB(SRAM_OEB), 
        .SRAM_CLK(SRAM_CLK), .SRAM_A(SRAM_A), .SRAM_D(SRAM_D), .SRAM_RDAT(
        xdat_o), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .RD_DET(RD_DET), .STB_OVP(
        1'b0), .TX_DAT(TX_DAT), .TX_EN(TX_EN), .OSC_STOP(OSC_STOP), .OSC_LOW(
        OSC_LOW), .SLEEP(SLEEP), .PWRDN(PWRDN), .OCDRV_ENZ(), .DAC1_V(DAC1), 
        .SAMPL_SEL(SAMPL_SEL), .DAC1_COMP(COMP_O), .CCI2C_EN(CCI2C_EN), 
        .ANA_TM(ANA_TM), .DM_FAULT(DN_FAULT), .DM_COMP(DN_COMP), .DP_COMP(
        DP_COMP), .DI_GPIO(DI_GPIO), .DO_GPIO(DO_GPIO), .OE_GPIO(OE_GPIO), 
        .GPIO_PU(PU_GPIO), .GPIO_PD(PD_GPIO), .GPIO_IE(IE_GPIO), .DO_TS(DO_TS), 
        .DI_TS(DI_TS), .REGTRM(REGTRM), .ANAOPT({ANAOPT[7:5], 
        SYNOPSYS_UNCONNECTED_24, ANAOPT[3:2], SYNOPSYS_UNCONNECTED_25, 
        ANAOPT[0]}), .DUMMY_IN(DUMMY_IN), .DAC3_V(DAC3_V), .i_clk(OSC_O), 
        .i_rstz(RSTB), .atpg_en(tm_atpg), .di_tst(DI_TST), .tm_atpg(tm_atpg)
         );
  BUFX12 U3 ( .A(PMEM_PGM), .Y(n1) );
endmodule


module core_a0 ( SRCI, XANAV, BCK_REGX, ANA_REGX, LFOSC_ENB, STB_RP, RD_ENB, 
        OCP_SEL, PWREN_HOLD, CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, CC1_DOB, 
        CC2_DOB, DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, XTM, DO_CVCTL, DO_CCTRX, 
        DO_SRCCTL, DO_CCCTL, DO_DAC0, DO_DPDN, DO_VOOC, DO_PWR_I, PMEM_A, 
        PMEM_Q0, PMEM_Q1, PMEM_TWLB, PMEM_SAP, PMEM_CLK, PMEM_CSB, PMEM_RE, 
        PMEM_PGM, VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, 
        SRAM_A, SRAM_D, SRAM_RDAT, RX_DAT, RX_SQL, RD_DET, STB_OVP, TX_DAT, 
        TX_EN, OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, DAC1_V, SAMPL_SEL, 
        DAC1_COMP, CCI2C_EN, ANA_TM, DM_FAULT, DM_COMP, DP_COMP, DI_GPIO, 
        DO_GPIO, OE_GPIO, GPIO_PU, GPIO_PD, GPIO_IE, DO_TS, DI_TS, REGTRM, 
        ANAOPT, DUMMY_IN, DAC3_V, i_clk, i_rstz, atpg_en, di_tst, tm_atpg );
  input [5:0] SRCI;
  input [4:0] XANAV;
  output [15:0] BCK_REGX;
  output [15:0] ANA_REGX;
  output [3:0] XTM;
  output [7:0] DO_CVCTL;
  output [7:0] DO_CCTRX;
  output [7:0] DO_SRCCTL;
  output [7:0] DO_CCCTL;
  output [10:0] DO_DAC0;
  output [5:0] DO_DPDN;
  output [3:0] DO_VOOC;
  output [7:0] DO_PWR_I;
  output [15:0] PMEM_A;
  input [7:0] PMEM_Q0;
  input [7:0] PMEM_Q1;
  output [1:0] PMEM_TWLB;
  output [1:0] PMEM_SAP;
  output [1:0] PMEM_CLK;
  output [10:0] SRAM_A;
  output [7:0] SRAM_D;
  input [7:0] SRAM_RDAT;
  output [9:0] DAC1_V;
  output [17:0] SAMPL_SEL;
  output [3:0] ANA_TM;
  input [6:0] DI_GPIO;
  output [6:0] DO_GPIO;
  output [6:0] OE_GPIO;
  output [6:0] GPIO_PU;
  output [6:0] GPIO_PD;
  output [1:0] GPIO_IE;
  output [3:0] DO_TS;
  output [55:0] REGTRM;
  output [7:0] ANAOPT;
  output [7:0] DUMMY_IN;
  output [5:0] DAC3_V;
  input CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, RX_DAT, RX_SQL, RD_DET, STB_OVP,
         DAC1_COMP, DM_FAULT, DM_COMP, DP_COMP, DI_TS, i_clk, i_rstz, atpg_en,
         di_tst;
  output LFOSC_ENB, STB_RP, RD_ENB, OCP_SEL, PWREN_HOLD, CC1_DOB, CC2_DOB,
         DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, PMEM_CSB, PMEM_RE, PMEM_PGM,
         VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, TX_DAT,
         TX_EN, OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, CCI2C_EN, tm_atpg;
  wire   N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, n638, n639, aswclk, detclk, tclk_sel, s_clk, aswkup, x_clk,
         t_di_gpio4, r_osc_gate, g_clk, xram_ce, iram_ce, sram_en, r_i2c_attr,
         esfrm_oe, esfrm_we, sfrack, ictlr_psrack, esfrm_rrdy, memwr, memrd,
         memrd_c, memack, o_cpurst, hit_xd, hit_xr, hit_ps, hit_ps_c,
         mcu_ram_r, mcu_ram_w, regx_re, iram_we, xram_we, regx_we, bist_en,
         bist_wr, srstz, prl_cany0w, prl_cany0r, mempsrd, r_bclk_sel,
         r_hold_mcu, t0_intr, fcp_intr, dpdm_urx, s0_rxdoe, mcuo_scl, mcuo_sda,
         mempsack, mempswr, mempsrd_c, sfr_w, sfr_r, ictlr_psack, ictlr_inc,
         set_hold, bkpt_hold, bkpt_ena, r_psrd, r_pswr, prl_cany0, prl_c0set,
         pmem_pgm, pmem_re, pmem_csb, we_twlb, r_otp_wpls, pwrdn_rst,
         r_otp_pwdn_en, ramacc, r_sleep, ps_pwrdn, r_pwrdn, r_ocdrv_enz,
         r_osc_stop, r_pwrv_upd, r_otpi_gate, r_fcpre, r_fortxdat, r_fortxrdy,
         r_fortxen, r_gpio_tm, pid_goidle, pid_gobusy, bus_idle, sse_idle,
         r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, r_unlock, r_first, r_last,
         r_fiforst, r_set_cpmsgid, r_txendk, r_txshrt, r_auto_discard,
         r_dat_portrole, r_dat_datarole, r_pshords, r_discard, r_strtch,
         r_i2c_ninc, r_i2c_fwnak, r_i2c_fwack, hwi2c_stretch, i2c_ev_6_,
         i2c_ev_3, i2c_ev_2, prl_discard, prl_GCTxDone, pff_obsd, pff_empty,
         pff_full, ptx_ack, clk_1500k, clk_500k, clk_500, prstz, sse_rdrdy,
         upd_rdrdy, sse_prefetch, slvo_sda, slvo_re, slvo_early, dm_comp,
         dp_comp, di_cc, ptx_cc, ptx_oe, sh_rst, sh_hold, fcp_oe, fcp_do,
         sdischg_duty, clk_100k, r_imp_osc, r_vpp_en, r_vpp0v_en, di_ts,
         r_xana_23, r_xana_19, r_xana_18, divff_8, divff_5, clk_50k, N449,
         N450, o_dodat0_15_, o_dodat5_2_, N570, N571, N572, N573, N574, N579,
         N580, N581, N582, N583, N584, N585, N586, N1483, N1488, N1493, N1498,
         net8831, n504, n505, n506, n507, n51, n52, n53, n110, n111, n112,
         n113, n114, n115, n116, n117, n8, n20, n21, n22, n132, n535, n632,
         n633, n634, n635, n636, n637, n672, n673, n674, n706, n761, n762,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n857, n858, n859, n860, n861, n862, n863, n869, n875,
         n899, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n955, n957, n958, n959, n960, n961, n962,
         n963, n964, n970, n972, n973, n979, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1086, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1, n2, n3, n4, n5, n6, n7,
         n9, n10, n11, n12, n13, n14, n16, n17, n18, n19, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100;
  wire   [9:0] aswclk_ps;
  wire   [9:0] detclk_ps;
  wire   [7:0] sse_wdat;
  wire   [7:0] prx_fifowdat;
  wire   [7:0] sse_adr;
  wire   [7:0] prl_cany0adr;
  wire   [7:0] esfrm_wdat;
  wire   [6:0] esfrm_adr;
  wire   [7:0] mcu_esfrrdat;
  wire   [7:0] delay_inst;
  wire   [7:0] esfrm_rdat;
  wire   [3:0] r_pg0_sel;
  wire   [15:0] memaddr;
  wire   [15:0] memaddr_c;
  wire   [7:0] memdatao;
  wire   [7:0] idat_adr;
  wire   [7:0] idat_wdat;
  wire   [10:0] iram_a;
  wire   [10:0] xram_a;
  wire   [7:0] iram_d;
  wire   [7:0] xram_d;
  wire   [1:0] sram_rdat;
  wire   [7:0] regx_rdat;
  wire   [10:0] bist_adr;
  wire   [7:0] bist_wdat;
  wire   [7:0] memdatai;
  wire   [7:0] ictlr_inst;
  wire   [15:0] mcu_pc;
  wire   [22:16] mcu_dbgpo;
  wire   [3:2] sfr_intr;
  wire   [7:0] exint;
  wire   [7:0] ff_p0;
  wire   [6:0] do_p0;
  wire   [7:0] sfr_rdat;
  wire   [7:0] sfr_wdat;
  wire   [6:0] sfr_adr;
  wire   [14:0] bkpt_pc;
  wire   [14:0] r_inst_ofs;
  wire   [1:0] pmem_clk;
  wire   [7:0] pmem_q0;
  wire   [7:0] pmem_q1;
  wire   [1:0] pmem_twlb;
  wire   [1:0] wd_twlb;
  wire   [1:0] r_sqlch;
  wire   [3:2] r_ccrx;
  wire   [1:0] r_rxdb_opt;
  wire   [7:4] r_pwrctl;
  wire   [5:0] di_pro;
  wire   [7:0] r_cvctl;
  wire   [7:0] r_srcctl;
  wire   [7:0] r_dpdmctl;
  wire   [11:0] r_fw_pwrv;
  wire   [5:0] r_cvcwr;
  wire   [15:0] r_cvofs;
  wire   [7:0] r_cctrx;
  wire   [7:0] r_ccctl;
  wire   [6:0] r_fcpwr;
  wire   [7:0] fcp_r_dat;
  wire   [7:0] fcp_r_sta;
  wire   [7:0] fcp_r_msk;
  wire   [7:0] fcp_r_ctl;
  wire   [7:0] fcp_r_crc;
  wire   [7:0] fcp_r_acc;
  wire   [7:0] fcp_r_tui;
  wire   [7:0] r_accctl;
  wire   [7:5] r_comp_opt;
  wire   [14:0] sfr_dacwr;
  wire   [17:0] r_dac_en;
  wire   [17:0] r_sar_en;
  wire   [7:0] r_isofs;
  wire   [7:0] r_adofs;
  wire   [7:0] dac_r_ctl;
  wire   [7:0] dac_r_cmpsta;
  wire   [17:0] dac_r_comp;
  wire   [143:0] dac_r_vs;
  wire   [5:0] x_daclsb;
  wire   [6:0] REVID;
  wire   [6:0] r_pu_gpio;
  wire   [6:0] r_pd_gpio;
  wire   [6:0] r_gpio_oe;
  wire   [1:0] r_gpio_ie;
  wire   [55:0] r_regtrm;
  wire   [3:0] r_ana_tm;
  wire   [7:0] i2c_ltbuf;
  wire   [7:0] i2c_lt_ofs;
  wire   [4:0] r_txnumk;
  wire   [1:0] r_auto_gdcrc;
  wire   [1:0] r_spec;
  wire   [1:0] r_dat_spec;
  wire   [6:0] r_txauto;
  wire   [6:0] r_rxords_ena;
  wire   [7:1] r_i2c_deva;
  wire   [2:0] prl_cpmsgid;
  wire   [1:0] pff_ack;
  wire   [7:0] pff_rdat;
  wire   [15:0] pff_rxpart;
  wire   [5:0] pff_ptr;
  wire   [6:0] prx_setsta;
  wire   [1:0] prx_rst;
  wire   [4:0] prx_rcvinf;
  wire   [5:0] prx_adpn;
  wire   [3:0] prx_fsm;
  wire   [2:0] ptx_fsm;
  wire   [3:0] prl_fsm;
  wire   [3:0] slvo_ev;
  wire   [1:0] r_i2cslv_route;
  wire   [5:4] r_i2crout;
  wire   [1:0] r_i2cmcu_route;
  wire   [18:17] upd_dbgpo;
  wire   [7:0] r_dacwdat;
  wire   [17:8] wr_dacv;
  wire   [10:7] r_dacwr;
  wire   [17:0] dacmux_sel;
  wire   [3:0] comp_smpl;
  wire   [7:0] r_cvcwdat;
  wire   [7:0] r_sdischg;
  wire   [7:0] r_vcomp;
  wire   [7:0] r_idacsh;
  wire   [7:0] r_cvofsx;
  wire   [7:0] r_xtm;
  wire   [6:0] bist_r_ctl;
  wire   [1:0] regx_hitbst;
  wire   [7:0] bist_r_dat;
  wire   [1:0] regx_wrpwm;
  wire   [15:0] r_pwm;
  wire   [1:0] r_sap;
  wire   [3:0] lt_gpi;
  wire   [6:0] r_do_ts;
  wire   [3:0] r_dpdo_sel;
  wire   [3:0] r_dndo_sel;
  wire   [4:0] di_aswk;
  wire   [15:8] r_xana;
  wire   [4:0] di_xanav;
  wire   [7:0] r_aopt;
  wire   [6:0] di_gpio;
  wire   [7:6] do_opt;
  wire   [1:0] pwm_o;
  wire   [15:0] d_dodat;
  wire   [3:0] r_lt_gpi;

  CKBUFX1 U0_ASWCLK_BUF_0_ ( .A(aswclk_ps[0]), .Y(aswclk_ps[1]) );
  CKBUFX1 U0_ASWCLK_BUF_1_ ( .A(aswclk_ps[1]), .Y(aswclk_ps[2]) );
  CKBUFX1 U0_ASWCLK_BUF_2_ ( .A(aswclk_ps[2]), .Y(aswclk_ps[3]) );
  CKBUFX1 U0_ASWCLK_BUF_3_ ( .A(aswclk_ps[3]), .Y(aswclk_ps[4]) );
  CKBUFX1 U0_ASWCLK_BUF_4_ ( .A(aswclk_ps[4]), .Y(aswclk_ps[5]) );
  CKBUFX1 U0_ASWCLK_BUF_5_ ( .A(aswclk_ps[5]), .Y(aswclk_ps[6]) );
  CKBUFX1 U0_ASWCLK_BUF_6_ ( .A(aswclk_ps[6]), .Y(aswclk_ps[7]) );
  CKBUFX1 U0_ASWCLK_BUF_7_ ( .A(aswclk_ps[7]), .Y(aswclk_ps[8]) );
  CKBUFX1 U0_ASWCLK_BUF_8_ ( .A(aswclk_ps[8]), .Y(aswclk_ps[9]) );
  CKBUFX1 U0_ASWCLK_BUF_9_ ( .A(aswclk_ps[9]), .Y(aswclk) );
  CKBUFX1 U0_DETCLK_BUF_0_ ( .A(detclk_ps[0]), .Y(detclk_ps[1]) );
  CKBUFX1 U0_DETCLK_BUF_1_ ( .A(detclk_ps[1]), .Y(detclk_ps[2]) );
  CKBUFX1 U0_DETCLK_BUF_2_ ( .A(detclk_ps[2]), .Y(detclk_ps[3]) );
  CKBUFX1 U0_DETCLK_BUF_3_ ( .A(detclk_ps[3]), .Y(detclk_ps[4]) );
  CKBUFX1 U0_DETCLK_BUF_4_ ( .A(detclk_ps[4]), .Y(detclk_ps[5]) );
  CKBUFX1 U0_DETCLK_BUF_5_ ( .A(detclk_ps[5]), .Y(detclk_ps[6]) );
  CKBUFX1 U0_DETCLK_BUF_6_ ( .A(detclk_ps[6]), .Y(detclk_ps[7]) );
  CKBUFX1 U0_DETCLK_BUF_7_ ( .A(detclk_ps[7]), .Y(detclk_ps[8]) );
  CKBUFX1 U0_DETCLK_BUF_8_ ( .A(detclk_ps[8]), .Y(detclk_ps[9]) );
  CKBUFX1 U0_DETCLK_BUF_9_ ( .A(detclk_ps[9]), .Y(detclk) );
  AND2X1 U0_SCAN_EN ( .A(DI_GPIO[2]), .B(n85), .Y(n8) );
  CKMUX2X1 U0_CLK_MUX ( .D0(i_clk), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(s_clk)
         );
  CKMUX2X1 U0_DCLKMUX ( .D0(RD_DET), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        detclk_ps[0]) );
  CKMUX2X1 U0_ACLKMUX ( .D0(aswkup), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        aswclk_ps[0]) );
  CKBUFX1 U0_MCK_BUF ( .A(i_clk), .Y(x_clk) );
  CKBUFX1 U0_TCK_BUF ( .A(DI_GPIO[4]), .Y(t_di_gpio4) );
  CLKDLX1 U0_MCLK_ICG ( .CK(s_clk), .E(n259), .SE(n78), .ECK(g_clk) );
  CLKDLX1 U0_SRAM_ICG ( .CK(g_clk), .E(sram_en), .SE(n86), .ECK(SRAM_CLK) );
  INVX1 U0_REVIDZ_0_ ( .A(1'b1), .Y(REVID[0]) );
  INVX1 U0_REVIDZ_1_ ( .A(1'b1), .Y(REVID[1]) );
  INVX1 U0_REVIDZ_2_ ( .A(1'b1), .Y(REVID[2]) );
  INVX1 U0_REVIDZ_3_ ( .A(1'b1), .Y(REVID[3]) );
  INVX1 U0_REVIDZ_4_ ( .A(1'b0), .Y(REVID[4]) );
  INVX1 U0_REVIDZ_5_ ( .A(1'b0), .Y(REVID[5]) );
  INVX1 U0_REVIDZ_6_ ( .A(1'b1), .Y(REVID[6]) );
  INVX1 U94 ( .A(n53), .Y(n51) );
  INVX1 U104 ( .A(n53), .Y(n52) );
  INVX1 U138 ( .A(srstz), .Y(n53) );
  MUX2X1 U987 ( .D0(n638), .D1(ANA_REGX[0]), .S(n8), .Y(DO_GPIO[6]) );
  MUX2X1 U988 ( .D0(n639), .D1(PMEM_A[15]), .S(n8), .Y(DO_GPIO[5]) );
  AND2X4 U246 ( .A(r_sap[1]), .B(n58), .Y(PMEM_SAP[1]) );
  AND2X4 U247 ( .A(r_sap[0]), .B(n58), .Y(PMEM_SAP[0]) );
  mpb_a0 u0_mpb ( .i_rd({prl_cany0r, n706}), .i_wr({prl_cany0w, i2c_ev_3}), 
        .wdat0(sse_wdat), .wdat1(prx_fifowdat), .addr0(sse_adr), .addr1(
        prl_cany0adr), .r_i2c_attr(r_i2c_attr), .esfrm_oe(esfrm_oe), 
        .esfrm_we(esfrm_we), .sfrack(sfrack), .esfrm_wdat(esfrm_wdat), 
        .esfrm_adr(esfrm_adr), .mcu_esfr_rdat(mcu_esfrrdat), .delay_rdat(
        delay_inst), .delay_rrdy(ictlr_psrack), .esfrm_rrdy(esfrm_rrdy), 
        .esfrm_rdat(esfrm_rdat), .channel_sel(1'b0), .r_pg0_sel(r_pg0_sel), 
        .dma_w(1'b0), .dma_r(1'b0), .dma_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_wdat({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_ack(), .memaddr(memaddr), 
        .memaddr_c({memaddr_c[15:7], n31, n28, memaddr_c[4], n1, n29, 
        memaddr_c[1:0]}), .memwr(memwr), .memrd(memrd), .memrd_c(memrd_c), 
        .cpurst(o_cpurst), .memdatao(memdatao), .memack(memack), .hit_xd(
        hit_xd), .hit_xr(hit_xr), .hit_ps(hit_ps), .hit_ps_c(hit_ps_c), 
        .idat_r(mcu_ram_r), .idat_w(mcu_ram_w), .idat_adr(idat_adr), 
        .idat_wdat(idat_wdat), .iram_ce(iram_ce), .xram_ce(xram_ce), .regx_re(
        regx_re), .iram_we(iram_we), .xram_we(xram_we), .regx_we(regx_we), 
        .iram_a(iram_a), .xram_a(xram_a), .iram_d(iram_d), .xram_d(xram_d), 
        .iram_rdat({n1123, n1120, n1119, n1116, n1118, n1121, sram_rdat}), 
        .xram_rdat({n1123, n1120, n1119, n1116, n1118, n1121, sram_rdat}), 
        .regx_rdat(regx_rdat), .bist_en(n10), .bist_wr(bist_wr), .bist_adr(
        bist_adr), .bist_wdat(bist_wdat), .bist_xram(1'b0), .mclk(g_clk), 
        .srstz(n51), .test_si(n535), .test_so(n132), .test_se(n8) );
  mcu51_a0 u0_mcu ( .bclki2c(r_bclk_sel), .pc_ini({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .slp2wakeup(1'b0), .r_hold_mcu(r_hold_mcu), .wdt_slow(1'b0), .wdtov({n535, 
        SYNOPSYS_UNCONNECTED_1}), .mdubsy(), .cs_run(), .t0_intr(t0_intr), 
        .clki2c(g_clk), .clkmdu(g_clk), .clkur0(g_clk), .clktm0(g_clk), 
        .clktm1(g_clk), .clkwdt(g_clk), .i2c_autoack(1'b0), .i2c_con_ens1(), 
        .clkcpu(g_clk), .clkper(g_clk), .reset(n53), .ro(o_cpurst), .port0i({
        n1110, di_gpio[6:4], n1117, di_gpio[2:0]}), .exint_9(fcp_intr), 
        .exint({exint[7:4], n674, n673, exint[1:0]}), .clkcpuen(), .clkperen(), 
        .port0o({SYNOPSYS_UNCONNECTED_2, do_p0}), .port0ff(ff_p0), .rxd0o(
        do_opt[7]), .txd0(do_opt[6]), .rxd0i(dpdm_urx), .rxd0oe(s0_rxdoe), 
        .scli(n505), .sdai(n507), .sclo(mcuo_scl), .sdao(mcuo_sda), 
        .waitstaten(), .mempsack(mempsack), .memack(memack), .memdatai(
        memdatai), .memdatao(memdatao), .memaddr(memaddr), .mempswr(mempswr), 
        .mempsrd(mempsrd), .memwr(memwr), .memrd(memrd), .memdatao_comb({
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10}), .memaddr_comb(
        memaddr_c), .mempswr_comb(), .mempsrd_comb(mempsrd_c), .memwr_comb(), 
        .memrd_comb(memrd_c), .ramdatai({n1123, n1120, n1119, n1116, n1118, 
        n1121, sram_rdat}), .ramdatao(idat_wdat), .ramaddr(idat_adr), .ramwe(
        mcu_ram_w), .ramoe(mcu_ram_r), .dbgpo({SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, mcu_dbgpo, mcu_pc}), 
        .sfrack(sfrack), .sfrdatai(sfr_rdat), .sfrdatao(sfr_wdat), .sfraddr(
        sfr_adr), .sfrwe(sfr_w), .sfroe(sfr_r), .esfrm_wrdata(esfrm_wdat), 
        .esfrm_addr(esfrm_adr), .esfrm_we(esfrm_we), .esfrm_oe(esfrm_oe), 
        .esfrm_rddata(mcu_esfrrdat), .test_si2(DI_GPIO[1]), .test_si1(n633), 
        .test_so1(n632), .test_se(n8) );
  ictlr_a0 u0_ictlr ( .bkpt_ena(bkpt_ena), .bkpt_pc(bkpt_pc), .memaddr_c({
        memaddr_c[14:7], n31, n28, memaddr_c[4], n1, n29, memaddr_c[1:0]}), 
        .memaddr(memaddr[14:0]), .mcu_psr_c(mempsrd_c), .mcu_psw(mempswr), 
        .hit_ps_c(hit_ps_c), .hit_ps(hit_ps), .mempsack(ictlr_psack), 
        .memdatao(memdatao), .o_set_hold(set_hold), .o_bkp_hold(bkpt_hold), 
        .o_ofs_inc(ictlr_inc), .o_inst(ictlr_inst), .d_inst(delay_inst), 
        .sfr_psrack(ictlr_psrack), .sfr_psofs(r_inst_ofs), .sfr_psr(r_psrd), 
        .sfr_psw(r_pswr), .dw_rst(prl_c0set), .dw_ena(n13), .sfr_wdat({n54, 
        n49, n47, n45, n42, n40, n38, n35}), .pmem_pgm(pmem_pgm), .pmem_re(
        pmem_re), .pmem_csb(pmem_csb), .pmem_clk(pmem_clk), .pmem_a(PMEM_A), 
        .pmem_q0(pmem_q0), .pmem_q1(pmem_q1), .pmem_twlb(pmem_twlb), .wd_twlb(
        wd_twlb), .we_twlb(we_twlb), .pwrdn_rst(pwrdn_rst), .r_pwdn_en(
        r_otp_pwdn_en), .r_multi(r_otp_wpls), .r_hold_mcu(r_hold_mcu), .clk(
        g_clk), .srst(o_cpurst), .test_si3(n632), .test_si2(slvo_sda), 
        .test_si1(n637), .test_so2(n633), .test_so1(n636), .test_se(n8) );
  regbank_a0 u0_regbank ( .srci({di_pro[5], n1108, n1112, n1113, n1111, 
        di_pro[0]}), .dm_fault(di_aswk[3]), .cc1_di(n1122), .cc2_di(n1115), 
        .di_rd_det(n1109), .di_stbovp(di_aswk[1]), .i_tmrf(t0_intr), 
        .i_vcbyval(r_xtm[4]), .dnchk_en(o_dodat5_2_), .r_pwrv_upd(r_pwrv_upd), 
        .aswkup(aswkup), .ps_pwrdn(ps_pwrdn), .r_sleep(r_sleep), .r_pwrdn(
        r_pwrdn), .r_ocdrv_enz(r_ocdrv_enz), .r_osc_stop(r_osc_stop), 
        .r_osc_lo(o_dodat0_15_), .r_osc_gate(r_osc_gate), .r_fw_pwrv(r_fw_pwrv), .r_cvcwr(r_cvcwr[1:0]), .r_cvofs(r_cvofs), .r_otpi_gate(r_otpi_gate), 
        .r_pwrctl(r_pwrctl), .r_pwr_i(DO_PWR_I), .r_cvctl(r_cvctl), .r_srcctl(
        r_srcctl), .r_dpdmctl(r_dpdmctl), .r_ccrx({r_sqlch, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, r_ccrx, r_rxdb_opt}), 
        .r_cctrx(r_cctrx), .r_ccctl(r_ccctl), .r_fcpwr(r_fcpwr), .r_fcpre(
        r_fcpre), .fcp_r_dat(fcp_r_dat), .fcp_r_sta(fcp_r_sta), .fcp_r_msk(
        fcp_r_msk), .fcp_r_ctl(fcp_r_ctl), .fcp_r_crc(fcp_r_crc), .fcp_r_acc(
        fcp_r_acc), .fcp_r_tui(fcp_r_tui), .r_accctl(r_accctl), .r_bclk_sel(
        r_bclk_sel), .r_dacwr(sfr_dacwr), .r_dac_en(r_dac_en[7:0]), .r_sar_en(
        r_sar_en[7:0]), .r_adofs(r_adofs), .r_isofs(r_isofs), .x_daclsb(
        x_daclsb), .r_comp_opt({r_comp_opt, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26}), .dac_r_ctl(
        dac_r_ctl), .dac_r_comp(dac_r_comp[7:0]), .dac_r_cmpsta(dac_r_cmpsta), 
        .dac_r_vs(dac_r_vs[63:0]), .REVID(REVID), .atpg_en(n85), .sfr_r(sfr_r), 
        .sfr_w(sfr_w), .set_hold(set_hold), .bkpt_hold(bkpt_hold), .cpurst(
        o_cpurst), .sfr_addr({1'b1, sfr_adr}), .sfr_wdat({n54, n49, n47, n44, 
        n42, n40, n37, n35}), .sfr_rdat(sfr_rdat), .ff_p0(ff_p0), .di_p0({
        n1110, di_gpio[6:4], n1117, di_gpio[2:0]}), .ictlr_idle(pmem_csb), 
        .ictlr_inc(ictlr_inc), .r_inst_ofs(r_inst_ofs), .r_psrd(r_psrd), 
        .r_pswr(r_pswr), .r_fortxdat(r_fortxdat), .r_fortxrdy(r_fortxrdy), 
        .r_fortxen(r_fortxen), .r_ana_tm(r_ana_tm), .r_gpio_tm(r_gpio_tm), 
        .r_gpio_ie(r_gpio_ie), .r_gpio_oe(r_gpio_oe), .r_gpio_pu(r_pu_gpio), 
        .r_gpio_pd(r_pd_gpio), .r_gpio_s0({N269, N268, N267}), .r_gpio_s1({
        N266, N265, N264}), .r_gpio_s2({N263, N262, N261}), .r_gpio_s3({N260, 
        N259, N258}), .r_regtrm(r_regtrm), .i_pc(mcu_pc), .i_goidle(pid_goidle), .i_gobusy(pid_gobusy), .i_i2c_idle(sse_idle), .bus_idle(bus_idle), 
        .i2c_stretch(hwi2c_stretch), .i_i2c_rwbuf(sse_wdat), .i_i2c_ltbuf(
        i2c_ltbuf), .i_i2c_ofs(i2c_lt_ofs), .o_intr({exint[6], sfr_intr, 
        exint[5:4]}), .r_auto_gdcrc(r_auto_gdcrc), .r_exist1st(r_exist1st), 
        .r_ordrs4(r_ordrs4), .r_fifopsh(r_fifopsh), .r_fifopop(r_fifopop), 
        .r_unlock(r_unlock), .r_first(r_first), .r_last(r_last), .r_fiforst(
        r_fiforst), .r_set_cpmsgid(r_set_cpmsgid), .r_txendk(r_txendk), 
        .r_txnumk(r_txnumk), .r_txshrt(r_txshrt), .r_auto_discard(
        r_auto_discard), .r_hold_mcu(r_hold_mcu), .r_txauto(r_txauto), 
        .r_rxords_ena(r_rxords_ena), .r_spec(r_spec), .r_dat_spec(r_dat_spec), 
        .r_dat_portrole(r_dat_portrole), .r_dat_datarole(r_dat_datarole), 
        .r_discard(r_discard), .r_pshords(r_pshords), .r_pg0_sel(r_pg0_sel), 
        .r_strtch(r_strtch), .r_i2c_attr(r_i2c_attr), .r_i2c_ninc(r_i2c_ninc), 
        .r_hwi2c_en(), .r_i2c_fwnak(r_i2c_fwnak), .r_i2c_fwack(r_i2c_fwack), 
        .r_i2c_deva(r_i2c_deva), .i2c_ev({n706, i2c_ev_6_, slvo_ev[3:2], 
        i2c_ev_3, i2c_ev_2, slvo_ev[1:0]}), .prl_c0set(prl_c0set), .prl_cany0(
        n12), .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), 
        .prl_cpmsgid(prl_cpmsgid), .pff_ack(pff_ack), .prx_rst(prx_rst), 
        .pff_obsd(pff_obsd), .pff_full(pff_full), .pff_empty(pff_empty), 
        .ptx_ack(ptx_ack), .pff_ptr(pff_ptr), .prx_adpn(prx_adpn), .pff_rdat(
        pff_rdat), .pff_rxpart(pff_rxpart), .prx_rcvinf(prx_rcvinf), .ptx_fsm(
        ptx_fsm), .prx_fsm(prx_fsm), .prl_fsm(prl_fsm), .prx_setsta(prx_setsta), .clk_1500k(clk_1500k), .clk_500k(clk_500k), .clk_500(clk_500), .clk(g_clk), 
        .xrstz(i_rstz), .xclk(s_clk), .dbgpo({SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58}), .srstz(srstz), .prstz(prstz), .test_si2(
        r_pwm[15]), .test_si1(n636), .test_so2(n22), .test_so1(n635), 
        .test_se(n8) );
  i2cslv_a0 u0_i2cslv ( .i_sda(n506), .i_scl(n504), .o_sda(slvo_sda), .i_deva(
        r_i2c_deva), .i_inc(n672), .i_fwnak(r_i2c_fwnak), .i_fwack(r_i2c_fwack), .o_we(i2c_ev_3), .o_re(slvo_re), .o_r_early(slvo_early), .o_idle(sse_idle), 
        .o_dec(), .o_busev(slvo_ev), .o_ofs(sse_adr), .o_lt_ofs(i2c_lt_ofs), 
        .o_wdat(sse_wdat), .o_lt_buf(i2c_ltbuf), .o_dbgpo({
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66}), .i_rdat(esfrm_rdat), .i_rd_mem(sse_rdrdy), .i_clk(g_clk), .i_rstz(n52), .i_prefetch(sse_prefetch), 
        .test_si(n634), .test_se(n8) );
  updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 u0_updphy ( .i_cc(di_cc), .i_cc_49(n1114), .i_sqlch(n1107), .r_sqlch(r_sqlch), .r_adprx_en(r_ccrx[3]), .r_adp2nd(
        r_ccrx[2]), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), .r_fifopsh(
        r_fifopsh), .r_fifopop(r_fifopop), .r_fiforst(r_fiforst), .r_unlock(
        r_unlock), .r_first(r_first), .r_last(r_last), .r_set_cpmsgid(
        r_set_cpmsgid), .r_rdy(upd_rdrdy), .r_wdat({n54, n49, n47, n44, n42, 
        n40, n37, n35}), .r_rdat(esfrm_rdat), .r_txnumk(r_txnumk), .r_txendk(
        r_txendk), .r_txshrt(r_txshrt), .r_auto_discard(r_auto_discard), 
        .r_txauto(r_txauto), .r_rxords_ena(r_rxords_ena), .r_spec(r_spec), 
        .r_dat_spec(r_dat_spec), .r_auto_gdcrc(r_auto_gdcrc), .r_rxdb_opt(
        r_rxdb_opt), .r_pshords(r_pshords), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_discard(r_discard), .pid_goidle(
        pid_goidle), .pid_gobusy(pid_gobusy), .pff_ack(pff_ack), .pff_rdat(
        pff_rdat), .pff_rxpart(pff_rxpart), .prx_rcvinf(prx_rcvinf), 
        .pff_obsd(pff_obsd), .pff_ptr(pff_ptr), .pff_empty(pff_empty), 
        .pff_full(pff_full), .ptx_ack(ptx_ack), .ptx_cc(ptx_cc), .ptx_oe(
        ptx_oe), .prx_setsta(prx_setsta), .prx_rst(prx_rst), .prl_c0set(
        prl_c0set), .prl_cany0(prl_cany0), .prl_cany0r(prl_cany0r), 
        .prl_cany0w(prl_cany0w), .prl_discard(prl_discard), .prl_GCTxDone(
        prl_GCTxDone), .prl_cany0adr(prl_cany0adr), .prl_cpmsgid(prl_cpmsgid), 
        .prx_fifowdat(prx_fifowdat), .ptx_fsm(ptx_fsm), .prl_fsm(prl_fsm), 
        .prx_fsm(prx_fsm), .prx_adpn(prx_adpn), .dbgpo({
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, upd_dbgpo, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .clk(g_clk), 
        .srstz(prstz), .test_si(bist_r_ctl[3]), .test_so(n20), .test_se(n8) );
  dacmux_a0 u0_dacmux ( .clk(g_clk), .srstz(n51), .i_comp(n1110), .r_comp_opt(
        r_comp_opt), .r_wdat(r_dacwdat), .r_adofs(r_adofs), .r_isofs(r_isofs), 
        .r_wr({r_dacwr, sfr_dacwr[14:8]}), .dacv_wr({wr_dacv, sfr_dacwr[7:0]}), 
        .o_dacv(dac_r_vs), .o_shrst(sh_rst), .o_hold(sh_hold), .o_dac1(DAC1_V), 
        .o_daci_sel(dacmux_sel), .o_dat(dac_r_comp), .r_dac_en(r_dac_en), 
        .r_sar_en(r_sar_en), .o_dactl(dac_r_ctl), .o_cmpsta(dac_r_cmpsta), 
        .x_daclsb(x_daclsb), .o_intr(exint[7]), .o_smpl({
        SYNOPSYS_UNCONNECTED_97, comp_smpl}), .test_si2(r_vcomp[7]), 
        .test_si1(DI_GPIO[0]), .test_so1(n637), .test_se(n8) );
  fcp_a0 u0_fcp ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(1'b0), .intr(
        fcp_intr), .tx_en(fcp_oe), .tx_dat(fcp_do), .r_dat(fcp_r_dat), .r_sta(
        fcp_r_sta), .r_ctl(fcp_r_ctl), .r_msk(fcp_r_msk), .r_crc(fcp_r_crc), 
        .r_acc(fcp_r_acc), .r_dpdmsta(r_accctl), .r_wdat({n54, n49, n47, n44, 
        n42, n40, n37, n34}), .r_wr(r_fcpwr), .r_re(r_fcpre), .clk(g_clk), 
        .srstz(n52), .r_tui(fcp_r_tui), .test_si(divff_5), .test_so(n634), 
        .test_se(n8) );
  cvctl_a0 u0_cvctl ( .r_cvcwr(r_cvcwr), .wdat(r_cvcwdat), .r_sdischg(
        r_sdischg), .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), .r_cvofsx(r_cvofsx), .r_cvofs(r_cvofs), .sdischg_duty(sdischg_duty), .r_hlsb_en(r_pwrctl[4]), 
        .r_hlsb_sel(r_pwrctl[5]), .r_hlsb_freq(r_xtm[5]), .r_hlsb_duty(
        r_xtm[6]), .r_fw_pwrv(r_fw_pwrv), .r_dac0(DO_DAC0), .r_dac3(DAC3_V), 
        .clk_100k(clk_100k), .clk(g_clk), .srstz(n52), .test_si(d_dodat[15]), 
        .test_se(n8) );
  regx_a0 u0_regx ( .regx_r(regx_re), .regx_w(regx_we), .di_drposc(di_aswk[0]), 
        .di_imposc(di_aswk[4]), .di_rd_det(n1109), .di_stbovp(di_aswk[1]), 
        .clk_500k(clk_500k), .r_imp_osc(r_imp_osc), .regx_addr(xram_a[6:0]), 
        .regx_wdat(xram_d), .regx_rdat(regx_rdat), .regx_hitbst(regx_hitbst), 
        .regx_wrpwm(regx_wrpwm), .regx_wrcvc({r_cvcwr[2], r_cvcwr[5:3]}), 
        .r_sdischg(r_sdischg), .r_bistctl(bist_r_ctl), .r_bistdat(bist_r_dat), 
        .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), .r_cvofsx(r_cvofsx), .r_pwm(
        r_pwm), .regx_wrdac({wr_dacv[17:16], r_dacwr[10:9], wr_dacv[15:8], 
        r_dacwr[8:7]}), .dac_r_vs(dac_r_vs[143:64]), .dac_comp(
        dac_r_comp[17:8]), .r_dac_en(r_dac_en[17:8]), .r_sar_en(r_sar_en[17:8]), .r_aopt(r_aopt), .r_xtm(r_xtm), .r_adummyi(DUMMY_IN), .r_bck0(BCK_REGX[7:0]), 
        .r_bck1(BCK_REGX[15:8]), .r_i2crout({r_i2crout, r_i2cmcu_route, 
        r_i2cslv_route}), .r_xana({r_xana_23, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, r_xana_19, 
        r_xana_18, OCP_SEL, PWREN_HOLD, r_xana, ANA_REGX[7:0]}), .di_xana(
        di_xanav), .lt_gpi(lt_gpi), .di_tst(di_tst), .bkpt_pc(bkpt_pc), 
        .bkpt_ena(bkpt_ena), .we_twlb(we_twlb), .r_vpp_en(r_vpp_en), 
        .r_vpp0v_en(r_vpp0v_en), .r_otp_pwdn_en(r_otp_pwdn_en), .r_otp_wpls(
        r_otp_wpls), .wd_twlb(wd_twlb), .r_sap(r_sap), .r_twlb(pmem_twlb), 
        .upd_pwrv(r_pwrv_upd), .ramacc(ramacc), .sse_idle(sse_idle), 
        .bus_idle(bus_idle), .r_do_ts(r_do_ts), .r_dpdo_sel(r_dpdo_sel), 
        .r_dndo_sel(r_dndo_sel), .di_ts(di_ts), .detclk(detclk), .aswclk(
        aswclk), .atpg_en(n81), .di_aswk({di_aswk[4:3], n1109, di_aswk[1:0]}), 
        .clk(g_clk), .rrstz(srstz), .test_si2(n20), .test_si1(n22), .test_so1(
        n21), .test_se(n8) );
  srambist_a0 u0_srambist ( .clk(g_clk), .srstz(n52), .reg_hit(regx_hitbst), 
        .reg_w(regx_we), .reg_r(regx_re), .reg_wdat(xram_d), .iram_rdat({n1123, 
        n1120, n1119, n1116, n1118, n1121, sram_rdat}), .xram_rdat({n1123, 
        n1120, n1119, n1116, n1118, n1121, sram_rdat}), .bist_en(bist_en), 
        .bist_xram(), .bist_wr(bist_wr), .bist_adr(bist_adr), .bist_wdat(
        bist_wdat), .o_bistctl(bist_r_ctl), .o_bistdat(bist_r_dat), .test_si(
        n21), .test_se(n8) );
  divclk_a0 u0_divclk ( .mclk(g_clk), .srstz(n52), .atpg_en(n78), .clk_1500k(
        clk_1500k), .clk_500k(clk_500k), .clk_100k(clk_100k), .clk_50k(clk_50k), .clk_500(clk_500), .divff_8(divff_8), .divff_5(divff_5), .test_si(
        r_sar_en[17]), .test_se(n8) );
  glpwm_a0_0 u0_pwm_0_ ( .clk(g_clk), .rstz(n52), .clk_base(clk_50k), .we(
        regx_wrpwm[0]), .wdat(xram_d), .r_pwm(r_pwm[7:0]), .pwm_o(pwm_o[0]), 
        .test_si(n132), .test_se(n8) );
  glpwm_a0_1 u0_pwm_1_ ( .clk(g_clk), .rstz(n51), .clk_base(clk_50k), .we(
        regx_wrpwm[1]), .wdat(xram_d), .r_pwm(r_pwm[15:8]), .pwm_o(pwm_o[1]), 
        .test_si(r_pwm[7]), .test_se(n8) );
  SNPS_CLOCK_GATE_HIGH_core_a0 clk_gate_d_dodat_reg ( .CLK(g_clk), .EN(N570), 
        .ENCLK(net8831), .TE(n8) );
  DLNQX1 r_lt_gpi_reg_3_ ( .D(DI_GPIO[0]), .XG(i_rstz), .Q(r_lt_gpi[3]) );
  DLNQX1 r_lt_gpi_reg_2_ ( .D(DI_GPIO[1]), .XG(i_rstz), .Q(r_lt_gpi[2]) );
  DLNQX1 r_lt_gpi_reg_0_ ( .D(DI_GPIO[3]), .XG(i_rstz), .Q(r_lt_gpi[0]) );
  DLNQX1 r_lt_gpi_reg_1_ ( .D(DI_GPIO[2]), .XG(i_rstz), .Q(r_lt_gpi[1]) );
  SDFFQX1 d_dodat_reg_15_ ( .D(N571), .SIN(d_dodat[14]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[15]) );
  SDFFQX1 d_dodat_reg_11_ ( .D(N1483), .SIN(d_dodat[10]), .SMC(n8), .C(net8831), .Q(d_dodat[11]) );
  SDFFQX1 d_dodat_reg_12_ ( .D(N574), .SIN(d_dodat[11]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[12]) );
  SDFFQX1 d_dodat_reg_8_ ( .D(N1498), .SIN(d_dodat[7]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[8]) );
  SDFFQX1 d_dodat_reg_10_ ( .D(N1488), .SIN(d_dodat[9]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[10]) );
  SDFFQX1 d_dodat_reg_9_ ( .D(N1493), .SIN(d_dodat[8]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[9]) );
  SDFFQX1 d_dodat_reg_13_ ( .D(N573), .SIN(d_dodat[12]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[13]) );
  SDFFQX1 d_dodat_reg_14_ ( .D(N572), .SIN(d_dodat[13]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[14]) );
  SDFFQX1 d_dodat_reg_4_ ( .D(N582), .SIN(d_dodat[3]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[4]) );
  SDFFQX1 d_dodat_reg_1_ ( .D(N585), .SIN(d_dodat[0]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[1]) );
  SDFFQX1 d_dodat_reg_0_ ( .D(N586), .SIN(n635), .SMC(n8), .C(net8831), .Q(
        d_dodat[0]) );
  SDFFQX1 d_dodat_reg_3_ ( .D(N583), .SIN(d_dodat[2]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[3]) );
  SDFFQX1 d_dodat_reg_5_ ( .D(N581), .SIN(d_dodat[4]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[5]) );
  SDFFQX1 d_dodat_reg_6_ ( .D(N580), .SIN(d_dodat[5]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[6]) );
  SDFFQX1 d_dodat_reg_2_ ( .D(N584), .SIN(d_dodat[1]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[2]) );
  SDFFQX1 d_dodat_reg_7_ ( .D(N579), .SIN(d_dodat[6]), .SMC(n8), .C(net8831), 
        .Q(d_dodat[7]) );
  MUX4X1 U596 ( .D0(n196), .D1(n207), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N267), 
        .S1(N268), .Y(n117) );
  MUX4X1 U595 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N267), .S1(N268), .Y(n116) );
  MUX2X1 U594 ( .D0(n117), .D1(n116), .S(N269), .Y(DO_GPIO[0]) );
  MUX4X1 U599 ( .D0(n196), .D1(n207), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N264), 
        .S1(N265), .Y(n115) );
  MUX4X1 U598 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N264), .S1(N265), .Y(n114) );
  MUX2X1 U597 ( .D0(n115), .D1(n114), .S(N266), .Y(DO_GPIO[1]) );
  MUX4X1 U587 ( .D0(n196), .D1(n207), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N261), 
        .S1(N262), .Y(n113) );
  MUX4X1 U586 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N261), .S1(N262), .Y(n112) );
  MUX2X1 U585 ( .D0(n113), .D1(n112), .S(N263), .Y(N450) );
  MUX4X1 U584 ( .D0(n196), .D1(n207), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N258), 
        .S1(N259), .Y(n111) );
  MUX4X1 U583 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N258), .S1(N259), .Y(n110) );
  MUX2X1 U582 ( .D0(n111), .D1(n110), .S(N260), .Y(N449) );
  INVX2 U3 ( .A(wr_dacv[11]), .Y(n90) );
  NOR8X1 U4 ( .A(n96), .B(wr_dacv[13]), .C(n95), .D(n94), .E(n93), .F(
        r_dacwr[7]), .G(n92), .H(n91), .Y(n97) );
  AND2X1 U5 ( .A(r_vpp0v_en), .B(ps_pwrdn), .Y(pwrdn_rst) );
  AND2X1 U6 ( .A(n98), .B(n99), .Y(sse_prefetch) );
  BUFX3 U7 ( .A(memaddr_c[2]), .Y(n29) );
  BUFX3 U8 ( .A(memaddr_c[3]), .Y(n1) );
  OA21X1 U9 ( .B(hit_xd), .C(hit_xr), .A(memrd), .Y(n2) );
  NAND2X2 U10 ( .A(pmem_pgm), .B(n59), .Y(n3) );
  INVXL U11 ( .A(n215), .Y(n4) );
  INVX8 U12 ( .A(n3), .Y(PMEM_PGM) );
  INVXL U13 ( .A(n2), .Y(n5) );
  INVXL U14 ( .A(n2), .Y(n6) );
  BUFX3 U15 ( .A(iram_ce), .Y(n7) );
  BUFX3 U16 ( .A(xram_ce), .Y(n9) );
  BUFX3 U17 ( .A(bist_en), .Y(n10) );
  INVX1 U18 ( .A(prl_cany0), .Y(n11) );
  INVX1 U19 ( .A(n11), .Y(n12) );
  INVX1 U20 ( .A(n11), .Y(n13) );
  BUFX3 U21 ( .A(n1096), .Y(n14) );
  INVXL U22 ( .A(n86), .Y(n59) );
  OR2X2 U23 ( .A(wr_dacv[10]), .B(wr_dacv[9]), .Y(n91) );
  OR2X2 U24 ( .A(wr_dacv[15]), .B(wr_dacv[14]), .Y(n96) );
  INVX1 U25 ( .A(memaddr_c[6]), .Y(n30) );
  MUX2XL U26 ( .D0(xram_d[2]), .D1(sfr_wdat[2]), .S(n33), .Y(r_dacwdat[2]) );
  MUX2XL U27 ( .D0(xram_d[1]), .D1(n38), .S(n33), .Y(r_dacwdat[1]) );
  AO22XL U28 ( .A(iram_a[3]), .B(iram_ce), .C(xram_a[3]), .D(xram_ce), .Y(
        SRAM_A[3]) );
  INVX1 U29 ( .A(fcp_oe), .Y(n228) );
  NAND21X1 U30 ( .B(r_cvctl[0]), .A(n56), .Y(DO_CVCTL[0]) );
  NAND21X1 U31 ( .B(r_cvctl[1]), .A(n56), .Y(DO_CVCTL[1]) );
  AND2X1 U32 ( .A(r_srcctl[7]), .B(n61), .Y(DO_SRCCTL[7]) );
  AND2X1 U33 ( .A(r_ccctl[1]), .B(n64), .Y(DO_CCCTL[1]) );
  AND2X1 U34 ( .A(r_ccctl[3]), .B(n64), .Y(DO_CCCTL[3]) );
  AND2X1 U35 ( .A(r_srcctl[6]), .B(n61), .Y(DO_SRCCTL[6]) );
  AND2X1 U36 ( .A(r_xana[12]), .B(n65), .Y(ANA_REGX[12]) );
  AND2X1 U37 ( .A(r_aopt[1]), .B(n57), .Y(ANAOPT[1]) );
  AND2X1 U38 ( .A(r_aopt[4]), .B(n66), .Y(ANAOPT[4]) );
  AND2X1 U39 ( .A(r_xana[8]), .B(n65), .Y(ANA_REGX[8]) );
  AND2X1 U40 ( .A(r_xana[9]), .B(n65), .Y(ANA_REGX[9]) );
  AND2X1 U41 ( .A(r_ccctl[2]), .B(n64), .Y(DO_CCCTL[2]) );
  AND2X1 U42 ( .A(r_cvctl[3]), .B(n63), .Y(DO_CVCTL[3]) );
  AND2X1 U43 ( .A(r_cvctl[4]), .B(n62), .Y(DO_CVCTL[4]) );
  OR2X1 U44 ( .A(wr_dacv[8]), .B(r_dacwr[8]), .Y(n93) );
  INVX1 U45 ( .A(n97), .Y(n32) );
  NAND21X1 U46 ( .B(wr_dacv[12]), .A(n90), .Y(n92) );
  NAND21X1 U47 ( .B(wr_dacv[17]), .A(n89), .Y(n95) );
  INVX1 U48 ( .A(wr_dacv[16]), .Y(n89) );
  INVX1 U49 ( .A(n43), .Y(n42) );
  NAND21X1 U50 ( .B(n182), .A(n56), .Y(SRAM_CEB) );
  NOR3XL U51 ( .A(r_cvcwr[4]), .B(r_cvcwr[3]), .C(r_cvcwr[5]), .Y(n16) );
  INVX1 U52 ( .A(n36), .Y(n35) );
  INVX1 U53 ( .A(n41), .Y(n40) );
  INVX1 U54 ( .A(n46), .Y(n44) );
  INVX1 U55 ( .A(n55), .Y(n54) );
  INVX1 U56 ( .A(n50), .Y(n49) );
  INVX1 U57 ( .A(n48), .Y(n47) );
  INVX1 U58 ( .A(n39), .Y(n37) );
  INVX1 U59 ( .A(n39), .Y(n38) );
  INVX1 U60 ( .A(n46), .Y(n45) );
  INVX1 U61 ( .A(n36), .Y(n34) );
  INVX1 U62 ( .A(n903), .Y(n188) );
  INVX1 U63 ( .A(n1092), .Y(n101) );
  INVX1 U64 ( .A(n927), .Y(n118) );
  INVX1 U65 ( .A(n905), .Y(n108) );
  INVX1 U66 ( .A(n85), .Y(n56) );
  INVX1 U67 ( .A(n85), .Y(n57) );
  INVX1 U68 ( .A(atpg_en), .Y(n71) );
  INVX1 U69 ( .A(n81), .Y(n70) );
  INVX1 U70 ( .A(n83), .Y(n68) );
  INVX1 U71 ( .A(n80), .Y(n69) );
  INVX1 U72 ( .A(n86), .Y(n60) );
  INVX1 U73 ( .A(n86), .Y(n58) );
  INVX1 U74 ( .A(n85), .Y(n67) );
  INVX1 U75 ( .A(n86), .Y(n66) );
  INVX1 U76 ( .A(n78), .Y(n65) );
  INVX1 U77 ( .A(n86), .Y(n64) );
  INVX1 U78 ( .A(n78), .Y(n63) );
  INVX1 U79 ( .A(n86), .Y(n62) );
  INVX1 U80 ( .A(n86), .Y(n61) );
  INVX1 U81 ( .A(n81), .Y(n72) );
  INVX1 U82 ( .A(atpg_en), .Y(n75) );
  INVX1 U83 ( .A(n80), .Y(n77) );
  INVX1 U84 ( .A(n84), .Y(n76) );
  INVX1 U85 ( .A(n83), .Y(n74) );
  INVX1 U86 ( .A(n85), .Y(n73) );
  OR2X1 U87 ( .A(r_dacwr[10]), .B(r_dacwr[9]), .Y(n94) );
  INVX1 U88 ( .A(sfr_wdat[3]), .Y(n43) );
  INVX1 U89 ( .A(SRAM_A[4]), .Y(n178) );
  INVX1 U90 ( .A(sram_en), .Y(n182) );
  INVX1 U91 ( .A(n849), .Y(SRAM_D[7]) );
  INVX1 U92 ( .A(sfr_wdat[0]), .Y(n36) );
  INVX1 U93 ( .A(n850), .Y(SRAM_D[0]) );
  INVX1 U95 ( .A(sfr_wdat[4]), .Y(n46) );
  INVX1 U96 ( .A(sfr_wdat[6]), .Y(n50) );
  INVX1 U97 ( .A(sfr_wdat[7]), .Y(n55) );
  INVX1 U98 ( .A(sfr_wdat[5]), .Y(n48) );
  INVX1 U99 ( .A(sfr_wdat[2]), .Y(n41) );
  INVX1 U100 ( .A(sfr_wdat[1]), .Y(n39) );
  OR2X1 U101 ( .A(iram_we), .B(xram_we), .Y(n963) );
  OAI21X1 U102 ( .B(xram_we), .C(iram_we), .A(n72), .Y(SRAM_WEB) );
  OR2X1 U103 ( .A(n924), .B(n929), .Y(n905) );
  OR2X1 U105 ( .A(n907), .B(n905), .Y(n1092) );
  NAND42X1 U106 ( .C(n911), .D(n908), .A(n1094), .B(n257), .Y(n991) );
  NOR4XL U107 ( .A(n1092), .B(n927), .C(n1086), .D(n188), .Y(n1094) );
  INVX1 U108 ( .A(n125), .Y(n186) );
  NAND21X1 U109 ( .B(n991), .A(n950), .Y(n125) );
  NAND42X1 U110 ( .C(n912), .D(n910), .A(n255), .B(n256), .Y(n1086) );
  XOR2X1 U111 ( .A(DO_DAC0[0]), .B(DAC3_V[5]), .Y(n165) );
  NOR2X1 U112 ( .A(n923), .B(n926), .Y(n903) );
  OR2X1 U113 ( .A(n913), .B(n899), .Y(n927) );
  INVX1 U114 ( .A(n972), .Y(n196) );
  INVX1 U115 ( .A(n1076), .Y(n255) );
  INVX1 U116 ( .A(n1079), .Y(n256) );
  NAND2X1 U117 ( .A(n950), .B(n991), .Y(n119) );
  INVX1 U118 ( .A(n906), .Y(n257) );
  OR3XL U119 ( .A(n926), .B(n899), .C(n1086), .Y(n1093) );
  OR2X1 U120 ( .A(n912), .B(n927), .Y(n1077) );
  AOI21BBXL U121 ( .B(n907), .C(n924), .A(n261), .Y(n1078) );
  INVX1 U122 ( .A(s0_rxdoe), .Y(n258) );
  INVX1 U123 ( .A(n911), .Y(n104) );
  NOR2X1 U124 ( .A(n209), .B(n205), .Y(n1000) );
  INVX1 U125 ( .A(n88), .Y(n86) );
  INVX1 U126 ( .A(n87), .Y(n85) );
  INVX1 U127 ( .A(n88), .Y(n82) );
  INVX1 U128 ( .A(n88), .Y(n81) );
  INVX1 U129 ( .A(n88), .Y(n83) );
  INVX1 U130 ( .A(n88), .Y(n84) );
  INVX1 U131 ( .A(n88), .Y(n79) );
  INVX1 U132 ( .A(n88), .Y(n80) );
  AOI21X1 U133 ( .B(n210), .C(n204), .A(n86), .Y(CCI2C_EN) );
  NAND2X1 U134 ( .A(n254), .B(n56), .Y(OCDRV_ENZ) );
  NAND2X1 U135 ( .A(n229), .B(n56), .Y(SH_HOLD) );
  NOR2X1 U136 ( .A(n83), .B(n191), .Y(OSC_LOW) );
  MUX2X2 U137 ( .D0(n35), .D1(xram_d[0]), .S(n32), .Y(r_dacwdat[0]) );
  MUX2BXL U139 ( .D0(xram_d[5]), .D1(n48), .S(n33), .Y(r_dacwdat[5]) );
  MUX2BXL U140 ( .D0(xram_d[6]), .D1(n50), .S(n33), .Y(r_dacwdat[6]) );
  MUX2X1 U141 ( .D0(xram_d[4]), .D1(n45), .S(n33), .Y(r_dacwdat[4]) );
  MUX2BXL U142 ( .D0(xram_d[7]), .D1(n55), .S(n33), .Y(r_dacwdat[7]) );
  MUX2BXL U143 ( .D0(xram_d[3]), .D1(n43), .S(n33), .Y(r_dacwdat[3]) );
  NAND32X1 U144 ( .B(n1091), .C(n106), .A(n105), .Y(DO_GPIO[2]) );
  AO22X1 U145 ( .A(n906), .B(n1122), .C(n923), .D(di_pro[5]), .Y(n1091) );
  OA22X1 U146 ( .A(n104), .B(n103), .C(n102), .D(n101), .Y(n105) );
  AO2222XL U147 ( .A(N450), .B(n119), .C(n908), .D(n100), .E(mcu_dbgpo[20]), 
        .F(n1093), .G(r_osc_stop), .H(n913), .Y(n106) );
  NOR2X1 U148 ( .A(n82), .B(n937), .Y(DO_TS[3]) );
  OAI2B11X1 U149 ( .D(regx_rdat[7]), .C(n814), .A(n815), .B(n816), .Y(
        memdatai[7]) );
  AOI22X1 U150 ( .A(n817), .B(n1123), .C(ictlr_inst[7]), .D(n6), .Y(n816) );
  XNOR2XL U151 ( .A(n986), .B(n987), .Y(N1483) );
  XNOR2XL U152 ( .A(DO_DAC0[6]), .B(n988), .Y(n987) );
  XNOR2XL U153 ( .A(n989), .B(n860), .Y(n986) );
  XNOR2XL U154 ( .A(n199), .B(dacmux_sel[11]), .Y(n988) );
  XNOR2XL U155 ( .A(DAC1_V[5]), .B(n849), .Y(n989) );
  AOI22X1 U156 ( .A(xram_d[7]), .B(xram_we), .C(iram_we), .D(iram_d[7]), .Y(
        n849) );
  OR2X1 U157 ( .A(slvo_early), .B(slvo_re), .Y(n706) );
  OAI2B11X1 U158 ( .D(regx_rdat[4]), .C(n814), .A(n815), .B(n821), .Y(
        memdatai[4]) );
  AOI22X1 U159 ( .A(n817), .B(n1116), .C(ictlr_inst[4]), .D(n6), .Y(n821) );
  OAI2B11X1 U160 ( .D(regx_rdat[2]), .C(n814), .A(n815), .B(n823), .Y(
        memdatai[2]) );
  AOI22X1 U161 ( .A(n817), .B(n1121), .C(ictlr_inst[2]), .D(n5), .Y(n823) );
  OAI2B11X1 U162 ( .D(regx_rdat[5]), .C(n814), .A(n815), .B(n820), .Y(
        memdatai[5]) );
  AOI22X1 U163 ( .A(n817), .B(n1119), .C(ictlr_inst[5]), .D(n5), .Y(n820) );
  OAI2B11X1 U164 ( .D(regx_rdat[1]), .C(n814), .A(n815), .B(n824), .Y(
        memdatai[1]) );
  AOI22X1 U165 ( .A(n817), .B(sram_rdat[1]), .C(ictlr_inst[1]), .D(n6), .Y(
        n824) );
  OR2X1 U166 ( .A(iram_ce), .B(xram_ce), .Y(sram_en) );
  AO22XL U167 ( .A(iram_a[4]), .B(iram_ce), .C(xram_a[4]), .D(xram_ce), .Y(
        SRAM_A[4]) );
  XOR2X1 U168 ( .A(n147), .B(n146), .Y(N579) );
  XNOR3X1 U169 ( .A(n145), .B(n144), .C(n143), .Y(n147) );
  XOR3X1 U170 ( .A(SRAM_A[7]), .B(SRAM_D[3]), .C(n937), .Y(n146) );
  INVX1 U171 ( .A(DAC1_V[1]), .Y(n144) );
  XNOR3X1 U172 ( .A(n17), .B(n18), .C(SRAM_A[9]), .Y(N1493) );
  XNOR3X1 U173 ( .A(DO_DAC0[4]), .B(dacmux_sel[9]), .C(DAC1_V[3]), .Y(n17) );
  XNOR2XL U174 ( .A(SRAM_D[5]), .B(n862), .Y(n18) );
  XNOR3X1 U175 ( .A(n19), .B(n23), .C(n861), .Y(N1488) );
  XNOR3X1 U176 ( .A(DO_DAC0[5]), .B(dacmux_sel[10]), .C(DAC1_V[4]), .Y(n19) );
  XNOR2XL U177 ( .A(SRAM_D[6]), .B(SRAM_A[10]), .Y(n23) );
  XNOR3X1 U178 ( .A(n24), .B(n25), .C(SRAM_A[8]), .Y(N1498) );
  XNOR3X1 U179 ( .A(DO_DAC0[3]), .B(dacmux_sel[8]), .C(DAC1_V[2]), .Y(n24) );
  XNOR2XL U180 ( .A(SRAM_D[4]), .B(n863), .Y(n25) );
  OAI2B11X1 U181 ( .D(regx_rdat[3]), .C(n814), .A(n815), .B(n822), .Y(
        memdatai[3]) );
  AOI22X1 U182 ( .A(n817), .B(n1118), .C(ictlr_inst[3]), .D(n5), .Y(n822) );
  AO22XL U183 ( .A(iram_a[0]), .B(iram_ce), .C(xram_a[0]), .D(xram_ce), .Y(
        SRAM_A[0]) );
  AO22XL U184 ( .A(iram_a[1]), .B(iram_ce), .C(xram_a[1]), .D(xram_ce), .Y(
        SRAM_A[1]) );
  AO22XL U185 ( .A(iram_a[2]), .B(iram_ce), .C(xram_a[2]), .D(xram_ce), .Y(
        SRAM_A[2]) );
  AO22XL U186 ( .A(iram_a[5]), .B(iram_ce), .C(xram_a[5]), .D(xram_ce), .Y(
        SRAM_A[5]) );
  XOR2X1 U187 ( .A(n149), .B(n148), .Y(N584) );
  XOR3X1 U188 ( .A(DAC3_V[2]), .B(dacmux_sel[2]), .C(DO_PWR_I[2]), .Y(n149) );
  XOR3X1 U189 ( .A(o_dodat5_2_), .B(SRAM_A[2]), .C(DO_GPIO[2]), .Y(n148) );
  XOR2X1 U190 ( .A(n157), .B(n156), .Y(N580) );
  XNOR3X1 U191 ( .A(n155), .B(dacmux_sel[6]), .C(n154), .Y(n156) );
  XOR3X1 U192 ( .A(SRAM_A[6]), .B(SRAM_D[2]), .C(n638), .Y(n157) );
  INVX1 U193 ( .A(DAC1_V[0]), .Y(n154) );
  XOR2X1 U194 ( .A(n167), .B(n166), .Y(N581) );
  XNOR3X1 U195 ( .A(n165), .B(n164), .C(n163), .Y(n167) );
  XOR3X1 U196 ( .A(SRAM_D[1]), .B(SRAM_A[5]), .C(n639), .Y(n166) );
  INVX1 U197 ( .A(DO_PWR_I[5]), .Y(n164) );
  XOR2X1 U198 ( .A(n169), .B(n168), .Y(N583) );
  XOR3X1 U199 ( .A(DAC3_V[3]), .B(dacmux_sel[3]), .C(DO_PWR_I[3]), .Y(n168) );
  XOR3X1 U200 ( .A(CC1_DOB), .B(DO_GPIO[3]), .C(SRAM_A[3]), .Y(n169) );
  XOR2X1 U201 ( .A(n172), .B(n171), .Y(N586) );
  XOR3X1 U202 ( .A(dacmux_sel[16]), .B(DO_PWR_I[0]), .C(n170), .Y(n171) );
  XOR3X1 U203 ( .A(dacmux_sel[0]), .B(n227), .C(SRAM_A[0]), .Y(n172) );
  XOR2X1 U204 ( .A(DAC3_V[0]), .B(DO_GPIO[0]), .Y(n170) );
  XOR2X1 U205 ( .A(n176), .B(n175), .Y(N585) );
  XOR3X1 U206 ( .A(dacmux_sel[17]), .B(DO_PWR_I[1]), .C(n174), .Y(n175) );
  XOR3X1 U207 ( .A(dacmux_sel[1]), .B(n173), .C(SRAM_A[1]), .Y(n176) );
  XOR2X1 U208 ( .A(DAC3_V[1]), .B(DO_GPIO[1]), .Y(n174) );
  XOR2X1 U209 ( .A(n180), .B(n179), .Y(N582) );
  XOR3X1 U210 ( .A(DO_PWR_I[4]), .B(DAC3_V[4]), .C(n177), .Y(n180) );
  XOR3X1 U211 ( .A(dacmux_sel[4]), .B(n26), .C(n178), .Y(n179) );
  XOR2X1 U212 ( .A(DO_GPIO[4]), .B(n850), .Y(n177) );
  XOR2X1 U213 ( .A(n185), .B(n184), .Y(N572) );
  XOR3X1 U214 ( .A(dacmux_sel[14]), .B(DAC1_V[8]), .C(n181), .Y(n185) );
  XOR3X1 U215 ( .A(n183), .B(n182), .C(n857), .Y(n184) );
  XOR2X1 U216 ( .A(DO_DAC0[9]), .B(TX_EN), .Y(n181) );
  OAI2B11X1 U217 ( .D(regx_rdat[0]), .C(n814), .A(n815), .B(n825), .Y(
        memdatai[0]) );
  AOI22X1 U218 ( .A(n817), .B(sram_rdat[0]), .C(ictlr_inst[0]), .D(n6), .Y(
        n825) );
  AO22X1 U219 ( .A(iram_d[6]), .B(iram_we), .C(xram_d[6]), .D(xram_we), .Y(
        SRAM_D[6]) );
  AO22X1 U220 ( .A(iram_d[5]), .B(iram_we), .C(xram_d[5]), .D(xram_we), .Y(
        SRAM_D[5]) );
  OAI2B11X1 U221 ( .D(regx_rdat[6]), .C(n814), .A(n815), .B(n819), .Y(
        memdatai[6]) );
  AOI22X1 U222 ( .A(n817), .B(n1120), .C(ictlr_inst[6]), .D(n5), .Y(n819) );
  MUX2X1 U223 ( .D0(xram_d[7]), .D1(n54), .S(n16), .Y(r_cvcwdat[7]) );
  MUX2X1 U224 ( .D0(xram_d[2]), .D1(n40), .S(n16), .Y(r_cvcwdat[2]) );
  MUX2X1 U225 ( .D0(xram_d[5]), .D1(n47), .S(n16), .Y(r_cvcwdat[5]) );
  MUX2X1 U226 ( .D0(xram_d[1]), .D1(n38), .S(n16), .Y(r_cvcwdat[1]) );
  MUX2X1 U227 ( .D0(xram_d[0]), .D1(n35), .S(n16), .Y(r_cvcwdat[0]) );
  MUX2X1 U228 ( .D0(xram_d[3]), .D1(n42), .S(n16), .Y(r_cvcwdat[3]) );
  MUX2X1 U229 ( .D0(xram_d[4]), .D1(n45), .S(n16), .Y(r_cvcwdat[4]) );
  MUX2X1 U230 ( .D0(xram_d[6]), .D1(n49), .S(n16), .Y(r_cvcwdat[6]) );
  AO22X1 U231 ( .A(iram_d[4]), .B(iram_we), .C(xram_d[4]), .D(xram_we), .Y(
        SRAM_D[4]) );
  AO22X1 U232 ( .A(iram_d[3]), .B(iram_we), .C(xram_d[3]), .D(xram_we), .Y(
        SRAM_D[3]) );
  AO22X1 U233 ( .A(iram_d[2]), .B(iram_we), .C(xram_d[2]), .D(xram_we), .Y(
        SRAM_D[2]) );
  NAND21X1 U234 ( .B(n5), .A(hit_xr), .Y(n814) );
  XNOR2XL U235 ( .A(n938), .B(n939), .Y(N574) );
  XNOR2XL U236 ( .A(DO_DAC0[7]), .B(n940), .Y(n939) );
  XNOR2XL U237 ( .A(n941), .B(n942), .Y(n938) );
  XNOR2XL U238 ( .A(r_xana_19), .B(n232), .Y(n940) );
  AOI22X1 U239 ( .A(xram_d[0]), .B(xram_we), .C(iram_d[0]), .D(iram_we), .Y(
        n850) );
  AO22X1 U240 ( .A(iram_d[1]), .B(iram_we), .C(xram_d[1]), .D(xram_we), .Y(
        SRAM_D[1]) );
  NOR2X1 U241 ( .A(n5), .B(hit_xr), .Y(n817) );
  AOI221XL U242 ( .A(n1047), .B(r_osc_stop), .C(r_ocdrv_enz), .D(n1045), .E(
        n1059), .Y(n1058) );
  OAI22X1 U243 ( .A(n198), .B(n219), .C(n259), .D(n218), .Y(n1059) );
  XNOR2XL U244 ( .A(DO_DAC0[8]), .B(n230), .Y(n946) );
  XNOR2XL U245 ( .A(o_dodat0_15_), .B(dacmux_sel[15]), .Y(n961) );
  XNOR2XL U248 ( .A(n944), .B(n945), .Y(N573) );
  XNOR2XL U249 ( .A(n947), .B(n948), .Y(n944) );
  XNOR2XL U250 ( .A(DAC1_V[7]), .B(n946), .Y(n945) );
  XNOR2XL U251 ( .A(n949), .B(n858), .Y(n947) );
  XNOR2XL U252 ( .A(n958), .B(n959), .Y(N571) );
  XNOR2XL U253 ( .A(n962), .B(n963), .Y(n958) );
  XNOR2XL U254 ( .A(n960), .B(n961), .Y(n959) );
  XNOR2XL U255 ( .A(n964), .B(n904), .Y(n962) );
  INVX1 U256 ( .A(dacmux_sel[7]), .Y(n143) );
  INVX1 U257 ( .A(dacmux_sel[5]), .Y(n163) );
  NOR2X1 U258 ( .A(n237), .B(n229), .Y(N570) );
  OAI31XL U259 ( .A(n1099), .B(n1103), .C(n1096), .D(n774), .Y(n924) );
  OAI31XL U260 ( .A(n1098), .B(n1103), .C(n1096), .D(n775), .Y(n929) );
  INVX1 U261 ( .A(pwm_o[1]), .Y(n197) );
  OAI31XL U262 ( .A(n1100), .B(n14), .C(n1099), .D(n781), .Y(n911) );
  OAI22X1 U263 ( .A(n212), .B(n995), .C(mcuo_scl), .D(n208), .Y(n972) );
  OAI31XL U264 ( .A(n1101), .B(n1096), .C(n1100), .D(n783), .Y(n1076) );
  OAI31XL U265 ( .A(n1097), .B(n1096), .C(n1100), .D(n784), .Y(n1079) );
  OAI31XL U266 ( .A(n1097), .B(n1096), .C(n1102), .D(n780), .Y(n908) );
  OAI32X1 U267 ( .A(n1102), .B(n14), .C(n1098), .D(n72), .E(n266), .Y(n899) );
  OAI31XL U268 ( .A(n1095), .B(n1096), .C(n1098), .D(n771), .Y(n926) );
  OAI31XL U269 ( .A(n1101), .B(n14), .C(n1095), .D(n772), .Y(n907) );
  OAI31XL U270 ( .A(n1099), .B(n1096), .C(n1102), .D(n778), .Y(n912) );
  OAI31XL U271 ( .A(n1095), .B(n1096), .C(n1099), .D(n770), .Y(n923) );
  OAI31XL U272 ( .A(n1101), .B(n1096), .C(n1102), .D(n779), .Y(n910) );
  OAI31XL U273 ( .A(n1100), .B(n14), .C(n1098), .D(n782), .Y(n913) );
  OAI31XL U274 ( .A(n1095), .B(n14), .C(n1097), .D(n773), .Y(n906) );
  NOR2X1 U275 ( .A(n81), .B(n860), .Y(OE_GPIO[3]) );
  NOR2X1 U276 ( .A(n81), .B(n861), .Y(OE_GPIO[2]) );
  NOR2X1 U277 ( .A(n81), .B(n859), .Y(OE_GPIO[4]) );
  NOR2X1 U278 ( .A(n83), .B(n862), .Y(OE_GPIO[1]) );
  NOR2X1 U279 ( .A(n83), .B(n863), .Y(OE_GPIO[0]) );
  NAND2X1 U280 ( .A(n858), .B(n57), .Y(OE_GPIO[5]) );
  NAND2X1 U281 ( .A(n857), .B(n56), .Y(OE_GPIO[6]) );
  AO22X1 U282 ( .A(n929), .B(di_cc), .C(n1110), .D(n907), .Y(n928) );
  OAI22X1 U283 ( .A(n255), .B(n192), .C(n256), .D(n239), .Y(n930) );
  OAI22X1 U284 ( .A(n260), .B(n903), .C(n256), .D(n904), .Y(n902) );
  NOR3XL U285 ( .A(n788), .B(n792), .C(n261), .Y(di_cc) );
  INVX1 U286 ( .A(n1114), .Y(n261) );
  ENOX1 U287 ( .A(n257), .B(n904), .C(n1108), .D(n926), .Y(n925) );
  INVX1 U288 ( .A(n973), .Y(n207) );
  INVX1 U289 ( .A(di_gpio[2]), .Y(n190) );
  INVX1 U290 ( .A(n791), .Y(n212) );
  INVX1 U291 ( .A(n786), .Y(n208) );
  AOI222XL U292 ( .A(n786), .B(n803), .C(n788), .D(n804), .E(n205), .F(n805), 
        .Y(n505) );
  AOI222XL U293 ( .A(n786), .B(n787), .C(n788), .D(n789), .E(n205), .F(n790), 
        .Y(n507) );
  OAI22AX1 U294 ( .D(n806), .C(n807), .A(di_gpio[0]), .B(n806), .Y(n803) );
  NAND2X1 U295 ( .A(n802), .B(n252), .Y(n806) );
  EORX1 U296 ( .A(n808), .B(n809), .C(n809), .D(di_gpio[1]), .Y(n807) );
  NAND2X1 U297 ( .A(n797), .B(n253), .Y(n809) );
  AOI222XL U298 ( .A(n791), .B(n787), .C(n792), .D(n789), .E(n209), .F(n790), 
        .Y(n506) );
  AOI222XL U299 ( .A(n791), .B(n803), .C(n792), .D(n804), .E(n209), .F(n805), 
        .Y(n504) );
  NOR2X1 U300 ( .A(n201), .B(n202), .Y(n1067) );
  INVX1 U301 ( .A(di_gpio[0]), .Y(n195) );
  INVX1 U302 ( .A(n1113), .Y(n260) );
  INVX1 U303 ( .A(n955), .Y(n187) );
  XOR2X1 U304 ( .A(DO_PWR_I[7]), .B(DO_DAC0[2]), .Y(n145) );
  XOR2X1 U305 ( .A(DO_PWR_I[6]), .B(DO_DAC0[1]), .Y(n155) );
  INVX1 U306 ( .A(n1110), .Y(n103) );
  INVX1 U307 ( .A(n1107), .Y(n102) );
  INVX1 U308 ( .A(n1068), .Y(n130) );
  XNOR2XL U309 ( .A(DO_DAC0[10]), .B(DAC1_V[9]), .Y(n960) );
  XOR2X1 U310 ( .A(DAC1_V[6]), .B(n859), .Y(n941) );
  INVX1 U311 ( .A(n957), .Y(n183) );
  OAI22X1 U312 ( .A(n197), .B(n219), .C(n218), .D(n245), .Y(n1051) );
  OAI22X1 U313 ( .A(n198), .B(n221), .C(n191), .D(n1013), .Y(n1012) );
  OAI22X1 U314 ( .A(n995), .B(n210), .C(mcuo_scl), .D(n204), .Y(n123) );
  AND2X1 U315 ( .A(n706), .B(n99), .Y(i2c_ev_6_) );
  INVX1 U316 ( .A(n26), .Y(CC2_DOB) );
  INVX1 U317 ( .A(n200), .Y(o_dodat5_2_) );
  OAI22X1 U318 ( .A(n995), .B(n1031), .C(mcuo_scl), .D(n1032), .Y(n999) );
  AOI222XL U319 ( .A(n1015), .B(r_xana_19), .C(n223), .D(di_aswk[0]), .E(n222), 
        .F(di_aswk[4]), .Y(n1017) );
  AOI222XL U320 ( .A(n1046), .B(n187), .C(n1047), .D(n1107), .E(n1045), .F(
        n1122), .Y(n1056) );
  INVX1 U321 ( .A(n904), .Y(TX_DAT) );
  AOI221XL U322 ( .A(n222), .B(o_dodat5_2_), .C(n1015), .D(n227), .E(n1018), 
        .Y(n1016) );
  OAI22AX1 U323 ( .D(n1011), .C(n875), .A(n1019), .B(n241), .Y(n1018) );
  AOI221XL U324 ( .A(n222), .B(n1112), .C(n1015), .D(di_pro[0]), .E(n1027), 
        .Y(n1026) );
  ENOX1 U325 ( .A(n260), .B(n1019), .C(n1111), .D(n1011), .Y(n1027) );
  INVX1 U326 ( .A(n1013), .Y(n222) );
  INVX1 U327 ( .A(n1019), .Y(n223) );
  INVX1 U328 ( .A(o_dodat0_15_), .Y(n191) );
  INVX1 U329 ( .A(n1036), .Y(n219) );
  INVX1 U330 ( .A(n1046), .Y(n218) );
  INVX1 U331 ( .A(n788), .Y(n204) );
  INVX1 U332 ( .A(n792), .Y(n210) );
  INVX1 U333 ( .A(n1015), .Y(n221) );
  NOR2X1 U334 ( .A(n225), .B(n217), .Y(n1045) );
  AOI222XL U335 ( .A(n1015), .B(n1108), .C(n1011), .D(di_pro[5]), .E(n222), 
        .F(di_aswk[3]), .Y(n1025) );
  INVX1 U336 ( .A(n869), .Y(n227) );
  INVX1 U337 ( .A(r_ocdrv_enz), .Y(n254) );
  INVX1 U338 ( .A(n949), .Y(n203) );
  INVX1 U339 ( .A(n1032), .Y(n205) );
  INVX1 U340 ( .A(n1031), .Y(n209) );
  NOR2X1 U341 ( .A(n955), .B(n82), .Y(TX_EN) );
  INVX1 U342 ( .A(n848), .Y(n246) );
  INVX1 U343 ( .A(n875), .Y(n173) );
  INVX1 U344 ( .A(sh_hold), .Y(n229) );
  NAND2X1 U345 ( .A(n761), .B(n931), .Y(n950) );
  NOR21XL U346 ( .B(r_pwrdn), .A(n81), .Y(PWRDN) );
  NOR21XL U347 ( .B(dacmux_sel[11]), .A(n78), .Y(SAMPL_SEL[11]) );
  NOR21XL U348 ( .B(n964), .A(n84), .Y(DO_VOOC[3]) );
  OR2X2 U349 ( .A(pmem_csb), .B(n80), .Y(PMEM_CSB) );
  INVX1 U350 ( .A(n88), .Y(n78) );
  INVX1 U351 ( .A(atpg_en), .Y(n88) );
  NAND2X1 U352 ( .A(n57), .B(n762), .Y(tclk_sel) );
  AND2X1 U353 ( .A(dacmux_sel[5]), .B(n67), .Y(SAMPL_SEL[5]) );
  AND2X1 U354 ( .A(dacmux_sel[7]), .B(n66), .Y(SAMPL_SEL[7]) );
  INVX1 U355 ( .A(n267), .Y(n139) );
  NAND2X1 U356 ( .A(n262), .B(n263), .Y(n1103) );
  AND2X1 U357 ( .A(n957), .B(n60), .Y(DO_VOOC[2]) );
  AND2X1 U358 ( .A(dacmux_sel[15]), .B(n67), .Y(SAMPL_SEL[15]) );
  AND2X1 U359 ( .A(dacmux_sel[6]), .B(n66), .Y(SAMPL_SEL[6]) );
  AND2X1 U360 ( .A(dacmux_sel[4]), .B(n67), .Y(SAMPL_SEL[4]) );
  AND2X1 U361 ( .A(dacmux_sel[1]), .B(n67), .Y(SAMPL_SEL[1]) );
  AND2X1 U362 ( .A(dacmux_sel[14]), .B(n67), .Y(SAMPL_SEL[14]) );
  AND2X1 U363 ( .A(dacmux_sel[16]), .B(n67), .Y(SAMPL_SEL[16]) );
  AND2X1 U364 ( .A(dacmux_sel[17]), .B(n67), .Y(SAMPL_SEL[17]) );
  AND2X1 U365 ( .A(dacmux_sel[0]), .B(n67), .Y(SAMPL_SEL[0]) );
  NAND2X1 U366 ( .A(n264), .B(n265), .Y(n1097) );
  AND2X1 U367 ( .A(r_xana_19), .B(n66), .Y(STB_RP) );
  INVX1 U368 ( .A(atpg_en), .Y(n87) );
  AND2X1 U369 ( .A(n948), .B(n61), .Y(DO_VOOC[1]) );
  AND2X1 U370 ( .A(r_srcctl[0]), .B(n62), .Y(DO_SRCCTL[0]) );
  AND2X1 U371 ( .A(n942), .B(n61), .Y(DO_VOOC[0]) );
  AND2X1 U372 ( .A(r_osc_stop), .B(n58), .Y(OSC_STOP) );
  NOR2X1 U373 ( .A(n83), .B(n263), .Y(lt_gpi[3]) );
  NOR2X1 U374 ( .A(n83), .B(n262), .Y(lt_gpi[2]) );
  NOR2X1 U375 ( .A(n82), .B(n264), .Y(lt_gpi[1]) );
  NOR2X1 U376 ( .A(n82), .B(n265), .Y(lt_gpi[0]) );
  NAND2X1 U377 ( .A(n199), .B(n57), .Y(RD_ENB) );
  NAND2X1 U378 ( .A(n245), .B(n57), .Y(SLEEP) );
  INVX1 U379 ( .A(n762), .Y(n158) );
  NOR2X1 U380 ( .A(n82), .B(n237), .Y(SH_RST) );
  NOR2X1 U381 ( .A(n84), .B(n192), .Y(DO_DPDN[0]) );
  NOR2X1 U382 ( .A(n85), .B(n241), .Y(DO_SRCCTL[5]) );
  NOR2X1 U383 ( .A(n83), .B(n242), .Y(DO_DPDN[3]) );
  NOR2X1 U384 ( .A(n85), .B(n239), .Y(DO_CCCTL[0]) );
  NOR2X1 U385 ( .A(n84), .B(n226), .Y(VPP_SEL) );
  NOR2X1 U386 ( .A(n81), .B(n233), .Y(SAMPL_SEL[9]) );
  INVX1 U387 ( .A(dacmux_sel[9]), .Y(n233) );
  NOR2X1 U388 ( .A(n79), .B(n234), .Y(SAMPL_SEL[8]) );
  INVX1 U389 ( .A(dacmux_sel[8]), .Y(n234) );
  NOR2X1 U390 ( .A(atpg_en), .B(n235), .Y(SAMPL_SEL[2]) );
  INVX1 U391 ( .A(dacmux_sel[2]), .Y(n235) );
  NOR2X1 U392 ( .A(n80), .B(n236), .Y(SAMPL_SEL[3]) );
  INVX1 U393 ( .A(dacmux_sel[3]), .Y(n236) );
  NOR2X1 U394 ( .A(n81), .B(n231), .Y(SAMPL_SEL[10]) );
  INVX1 U395 ( .A(dacmux_sel[10]), .Y(n231) );
  NOR2X1 U396 ( .A(n82), .B(n232), .Y(SAMPL_SEL[12]) );
  NOR2X1 U397 ( .A(n84), .B(n230), .Y(SAMPL_SEL[13]) );
  NOR2X1 U398 ( .A(n84), .B(n200), .Y(ANAOPT[3]) );
  NOR2X1 U399 ( .A(n82), .B(n949), .Y(ANAOPT[5]) );
  NOR2X1 U400 ( .A(n84), .B(n875), .Y(DO_SRCCTL[4]) );
  NOR2X1 U401 ( .A(n84), .B(n869), .Y(DO_SRCCTL[1]) );
  BUFX3 U402 ( .A(memaddr_c[5]), .Y(n28) );
  AO222X1 U403 ( .A(n1076), .B(r_dpdmctl[4]), .C(n908), .D(pmem_csb), .E(n910), 
        .F(dm_comp), .Y(n1075) );
  NAND3X1 U404 ( .A(n1072), .B(n1073), .C(n1074), .Y(DO_GPIO[4]) );
  AOI221XL U405 ( .A(n188), .B(n1111), .C(mcu_dbgpo[18]), .D(n1077), .E(n1078), 
        .Y(n1073) );
  AOI222XL U406 ( .A(upd_dbgpo[18]), .B(n929), .C(n187), .D(n1079), .E(n186), 
        .F(n1080), .Y(n1072) );
  AOI221XL U407 ( .A(slvo_sda), .B(n906), .C(comp_smpl[1]), .D(n911), .E(n1075), .Y(n1074) );
  MUX3X1 U408 ( .D0(n1064), .D1(n1063), .D2(n133), .S0(r_do_ts[6]), .S1(
        r_do_ts[3]), .Y(n937) );
  AOI222XL U409 ( .A(divff_5), .B(n1065), .C(n1066), .D(dp_comp), .E(n1067), 
        .F(n1122), .Y(n1064) );
  AOI222XL U410 ( .A(n1065), .B(di_xanav[1]), .C(n1068), .D(di_xanav[0]), .E(
        n1066), .F(n1108), .Y(n1063) );
  OA21X1 U411 ( .B(n131), .C(n130), .A(n129), .Y(n133) );
  OR2X1 U412 ( .A(pmem_clk[0]), .B(pmem_clk[1]), .Y(n100) );
  INVX1 U413 ( .A(pmem_clk[0]), .Y(n131) );
  AO22X1 U414 ( .A(iram_a[9]), .B(n7), .C(xram_a[9]), .D(n9), .Y(SRAM_A[9]) );
  AO22X1 U415 ( .A(iram_a[8]), .B(n7), .C(xram_a[8]), .D(n9), .Y(SRAM_A[8]) );
  AO22X1 U416 ( .A(iram_a[7]), .B(n7), .C(xram_a[7]), .D(n9), .Y(SRAM_A[7]) );
  AO22X1 U417 ( .A(iram_a[10]), .B(iram_ce), .C(xram_a[10]), .D(xram_ce), .Y(
        SRAM_A[10]) );
  NAND42X1 U418 ( .C(r_pg0_sel[1]), .D(r_pg0_sel[0]), .A(r_pg0_sel[3]), .B(
        r_pg0_sel[2]), .Y(n98) );
  INVX1 U419 ( .A(sse_adr[7]), .Y(n99) );
  OAI31XL U420 ( .A(n812), .B(o_cpurst), .C(hit_ps), .D(n813), .Y(mempsack) );
  NOR2X1 U421 ( .A(mempsrd), .B(mempswr), .Y(n812) );
  NAND2X1 U422 ( .A(ictlr_psack), .B(hit_ps), .Y(n813) );
  OAI21BBX1 U423 ( .A(SRAM_RDAT[7]), .B(n76), .C(n770), .Y(n1123) );
  NAND32X1 U424 ( .B(n153), .C(n152), .A(n151), .Y(n638) );
  NAND43X1 U425 ( .B(n928), .C(n925), .D(n930), .A(n150), .Y(n152) );
  AO222X1 U426 ( .A(mcu_dbgpo[17]), .B(n927), .C(n912), .D(mcu_dbgpo[16]), .E(
        fcp_oe), .F(n910), .Y(n153) );
  AOI222XL U427 ( .A(pmem_pgm), .B(n908), .C(do_p0[6]), .D(n186), .E(
        comp_smpl[3]), .F(n911), .Y(n151) );
  OAI21BBX1 U428 ( .A(SRAM_RDAT[4]), .B(n76), .C(n773), .Y(n1116) );
  OAI21BBX1 U429 ( .A(SRAM_RDAT[5]), .B(n76), .C(n772), .Y(n1119) );
  OAI21BBX1 U430 ( .A(SRAM_RDAT[6]), .B(n76), .C(n771), .Y(n1120) );
  OAI21BBX1 U431 ( .A(SRAM_RDAT[2]), .B(n76), .C(n775), .Y(n1121) );
  OAI21BBX1 U432 ( .A(SRAM_RDAT[0]), .B(n75), .C(n777), .Y(sram_rdat[0]) );
  OAI21BBX1 U433 ( .A(SRAM_RDAT[1]), .B(n75), .C(n776), .Y(sram_rdat[1]) );
  AO222X1 U434 ( .A(comp_smpl[2]), .B(n911), .C(n901), .D(n186), .E(
        upd_dbgpo[17]), .F(n905), .Y(n161) );
  XNOR2XL U435 ( .A(do_p0[5]), .B(n197), .Y(n901) );
  NAND43X1 U436 ( .B(n162), .C(n161), .D(n160), .A(n159), .Y(n639) );
  AOI211X1 U437 ( .C(n906), .D(n187), .A(n909), .B(n902), .Y(n159) );
  AO222X1 U438 ( .A(pmem_re), .B(n908), .C(o_dodat0_15_), .D(n913), .E(
        mcu_dbgpo[19]), .F(n899), .Y(n162) );
  AO222X1 U439 ( .A(i_rstz), .B(n158), .C(mcu_dbgpo[22]), .D(n912), .E(dp_comp), .F(n907), .Y(n160) );
  OAI21BBX1 U440 ( .A(SRAM_RDAT[3]), .B(n76), .C(n774), .Y(n1118) );
  NAND32X1 U441 ( .B(n122), .C(n121), .A(n120), .Y(DO_GPIO[3]) );
  OAI22X1 U442 ( .A(n118), .B(n109), .C(n108), .D(n107), .Y(n122) );
  AO2222XL U443 ( .A(n907), .B(n1114), .C(mcu_dbgpo[21]), .D(n1086), .E(n906), 
        .F(n1115), .G(di_pro[0]), .H(n188), .Y(n121) );
  AOI222XL U444 ( .A(comp_smpl[0]), .B(n911), .C(N449), .D(n119), .E(r_vpp_en), 
        .F(n908), .Y(n120) );
  OAI21BBX1 U445 ( .A(hit_ps), .B(mempsrd), .C(n6), .Y(n815) );
  OAI221X1 U446 ( .A(r_dpdmctl[0]), .B(n1033), .C(n1034), .D(n243), .E(n1035), 
        .Y(n942) );
  INVX1 U447 ( .A(r_dpdmctl[0]), .Y(n243) );
  OAI211X1 U448 ( .C(fcp_do), .D(n228), .A(n1036), .B(n1037), .Y(n1035) );
  AOI22X1 U449 ( .A(r_dndo_sel[3]), .B(n1041), .C(n1042), .D(n220), .Y(n1034)
         );
  AOI22X1 U450 ( .A(r_dndo_sel[3]), .B(n1053), .C(n1054), .D(n220), .Y(n1033)
         );
  OAI22X1 U451 ( .A(n1055), .B(n224), .C(r_dndo_sel[2]), .D(n1056), .Y(n1054)
         );
  OAI22X1 U452 ( .A(n1057), .B(n224), .C(r_dndo_sel[2]), .D(n1058), .Y(n1053)
         );
  AOI222XL U453 ( .A(n1036), .B(di_pro[0]), .C(n1047), .D(n1113), .E(n203), 
        .F(n1045), .Y(n1055) );
  INVX1 U454 ( .A(r_osc_gate), .Y(n259) );
  AND2X1 U455 ( .A(bist_r_ctl[5]), .B(n66), .Y(SRAM_OEB) );
  NAND2X1 U456 ( .A(d_dodat[7]), .B(n80), .Y(n770) );
  INVX1 U457 ( .A(dacmux_sel[13]), .Y(n230) );
  INVX1 U458 ( .A(dacmux_sel[12]), .Y(n232) );
  NOR21XL U459 ( .B(esfrm_rrdy), .A(n13), .Y(sse_rdrdy) );
  NAND2X1 U460 ( .A(d_dodat[3]), .B(atpg_en), .Y(n774) );
  NAND2X1 U461 ( .A(d_dodat[2]), .B(n80), .Y(n775) );
  NAND2X1 U462 ( .A(d_dodat[4]), .B(n80), .Y(n773) );
  NAND2X1 U463 ( .A(d_dodat[6]), .B(n79), .Y(n771) );
  NAND2X1 U464 ( .A(d_dodat[5]), .B(n79), .Y(n772) );
  NAND2X1 U465 ( .A(d_dodat[0]), .B(atpg_en), .Y(n777) );
  NAND2X1 U466 ( .A(d_dodat[1]), .B(n79), .Y(n776) );
  INVX1 U467 ( .A(sh_rst), .Y(n237) );
  OAI211X1 U468 ( .C(r_gpio_tm), .D(di_tst), .A(n72), .B(i_rstz), .Y(n1096) );
  AND2X1 U469 ( .A(esfrm_rrdy), .B(n13), .Y(upd_rdrdy) );
  XNOR2XL U470 ( .A(do_p0[4]), .B(n198), .Y(n1080) );
  OR2X1 U471 ( .A(mcu_ram_r), .B(mcu_ram_w), .Y(ramacc) );
  OAI21X1 U472 ( .B(pmem_pgm), .C(hwi2c_stretch), .A(r_strtch), .Y(n995) );
  INVX1 U473 ( .A(pwm_o[0]), .Y(n198) );
  NOR32XL U474 ( .B(n943), .C(n950), .A(r_gpio_oe[5]), .Y(n858) );
  NAND2X1 U475 ( .A(n991), .B(i_rstz), .Y(n943) );
  AO21X1 U476 ( .B(n140), .C(n943), .A(n139), .Y(n861) );
  OAI221X1 U477 ( .A(n848), .B(s0_rxdoe), .C(n801), .D(n985), .E(r_gpio_oe[2]), 
        .Y(n140) );
  AOI22X1 U478 ( .A(n207), .B(N261), .C(n196), .D(n249), .Y(n985) );
  NOR21XL U479 ( .B(n943), .A(r_gpio_oe[4]), .Y(n859) );
  NAND32X1 U480 ( .B(n139), .C(n138), .A(r_gpio_oe[1]), .Y(n862) );
  AO22X1 U481 ( .A(n797), .B(n979), .C(n137), .D(n258), .Y(n138) );
  INVX1 U482 ( .A(n845), .Y(n137) );
  OAI22X1 U483 ( .A(N264), .B(n972), .C(n253), .D(n973), .Y(n979) );
  NAND32X1 U484 ( .B(n139), .C(n136), .A(r_gpio_oe[0]), .Y(n863) );
  AO22X1 U485 ( .A(n802), .B(n970), .C(n135), .D(n258), .Y(n136) );
  INVX1 U486 ( .A(n844), .Y(n135) );
  OAI22X1 U487 ( .A(N267), .B(n972), .C(n252), .D(n973), .Y(n970) );
  INVX1 U488 ( .A(n142), .Y(n857) );
  NAND32X1 U489 ( .B(n141), .C(r_gpio_oe[6]), .A(n950), .Y(n142) );
  INVX1 U490 ( .A(n943), .Y(n141) );
  NAND2X1 U491 ( .A(d_dodat[13]), .B(atpg_en), .Y(n779) );
  NAND2X1 U492 ( .A(d_dodat[11]), .B(n79), .Y(n781) );
  NAND2X1 U493 ( .A(d_dodat[12]), .B(n82), .Y(n780) );
  AOI22X1 U494 ( .A(n207), .B(N258), .C(n196), .D(n250), .Y(n992) );
  NAND2X1 U495 ( .A(d_dodat[9]), .B(n78), .Y(n783) );
  NAND2X1 U496 ( .A(d_dodat[15]), .B(n79), .Y(n778) );
  NAND2X1 U497 ( .A(d_dodat[8]), .B(n80), .Y(n784) );
  OAI21BBX1 U498 ( .A(n990), .B(n943), .C(n267), .Y(n860) );
  OAI211X1 U499 ( .C(n992), .D(n993), .A(n994), .B(r_gpio_oe[3]), .Y(n990) );
  NAND21X1 U500 ( .B(N259), .A(n248), .Y(n993) );
  NAND4X1 U501 ( .A(N259), .B(N260), .C(N258), .D(n258), .Y(n994) );
  NAND2X1 U502 ( .A(d_dodat[10]), .B(n79), .Y(n782) );
  INVX1 U503 ( .A(d_dodat[14]), .Y(n266) );
  OAI22AX1 U504 ( .D(r_fortxrdy), .C(r_fortxdat), .A(r_fortxrdy), .B(ptx_cc), 
        .Y(n904) );
  OAI21BBX1 U505 ( .A(RX_DAT), .B(n74), .C(n783), .Y(n1114) );
  OAI21BBX1 U506 ( .A(DI_GPIO[2]), .B(n74), .C(n775), .Y(di_gpio[2]) );
  OAI22X1 U507 ( .A(slvo_sda), .B(n212), .C(mcuo_sda), .D(n208), .Y(n973) );
  MUX2BXL U508 ( .D0(n1070), .D1(n1069), .S(r_do_ts[6]), .Y(n129) );
  AO222X1 U509 ( .A(di_aswk[3]), .B(n1067), .C(di_pro[5]), .D(n1066), .E(n1112), .F(n1065), .Y(n1069) );
  AOI211X1 U510 ( .C(n1115), .D(n1067), .A(n1068), .B(n1071), .Y(n1070) );
  AO22X1 U511 ( .A(divff_8), .B(n1065), .C(dm_comp), .D(n201), .Y(n1071) );
  OAI21BBX1 U512 ( .A(SRCI[5]), .B(n73), .C(n780), .Y(di_pro[5]) );
  OAI21BBX1 U513 ( .A(DI_GPIO[3]), .B(n75), .C(n774), .Y(n1117) );
  OAI21BBX1 U514 ( .A(SRCI[3]), .B(n73), .C(n782), .Y(n1112) );
  NOR2X1 U515 ( .A(n216), .B(r_i2cmcu_route[1]), .Y(n788) );
  NOR2X1 U516 ( .A(n211), .B(r_i2cslv_route[1]), .Y(n792) );
  NOR2X1 U517 ( .A(r_i2cmcu_route[0]), .B(r_i2cmcu_route[1]), .Y(n786) );
  NOR2X1 U518 ( .A(r_i2cslv_route[0]), .B(r_i2cslv_route[1]), .Y(n791) );
  OAI21BBX1 U519 ( .A(DM_FAULT), .B(n73), .C(n778), .Y(di_aswk[3]) );
  AOI222XL U520 ( .A(x_clk), .B(n158), .C(n924), .D(n1114), .E(n923), .F(n1112), .Y(n150) );
  OAI21BBX1 U521 ( .A(DP_COMP), .B(n74), .C(n779), .Y(dp_comp) );
  OAI21BBX1 U522 ( .A(DM_COMP), .B(n73), .C(n780), .Y(dm_comp) );
  OAI21BBX1 U523 ( .A(SRCI[4]), .B(n73), .C(n781), .Y(n1108) );
  OAI22AX1 U524 ( .D(n826), .C(n827), .A(n195), .B(n826), .Y(exint[1]) );
  NAND2X1 U525 ( .A(n833), .B(N267), .Y(n826) );
  OAI22AX1 U526 ( .D(n828), .C(n829), .A(di_gpio[1]), .B(n828), .Y(n827) );
  NAND3X1 U527 ( .A(N264), .B(n251), .C(N266), .Y(n828) );
  OAI22AX1 U528 ( .D(n834), .C(n835), .A(n195), .B(n834), .Y(exint[0]) );
  NAND2X1 U529 ( .A(n833), .B(n252), .Y(n834) );
  OAI22AX1 U530 ( .D(n836), .C(n837), .A(di_gpio[1]), .B(n836), .Y(n835) );
  NAND3X1 U531 ( .A(n253), .B(n251), .C(N266), .Y(n836) );
  NOR2X1 U532 ( .A(n1117), .B(N259), .Y(n800) );
  INVX1 U533 ( .A(r_do_ts[4]), .Y(n201) );
  AOI32X1 U534 ( .A(n800), .B(n830), .C(n831), .D(n247), .E(n190), .Y(n829) );
  NOR2X1 U535 ( .A(n250), .B(n248), .Y(n831) );
  INVX1 U536 ( .A(n830), .Y(n247) );
  NAND2X1 U537 ( .A(n832), .B(N261), .Y(n830) );
  AOI32X1 U538 ( .A(N260), .B(n800), .C(n838), .D(n839), .E(n190), .Y(n837) );
  NOR2X1 U539 ( .A(N258), .B(n839), .Y(n838) );
  AND2X1 U540 ( .A(n832), .B(n249), .Y(n839) );
  NOR2X1 U541 ( .A(n201), .B(r_do_ts[5]), .Y(n1065) );
  INVX1 U542 ( .A(r_do_ts[5]), .Y(n202) );
  INVX1 U543 ( .A(r_i2cmcu_route[0]), .Y(n216) );
  INVX1 U544 ( .A(r_i2cslv_route[0]), .Y(n211) );
  ENOX1 U545 ( .A(n255), .B(n242), .C(n910), .D(fcp_do), .Y(n909) );
  NOR2X1 U546 ( .A(n202), .B(r_do_ts[4]), .Y(n1066) );
  NAND3X1 U547 ( .A(N266), .B(N265), .C(N264), .Y(n845) );
  NAND3X1 U548 ( .A(N269), .B(N268), .C(N267), .Y(n844) );
  OAI21BBX1 U549 ( .A(DAC1_COMP), .B(n74), .C(n784), .Y(n1110) );
  OAI21BBX1 U550 ( .A(DI_GPIO[0]), .B(n74), .C(n777), .Y(di_gpio[0]) );
  OAI21BBX1 U551 ( .A(SRCI[2]), .B(n73), .C(n783), .Y(n1113) );
  OAI21BBX1 U552 ( .A(DI_GPIO[1]), .B(n74), .C(n776), .Y(di_gpio[1]) );
  OAI21BBX1 U553 ( .A(CC1_DI), .B(n73), .C(n770), .Y(n1122) );
  OAI21BBX1 U554 ( .A(CC2_DI), .B(n73), .C(n778), .Y(n1115) );
  NOR2X1 U555 ( .A(r_fortxen), .B(ptx_oe), .Y(n955) );
  OAI22X1 U556 ( .A(n840), .B(n215), .C(n4), .D(n841), .Y(dpdm_urx) );
  AOI22AXL U557 ( .A(r_pwrctl[7]), .B(n214), .D(r_pwrctl[7]), .C(n842), .Y(
        n840) );
  AOI22X1 U558 ( .A(n842), .B(n240), .C(r_pwrctl[6]), .D(n214), .Y(n841) );
  INVX1 U559 ( .A(n805), .Y(n214) );
  NOR2X1 U560 ( .A(r_do_ts[4]), .B(r_do_ts[5]), .Y(n1068) );
  NAND3X1 U561 ( .A(N263), .B(N261), .C(N262), .Y(n848) );
  INVX1 U562 ( .A(N261), .Y(n249) );
  OAI22AX1 U563 ( .D(n793), .C(n794), .A(di_gpio[0]), .B(n793), .Y(n787) );
  NAND2X1 U564 ( .A(N267), .B(n802), .Y(n793) );
  EORX1 U565 ( .A(n795), .B(n796), .C(n796), .D(di_gpio[1]), .Y(n794) );
  NAND2X1 U566 ( .A(N264), .B(n797), .Y(n796) );
  EORX1 U567 ( .A(n843), .B(n844), .C(n844), .D(di_gpio[0]), .Y(n842) );
  OAI22AX1 U568 ( .D(n845), .C(n846), .A(di_gpio[1]), .B(n845), .Y(n843) );
  AOI32X1 U569 ( .A(N259), .B(N260), .C(n847), .D(n246), .E(n190), .Y(n846) );
  NOR3XL U570 ( .A(n250), .B(n1117), .C(n246), .Y(n847) );
  OAI21BBX1 U571 ( .A(XANAV[1]), .B(n74), .C(n776), .Y(di_xanav[1]) );
  OAI21BBX1 U572 ( .A(XANAV[0]), .B(n73), .C(n777), .Y(di_xanav[0]) );
  AOI21X1 U573 ( .B(n798), .C(di_gpio[2]), .A(n799), .Y(n795) );
  AOI31X1 U574 ( .A(n800), .B(n248), .C(N258), .D(n798), .Y(n799) );
  NOR2X1 U575 ( .A(n249), .B(n801), .Y(n798) );
  AOI21X1 U576 ( .B(n810), .C(di_gpio[2]), .A(n811), .Y(n808) );
  AOI31X1 U577 ( .A(n250), .B(n248), .C(n800), .D(n810), .Y(n811) );
  NOR2X1 U578 ( .A(n801), .B(N261), .Y(n810) );
  INVX1 U579 ( .A(r_ccctl[0]), .Y(n239) );
  INVX1 U580 ( .A(r_accctl[4]), .Y(n192) );
  OAI21BBX1 U581 ( .A(RX_SQL), .B(n74), .C(n781), .Y(n1107) );
  OAI21BBX1 U588 ( .A(SRCI[0]), .B(n74), .C(n770), .Y(di_pro[0]) );
  OAI21BBX1 U589 ( .A(SRCI[1]), .B(n74), .C(n784), .Y(n1111) );
  INVX1 U590 ( .A(N267), .Y(n252) );
  INVX1 U591 ( .A(prx_rcvinf[4]), .Y(n107) );
  INVX1 U592 ( .A(N260), .Y(n248) );
  INVX1 U593 ( .A(N264), .Y(n253) );
  INVX1 U600 ( .A(N258), .Y(n250) );
  NOR2X1 U601 ( .A(N266), .B(N265), .Y(n797) );
  NOR2X1 U602 ( .A(N269), .B(N268), .Y(n802) );
  OR2X1 U603 ( .A(N263), .B(N262), .Y(n801) );
  INVX1 U604 ( .A(r_dpdmctl[6]), .Y(n242) );
  AND2X1 U605 ( .A(r_do_ts[2]), .B(n61), .Y(DO_TS[2]) );
  INVX1 U606 ( .A(mcu_dbgpo[16]), .Y(n109) );
  OAI21BBX1 U607 ( .A(DI_GPIO[5]), .B(n75), .C(n772), .Y(di_gpio[5]) );
  OAI21BBX1 U608 ( .A(DI_GPIO[6]), .B(n75), .C(n771), .Y(di_gpio[6]) );
  OAI21BBX1 U609 ( .A(DI_TS), .B(n75), .C(n781), .Y(di_ts) );
  MUX4X1 U610 ( .D0(n134), .D1(n1008), .D2(n1020), .D3(n1007), .S0(
        r_dpdo_sel[3]), .S1(r_dpdo_sel[2]), .Y(n957) );
  OAI22X1 U611 ( .A(n1025), .B(n189), .C(r_dpdo_sel[1]), .D(n1026), .Y(n1020)
         );
  OAI22X1 U612 ( .A(n1016), .B(n189), .C(r_dpdo_sel[1]), .D(n1017), .Y(n1007)
         );
  AO21X1 U613 ( .B(n1004), .C(n189), .A(n1021), .Y(n134) );
  OAI22X1 U614 ( .A(n1009), .B(n189), .C(r_dpdo_sel[1]), .D(n1010), .Y(n1008)
         );
  AOI221XL U615 ( .A(n1011), .B(di_aswk[1]), .C(n223), .D(r_ocdrv_enz), .E(
        n1014), .Y(n1009) );
  AOI221XL U616 ( .A(n1011), .B(pwm_o[1]), .C(n223), .D(r_osc_stop), .E(n1012), 
        .Y(n1010) );
  ENOX1 U617 ( .A(n1013), .B(n199), .C(n1109), .D(n1015), .Y(n1014) );
  OAI22X1 U618 ( .A(n1049), .B(n224), .C(r_dndo_sel[2]), .D(n1050), .Y(n1041)
         );
  AOI221XL U619 ( .A(r_xana[12]), .B(n1047), .C(n1045), .D(CC2_DOB), .E(n1052), 
        .Y(n1049) );
  AOI221XL U620 ( .A(n1047), .B(o_dodat0_15_), .C(n1045), .D(r_pwrdn), .E(
        n1051), .Y(n1050) );
  OAI22X1 U621 ( .A(n226), .B(n219), .C(n875), .D(n218), .Y(n1052) );
  MUX2IX1 U622 ( .D0(n123), .D1(n124), .S(r_i2crout[4]), .Y(n26) );
  MUX2X1 U623 ( .D0(n124), .D1(n123), .S(r_i2crout[4]), .Y(CC1_DOB) );
  OAI21BBX1 U624 ( .A(DRP_OSC), .B(n72), .C(n779), .Y(di_aswk[0]) );
  INVX1 U625 ( .A(r_xana_18), .Y(n199) );
  OAI22X1 U626 ( .A(n1022), .B(n189), .C(r_dpdo_sel[1]), .D(n1023), .Y(n1021)
         );
  AOI22X1 U627 ( .A(n223), .B(n1107), .C(n222), .D(n1114), .Y(n1023) );
  AOI221XL U628 ( .A(n1011), .B(TX_DAT), .C(n223), .D(n1122), .E(n1024), .Y(
        n1022) );
  ENOX1 U629 ( .A(n955), .B(n221), .C(n1115), .D(n222), .Y(n1024) );
  AOI221XL U630 ( .A(n1045), .B(CC1_DOB), .C(n1046), .D(n227), .E(n193), .Y(
        n1057) );
  INVX1 U631 ( .A(n1060), .Y(n193) );
  AOI32X1 U632 ( .A(n1036), .B(r_vpp0v_en), .C(r_pwrdn), .D(n1047), .E(
        r_srcctl[0]), .Y(n1060) );
  INVX1 U633 ( .A(sfr_intr[2]), .Y(n673) );
  NOR21XL U634 ( .B(i2c_ev_3), .A(sse_adr[7]), .Y(i2c_ev_2) );
  NOR21XL U635 ( .B(N263), .A(N262), .Y(n832) );
  OAI211X1 U636 ( .C(sdischg_duty), .D(n128), .A(r_srcctl[4]), .B(n127), .Y(
        n875) );
  INVX1 U637 ( .A(r_sdischg[6]), .Y(n128) );
  NOR2X1 U638 ( .A(r_dpdo_sel[0]), .B(r_dpdmctl[2]), .Y(n1015) );
  NOR2X1 U639 ( .A(r_dndo_sel[0]), .B(r_dndo_sel[1]), .Y(n1036) );
  NOR2X1 U640 ( .A(n225), .B(r_dndo_sel[0]), .Y(n1046) );
  OAI221X1 U641 ( .A(r_pwrctl[7]), .B(n996), .C(r_i2crout[5]), .D(n206), .E(
        n997), .Y(n964) );
  OAI21X1 U642 ( .B(s0_rxdoe), .C(n215), .A(r_pwrctl[7]), .Y(n997) );
  INVX1 U643 ( .A(n998), .Y(n206) );
  AOI22X1 U644 ( .A(r_i2crout[5]), .B(n999), .C(r_dpdmctl[3]), .D(n1000), .Y(
        n996) );
  OAI21BBX1 U645 ( .A(IMP_OSC), .B(n77), .C(n779), .Y(di_aswk[4]) );
  NOR2X1 U646 ( .A(n217), .B(r_dndo_sel[1]), .Y(n1047) );
  NAND2X1 U647 ( .A(r_dpdo_sel[0]), .B(n244), .Y(n1019) );
  OAI21BBX1 U648 ( .A(RD_DET), .B(n73), .C(n780), .Y(n1109) );
  NAND2X1 U649 ( .A(r_dpdo_sel[0]), .B(r_dpdmctl[2]), .Y(n1013) );
  OAI22X1 U650 ( .A(mcuo_sda), .B(n204), .C(slvo_sda), .D(n210), .Y(n124) );
  NOR2X1 U651 ( .A(n244), .B(r_dpdo_sel[0]), .Y(n1011) );
  XOR2X1 U652 ( .A(r_aopt[3]), .B(n27), .Y(n200) );
  NAND2X1 U653 ( .A(di_aswk[4]), .B(r_imp_osc), .Y(n27) );
  INVX1 U654 ( .A(r_dpdmctl[2]), .Y(n244) );
  OAI22X1 U655 ( .A(n1043), .B(n224), .C(r_dndo_sel[2]), .D(n1044), .Y(n1042)
         );
  AOI221XL U656 ( .A(n1046), .B(n1110), .C(n1036), .D(n1111), .E(n1048), .Y(
        n1043) );
  AOI222XL U657 ( .A(n1045), .B(n1115), .C(n1046), .D(TX_DAT), .E(n1047), .F(
        n1114), .Y(n1044) );
  AO22X1 U658 ( .A(di_pro[5]), .B(n1045), .C(n1112), .D(n1047), .Y(n1048) );
  AOI211X1 U659 ( .C(n1038), .D(n228), .A(r_dndo_sel[3]), .B(r_dndo_sel[2]), 
        .Y(n1037) );
  OAI21BBX1 U660 ( .A(n1039), .B(r_pwrctl[6]), .C(n1040), .Y(n1038) );
  OAI22X1 U661 ( .A(n215), .B(do_opt[6]), .C(do_opt[7]), .D(r_i2crout[5]), .Y(
        n1039) );
  OAI21BBX1 U662 ( .A(n1000), .B(r_dpdmctl[0]), .C(n240), .Y(n1040) );
  INVX1 U663 ( .A(r_dndo_sel[0]), .Y(n217) );
  INVX1 U664 ( .A(r_otpi_gate), .Y(n127) );
  ENOX1 U665 ( .A(n87), .B(n266), .C(PMEM_Q0[6]), .D(n87), .Y(pmem_q0[6]) );
  OAI21BBX1 U666 ( .A(PMEM_Q1[6]), .B(n88), .C(n771), .Y(pmem_q1[6]) );
  NOR21XL U667 ( .B(N269), .A(N268), .Y(n833) );
  OAI21BBX1 U668 ( .A(PMEM_Q0[7]), .B(n77), .C(n778), .Y(pmem_q0[7]) );
  OAI21BBX1 U669 ( .A(PMEM_Q1[7]), .B(n87), .C(n770), .Y(pmem_q1[7]) );
  OAI21BBX1 U670 ( .A(PMEM_Q1[1]), .B(n77), .C(n776), .Y(pmem_q1[1]) );
  OAI21BBX1 U671 ( .A(PMEM_Q0[1]), .B(n76), .C(n783), .Y(pmem_q0[1]) );
  OAI21BBX1 U672 ( .A(PMEM_Q1[5]), .B(n77), .C(n772), .Y(pmem_q1[5]) );
  OAI21BBX1 U673 ( .A(PMEM_Q0[5]), .B(n77), .C(n779), .Y(pmem_q0[5]) );
  OAI21BBX1 U674 ( .A(PMEM_Q1[3]), .B(n77), .C(n774), .Y(pmem_q1[3]) );
  OAI21BBX1 U675 ( .A(PMEM_Q0[3]), .B(n76), .C(n781), .Y(pmem_q0[3]) );
  OAI21BBX1 U676 ( .A(PMEM_Q0[2]), .B(n76), .C(n782), .Y(pmem_q0[2]) );
  OAI21BBX1 U677 ( .A(PMEM_Q1[2]), .B(n77), .C(n775), .Y(pmem_q1[2]) );
  OAI21BBX1 U678 ( .A(r_xtm[7]), .B(n254), .C(r_aopt[5]), .Y(n949) );
  OAI211X1 U679 ( .C(sdischg_duty), .D(n126), .A(r_srcctl[1]), .B(n127), .Y(
        n869) );
  INVX1 U680 ( .A(r_sdischg[5]), .Y(n126) );
  INVX1 U681 ( .A(r_i2crout[5]), .Y(n215) );
  OAI21BBX1 U682 ( .A(STB_OVP), .B(n72), .C(n779), .Y(di_aswk[1]) );
  NAND2X1 U683 ( .A(r_i2cmcu_route[1]), .B(n216), .Y(n1032) );
  NAND2X1 U684 ( .A(r_i2cslv_route[1]), .B(n211), .Y(n1031) );
  OAI211X1 U685 ( .C(r_pwrctl[6]), .D(n1028), .A(n228), .B(n1029), .Y(n948) );
  AOI22X1 U686 ( .A(r_pwrctl[6]), .B(n1030), .C(r_i2crout[5]), .D(n998), .Y(
        n1029) );
  AOI22X1 U687 ( .A(n999), .B(n215), .C(r_dpdmctl[1]), .D(n1000), .Y(n1028) );
  NAND2X1 U688 ( .A(n258), .B(n215), .Y(n1030) );
  INVX1 U689 ( .A(N265), .Y(n251) );
  INVX1 U690 ( .A(r_i2c_ninc), .Y(n672) );
  AOI211X1 U691 ( .C(r_pwrctl[7]), .D(n1005), .A(r_dpdo_sel[0]), .B(n1006), 
        .Y(n1004) );
  OAI22X1 U692 ( .A(do_opt[7]), .B(n215), .C(r_i2crout[5]), .D(do_opt[6]), .Y(
        n1005) );
  AOI21X1 U693 ( .B(r_dpdmctl[2]), .C(n1000), .A(r_pwrctl[7]), .Y(n1006) );
  INVX1 U694 ( .A(r_dndo_sel[1]), .Y(n225) );
  INVX1 U695 ( .A(r_vpp_en), .Y(n226) );
  INVX1 U696 ( .A(r_srcctl[5]), .Y(n241) );
  INVX1 U697 ( .A(r_sleep), .Y(n245) );
  OAI22X1 U698 ( .A(slvo_sda), .B(n1031), .C(mcuo_sda), .D(n1032), .Y(n998) );
  OAI21BBX1 U699 ( .A(PMEM_Q0[0]), .B(n76), .C(n784), .Y(pmem_q0[0]) );
  OAI21BBX1 U700 ( .A(PMEM_Q1[0]), .B(n77), .C(n777), .Y(pmem_q1[0]) );
  OAI21BBX1 U701 ( .A(PMEM_Q0[4]), .B(n77), .C(n780), .Y(pmem_q0[4]) );
  OAI21BBX1 U702 ( .A(PMEM_Q1[4]), .B(n77), .C(n773), .Y(pmem_q1[4]) );
  INVX1 U703 ( .A(r_dpdo_sel[1]), .Y(n189) );
  INVX1 U704 ( .A(r_dndo_sel[2]), .Y(n224) );
  INVX1 U705 ( .A(r_pwrctl[6]), .Y(n240) );
  INVX1 U706 ( .A(sfr_intr[3]), .Y(n674) );
  OAI22X1 U707 ( .A(dp_comp), .B(n215), .C(r_i2crout[5]), .D(dm_comp), .Y(n805) );
  OAI22X1 U708 ( .A(n4), .B(dp_comp), .C(dm_comp), .D(n215), .Y(n790) );
  OAI22X1 U709 ( .A(r_i2crout[4]), .B(n1122), .C(n1115), .D(n213), .Y(n789) );
  OAI22X1 U710 ( .A(n1122), .B(n213), .C(r_i2crout[4]), .D(n1115), .Y(n804) );
  INVX1 U711 ( .A(r_dndo_sel[3]), .Y(n220) );
  INVX1 U712 ( .A(r_i2crout[4]), .Y(n213) );
  OAI21BBX1 U713 ( .A(t_di_gpio4), .B(n75), .C(n773), .Y(di_gpio[4]) );
  OAI21BBX1 U714 ( .A(XANAV[2]), .B(n75), .C(n775), .Y(di_xanav[2]) );
  OAI21BBX1 U715 ( .A(XANAV[3]), .B(n75), .C(n774), .Y(di_xanav[3]) );
  OAI21BBX1 U716 ( .A(XANAV[4]), .B(n75), .C(n773), .Y(di_xanav[4]) );
  NAND21X1 U717 ( .B(r_gpio_ie[0]), .A(n56), .Y(GPIO_IE[0]) );
  AND2X2 U718 ( .A(pmem_twlb[1]), .B(n58), .Y(PMEM_TWLB[1]) );
  AND2X2 U719 ( .A(pmem_twlb[0]), .B(n59), .Y(PMEM_TWLB[0]) );
  NAND21X1 U720 ( .B(i_rstz), .A(di_tst), .Y(n267) );
  NAND21X1 U721 ( .B(r_gpio_ie[1]), .A(n56), .Y(GPIO_IE[1]) );
  AND3X1 U722 ( .A(di_tst), .B(n761), .C(n265), .Y(tm_atpg) );
  AND2X1 U723 ( .A(pmem_re), .B(n58), .Y(PMEM_RE) );
  AND2X1 U724 ( .A(pmem_clk[0]), .B(n58), .Y(PMEM_CLK[0]) );
  AND2X1 U725 ( .A(pmem_clk[1]), .B(n58), .Y(PMEM_CLK[1]) );
  NOR2X1 U726 ( .A(n1103), .B(r_lt_gpi[1]), .Y(n761) );
  AND2X1 U727 ( .A(di_tst), .B(n62), .Y(n931) );
  NAND3X1 U728 ( .A(r_lt_gpi[0]), .B(n761), .C(n931), .Y(n762) );
  NAND21X1 U729 ( .B(r_cctrx[2]), .A(n56), .Y(DO_CCTRX[2]) );
  NAND21X1 U730 ( .B(r_cctrx[1]), .A(n56), .Y(DO_CCTRX[1]) );
  AND2X1 U731 ( .A(r_pu_gpio[1]), .B(n60), .Y(GPIO_PU[1]) );
  AND2X1 U732 ( .A(r_pd_gpio[6]), .B(n60), .Y(GPIO_PD[6]) );
  AND2X1 U733 ( .A(r_pd_gpio[5]), .B(n60), .Y(GPIO_PD[5]) );
  AND2X1 U734 ( .A(r_pd_gpio[4]), .B(n60), .Y(GPIO_PD[4]) );
  AND2X1 U735 ( .A(r_pu_gpio[3]), .B(n59), .Y(GPIO_PU[3]) );
  AND2X1 U736 ( .A(r_pu_gpio[2]), .B(n59), .Y(GPIO_PU[2]) );
  AND2X1 U737 ( .A(r_pu_gpio[0]), .B(n60), .Y(GPIO_PU[0]) );
  AND2X1 U738 ( .A(r_pd_gpio[2]), .B(n60), .Y(GPIO_PD[2]) );
  AND2X1 U739 ( .A(r_do_ts[1]), .B(n61), .Y(DO_TS[1]) );
  AND2X1 U740 ( .A(r_do_ts[0]), .B(n61), .Y(DO_TS[0]) );
  AND2X1 U741 ( .A(r_pu_gpio[6]), .B(n59), .Y(GPIO_PU[6]) );
  AND2X1 U742 ( .A(r_pu_gpio[5]), .B(n59), .Y(GPIO_PU[5]) );
  AND2X1 U743 ( .A(r_pu_gpio[4]), .B(n59), .Y(GPIO_PU[4]) );
  AND2X1 U744 ( .A(r_pd_gpio[3]), .B(n60), .Y(GPIO_PD[3]) );
  AND2X1 U745 ( .A(r_pd_gpio[1]), .B(n60), .Y(GPIO_PD[1]) );
  AND2X1 U746 ( .A(r_pd_gpio[0]), .B(n60), .Y(GPIO_PD[0]) );
  INVX1 U747 ( .A(r_lt_gpi[0]), .Y(n265) );
  INVX1 U748 ( .A(r_lt_gpi[1]), .Y(n264) );
  INVX1 U749 ( .A(r_lt_gpi[3]), .Y(n263) );
  INVX1 U750 ( .A(r_lt_gpi[2]), .Y(n262) );
  NAND2X1 U751 ( .A(r_lt_gpi[2]), .B(n263), .Y(n1095) );
  NAND2X1 U752 ( .A(r_lt_gpi[1]), .B(r_lt_gpi[0]), .Y(n1099) );
  NAND2X1 U753 ( .A(r_lt_gpi[3]), .B(n262), .Y(n1100) );
  NAND2X1 U754 ( .A(r_lt_gpi[1]), .B(n265), .Y(n1098) );
  NAND2X1 U755 ( .A(r_lt_gpi[3]), .B(r_lt_gpi[2]), .Y(n1102) );
  NAND2X1 U756 ( .A(r_lt_gpi[0]), .B(n264), .Y(n1101) );
  AND2X1 U757 ( .A(PWRDN), .B(r_vpp0v_en), .Y(VPP_0V) );
  AND2X1 U758 ( .A(r_regtrm[0]), .B(n58), .Y(REGTRM[0]) );
  AND2X1 U759 ( .A(r_regtrm[1]), .B(n72), .Y(REGTRM[1]) );
  AND2X1 U760 ( .A(r_regtrm[2]), .B(n71), .Y(REGTRM[2]) );
  AND2X1 U761 ( .A(r_regtrm[3]), .B(n70), .Y(REGTRM[3]) );
  AND2X1 U762 ( .A(r_regtrm[4]), .B(n68), .Y(REGTRM[4]) );
  AND2X1 U763 ( .A(r_regtrm[5]), .B(n68), .Y(REGTRM[5]) );
  AND2X1 U764 ( .A(r_regtrm[6]), .B(n68), .Y(REGTRM[6]) );
  AND2X1 U765 ( .A(r_regtrm[7]), .B(n68), .Y(REGTRM[7]) );
  AND2X1 U766 ( .A(r_regtrm[8]), .B(n67), .Y(REGTRM[8]) );
  AND2X1 U767 ( .A(r_regtrm[9]), .B(n67), .Y(REGTRM[9]) );
  AND2X1 U768 ( .A(r_regtrm[11]), .B(n57), .Y(REGTRM[11]) );
  AND2X1 U769 ( .A(r_regtrm[13]), .B(n57), .Y(REGTRM[13]) );
  AND2X1 U770 ( .A(r_regtrm[14]), .B(n58), .Y(REGTRM[14]) );
  AND2X1 U771 ( .A(r_regtrm[15]), .B(n57), .Y(REGTRM[15]) );
  AND2X1 U772 ( .A(r_regtrm[16]), .B(n59), .Y(REGTRM[16]) );
  AND2X1 U773 ( .A(r_regtrm[17]), .B(n57), .Y(REGTRM[17]) );
  AND2X1 U774 ( .A(r_regtrm[19]), .B(n72), .Y(REGTRM[19]) );
  AND2X1 U775 ( .A(r_regtrm[21]), .B(n71), .Y(REGTRM[21]) );
  AND2X1 U776 ( .A(r_regtrm[22]), .B(n72), .Y(REGTRM[22]) );
  AND2X1 U777 ( .A(r_regtrm[23]), .B(n72), .Y(REGTRM[23]) );
  AND2X1 U778 ( .A(r_regtrm[40]), .B(n70), .Y(REGTRM[40]) );
  AND2X1 U779 ( .A(r_regtrm[41]), .B(n69), .Y(REGTRM[41]) );
  AND2X1 U780 ( .A(r_regtrm[43]), .B(n69), .Y(REGTRM[43]) );
  AND2X1 U781 ( .A(r_regtrm[44]), .B(n69), .Y(REGTRM[44]) );
  AND2X1 U782 ( .A(r_regtrm[45]), .B(n69), .Y(REGTRM[45]) );
  AND2X1 U783 ( .A(r_regtrm[46]), .B(n69), .Y(REGTRM[46]) );
  AND2X1 U784 ( .A(r_regtrm[47]), .B(n69), .Y(REGTRM[47]) );
  AND2X1 U785 ( .A(r_regtrm[48]), .B(n69), .Y(REGTRM[48]) );
  AND2X1 U786 ( .A(r_regtrm[49]), .B(n69), .Y(REGTRM[49]) );
  AND2X1 U787 ( .A(r_regtrm[51]), .B(n68), .Y(REGTRM[51]) );
  AND2X1 U788 ( .A(r_regtrm[52]), .B(n68), .Y(REGTRM[52]) );
  AND2X1 U789 ( .A(r_regtrm[53]), .B(n68), .Y(REGTRM[53]) );
  AND2X1 U790 ( .A(r_regtrm[54]), .B(n68), .Y(REGTRM[54]) );
  AND2X1 U791 ( .A(r_regtrm[55]), .B(n68), .Y(REGTRM[55]) );
  AND2X1 U792 ( .A(r_sdischg[7]), .B(n59), .Y(LDO3P9V) );
  AND2X1 U793 ( .A(r_dpdmctl[7]), .B(n62), .Y(DO_DPDN[4]) );
  AND2X1 U794 ( .A(r_xtm[0]), .B(n66), .Y(XTM[0]) );
  AND2X1 U795 ( .A(r_xtm[1]), .B(n66), .Y(XTM[1]) );
  AND2X1 U796 ( .A(r_ccctl[7]), .B(n63), .Y(DO_CCCTL[7]) );
  AND2X1 U797 ( .A(r_ccctl[6]), .B(n63), .Y(DO_CCCTL[6]) );
  AND2X1 U798 ( .A(r_ccctl[4]), .B(n64), .Y(DO_CCCTL[4]) );
  AND2X1 U799 ( .A(r_ccctl[5]), .B(n64), .Y(DO_CCCTL[5]) );
  AND2X1 U800 ( .A(r_srcctl[3]), .B(n61), .Y(DO_SRCCTL[3]) );
  AND2X1 U801 ( .A(r_srcctl[2]), .B(n61), .Y(DO_SRCCTL[2]) );
  AND2X1 U802 ( .A(r_dpdmctl[4]), .B(n62), .Y(DO_DPDN[1]) );
  AND2X1 U803 ( .A(x_daclsb[2]), .B(n64), .Y(DAC1_EN) );
  AND2X1 U804 ( .A(r_regtrm[12]), .B(n57), .Y(REGTRM[12]) );
  AND2X1 U805 ( .A(r_xana[15]), .B(n65), .Y(ANA_REGX[15]) );
  AND2X1 U806 ( .A(r_xana[13]), .B(n65), .Y(ANA_REGX[13]) );
  AND2X1 U807 ( .A(r_xana[14]), .B(n65), .Y(ANA_REGX[14]) );
  AND2X1 U808 ( .A(r_regtrm[10]), .B(n58), .Y(REGTRM[10]) );
  AND2X1 U809 ( .A(r_regtrm[18]), .B(n61), .Y(REGTRM[18]) );
  AND2X1 U810 ( .A(r_regtrm[20]), .B(n71), .Y(REGTRM[20]) );
  AND2X1 U811 ( .A(r_regtrm[25]), .B(n71), .Y(REGTRM[25]) );
  AND2X1 U812 ( .A(r_regtrm[26]), .B(n71), .Y(REGTRM[26]) );
  AND2X1 U813 ( .A(r_regtrm[27]), .B(n71), .Y(REGTRM[27]) );
  AND2X1 U814 ( .A(r_regtrm[28]), .B(n71), .Y(REGTRM[28]) );
  AND2X1 U815 ( .A(r_regtrm[29]), .B(n71), .Y(REGTRM[29]) );
  AND2X1 U816 ( .A(r_regtrm[30]), .B(n71), .Y(REGTRM[30]) );
  AND2X1 U817 ( .A(r_regtrm[31]), .B(n70), .Y(REGTRM[31]) );
  AND2X1 U818 ( .A(r_regtrm[32]), .B(n70), .Y(REGTRM[32]) );
  AND2X1 U819 ( .A(r_regtrm[33]), .B(n71), .Y(REGTRM[33]) );
  AND2X1 U820 ( .A(r_regtrm[34]), .B(n70), .Y(REGTRM[34]) );
  AND2X1 U821 ( .A(r_regtrm[35]), .B(n70), .Y(REGTRM[35]) );
  AND2X1 U822 ( .A(r_regtrm[36]), .B(n70), .Y(REGTRM[36]) );
  AND2X1 U823 ( .A(r_regtrm[37]), .B(n70), .Y(REGTRM[37]) );
  AND2X1 U824 ( .A(r_regtrm[38]), .B(n70), .Y(REGTRM[38]) );
  AND2X1 U825 ( .A(r_regtrm[39]), .B(n70), .Y(REGTRM[39]) );
  AND2X1 U826 ( .A(r_regtrm[42]), .B(n69), .Y(REGTRM[42]) );
  AND2X1 U827 ( .A(r_regtrm[50]), .B(n68), .Y(REGTRM[50]) );
  AND2X1 U828 ( .A(r_aopt[0]), .B(n69), .Y(ANAOPT[0]) );
  AND2X1 U829 ( .A(r_aopt[2]), .B(n66), .Y(ANAOPT[2]) );
  AND2X1 U830 ( .A(r_aopt[6]), .B(n65), .Y(ANAOPT[6]) );
  AND2X1 U831 ( .A(r_aopt[7]), .B(n65), .Y(ANAOPT[7]) );
  AND2X1 U832 ( .A(r_accctl[3]), .B(n62), .Y(DO_DPDN[5]) );
  AND2X1 U833 ( .A(r_cvctl[6]), .B(n62), .Y(DO_CVCTL[6]) );
  AND2X1 U836 ( .A(r_cvctl[7]), .B(n62), .Y(DO_CVCTL[7]) );
  AND2X1 U837 ( .A(r_cvctl[5]), .B(n62), .Y(DO_CVCTL[5]) );
  AND2X1 U838 ( .A(r_ana_tm[0]), .B(n64), .Y(ANA_TM[0]) );
  AND2X1 U839 ( .A(r_ana_tm[1]), .B(n64), .Y(ANA_TM[1]) );
  AND2X1 U840 ( .A(r_ana_tm[2]), .B(n64), .Y(ANA_TM[2]) );
  AND2X1 U841 ( .A(r_ana_tm[3]), .B(n64), .Y(ANA_TM[3]) );
  AND2X1 U842 ( .A(r_cctrx[3]), .B(n63), .Y(DO_CCTRX[3]) );
  AND2X1 U843 ( .A(r_cvctl[2]), .B(n63), .Y(DO_CVCTL[2]) );
  AND2X1 U844 ( .A(r_xana_23), .B(n59), .Y(LFOSC_ENB) );
  AND2X1 U845 ( .A(r_dpdmctl[5]), .B(n62), .Y(DO_DPDN[2]) );
  AND2X1 U846 ( .A(r_xana[10]), .B(n65), .Y(ANA_REGX[10]) );
  AND2X1 U847 ( .A(r_xana[11]), .B(n65), .Y(ANA_REGX[11]) );
  AND2X1 U848 ( .A(r_cctrx[7]), .B(n63), .Y(DO_CCTRX[7]) );
  AND2X1 U849 ( .A(r_cctrx[6]), .B(n63), .Y(DO_CCTRX[6]) );
  AND2X1 U850 ( .A(r_cctrx[5]), .B(n63), .Y(DO_CCTRX[5]) );
  AND2X1 U851 ( .A(r_cctrx[4]), .B(n63), .Y(DO_CCTRX[4]) );
  AND2X1 U852 ( .A(r_xtm[2]), .B(n66), .Y(XTM[2]) );
  AND2X1 U853 ( .A(r_xtm[3]), .B(n66), .Y(XTM[3]) );
  AND2X1 U854 ( .A(r_cctrx[0]), .B(n63), .Y(DO_CCTRX[0]) );
  AND2X1 U855 ( .A(r_regtrm[24]), .B(n72), .Y(REGTRM[24]) );
  INVX3 U856 ( .A(n30), .Y(n31) );
  AO22XL U857 ( .A(iram_a[6]), .B(iram_ce), .C(xram_a[6]), .D(xram_ce), .Y(
        SRAM_A[6]) );
  INVXL U858 ( .A(n32), .Y(n33) );
endmodule


module SNPS_CLOCK_GATE_HIGH_core_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_1 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o, test_si, 
        test_se );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we, test_si, test_se;
  output pwm_o;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, net8849, n1, n2, n3, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n29, n30, n31, n32, n33, n34,
         n35;
  wire   [6:0] pwmcnt;

  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  glreg_a0_1 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm), .test_si(pwmcnt[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8849), .TE(test_se) );
  SDFFSQX1 pwmcnt_reg_6_ ( .D(N20), .SIN(pwmcnt[5]), .SMC(test_se), .C(net8849), .XS(n2), .Q(pwmcnt[6]) );
  SDFFSQX1 pwmcnt_reg_4_ ( .D(N18), .SIN(pwmcnt[3]), .SMC(test_se), .C(net8849), .XS(n2), .Q(pwmcnt[4]) );
  SDFFSQX1 pwmcnt_reg_5_ ( .D(N19), .SIN(pwmcnt[4]), .SMC(test_se), .C(net8849), .XS(n2), .Q(pwmcnt[5]) );
  SDFFSQX1 pwmcnt_reg_2_ ( .D(N16), .SIN(pwmcnt[1]), .SMC(test_se), .C(net8849), .XS(n2), .Q(pwmcnt[2]) );
  SDFFSQX1 pwmcnt_reg_3_ ( .D(N17), .SIN(pwmcnt[2]), .SMC(test_se), .C(net8849), .XS(n2), .Q(pwmcnt[3]) );
  SDFFSQX1 pwmcnt_reg_1_ ( .D(N15), .SIN(pwmcnt[0]), .SMC(test_se), .C(net8849), .XS(n1), .Q(pwmcnt[1]) );
  SDFFSQX1 pwmcnt_reg_0_ ( .D(N14), .SIN(test_si), .SMC(test_se), .C(net8849), 
        .XS(n1), .Q(pwmcnt[0]) );
  INVX1 U6 ( .A(n4), .Y(n14) );
  NAND21X1 U7 ( .B(wdat[7]), .A(we), .Y(n4) );
  INVX1 U8 ( .A(n27), .Y(n18) );
  INVX1 U9 ( .A(n30), .Y(n10) );
  INVX1 U10 ( .A(n8), .Y(n9) );
  INVX1 U11 ( .A(n12), .Y(n7) );
  INVX1 U12 ( .A(n6), .Y(n11) );
  GEN2XL U13 ( .D(pwmcnt[0]), .E(pwmcnt[1]), .C(n10), .B(r_pwm[7]), .A(n14), 
        .Y(N15) );
  GEN2XL U14 ( .D(pwmcnt[5]), .E(n6), .C(n13), .B(r_pwm[7]), .A(n14), .Y(N19)
         );
  GEN2XL U15 ( .D(pwmcnt[3]), .E(n8), .C(n7), .B(r_pwm[7]), .A(n14), .Y(N17)
         );
  GEN2XL U16 ( .D(pwmcnt[4]), .E(n12), .C(n11), .B(r_pwm[7]), .A(n14), .Y(N18)
         );
  GEN2XL U17 ( .D(pwmcnt[2]), .E(n30), .C(n9), .B(r_pwm[7]), .A(n14), .Y(N16)
         );
  AO21X1 U18 ( .B(r_pwm[7]), .C(n29), .A(n14), .Y(N14) );
  AO21X1 U19 ( .B(r_pwm[7]), .C(n15), .A(n14), .Y(N20) );
  XOR2X1 U20 ( .A(pwmcnt[6]), .B(n13), .Y(n15) );
  OR2X1 U21 ( .A(n14), .B(r_pwm[7]), .Y(N13) );
  OR2X1 U22 ( .A(pwmcnt[0]), .B(pwmcnt[1]), .Y(n30) );
  OAI221X1 U23 ( .A(n19), .B(n20), .C(pwmcnt[6]), .D(n16), .E(n21), .Y(pwm_o)
         );
  AOI32X1 U24 ( .A(n22), .B(n31), .C(r_pwm[4]), .D(r_pwm[5]), .E(n35), .Y(n20)
         );
  OAI211X1 U25 ( .C(r_pwm[4]), .D(n31), .A(n22), .B(n23), .Y(n21) );
  INVX1 U26 ( .A(pwmcnt[4]), .Y(n31) );
  NOR2X1 U27 ( .A(n34), .B(r_pwm[3]), .Y(n27) );
  AOI211X1 U28 ( .C(n30), .D(n17), .A(n27), .B(n28), .Y(n26) );
  INVX1 U29 ( .A(r_pwm[1]), .Y(n17) );
  AOI21X1 U30 ( .B(r_pwm[1]), .C(n32), .A(r_pwm[0]), .Y(n28) );
  AOI21X1 U31 ( .B(n24), .C(n25), .A(n19), .Y(n23) );
  AOI32X1 U32 ( .A(n18), .B(n33), .C(r_pwm[2]), .D(r_pwm[3]), .E(n34), .Y(n24)
         );
  OAI221X1 U33 ( .A(n29), .B(n32), .C(r_pwm[2]), .D(n33), .E(n26), .Y(n25) );
  INVX1 U34 ( .A(pwmcnt[2]), .Y(n33) );
  INVX1 U35 ( .A(pwmcnt[1]), .Y(n32) );
  INVX1 U36 ( .A(pwmcnt[3]), .Y(n34) );
  AND2X1 U37 ( .A(pwmcnt[6]), .B(n16), .Y(n19) );
  INVX1 U38 ( .A(pwmcnt[0]), .Y(n29) );
  INVX1 U39 ( .A(r_pwm[6]), .Y(n16) );
  NAND21X1 U40 ( .B(r_pwm[5]), .A(pwmcnt[5]), .Y(n22) );
  INVX1 U41 ( .A(pwmcnt[5]), .Y(n35) );
  NAND21X1 U42 ( .B(pwmcnt[2]), .A(n10), .Y(n8) );
  NAND21X1 U43 ( .B(pwmcnt[3]), .A(n9), .Y(n12) );
  NAND21X1 U44 ( .B(pwmcnt[4]), .A(n7), .Y(n6) );
  INVX1 U45 ( .A(n5), .Y(n13) );
  NAND21X1 U46 ( .B(pwmcnt[5]), .A(n11), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8867;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8867), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8867), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8867), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8867), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8867), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8867), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8867), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8867), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8867), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_0 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o, test_si, 
        test_se );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we, test_si, test_se;
  output pwm_o;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, net8885, n1, n2, n3, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n29, n30, n31, n32, n33, n34,
         n35;
  wire   [6:0] pwmcnt;

  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  glreg_a0_0 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm), .test_si(pwmcnt[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8885), .TE(test_se) );
  SDFFSQX1 pwmcnt_reg_6_ ( .D(N20), .SIN(pwmcnt[5]), .SMC(test_se), .C(net8885), .XS(n2), .Q(pwmcnt[6]) );
  SDFFSQX1 pwmcnt_reg_4_ ( .D(N18), .SIN(pwmcnt[3]), .SMC(test_se), .C(net8885), .XS(n2), .Q(pwmcnt[4]) );
  SDFFSQX1 pwmcnt_reg_5_ ( .D(N19), .SIN(pwmcnt[4]), .SMC(test_se), .C(net8885), .XS(n2), .Q(pwmcnt[5]) );
  SDFFSQX1 pwmcnt_reg_2_ ( .D(N16), .SIN(pwmcnt[1]), .SMC(test_se), .C(net8885), .XS(n2), .Q(pwmcnt[2]) );
  SDFFSQX1 pwmcnt_reg_3_ ( .D(N17), .SIN(pwmcnt[2]), .SMC(test_se), .C(net8885), .XS(n2), .Q(pwmcnt[3]) );
  SDFFSQX1 pwmcnt_reg_1_ ( .D(N15), .SIN(pwmcnt[0]), .SMC(test_se), .C(net8885), .XS(n1), .Q(pwmcnt[1]) );
  SDFFSQX1 pwmcnt_reg_0_ ( .D(N14), .SIN(test_si), .SMC(test_se), .C(net8885), 
        .XS(n1), .Q(pwmcnt[0]) );
  INVX1 U6 ( .A(n4), .Y(n14) );
  NAND21X1 U7 ( .B(wdat[7]), .A(we), .Y(n4) );
  INVX1 U8 ( .A(n27), .Y(n18) );
  INVX1 U9 ( .A(n30), .Y(n10) );
  INVX1 U10 ( .A(n8), .Y(n9) );
  INVX1 U11 ( .A(n12), .Y(n7) );
  INVX1 U12 ( .A(n6), .Y(n11) );
  GEN2XL U13 ( .D(pwmcnt[0]), .E(pwmcnt[1]), .C(n10), .B(r_pwm[7]), .A(n14), 
        .Y(N15) );
  GEN2XL U14 ( .D(pwmcnt[5]), .E(n6), .C(n13), .B(r_pwm[7]), .A(n14), .Y(N19)
         );
  GEN2XL U15 ( .D(pwmcnt[3]), .E(n8), .C(n7), .B(r_pwm[7]), .A(n14), .Y(N17)
         );
  GEN2XL U16 ( .D(pwmcnt[4]), .E(n12), .C(n11), .B(r_pwm[7]), .A(n14), .Y(N18)
         );
  GEN2XL U17 ( .D(pwmcnt[2]), .E(n30), .C(n9), .B(r_pwm[7]), .A(n14), .Y(N16)
         );
  AO21X1 U18 ( .B(r_pwm[7]), .C(n29), .A(n14), .Y(N14) );
  AO21X1 U19 ( .B(r_pwm[7]), .C(n15), .A(n14), .Y(N20) );
  XOR2X1 U20 ( .A(pwmcnt[6]), .B(n13), .Y(n15) );
  OR2X1 U21 ( .A(n14), .B(r_pwm[7]), .Y(N13) );
  OR2X1 U22 ( .A(pwmcnt[0]), .B(pwmcnt[1]), .Y(n30) );
  NOR2X1 U23 ( .A(n34), .B(r_pwm[3]), .Y(n27) );
  AOI211X1 U24 ( .C(n30), .D(n17), .A(n27), .B(n28), .Y(n26) );
  INVX1 U25 ( .A(r_pwm[1]), .Y(n17) );
  AOI21X1 U26 ( .B(r_pwm[1]), .C(n32), .A(r_pwm[0]), .Y(n28) );
  AOI21X1 U27 ( .B(n24), .C(n25), .A(n19), .Y(n23) );
  AOI32X1 U28 ( .A(n18), .B(n33), .C(r_pwm[2]), .D(r_pwm[3]), .E(n34), .Y(n24)
         );
  OAI221X1 U29 ( .A(n29), .B(n32), .C(r_pwm[2]), .D(n33), .E(n26), .Y(n25) );
  INVX1 U30 ( .A(pwmcnt[2]), .Y(n33) );
  INVX1 U31 ( .A(pwmcnt[1]), .Y(n32) );
  OAI221X1 U32 ( .A(n19), .B(n20), .C(pwmcnt[6]), .D(n16), .E(n21), .Y(pwm_o)
         );
  AOI32X1 U33 ( .A(n22), .B(n31), .C(r_pwm[4]), .D(r_pwm[5]), .E(n35), .Y(n20)
         );
  OAI211X1 U34 ( .C(r_pwm[4]), .D(n31), .A(n22), .B(n23), .Y(n21) );
  INVX1 U35 ( .A(pwmcnt[3]), .Y(n34) );
  AND2X1 U36 ( .A(pwmcnt[6]), .B(n16), .Y(n19) );
  INVX1 U37 ( .A(pwmcnt[0]), .Y(n29) );
  INVX1 U38 ( .A(r_pwm[6]), .Y(n16) );
  NAND21X1 U39 ( .B(r_pwm[5]), .A(pwmcnt[5]), .Y(n22) );
  INVX1 U40 ( .A(pwmcnt[5]), .Y(n35) );
  INVX1 U41 ( .A(pwmcnt[4]), .Y(n31) );
  NAND21X1 U42 ( .B(pwmcnt[2]), .A(n10), .Y(n8) );
  NAND21X1 U43 ( .B(pwmcnt[3]), .A(n9), .Y(n12) );
  NAND21X1 U44 ( .B(pwmcnt[4]), .A(n7), .Y(n6) );
  INVX1 U45 ( .A(n5), .Y(n13) );
  NAND21X1 U46 ( .B(pwmcnt[5]), .A(n11), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8903;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8903), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8903), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8903), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8903), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8903), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8903), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8903), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8903), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8903), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module divclk_a0 ( mclk, srstz, atpg_en, clk_1500k, clk_500k, clk_100k, 
        clk_50k, clk_500, divff_8, divff_5, test_si, test_se );
  input mclk, srstz, atpg_en, test_si, test_se;
  output clk_1500k, clk_500k, clk_100k, clk_50k, clk_500, divff_8, divff_5;
  wire   div100k_2, N11, N12, N17, N18, N24, N25, N26, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, n7, n8, n9, n10, n1, n2,
         n3, n11, n12, n13, n4, n5, n6;
  wire   [1:0] div8;
  wire   [1:0] div500k_5;
  wire   [1:0] div1p5m_3;
  wire   [6:0] div50k_100;

  CLKDLX1 U0_D1P5M_ICG ( .CK(mclk), .E(n7), .SE(atpg_en), .ECK(clk_1500k) );
  CLKDLX1 U0_D500K_ICG ( .CK(clk_1500k), .E(n8), .SE(atpg_en), .ECK(clk_500k)
         );
  CLKDLX1 U0_D100K_ICG ( .CK(clk_500k), .E(n9), .SE(atpg_en), .ECK(clk_100k)
         );
  CLKDLX1 U0_D50K_ICG ( .CK(clk_100k), .E(div100k_2), .SE(atpg_en), .ECK(
        clk_50k) );
  CLKDLX1 U0_D0P5K_ICG ( .CK(clk_50k), .E(n10), .SE(atpg_en), .ECK(clk_500) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(srstz), .Y(n3) );
  divclk_a0_DW01_inc_0 add_48 ( .A(div50k_100), .SUM({N39, N38, N37, N36, N35, 
        N34, N33}) );
  SDFFRQX1 div1p5m_3_reg_1_ ( .D(N18), .SIN(div1p5m_3[0]), .SMC(test_se), .C(
        clk_1500k), .XR(n1), .Q(div1p5m_3[1]) );
  SDFFRQX1 div1p5m_3_reg_0_ ( .D(N17), .SIN(test_si), .SMC(test_se), .C(
        clk_1500k), .XR(n1), .Q(div1p5m_3[0]) );
  SDFFRQX1 div100k_2_reg ( .D(n4), .SIN(div50k_100[6]), .SMC(test_se), .C(
        clk_100k), .XR(n1), .Q(div100k_2) );
  SDFFRQX1 div50k_100_reg_6_ ( .D(N46), .SIN(div50k_100[5]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[6]) );
  SDFFRQX1 div50k_100_reg_5_ ( .D(N45), .SIN(div50k_100[4]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[5]) );
  SDFFRQX1 div50k_100_reg_4_ ( .D(N44), .SIN(div50k_100[3]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[4]) );
  SDFFRQX1 div50k_100_reg_3_ ( .D(N43), .SIN(div50k_100[2]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[3]) );
  SDFFRQX1 div500k_5_reg_0_ ( .D(N24), .SIN(div100k_2), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(div500k_5[0]) );
  SDFFRQX1 div8_reg_1_ ( .D(N11), .SIN(div8[0]), .SMC(test_se), .C(mclk), .XR(
        n1), .Q(div8[1]) );
  SDFFRQX1 div500k_5_reg_1_ ( .D(N25), .SIN(div500k_5[0]), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(div500k_5[1]) );
  SDFFRQX1 div8_reg_0_ ( .D(n5), .SIN(div1p5m_3[1]), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(div8[0]) );
  SDFFRQX1 div50k_100_reg_1_ ( .D(N41), .SIN(div50k_100[0]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[1]) );
  SDFFRQX1 div50k_100_reg_2_ ( .D(N42), .SIN(div50k_100[1]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[2]) );
  SDFFRQX1 div50k_100_reg_0_ ( .D(N40), .SIN(divff_8), .SMC(test_se), .C(
        clk_50k), .XR(n1), .Q(div50k_100[0]) );
  SDFFRQX1 div500k_5_reg_2_ ( .D(N26), .SIN(div500k_5[1]), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(divff_5) );
  SDFFRQX1 div8_reg_2_ ( .D(N12), .SIN(div8[1]), .SMC(test_se), .C(mclk), .XR(
        n1), .Q(divff_8) );
  NOR21XL U6 ( .B(N35), .A(n10), .Y(N42) );
  NOR21XL U7 ( .B(N36), .A(n10), .Y(N43) );
  NOR21XL U8 ( .B(N34), .A(n10), .Y(N41) );
  NOR21XL U9 ( .B(N37), .A(n10), .Y(N44) );
  NOR21XL U10 ( .B(N38), .A(n10), .Y(N45) );
  AND4X1 U11 ( .A(div50k_100[5]), .B(div50k_100[1]), .C(div50k_100[6]), .D(n12), .Y(n10) );
  NOR41XL U12 ( .D(div50k_100[0]), .A(div50k_100[4]), .B(div50k_100[3]), .C(
        div50k_100[2]), .Y(n12) );
  NOR21XL U13 ( .B(N33), .A(n10), .Y(N40) );
  NOR21XL U14 ( .B(N39), .A(n10), .Y(N46) );
  XNOR2XL U15 ( .A(n6), .B(div500k_5[0]), .Y(N25) );
  XNOR2XL U16 ( .A(divff_8), .B(n13), .Y(N12) );
  NAND2X1 U17 ( .A(div8[1]), .B(div8[0]), .Y(n13) );
  ENOX1 U18 ( .A(divff_5), .B(n11), .C(N25), .D(divff_5), .Y(N26) );
  INVX1 U19 ( .A(div500k_5[1]), .Y(n6) );
  NOR32XL U20 ( .B(divff_5), .C(n11), .A(N25), .Y(n9) );
  NOR32XL U21 ( .B(divff_8), .C(n5), .A(div8[1]), .Y(n7) );
  NOR21XL U22 ( .B(div1p5m_3[0]), .A(div1p5m_3[1]), .Y(N18) );
  NOR21XL U23 ( .B(div1p5m_3[1]), .A(div1p5m_3[0]), .Y(n8) );
  XNOR2XL U24 ( .A(n5), .B(div8[1]), .Y(N11) );
  AOI21X1 U25 ( .B(divff_5), .C(n6), .A(div500k_5[0]), .Y(N24) );
  INVX1 U26 ( .A(div8[0]), .Y(n5) );
  NAND2X1 U27 ( .A(div500k_5[1]), .B(div500k_5[0]), .Y(n11) );
  NOR2X1 U28 ( .A(div1p5m_3[1]), .B(div1p5m_3[0]), .Y(N17) );
  INVX1 U29 ( .A(div100k_2), .Y(n4) );
endmodule


module divclk_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module srambist_a0 ( clk, srstz, reg_hit, reg_w, reg_r, reg_wdat, iram_rdat, 
        xram_rdat, bist_en, bist_xram, bist_wr, bist_adr, bist_wdat, o_bistctl, 
        o_bistdat, test_si, test_se );
  input [1:0] reg_hit;
  input [7:0] reg_wdat;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  output [10:0] bist_adr;
  output [7:0] bist_wdat;
  output [6:0] o_bistctl;
  output [7:0] o_bistdat;
  input clk, srstz, reg_w, reg_r, test_si, test_se;
  output bist_en, bist_xram, bist_wr;
  wire   we_1_, bistctl_re, N21, busy_dly, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, r_bistfault, upd_fault, wd_fault, net8921, n110, n111, n10,
         n11, n12, n13, n28, n29, n30, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n87, n88, n3, n4, n6, n7, n9, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n31, n32, n86, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140;
  wire   [1:0] rw_sta;

  INVX1 U11 ( .A(n13), .Y(n11) );
  INVX1 U12 ( .A(n13), .Y(n12) );
  INVX1 U13 ( .A(n13), .Y(n10) );
  INVX1 U14 ( .A(srstz), .Y(n13) );
  INVX8 U151 ( .A(n11), .Y(n28) );
  INVX8 U152 ( .A(n10), .Y(n29) );
  glreg_WIDTH1_0 u0_bistfault ( .clk(clk), .arstz(n11), .we(upd_fault), .wdat(
        wd_fault), .rdat(o_bistctl[3]), .test_si(o_bistdat[7]), .test_se(
        test_se) );
  glreg_WIDTH5_1 u0_bistctl ( .clk(clk), .arstz(n11), .we(n30), .wdat({
        reg_wdat[6:4], reg_wdat[2], n9}), .rdat({o_bistctl[6:4], 
        o_bistctl[2:1]}), .test_si(rw_sta[1]), .test_se(test_se) );
  glreg_a0_6 u0_bistdat ( .clk(clk), .arstz(n10), .we(we_1_), .wdat({
        reg_wdat[7:2], n9, reg_wdat[0]}), .rdat(o_bistdat), .test_si(
        o_bistctl[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_srambist_a0 clk_gate_adr_reg ( .CLK(clk), .EN(N86), 
        .ENCLK(net8921), .TE(test_se) );
  srambist_a0_DW01_inc_0 add_65 ( .A(bist_adr), .SUM({N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64}) );
  SDFFQX1 busy_dly_reg ( .D(o_bistctl[0]), .SIN(bistctl_re), .SMC(test_se), 
        .C(clk), .Q(busy_dly) );
  SDFFQX1 r_bistfault_reg ( .D(n110), .SIN(busy_dly), .SMC(test_se), .C(clk), 
        .Q(r_bistfault) );
  SDFFRQX1 bistctl_re_reg ( .D(N21), .SIN(bist_adr[10]), .SMC(test_se), .C(clk), .XR(n11), .Q(bistctl_re) );
  SDFFQX1 rw_sta_reg_1_ ( .D(n135), .SIN(rw_sta[0]), .SMC(test_se), .C(clk), 
        .Q(rw_sta[1]) );
  SDFFQX1 rw_sta_reg_0_ ( .D(n111), .SIN(r_bistfault), .SMC(test_se), .C(clk), 
        .Q(rw_sta[0]) );
  SDFFQX1 adr_reg_10_ ( .D(N97), .SIN(bist_adr[9]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[10]) );
  SDFFQX1 adr_reg_9_ ( .D(N96), .SIN(bist_adr[8]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[9]) );
  SDFFQX1 adr_reg_8_ ( .D(N95), .SIN(bist_adr[7]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[8]) );
  SDFFQX1 adr_reg_7_ ( .D(N94), .SIN(bist_adr[6]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[7]) );
  SDFFQX1 adr_reg_6_ ( .D(N93), .SIN(bist_adr[5]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[6]) );
  SDFFQX1 adr_reg_5_ ( .D(N92), .SIN(bist_adr[4]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[5]) );
  SDFFQX1 adr_reg_4_ ( .D(N91), .SIN(bist_adr[3]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[4]) );
  SDFFQX1 adr_reg_2_ ( .D(N89), .SIN(bist_adr[1]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[2]) );
  SDFFQX1 adr_reg_3_ ( .D(N90), .SIN(bist_adr[2]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[3]) );
  SDFFQX1 adr_reg_1_ ( .D(N88), .SIN(bist_adr[0]), .SMC(test_se), .C(net8921), 
        .Q(bist_adr[1]) );
  SDFFQX1 adr_reg_0_ ( .D(N87), .SIN(test_si), .SMC(test_se), .C(net8921), .Q(
        bist_adr[0]) );
  INVX1 U3 ( .A(1'b1), .Y(bist_xram) );
  NAND2X1 U5 ( .A(n24), .B(n21), .Y(n7) );
  INVX1 U6 ( .A(n7), .Y(n3) );
  INVX1 U7 ( .A(n7), .Y(n4) );
  INVX1 U8 ( .A(n138), .Y(bist_en) );
  INVX1 U9 ( .A(n22), .Y(n6) );
  INVX1 U10 ( .A(n19), .Y(n30) );
  NAND2X1 U15 ( .A(reg_hit[0]), .B(reg_w), .Y(n19) );
  AND2X1 U16 ( .A(reg_w), .B(reg_hit[1]), .Y(we_1_) );
  INVX1 U17 ( .A(n14), .Y(n9) );
  INVX1 U18 ( .A(n54), .Y(n128) );
  NAND21X1 U19 ( .B(n24), .A(n23), .Y(n106) );
  INVX1 U20 ( .A(n20), .Y(n21) );
  INVX1 U21 ( .A(n22), .Y(n116) );
  NAND21X1 U22 ( .B(n24), .A(n21), .Y(n22) );
  AND2X1 U23 ( .A(reg_r), .B(reg_hit[0]), .Y(N21) );
  INVX1 U24 ( .A(n118), .Y(n120) );
  INVX1 U25 ( .A(n94), .Y(n91) );
  INVX1 U26 ( .A(n26), .Y(n31) );
  INVX1 U27 ( .A(n104), .Y(n25) );
  INVX1 U28 ( .A(n100), .Y(n103) );
  INVX1 U29 ( .A(n107), .Y(n99) );
  INVX1 U30 ( .A(n32), .Y(n96) );
  INVX1 U31 ( .A(n97), .Y(n93) );
  INVX1 U32 ( .A(reg_wdat[1]), .Y(n14) );
  OAI21X1 U33 ( .B(n132), .C(n127), .A(n77), .Y(bist_wdat[0]) );
  NAND2X1 U34 ( .A(n132), .B(n127), .Y(n77) );
  INVX1 U35 ( .A(n82), .Y(n127) );
  XNOR2XL U36 ( .A(n132), .B(n84), .Y(bist_wdat[1]) );
  AOI21X1 U37 ( .B(n80), .C(n79), .A(n82), .Y(n84) );
  XNOR2XL U38 ( .A(iram_rdat[2]), .B(n56), .Y(n49) );
  AOI21X1 U39 ( .B(n54), .C(n129), .A(n55), .Y(n56) );
  NAND2X1 U40 ( .A(n79), .B(n125), .Y(n80) );
  AOI31X1 U41 ( .A(iram_rdat[7]), .B(n47), .C(n48), .D(n133), .Y(n43) );
  AOI21X1 U42 ( .B(n128), .C(n140), .A(n49), .Y(n48) );
  INVX1 U43 ( .A(n78), .Y(n125) );
  INVX1 U44 ( .A(o_bistctl[0]), .Y(n138) );
  XOR2X1 U45 ( .A(iram_rdat[1]), .B(n53), .Y(n47) );
  AOI21X1 U46 ( .B(n54), .C(n46), .A(n55), .Y(n53) );
  XNOR2XL U47 ( .A(n132), .B(n83), .Y(bist_wdat[2]) );
  AOI21X1 U48 ( .B(n80), .C(n125), .A(n82), .Y(n83) );
  XOR2X1 U49 ( .A(bist_wdat[3]), .B(iram_rdat[3]), .Y(n72) );
  XOR2X1 U50 ( .A(bist_wdat[2]), .B(iram_rdat[2]), .Y(n76) );
  OAI22AX1 U51 ( .D(n80), .C(n77), .A(n132), .B(n80), .Y(bist_wdat[4]) );
  XNOR2XL U52 ( .A(iram_rdat[6]), .B(n65), .Y(n57) );
  OAI22X1 U53 ( .A(n131), .B(n129), .C(n66), .D(n133), .Y(n65) );
  XNOR2XL U54 ( .A(iram_rdat[0]), .B(n64), .Y(n58) );
  NAND2X1 U55 ( .A(n131), .B(n62), .Y(n64) );
  INVX1 U56 ( .A(iram_rdat[4]), .Y(n140) );
  INVX1 U57 ( .A(iram_rdat[5]), .Y(n139) );
  NOR4XL U58 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(n68) );
  XOR2X1 U59 ( .A(bist_wdat[0]), .B(iram_rdat[0]), .Y(n70) );
  XNOR2XL U60 ( .A(bist_wdat[5]), .B(n139), .Y(n69) );
  XOR2X1 U61 ( .A(bist_wdat[6]), .B(iram_rdat[6]), .Y(n71) );
  NOR4XL U62 ( .A(n73), .B(n74), .C(n75), .D(n76), .Y(n67) );
  XNOR2XL U63 ( .A(n140), .B(bist_wdat[4]), .Y(n73) );
  XOR2X1 U64 ( .A(bist_wdat[1]), .B(iram_rdat[1]), .Y(n75) );
  XNOR2XL U65 ( .A(n132), .B(iram_rdat[7]), .Y(n74) );
  OAI22X1 U66 ( .A(n77), .B(n80), .C(n81), .D(n132), .Y(bist_wdat[3]) );
  NOR2X1 U67 ( .A(n82), .B(n80), .Y(n81) );
  OAI22X1 U68 ( .A(n77), .B(n125), .C(n78), .D(n132), .Y(bist_wdat[6]) );
  NAND2X1 U69 ( .A(n46), .B(n129), .Y(n54) );
  INVX1 U70 ( .A(n35), .Y(n136) );
  INVX1 U71 ( .A(n66), .Y(n129) );
  INVX1 U72 ( .A(n63), .Y(n131) );
  NAND31X1 U73 ( .C(n23), .A(n17), .B(n34), .Y(n20) );
  MUX2IX1 U74 ( .D0(rw_sta[1]), .D1(rw_sta[0]), .S(o_bistctl[2]), .Y(n17) );
  MUX2AXL U75 ( .D0(o_bistctl[1]), .D1(n14), .S(n30), .Y(n24) );
  NAND2X1 U76 ( .A(n106), .B(n12), .Y(n102) );
  AO21X1 U77 ( .B(N68), .C(n4), .A(n86), .Y(N91) );
  GEN2XL U78 ( .D(n32), .E(bist_adr[4]), .C(n31), .B(n116), .A(n102), .Y(n86)
         );
  AO21X1 U79 ( .B(N65), .C(n4), .A(n92), .Y(N88) );
  GEN2XL U80 ( .D(bist_adr[0]), .E(bist_adr[1]), .C(n91), .B(n116), .A(n102), 
        .Y(n92) );
  AO21X1 U81 ( .B(N67), .C(n4), .A(n98), .Y(N90) );
  GEN2XL U82 ( .D(n97), .E(bist_adr[3]), .C(n96), .B(n116), .A(n102), .Y(n98)
         );
  AO21X1 U83 ( .B(n116), .C(n90), .A(n89), .Y(N87) );
  INVX1 U84 ( .A(bist_adr[0]), .Y(n90) );
  AO21X1 U85 ( .B(N64), .C(n3), .A(n102), .Y(n89) );
  AO21X1 U86 ( .B(N74), .C(n4), .A(n114), .Y(N97) );
  AO21X1 U87 ( .B(n113), .C(n116), .A(n112), .Y(n114) );
  XOR2X1 U88 ( .A(bist_adr[10]), .B(n117), .Y(n113) );
  AO21X1 U89 ( .B(N69), .C(n4), .A(n27), .Y(N92) );
  GEN2XL U90 ( .D(bist_adr[5]), .E(n26), .C(n25), .B(n116), .A(n102), .Y(n27)
         );
  AO21X1 U91 ( .B(N66), .C(n4), .A(n95), .Y(N89) );
  GEN2XL U92 ( .D(bist_adr[2]), .E(n94), .C(n93), .B(n6), .A(n102), .Y(n95) );
  AO21X1 U93 ( .B(N71), .C(n4), .A(n101), .Y(N94) );
  GEN2XL U94 ( .D(bist_adr[7]), .E(n100), .C(n99), .B(n116), .A(n102), .Y(n101) );
  AO21X1 U95 ( .B(N70), .C(n4), .A(n105), .Y(N93) );
  GEN2XL U96 ( .D(bist_adr[6]), .E(n104), .C(n103), .B(n116), .A(n102), .Y(
        n105) );
  AO21X1 U97 ( .B(N72), .C(n4), .A(n108), .Y(N95) );
  GEN2XL U98 ( .D(bist_adr[8]), .E(n107), .C(n120), .B(n116), .A(n112), .Y(
        n108) );
  AO21X1 U99 ( .B(N73), .C(n4), .A(n119), .Y(N96) );
  GEN2XL U100 ( .D(bist_adr[9]), .E(n118), .C(n117), .B(n116), .A(n115), .Y(
        n119) );
  INVX1 U101 ( .A(n16), .Y(n23) );
  NAND43X1 U102 ( .B(o_bistdat[6]), .C(n19), .D(n15), .A(o_bistdat[7]), .Y(n16) );
  INVX1 U103 ( .A(reg_wdat[0]), .Y(n15) );
  NAND21X1 U104 ( .B(n29), .A(n106), .Y(n112) );
  NAND32X1 U105 ( .B(n23), .C(n18), .A(n20), .Y(N86) );
  NOR4XL U106 ( .A(n87), .B(n88), .C(n123), .D(n124), .Y(n85) );
  INVX1 U107 ( .A(bist_adr[3]), .Y(n123) );
  INVX1 U108 ( .A(bist_adr[4]), .Y(n124) );
  OR2X1 U109 ( .A(bist_adr[0]), .B(bist_adr[1]), .Y(n94) );
  NAND21X1 U110 ( .B(bist_adr[4]), .A(n96), .Y(n26) );
  NAND21X1 U111 ( .B(bist_adr[3]), .A(n93), .Y(n32) );
  NAND21X1 U112 ( .B(bist_adr[8]), .A(n99), .Y(n118) );
  NAND21X1 U113 ( .B(bist_adr[5]), .A(n31), .Y(n104) );
  NAND21X1 U114 ( .B(bist_adr[6]), .A(n25), .Y(n100) );
  NAND21X1 U115 ( .B(bist_adr[7]), .A(n103), .Y(n107) );
  NAND21X1 U116 ( .B(bist_adr[2]), .A(n91), .Y(n97) );
  NAND4X1 U117 ( .A(bist_adr[8]), .B(bist_adr[7]), .C(bist_adr[6]), .D(
        bist_adr[5]), .Y(n87) );
  NAND3X1 U118 ( .A(bist_adr[1]), .B(bist_adr[0]), .C(bist_adr[2]), .Y(n88) );
  NOR2X1 U119 ( .A(o_bistdat[2]), .B(o_bistdat[3]), .Y(n82) );
  INVX1 U120 ( .A(o_bistdat[5]), .Y(n132) );
  NOR2X1 U121 ( .A(n126), .B(o_bistdat[3]), .Y(n78) );
  OAI22X1 U122 ( .A(o_bistdat[4]), .B(n50), .C(n128), .D(n51), .Y(n42) );
  XNOR2XL U123 ( .A(n131), .B(n140), .Y(n51) );
  NOR32XL U124 ( .B(n52), .C(n49), .A(n47), .Y(n50) );
  AOI21X1 U125 ( .B(iram_rdat[4]), .C(n128), .A(iram_rdat[7]), .Y(n52) );
  NOR42XL U126 ( .C(n122), .D(n12), .A(n121), .B(n40), .Y(n39) );
  NOR4XL U127 ( .A(n41), .B(n42), .C(n43), .D(n44), .Y(n40) );
  XNOR2XL U128 ( .A(n45), .B(n139), .Y(n44) );
  NAND3X1 U129 ( .A(n57), .B(n58), .C(n59), .Y(n41) );
  INVX1 U130 ( .A(o_bistdat[2]), .Y(n126) );
  NAND2X1 U131 ( .A(o_bistdat[3]), .B(n126), .Y(n79) );
  ENOX1 U132 ( .A(bistctl_re), .B(n37), .C(wd_fault), .D(srstz), .Y(n110) );
  AOI31X1 U133 ( .A(busy_dly), .B(n137), .C(n38), .D(n39), .Y(n37) );
  INVX1 U134 ( .A(n34), .Y(n137) );
  AOI211X1 U135 ( .C(n67), .D(n68), .A(n134), .B(n28), .Y(n38) );
  NOR3XL U136 ( .A(n138), .B(rw_sta[1]), .C(n121), .Y(bist_wr) );
  XNOR2XL U137 ( .A(iram_rdat[3]), .B(n60), .Y(n59) );
  NAND2X1 U138 ( .A(n61), .B(n62), .Y(n60) );
  OAI22X1 U139 ( .A(o_bistdat[4]), .B(n128), .C(n63), .D(n54), .Y(n61) );
  ENOX1 U140 ( .A(n77), .B(n79), .C(n79), .D(o_bistdat[5]), .Y(bist_wdat[5])
         );
  OAI21X1 U141 ( .B(n138), .C(n36), .A(n12), .Y(n35) );
  NOR2X1 U142 ( .A(n121), .B(n122), .Y(n36) );
  NOR2X1 U143 ( .A(n130), .B(o_bistdat[1]), .Y(n66) );
  INVX1 U144 ( .A(rw_sta[0]), .Y(n121) );
  INVX1 U145 ( .A(o_bistdat[0]), .Y(n130) );
  NAND2X1 U146 ( .A(o_bistdat[1]), .B(n130), .Y(n46) );
  INVX1 U147 ( .A(n33), .Y(n135) );
  AOI32X1 U148 ( .A(o_bistctl[2]), .B(bist_wr), .C(n11), .D(rw_sta[1]), .E(
        n136), .Y(n33) );
  NOR2X1 U149 ( .A(n55), .B(o_bistdat[4]), .Y(n63) );
  NOR2X1 U150 ( .A(o_bistdat[0]), .B(o_bistdat[1]), .Y(n55) );
  OAI32X1 U153 ( .A(n34), .B(n136), .C(n28), .D(n121), .E(n35), .Y(n111) );
  ENOX1 U154 ( .A(n131), .B(n46), .C(n46), .D(o_bistdat[4]), .Y(n45) );
  NAND2X1 U155 ( .A(n55), .B(o_bistdat[4]), .Y(n62) );
  INVX1 U157 ( .A(n109), .Y(n117) );
  NAND21X1 U158 ( .B(bist_adr[9]), .A(n120), .Y(n109) );
  INVX1 U159 ( .A(o_bistdat[4]), .Y(n133) );
  NAND21X1 U160 ( .B(rw_sta[1]), .A(n121), .Y(n34) );
  OR2X1 U161 ( .A(bistctl_re), .B(r_bistfault), .Y(upd_fault) );
  INVX1 U162 ( .A(o_bistctl[2]), .Y(n134) );
  INVX1 U163 ( .A(rw_sta[1]), .Y(n122) );
  NOR21XL U164 ( .B(r_bistfault), .A(bistctl_re), .Y(wd_fault) );
  OAI211X1 U165 ( .C(n85), .D(n120), .A(bist_adr[10]), .B(bist_adr[9]), .Y(
        o_bistctl[0]) );
  BUFX3 U166 ( .A(o_bistdat[5]), .Y(bist_wdat[7]) );
  INVX8 U167 ( .A(n11), .Y(n18) );
  INVX8 U168 ( .A(srstz), .Y(n115) );
endmodule


module srambist_a0_DW01_inc_0 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_srambist_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_6 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8939;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8939), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8939), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8939), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8939), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8939), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8939), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8939), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8939), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8939), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8957;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8957), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8957), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8957), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8957), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8957), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8957), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module regx_a0 ( regx_r, regx_w, di_drposc, di_imposc, di_rd_det, di_stbovp, 
        clk_500k, r_imp_osc, regx_addr, regx_wdat, regx_rdat, regx_hitbst, 
        regx_wrpwm, regx_wrcvc, r_sdischg, r_bistctl, r_bistdat, r_vcomp, 
        r_idacsh, r_cvofsx, r_pwm, regx_wrdac, dac_r_vs, dac_comp, r_dac_en, 
        r_sar_en, r_aopt, r_xtm, r_adummyi, r_bck0, r_bck1, r_i2crout, r_xana, 
        di_xana, lt_gpi, di_tst, bkpt_pc, bkpt_ena, we_twlb, r_vpp_en, 
        r_vpp0v_en, r_otp_pwdn_en, r_otp_wpls, wd_twlb, r_sap, r_twlb, 
        upd_pwrv, ramacc, sse_idle, bus_idle, r_do_ts, r_dpdo_sel, r_dndo_sel, 
        di_ts, detclk, aswclk, atpg_en, di_aswk, clk, rrstz, test_si2, 
        test_si1, test_so1, test_se );
  input [6:0] regx_addr;
  input [7:0] regx_wdat;
  output [7:0] regx_rdat;
  output [1:0] regx_hitbst;
  output [1:0] regx_wrpwm;
  output [3:0] regx_wrcvc;
  input [7:0] r_sdischg;
  input [6:0] r_bistctl;
  input [7:0] r_bistdat;
  input [7:0] r_vcomp;
  input [7:0] r_idacsh;
  input [7:0] r_cvofsx;
  input [15:0] r_pwm;
  output [13:0] regx_wrdac;
  input [79:0] dac_r_vs;
  input [9:0] dac_comp;
  input [9:0] r_dac_en;
  input [9:0] r_sar_en;
  output [7:0] r_aopt;
  output [7:0] r_xtm;
  output [7:0] r_adummyi;
  output [7:0] r_bck0;
  output [7:0] r_bck1;
  output [5:0] r_i2crout;
  output [23:0] r_xana;
  input [4:0] di_xana;
  input [3:0] lt_gpi;
  output [14:0] bkpt_pc;
  output [1:0] wd_twlb;
  output [1:0] r_sap;
  input [1:0] r_twlb;
  output [6:0] r_do_ts;
  output [3:0] r_dpdo_sel;
  output [3:0] r_dndo_sel;
  input [4:0] di_aswk;
  input regx_r, regx_w, di_drposc, di_imposc, di_rd_det, di_stbovp, clk_500k,
         di_tst, upd_pwrv, ramacc, sse_idle, bus_idle, di_ts, detclk, aswclk,
         atpg_en, clk, rrstz, test_si2, test_si1, test_se;
  output r_imp_osc, bkpt_ena, we_twlb, r_vpp_en, r_vpp0v_en, r_otp_pwdn_en,
         r_otp_wpls, test_so1;
  wire   we_19, we_7, we_5, we_4, reg1F_7, reg1F_6, reg1B_3_, reg10_7_, lt_drp,
         i2c_mode_upd, N8, d_we16, lt_reg1C_0, net8975, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n61, n74, n75, n76, n1, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151,
         SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153,
         SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155,
         SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157,
         SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159,
         SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161,
         SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163,
         SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165,
         SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167,
         SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169,
         SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171,
         SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173,
         SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175,
         SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177,
         SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179,
         SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181,
         SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183,
         SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185,
         SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187,
         SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189,
         SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191,
         SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193,
         SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195,
         SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197,
         SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199,
         SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201,
         SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203,
         SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205,
         SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207,
         SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209,
         SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211,
         SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213,
         SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215,
         SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217,
         SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219,
         SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221,
         SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223,
         SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225,
         SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227,
         SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229,
         SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231,
         SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233,
         SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235,
         SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237,
         SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239,
         SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241,
         SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243,
         SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245,
         SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247,
         SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249,
         SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251,
         SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253,
         SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255,
         SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257,
         SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259,
         SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261,
         SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263,
         SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265,
         SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267,
         SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269,
         SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271,
         SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273,
         SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275,
         SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277,
         SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279,
         SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281,
         SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283,
         SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285,
         SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287,
         SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289,
         SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291,
         SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293,
         SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295,
         SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297,
         SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299,
         SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301,
         SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303,
         SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305,
         SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307,
         SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309,
         SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311,
         SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313,
         SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315,
         SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317,
         SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319,
         SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321,
         SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323,
         SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325,
         SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327,
         SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329,
         SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331,
         SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333,
         SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335,
         SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337,
         SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339,
         SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341,
         SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343,
         SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345,
         SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347,
         SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349,
         SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351,
         SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353,
         SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355,
         SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357,
         SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359,
         SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361,
         SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363,
         SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365,
         SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367,
         SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369,
         SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371,
         SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373,
         SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375,
         SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377,
         SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379,
         SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381,
         SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383,
         SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385,
         SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387,
         SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389,
         SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391,
         SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393,
         SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395,
         SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397,
         SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399,
         SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401,
         SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403,
         SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405,
         SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407,
         SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409,
         SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411,
         SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413,
         SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415,
         SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417,
         SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419,
         SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421,
         SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423,
         SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425,
         SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427,
         SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429,
         SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431,
         SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433,
         SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435,
         SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437,
         SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439,
         SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441,
         SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443,
         SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445,
         SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447,
         SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449,
         SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451,
         SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453,
         SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455,
         SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457,
         SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459,
         SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461,
         SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463,
         SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465,
         SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467,
         SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469,
         SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471,
         SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473,
         SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475,
         SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477,
         SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479,
         SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481,
         SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483,
         SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485,
         SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487,
         SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489,
         SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491,
         SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493,
         SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495,
         SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497,
         SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499,
         SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501,
         SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503,
         SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505,
         SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507,
         SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509,
         SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511,
         SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513,
         SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515,
         SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517,
         SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519,
         SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521,
         SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523,
         SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525,
         SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527,
         SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529,
         SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531,
         SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533,
         SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535,
         SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537,
         SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539,
         SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541,
         SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543,
         SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545,
         SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547,
         SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549,
         SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551,
         SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553,
         SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555,
         SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557,
         SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559,
         SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561,
         SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563,
         SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565,
         SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567,
         SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569,
         SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571,
         SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573,
         SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575,
         SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577,
         SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579,
         SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581,
         SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583,
         SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585,
         SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587,
         SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589,
         SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591,
         SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593,
         SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595,
         SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597,
         SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599,
         SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601,
         SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603,
         SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605,
         SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607,
         SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609,
         SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611,
         SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613,
         SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615,
         SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617,
         SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619,
         SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621,
         SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623,
         SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625,
         SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627,
         SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629,
         SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631,
         SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633,
         SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635,
         SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637,
         SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639,
         SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641,
         SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643,
         SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645,
         SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647,
         SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649,
         SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651,
         SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653,
         SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655,
         SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657,
         SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659,
         SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661,
         SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663,
         SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665,
         SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667,
         SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669,
         SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671,
         SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673,
         SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675,
         SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677,
         SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679,
         SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681,
         SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683,
         SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685,
         SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687,
         SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689,
         SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691,
         SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693,
         SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695,
         SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697,
         SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699,
         SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701,
         SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703,
         SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705,
         SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707,
         SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709,
         SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711,
         SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713,
         SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715,
         SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717,
         SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719,
         SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721,
         SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723,
         SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725,
         SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727,
         SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729,
         SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731,
         SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733,
         SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735,
         SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737,
         SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739,
         SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741,
         SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743,
         SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745,
         SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747,
         SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749,
         SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751,
         SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753,
         SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755,
         SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757,
         SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759,
         SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761,
         SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763,
         SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765,
         SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767,
         SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769,
         SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771,
         SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773,
         SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775,
         SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777,
         SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779,
         SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781,
         SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783,
         SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785,
         SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787,
         SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789,
         SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791,
         SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793,
         SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795,
         SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797,
         SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799,
         SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801,
         SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803,
         SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805,
         SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807,
         SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809,
         SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811,
         SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813,
         SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815,
         SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817,
         SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819,
         SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821,
         SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823,
         SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825,
         SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827,
         SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829,
         SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831,
         SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833,
         SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835,
         SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837,
         SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839,
         SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841,
         SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843,
         SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845,
         SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847,
         SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849,
         SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851,
         SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853,
         SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855,
         SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857,
         SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859,
         SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861,
         SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863,
         SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865,
         SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867,
         SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869,
         SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871,
         SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873,
         SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875,
         SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877,
         SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879,
         SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881,
         SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883,
         SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885,
         SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887,
         SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889,
         SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891,
         SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893,
         SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895,
         SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897,
         SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899,
         SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901,
         SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903,
         SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905,
         SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907,
         SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909,
         SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911,
         SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913,
         SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915,
         SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917,
         SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919,
         SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921,
         SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923,
         SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925,
         SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927,
         SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929,
         SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931,
         SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933,
         SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935,
         SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937,
         SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939,
         SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941,
         SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943,
         SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945,
         SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947,
         SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949,
         SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951,
         SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953,
         SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955,
         SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957,
         SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959,
         SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961,
         SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963,
         SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965,
         SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967,
         SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969,
         SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971,
         SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973,
         SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975,
         SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977,
         SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979,
         SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981,
         SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983,
         SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985,
         SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987,
         SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989,
         SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991,
         SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993,
         SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995,
         SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997,
         SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999,
         SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001,
         SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003,
         SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005,
         SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007,
         SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009,
         SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011,
         SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013,
         SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015,
         SYNOPSYS_UNCONNECTED_1016;
  wire   [30:23] we;
  wire   [6:0] d_regx_addr;
  wire   [4:0] reg1F;
  wire   [3:2] reg1E;
  wire   [3:0] reg14;
  wire   [3:0] d_lt_gpi;
  wire   [5:0] lt_reg15_5_0;
  wire   [5:0] i2c_mode_wdat;
  wire   [5:0] d_lt_aswk;
  wire   [5:0] lt_aswk;
  wire   [7:0] wd18;

  INVX1 U73 ( .A(n58), .Y(n55) );
  INVX1 U74 ( .A(n58), .Y(n57) );
  INVX1 U75 ( .A(n59), .Y(n56) );
  INVX1 U76 ( .A(n58), .Y(n48) );
  INVX1 U77 ( .A(n59), .Y(n47) );
  INVX1 U78 ( .A(n58), .Y(n49) );
  INVX1 U79 ( .A(n59), .Y(n46) );
  INVX1 U80 ( .A(n59), .Y(n45) );
  INVX1 U81 ( .A(n58), .Y(n44) );
  INVX1 U82 ( .A(n59), .Y(n43) );
  INVX1 U83 ( .A(n60), .Y(n42) );
  INVX1 U84 ( .A(n58), .Y(n41) );
  INVX1 U85 ( .A(n59), .Y(n40) );
  INVX1 U86 ( .A(n58), .Y(n39) );
  INVX1 U87 ( .A(n60), .Y(n38) );
  INVX1 U88 ( .A(n58), .Y(n50) );
  INVX1 U89 ( .A(n58), .Y(n51) );
  INVX1 U90 ( .A(n59), .Y(n53) );
  INVX1 U91 ( .A(n58), .Y(n52) );
  INVX1 U92 ( .A(n59), .Y(n54) );
  INVX1 U94 ( .A(rrstz), .Y(n60) );
  INVX1 U95 ( .A(rrstz), .Y(n58) );
  INVX1 U96 ( .A(rrstz), .Y(n59) );
  glreg_a0_18 u0_reg04 ( .clk(clk), .arstz(n38), .we(we_4), .wdat({n13, n10, 
        n25, n22, n7, n19, wd_twlb[1], n16}), .rdat(r_bck0), .test_si(
        r_xana[23]), .test_se(test_se) );
  glreg_a0_17 u0_reg05 ( .clk(clk), .arstz(n39), .we(we_5), .wdat({n12, n10, 
        n25, n22, n7, n19, wd_twlb[1], n16}), .rdat(r_bck1), .test_si(
        r_bck0[7]), .test_se(test_se) );
  glreg_a0_16 u0_reg07 ( .clk(clk), .arstz(n40), .we(we_7), .wdat({n12, n9, 
        regx_wdat[5:4], n6, regx_wdat[2], wd_twlb[1], regx_wdat[0]}), .rdat(
        r_adummyi), .test_si(r_bck1[7]), .test_se(test_se) );
  glreg_WIDTH1_2 u0_reg10 ( .clk(clk), .arstz(n42), .we(1'b1), .wdat(ramacc), 
        .rdat(reg10_7_), .test_si(r_adummyi[7]), .test_se(test_se) );
  glreg_6_00000002 u0_reg12 ( .clk(clk), .arstz(n51), .we(we_twlb), .wdat({n13, 
        n10, n24, n21, n7, n18}), .rdat({r_vpp_en, r_vpp0v_en, r_otp_pwdn_en, 
        r_otp_wpls, r_sap}), .test_si(reg10_7_), .test_se(test_se) );
  glreg_a0_15 u0_reg13 ( .clk(clk), .arstz(n41), .we(we_19), .wdat({n13, n10, 
        n25, n22, n7, n19, wd_twlb}), .rdat({r_dpdo_sel, r_dndo_sel}), 
        .test_si(r_vpp_en), .test_se(test_se) );
  glreg_WIDTH6_1 u0_reg15 ( .clk(clk), .arstz(n55), .we(n76), .wdat({n25, n22, 
        n7, n19, wd_twlb[1], n16}), .rdat(lt_reg15_5_0), .test_si(
        r_dpdo_sel[3]), .test_se(test_se) );
  glreg_WIDTH6_0 u1_reg15 ( .clk(clk), .arstz(n54), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat(r_i2crout), .test_si(n114), .test_se(test_se) );
  glreg_a0_14 u0_reg17 ( .clk(clk), .arstz(n42), .we(we[23]), .wdat({n13, n10, 
        regx_wdat[5], n21, n7, regx_wdat[2], wd_twlb[1], n16}), .rdat(r_aopt), 
        .test_si(lt_reg15_5_0[5]), .test_se(test_se) );
  glreg_a0_13 u0_tmp18 ( .clk(clk), .arstz(n43), .we(we[24]), .wdat({n12, n9, 
        n24, n21, n6, n18, n63, wd_twlb[0]}), .rdat(wd18), .test_si(n116), 
        .test_se(test_se) );
  glreg_a0_12 u0_reg18 ( .clk(clk), .arstz(n44), .we(n75), .wdat(wd18), .rdat(
        bkpt_pc[7:0]), .test_si(r_aopt[7]), .test_se(test_se) );
  glreg_a0_11 u0_reg19 ( .clk(clk), .arstz(n45), .we(n75), .wdat({n13, n10, 
        n25, n22, n7, n19, n63, wd_twlb[0]}), .rdat({bkpt_ena, bkpt_pc[14:8]}), 
        .test_si(bkpt_pc[7]), .test_se(test_se) );
  glreg_a0_10 u0_reg1A ( .clk(clk), .arstz(n46), .we(we[26]), .wdat({n13, n10, 
        n25, n22, n7, n19, n63, n16}), .rdat(r_xtm), .test_si(n117), .test_se(
        test_se) );
  dbnc_WIDTH2_TIMEOUT2_7 u0_ts_db ( .o_dbc(reg1B_3_), .o_chg(), .i_org(di_ts), 
        .clk(clk), .rstz(n57), .test_si(wd18[7]), .test_so(n115), .test_se(
        test_se) );
  glreg_WIDTH7_0 u0_reg1B ( .clk(clk), .arstz(n50), .we(we[27]), .wdat({n13, 
        n10, n24, n22, n18, n63, n16}), .rdat(r_do_ts), .test_si(r_xtm[7]), 
        .test_se(test_se) );
  glreg_WIDTH1_1 u1_reg1C ( .clk(clk), .arstz(n38), .we(upd_pwrv), .wdat(
        lt_reg1C_0), .rdat(r_xana[0]), .test_si(test_si2), .test_se(test_se)
         );
  glreg_a0_9 u0_reg1C ( .clk(clk), .arstz(n49), .we(we[28]), .wdat({n12, n9, 
        n24, n21, n6, n18, n63, n16}), .rdat({r_xana[7:1], lt_reg1C_0}), 
        .test_si(r_do_ts[6]), .test_se(test_se) );
  glreg_a0_8 u0_reg1D ( .clk(clk), .arstz(n47), .we(we[29]), .wdat({n13, n10, 
        n25, n22, n6, n19, wd_twlb}), .rdat(r_xana[15:8]), .test_si(r_xana[7]), 
        .test_se(test_se) );
  glreg_a0_7 u0_reg1E ( .clk(clk), .arstz(n48), .we(we[30]), .wdat({n13, n10, 
        n25, n22, n7, n19, wd_twlb[1], n16}), .rdat({r_xana[23], r_imp_osc, 
        r_xana[21:20], reg1E, r_xana[17:16]}), .test_si(r_xana[15]), .test_se(
        test_se) );
  dbnc_WIDTH2_TIMEOUT2_6 u0_dosc_db ( .o_dbc(reg14[1]), .o_chg(), .i_org(
        di_imposc), .clk(clk), .rstz(n54), .test_si(lt_drp), .test_so(n119), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_5 u0_iosc_db ( .o_dbc(reg14[2]), .o_chg(), .i_org(
        di_drposc), .clk(clk), .rstz(n56), .test_si(n119), .test_so(n118), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_4 u0_xana_db ( .o_dbc(reg1F[0]), .o_chg(), .i_org(
        di_xana[0]), .clk(clk), .rstz(n57), .test_si(n115), .test_so(n114), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_3 u1_xana_db ( .o_dbc(reg1F[1]), .o_chg(), .i_org(
        di_xana[1]), .clk(clk), .rstz(rrstz), .test_si(r_i2crout[5]), 
        .test_so(n113), .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_2 u2_xana_db ( .o_dbc(reg1F[2]), .o_chg(), .i_org(
        di_xana[2]), .clk(clk), .rstz(n55), .test_si(n113), .test_so(n112), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_1 u3_xana_db ( .o_dbc(reg1F[3]), .o_chg(), .i_org(
        di_xana[3]), .clk(clk), .rstz(n56), .test_si(n112), .test_so(n111), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_0 u4_xana_db ( .o_dbc(reg1F[4]), .o_chg(), .i_org(
        di_xana[4]), .clk(clk), .rstz(n51), .test_si(n111), .test_so(test_so1), 
        .test_se(test_se) );
  dbnc_a0_1 u0_sbov_db ( .o_dbc(reg1F_6), .o_chg(), .i_org(di_stbovp), .clk(
        clk_500k), .rstz(n52), .test_si(bkpt_ena), .test_so(n116), .test_se(
        test_se) );
  dbnc_a0_0 u0_rdet_db ( .o_dbc(reg1F_7), .o_chg(), .i_org(di_rd_det), .clk(
        clk_500k), .rstz(n53), .test_si(n118), .test_so(n117), .test_se(
        test_se) );
  SNPS_CLOCK_GATE_HIGH_regx_a0 clk_gate_d_lt_gpi_reg ( .CLK(clk), .EN(n60), 
        .ENCLK(net8975), .TE(test_se) );
  regx_a0_DW_rightsh_0 srl_66 ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        dac_comp[9:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_sar_en[9:8], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_dac_en[9:8], 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_comp[7:0], r_sar_en[7:0], r_dac_en[7:0], dac_r_vs[63:0], 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_r_vs[79:64], reg1F_7, reg1F_6, 1'b0, reg1F, r_xana[23], r_imp_osc, 
        r_xana[21:20], reg1E, r_xana[17:0], r_do_ts[6:3], reg1B_3_, 
        r_do_ts[2:0], r_xtm, bkpt_ena, bkpt_pc, r_aopt, 1'b0, 1'b0, d_lt_aswk, 
        sse_idle, 1'b0, r_i2crout, d_lt_gpi, reg14, r_dpdo_sel, r_dndo_sel, 
        r_vpp_en, r_vpp0v_en, r_otp_pwdn_en, r_otp_wpls, r_sap, r_twlb, 
        r_bistdat, reg10_7_, r_bistctl, r_sdischg, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_pwm, r_adummyi, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_bck1, r_bck0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_cvofsx, r_idacsh, r_vcomp}), .DATA_TC(1'b0), .SH({d_regx_addr[6:4], 
        n29, n27, d_regx_addr[1:0], 1'b0, 1'b0, 1'b0}), .B({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, 
        SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, 
        SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, 
        SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, 
        SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, 
        SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, 
        SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, 
        SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, 
        SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, 
        SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, 
        SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, 
        SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, 
        SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, 
        SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, 
        SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, 
        SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, 
        SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, 
        SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, 
        SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, 
        SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, 
        SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, 
        SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, 
        SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, 
        SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, 
        SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, 
        SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, 
        SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, 
        SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, 
        SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, 
        SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, 
        SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, 
        SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, 
        SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, 
        SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, 
        SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, 
        SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, 
        SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, 
        SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, 
        SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, 
        SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, 
        SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, 
        SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, 
        SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, 
        SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, 
        SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, 
        SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, 
        SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, 
        SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, 
        SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, 
        SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, 
        SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, 
        SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, 
        SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, 
        SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, 
        SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, 
        SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, 
        SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, 
        SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, 
        SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, 
        SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, 
        SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, 
        SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, 
        SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, 
        SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, 
        SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, 
        SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, 
        SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, 
        SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, 
        SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, 
        SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, 
        SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, 
        SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, 
        SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, 
        SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, 
        SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, 
        SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, 
        SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, 
        SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, 
        SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, 
        SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, 
        SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, 
        SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, 
        SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, 
        SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, 
        SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, 
        SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, 
        SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, 
        SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, 
        SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, 
        SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, 
        SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, 
        SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, 
        SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, 
        SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, 
        SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, 
        SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, 
        SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, 
        SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, 
        SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, 
        SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, 
        SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, 
        SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, 
        SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, 
        SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, 
        SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, 
        SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, 
        SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, 
        SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, 
        SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, 
        SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, 
        SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, 
        SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, 
        SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, 
        SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, 
        SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, 
        SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, 
        SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, 
        SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, 
        SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, 
        SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, 
        SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, 
        SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, 
        SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, 
        SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, 
        SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, 
        SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, 
        SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, 
        SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, 
        SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, 
        SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, 
        SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, 
        SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, 
        SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, 
        SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, 
        SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, 
        SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, 
        SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, 
        SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, 
        SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, 
        SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, 
        SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, 
        SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, 
        SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, 
        SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, 
        SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, 
        SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, 
        SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, 
        SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, 
        SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, 
        SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, 
        SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, 
        SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, 
        SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, 
        SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, 
        SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, 
        SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, 
        SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, 
        SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, 
        SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, 
        SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, 
        SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, 
        SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, 
        SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, 
        SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, 
        SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, 
        SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, 
        SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, 
        SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, 
        SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, 
        SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, 
        SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, 
        SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, 
        SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, 
        SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, 
        SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, 
        SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, 
        SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, 
        SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, 
        SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, 
        SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, 
        SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, 
        SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, 
        SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, 
        SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, 
        SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, 
        SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, 
        SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, 
        SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, 
        SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, 
        SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, 
        SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, 
        SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, 
        SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, 
        SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, 
        SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, 
        SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, 
        SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, 
        SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, 
        SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, 
        SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, 
        SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, 
        SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, 
        SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, 
        SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, 
        SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, 
        SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, 
        SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, 
        SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, 
        SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, 
        SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, 
        SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, 
        SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, 
        SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, 
        SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, 
        SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, 
        SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, 
        SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, 
        SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, 
        SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, 
        SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, 
        SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, 
        SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, 
        SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, 
        SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, 
        SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, 
        SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, 
        SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, 
        SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, 
        SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, 
        SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, 
        SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, 
        SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, 
        SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, 
        SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, 
        SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, 
        SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, 
        SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, 
        SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, 
        SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, 
        SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, 
        SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, 
        SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, 
        SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, 
        SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, 
        SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, 
        SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, 
        SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, 
        SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, 
        SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, 
        SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, 
        SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, 
        SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, 
        SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, 
        SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, 
        SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, 
        SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, 
        SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, 
        SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, 
        SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, 
        SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, 
        SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, 
        SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, 
        SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, 
        SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, 
        SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, 
        SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, 
        SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, 
        SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, 
        SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, 
        SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, 
        SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, 
        SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, 
        SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, 
        SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, 
        SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, 
        SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, 
        SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, 
        SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, 
        SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, 
        SYNOPSYS_UNCONNECTED_1016, regx_rdat}) );
  SDFFQX1 d_we16_reg ( .D(N8), .SIN(d_regx_addr[6]), .SMC(test_se), .C(clk), 
        .Q(d_we16) );
  SDFFQX1 d_lt_gpi_reg_2_ ( .D(lt_gpi[2]), .SIN(d_lt_gpi[1]), .SMC(test_se), 
        .C(net8975), .Q(d_lt_gpi[2]) );
  SDFFQX1 d_lt_drp_reg ( .D(lt_drp), .SIN(d_lt_aswk[5]), .SMC(test_se), .C(clk), .Q(reg14[0]) );
  SDFFQX1 d_lt_aswk_reg_0_ ( .D(lt_aswk[0]), .SIN(reg14[3]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[0]) );
  SDFFQX1 d_regx_addr_reg_4_ ( .D(regx_addr[4]), .SIN(d_regx_addr[3]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[4]) );
  SDFFQX1 d_di_tst_reg ( .D(di_tst), .SIN(test_si1), .SMC(test_se), .C(clk), 
        .Q(reg14[3]) );
  SDFFQX1 d_lt_gpi_reg_1_ ( .D(lt_gpi[1]), .SIN(d_lt_gpi[0]), .SMC(test_se), 
        .C(net8975), .Q(d_lt_gpi[1]) );
  SDFFQX1 d_lt_gpi_reg_0_ ( .D(lt_gpi[0]), .SIN(reg14[0]), .SMC(test_se), .C(
        net8975), .Q(d_lt_gpi[0]) );
  SDFFQX1 d_lt_aswk_reg_5_ ( .D(lt_aswk[5]), .SIN(d_lt_aswk[4]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[5]) );
  SDFFQX1 d_lt_aswk_reg_4_ ( .D(lt_aswk[4]), .SIN(d_lt_aswk[3]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[4]) );
  SDFFQX1 d_lt_aswk_reg_3_ ( .D(lt_aswk[3]), .SIN(d_lt_aswk[2]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[3]) );
  SDFFQX1 d_lt_aswk_reg_2_ ( .D(lt_aswk[2]), .SIN(d_lt_aswk[1]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[2]) );
  SDFFQX1 d_lt_aswk_reg_1_ ( .D(lt_aswk[1]), .SIN(d_lt_aswk[0]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[1]) );
  SDFFQX1 d_regx_addr_reg_2_ ( .D(regx_addr[2]), .SIN(d_regx_addr[1]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[2]) );
  SDFFQX1 d_regx_addr_reg_3_ ( .D(regx_addr[3]), .SIN(d_regx_addr[2]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[3]) );
  SDFFQX1 d_lt_gpi_reg_3_ ( .D(lt_gpi[3]), .SIN(d_lt_gpi[2]), .SMC(test_se), 
        .C(net8975), .Q(d_lt_gpi[3]) );
  SDFFQX1 d_regx_addr_reg_1_ ( .D(regx_addr[1]), .SIN(d_regx_addr[0]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[1]) );
  SDFFQX1 d_regx_addr_reg_0_ ( .D(regx_addr[0]), .SIN(d_lt_gpi[3]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[0]) );
  SDFFQX1 d_regx_addr_reg_6_ ( .D(regx_addr[6]), .SIN(d_regx_addr[5]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[6]) );
  SDFFQX1 d_regx_addr_reg_5_ ( .D(regx_addr[5]), .SIN(d_regx_addr[4]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[5]) );
  SDFFRQX1 lt_drp_reg ( .D(di_drposc), .SIN(lt_aswk[5]), .SMC(test_se), .C(
        detclk), .XR(n52), .Q(lt_drp) );
  SDFFRQX1 lt_aswk_reg_5_ ( .D(1'b1), .SIN(lt_aswk[4]), .SMC(test_se), .C(
        aswclk), .XR(n74), .Q(lt_aswk[5]) );
  SDFFRQX1 lt_aswk_reg_4_ ( .D(di_aswk[4]), .SIN(lt_aswk[3]), .SMC(test_se), 
        .C(aswclk), .XR(n74), .Q(lt_aswk[4]) );
  SDFFRQX1 lt_aswk_reg_3_ ( .D(di_aswk[3]), .SIN(lt_aswk[2]), .SMC(test_se), 
        .C(aswclk), .XR(n74), .Q(lt_aswk[3]) );
  SDFFRQX1 lt_aswk_reg_2_ ( .D(di_aswk[2]), .SIN(lt_aswk[1]), .SMC(test_se), 
        .C(aswclk), .XR(n74), .Q(lt_aswk[2]) );
  SDFFRQX1 lt_aswk_reg_1_ ( .D(di_aswk[1]), .SIN(lt_aswk[0]), .SMC(test_se), 
        .C(aswclk), .XR(n74), .Q(lt_aswk[1]) );
  SDFFRQX1 lt_aswk_reg_0_ ( .D(di_aswk[0]), .SIN(d_we16), .SMC(test_se), .C(
        aswclk), .XR(n74), .Q(lt_aswk[0]) );
  INVX1 U4 ( .A(regx_addr[4]), .Y(n100) );
  INVX2 U7 ( .A(regx_addr[2]), .Y(n77) );
  AND2XL U8 ( .A(n120), .B(n127), .Y(regx_wrdac[2]) );
  NOR31X1 U9 ( .C(n34), .A(n100), .B(n122), .Y(n33) );
  INVX1 U10 ( .A(n130), .Y(n110) );
  INVX1 U11 ( .A(n70), .Y(n106) );
  INVX1 U12 ( .A(n73), .Y(n123) );
  INVX2 U13 ( .A(n101), .Y(n129) );
  INVX1 U14 ( .A(n79), .Y(n127) );
  INVX1 U15 ( .A(regx_addr[3]), .Y(n102) );
  AND3X1 U16 ( .A(regx_addr[3]), .B(n127), .C(n33), .Y(regx_wrdac[10]) );
  NAND21X1 U17 ( .B(regx_addr[0]), .A(n67), .Y(n130) );
  INVX1 U18 ( .A(n81), .Y(n67) );
  OR2X1 U19 ( .A(n122), .B(regx_addr[6]), .Y(n1) );
  INVX1 U20 ( .A(regx_addr[1]), .Y(n72) );
  INVXL U21 ( .A(regx_wdat[3]), .Y(n5) );
  INVXL U22 ( .A(n5), .Y(n6) );
  INVXL U23 ( .A(n5), .Y(n7) );
  INVXL U24 ( .A(regx_wdat[6]), .Y(n8) );
  INVXL U25 ( .A(n8), .Y(n9) );
  INVXL U26 ( .A(n8), .Y(n10) );
  INVXL U27 ( .A(regx_wdat[7]), .Y(n11) );
  INVXL U28 ( .A(n11), .Y(n12) );
  INVXL U29 ( .A(n11), .Y(n13) );
  INVXL U30 ( .A(regx_wdat[0]), .Y(n14) );
  INVXL U31 ( .A(n14), .Y(wd_twlb[0]) );
  INVXL U32 ( .A(n14), .Y(n16) );
  INVXL U33 ( .A(regx_wdat[2]), .Y(n17) );
  INVXL U34 ( .A(n17), .Y(n18) );
  INVXL U35 ( .A(n17), .Y(n19) );
  INVXL U36 ( .A(regx_wdat[4]), .Y(n20) );
  INVXL U37 ( .A(n20), .Y(n21) );
  INVXL U38 ( .A(n20), .Y(n22) );
  INVXL U39 ( .A(regx_wdat[5]), .Y(n23) );
  INVXL U40 ( .A(n23), .Y(n24) );
  INVXL U41 ( .A(n23), .Y(n25) );
  INVXL U42 ( .A(d_regx_addr[2]), .Y(n26) );
  INVXL U43 ( .A(n26), .Y(n27) );
  INVX1 U44 ( .A(d_regx_addr[3]), .Y(n28) );
  INVX1 U45 ( .A(n28), .Y(n29) );
  BUFX3 U46 ( .A(r_imp_osc), .Y(r_xana[22]) );
  AND3XL U47 ( .A(regx_addr[3]), .B(n129), .C(n33), .Y(regx_wrdac[11]) );
  AND3XL U48 ( .A(n33), .B(n129), .C(n102), .Y(regx_wrdac[1]) );
  NAND21XL U49 ( .B(regx_addr[3]), .A(n100), .Y(n98) );
  AND2XL U50 ( .A(n120), .B(n31), .Y(regx_wrdac[9]) );
  NOR2X2 U51 ( .A(n98), .B(n1), .Y(n35) );
  NAND21X1 U52 ( .B(n104), .A(regx_addr[5]), .Y(n122) );
  AND2X2 U53 ( .A(n35), .B(n129), .Y(regx_wrdac[13]) );
  AND3XL U54 ( .A(n33), .B(n127), .C(n102), .Y(regx_wrdac[0]) );
  INVXL U55 ( .A(regx_addr[6]), .Y(n34) );
  INVX1 U56 ( .A(n69), .Y(n108) );
  NOR2X1 U57 ( .A(regx_addr[0]), .B(regx_addr[1]), .Y(n30) );
  AND2XL U58 ( .A(n80), .B(n110), .Y(we[30]) );
  AND2X2 U59 ( .A(n35), .B(n127), .Y(regx_wrdac[12]) );
  INVXL U60 ( .A(n68), .Y(n109) );
  AND2XL U61 ( .A(n127), .B(n128), .Y(regx_hitbst[0]) );
  AND2XL U62 ( .A(n36), .B(n127), .Y(regx_wrcvc[0]) );
  AND2XL U63 ( .A(n126), .B(n127), .Y(regx_wrpwm[0]) );
  NAND21XL U64 ( .B(n101), .A(n80), .Y(n78) );
  AND2XL U65 ( .A(n31), .B(n126), .Y(regx_wrcvc[3]) );
  AND2XL U66 ( .A(n36), .B(n31), .Y(we_7) );
  AND2XL U67 ( .A(n80), .B(n127), .Y(we[24]) );
  AND2XL U68 ( .A(n71), .B(n106), .Y(we[27]) );
  AND2XL U69 ( .A(n106), .B(n128), .Y(we_19) );
  INVX1 U70 ( .A(n98), .Y(n121) );
  INVXL U71 ( .A(regx_addr[0]), .Y(n32) );
  NOR2XL U72 ( .A(regx_addr[3]), .B(n124), .Y(n36) );
  NAND21XL U93 ( .B(n124), .A(regx_addr[3]), .Y(n125) );
  NOR42XL U97 ( .C(n135), .D(n16), .A(n130), .B(n134), .Y(N8) );
  INVX1 U98 ( .A(n92), .Y(n76) );
  AND2XL U99 ( .A(n109), .B(n120), .Y(regx_wrdac[7]) );
  AND2XL U100 ( .A(n120), .B(n129), .Y(regx_wrdac[3]) );
  AND2XL U101 ( .A(n120), .B(n110), .Y(regx_wrdac[8]) );
  INVX1 U102 ( .A(n95), .Y(n128) );
  NAND21X1 U103 ( .B(n133), .A(n109), .Y(n92) );
  INVX1 U104 ( .A(n66), .Y(n80) );
  NAND21X1 U105 ( .B(n104), .A(n71), .Y(n66) );
  AND2X1 U106 ( .A(n71), .B(n108), .Y(we[28]) );
  AND2X1 U107 ( .A(n80), .B(n109), .Y(we[29]) );
  AND2X2 U108 ( .A(n120), .B(n123), .Y(regx_wrdac[4]) );
  NAND32XL U109 ( .B(n77), .C(n32), .A(n72), .Y(n68) );
  NAND32XL U110 ( .B(n77), .C(n104), .A(n30), .Y(n69) );
  NAND32X1 U111 ( .B(n97), .C(n100), .A(n102), .Y(n95) );
  NAND21X1 U112 ( .B(n95), .A(regx_w), .Y(n133) );
  INVX1 U113 ( .A(n96), .Y(we_twlb) );
  NAND21X1 U114 ( .B(n133), .A(n123), .Y(n96) );
  NAND32X1 U115 ( .B(n97), .C(n104), .A(n100), .Y(n124) );
  AND2X1 U116 ( .A(n123), .B(n36), .Y(regx_wrcvc[2]) );
  AND2XL U117 ( .A(n126), .B(n129), .Y(regx_wrpwm[1]) );
  AND2XL U118 ( .A(n36), .B(n129), .Y(regx_wrcvc[1]) );
  AND2XL U119 ( .A(n129), .B(n128), .Y(regx_hitbst[1]) );
  AND2XL U120 ( .A(n109), .B(n36), .Y(we_5) );
  NOR21XL U121 ( .B(n31), .A(n133), .Y(we[23]) );
  INVX1 U122 ( .A(n78), .Y(n75) );
  INVX1 U123 ( .A(n65), .Y(n71) );
  NAND32X1 U124 ( .B(n100), .C(n102), .A(n99), .Y(n65) );
  INVX1 U125 ( .A(regx_w), .Y(n104) );
  AND3XL U126 ( .A(n108), .B(n99), .C(n121), .Y(we_4) );
  INVX1 U127 ( .A(n97), .Y(n99) );
  AND2X1 U128 ( .A(n80), .B(n123), .Y(we[26]) );
  INVX1 U129 ( .A(n64), .Y(wd_twlb[1]) );
  INVX1 U130 ( .A(n64), .Y(n63) );
  NAND32X1 U131 ( .B(regx_addr[1]), .C(n32), .A(n77), .Y(n101) );
  NAND32XL U132 ( .B(regx_addr[0]), .C(n72), .A(n77), .Y(n73) );
  NOR2XL U133 ( .A(n81), .B(n32), .Y(n31) );
  NAND21X1 U134 ( .B(regx_addr[2]), .A(n30), .Y(n79) );
  NAND43X1 U135 ( .B(regx_addr[2]), .C(n32), .D(n72), .A(regx_w), .Y(n70) );
  OR2XL U136 ( .A(regx_addr[5]), .B(regx_addr[6]), .Y(n97) );
  INVX1 U137 ( .A(n125), .Y(n126) );
  AO21X1 U138 ( .B(bus_idle), .C(n94), .A(n93), .Y(i2c_mode_upd) );
  AND3X1 U139 ( .A(n76), .B(n13), .C(n8), .Y(n93) );
  NAND43X1 U140 ( .B(n91), .C(n90), .D(n89), .A(n88), .Y(n94) );
  AND2X1 U141 ( .A(n12), .B(n9), .Y(n135) );
  NAND42X1 U142 ( .C(n6), .D(n133), .A(n132), .B(n131), .Y(n134) );
  NOR2X1 U143 ( .A(n18), .B(wd_twlb[1]), .Y(n132) );
  NOR2X1 U144 ( .A(n24), .B(n21), .Y(n131) );
  INVX1 U145 ( .A(regx_wdat[1]), .Y(n64) );
  AND4X1 U146 ( .A(n87), .B(n92), .C(n86), .D(n85), .Y(n88) );
  XOR2X1 U147 ( .A(n82), .B(r_i2crout[2]), .Y(n87) );
  XOR2X1 U148 ( .A(n83), .B(r_i2crout[1]), .Y(n86) );
  XOR2X1 U149 ( .A(n84), .B(r_i2crout[0]), .Y(n85) );
  MUX2X1 U150 ( .D0(lt_reg15_5_0[2]), .D1(n19), .S(n76), .Y(i2c_mode_wdat[2])
         );
  MUX2X1 U151 ( .D0(lt_reg15_5_0[5]), .D1(n25), .S(n76), .Y(i2c_mode_wdat[5])
         );
  MUX2X1 U152 ( .D0(lt_reg15_5_0[4]), .D1(n22), .S(n76), .Y(i2c_mode_wdat[4])
         );
  MUX2X1 U153 ( .D0(lt_reg15_5_0[0]), .D1(n16), .S(n76), .Y(i2c_mode_wdat[0])
         );
  MUX2X1 U154 ( .D0(lt_reg15_5_0[3]), .D1(n7), .S(n76), .Y(i2c_mode_wdat[3])
         );
  MUX2X1 U155 ( .D0(lt_reg15_5_0[1]), .D1(n63), .S(n76), .Y(i2c_mode_wdat[1])
         );
  XNOR2XL U156 ( .A(reg1E[2]), .B(n61), .Y(r_xana[18]) );
  NAND2X1 U157 ( .A(r_xana[20]), .B(di_drposc), .Y(n61) );
  XNOR2XL U158 ( .A(reg1E[3]), .B(n61), .Y(r_xana[19]) );
  XOR2X1 U159 ( .A(r_i2crout[4]), .B(lt_reg15_5_0[4]), .Y(n91) );
  XOR2X1 U160 ( .A(r_i2crout[5]), .B(lt_reg15_5_0[5]), .Y(n90) );
  XOR2X1 U161 ( .A(r_i2crout[3]), .B(lt_reg15_5_0[3]), .Y(n89) );
  INVX1 U162 ( .A(lt_reg15_5_0[0]), .Y(n84) );
  INVX1 U163 ( .A(lt_reg15_5_0[1]), .Y(n83) );
  INVX1 U164 ( .A(lt_reg15_5_0[2]), .Y(n82) );
  OA21X1 U165 ( .B(n136), .C(atpg_en), .A(n53), .Y(n74) );
  INVX1 U166 ( .A(d_we16), .Y(n136) );
  NAND21X1 U167 ( .B(n77), .A(regx_addr[1]), .Y(n81) );
  INVX2 U168 ( .A(n103), .Y(n107) );
  NAND43X1 U169 ( .B(regx_addr[6]), .C(regx_addr[4]), .D(n102), .A(
        regx_addr[5]), .Y(n103) );
  INVX4 U170 ( .A(n105), .Y(n120) );
  NAND21X4 U171 ( .B(n104), .A(n107), .Y(n105) );
  AND2X4 U172 ( .A(n106), .B(n107), .Y(regx_wrdac[5]) );
  AND2X4 U173 ( .A(n108), .B(n107), .Y(regx_wrdac[6]) );
endmodule


module regx_a0_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718;

  BUFXL U2125 ( .A(SH[5]), .Y(n3633) );
  BUFX3 U2126 ( .A(SH[6]), .Y(n3634) );
  INVX1 U2127 ( .A(n3676), .Y(n3665) );
  INVX1 U2128 ( .A(n3677), .Y(n3664) );
  INVX1 U2129 ( .A(n3712), .Y(n3694) );
  INVX1 U2130 ( .A(n3712), .Y(n3693) );
  INVX1 U2131 ( .A(n3712), .Y(n3692) );
  INVX1 U2132 ( .A(n3675), .Y(n3668) );
  INVX1 U2133 ( .A(n3674), .Y(n3672) );
  INVX1 U2134 ( .A(n3711), .Y(n3706) );
  INVX1 U2135 ( .A(n3713), .Y(n3697) );
  INVX1 U2136 ( .A(n3714), .Y(n3703) );
  INVX1 U2137 ( .A(n3713), .Y(n3707) );
  INVX1 U2138 ( .A(n3711), .Y(n3708) );
  INVX1 U2139 ( .A(n3714), .Y(n3710) );
  INVX1 U2140 ( .A(n3674), .Y(n3673) );
  INVX1 U2141 ( .A(n3713), .Y(n3695) );
  INVX1 U2142 ( .A(n3713), .Y(n3696) );
  INVX1 U2143 ( .A(n3676), .Y(n3667) );
  INVX1 U2144 ( .A(n3714), .Y(n3709) );
  INVX1 U2145 ( .A(n3678), .Y(n3661) );
  INVX1 U2146 ( .A(n3678), .Y(n3660) );
  INVX1 U2147 ( .A(n3677), .Y(n3662) );
  INVX1 U2148 ( .A(n3677), .Y(n3663) );
  INVX1 U2149 ( .A(n3678), .Y(n3659) );
  INVX1 U2150 ( .A(n3676), .Y(n3666) );
  INVX1 U2151 ( .A(n3679), .Y(n3671) );
  INVX1 U2152 ( .A(n3679), .Y(n3670) );
  INVX1 U2153 ( .A(n3679), .Y(n3669) );
  INVX1 U2154 ( .A(n3712), .Y(n3700) );
  INVX1 U2155 ( .A(n3714), .Y(n3704) );
  INVX1 U2156 ( .A(n3714), .Y(n3705) );
  INVX1 U2157 ( .A(n3714), .Y(n3702) );
  INVX1 U2158 ( .A(n3711), .Y(n3701) );
  INVX1 U2159 ( .A(n3718), .Y(n3699) );
  INVX1 U2160 ( .A(n3718), .Y(n3698) );
  INVX1 U2161 ( .A(n3715), .Y(n3714) );
  INVX1 U2162 ( .A(n3716), .Y(n3712) );
  INVX1 U2163 ( .A(n3716), .Y(n3713) );
  INVX1 U2164 ( .A(n3687), .Y(n3676) );
  INVX1 U2165 ( .A(n3687), .Y(n3677) );
  INVX1 U2166 ( .A(n3688), .Y(n3675) );
  INVX1 U2167 ( .A(n3688), .Y(n3674) );
  INVX1 U2168 ( .A(n3642), .Y(n3635) );
  INVX1 U2169 ( .A(n3644), .Y(n3636) );
  INVX1 U2170 ( .A(n3643), .Y(n3637) );
  INVX1 U2171 ( .A(n3648), .Y(n3639) );
  INVX1 U2172 ( .A(n3649), .Y(n3640) );
  INVX1 U2173 ( .A(n3717), .Y(n3711) );
  INVX1 U2174 ( .A(n3686), .Y(n3680) );
  INVX1 U2175 ( .A(n3686), .Y(n3681) );
  INVX1 U2176 ( .A(n3646), .Y(n3641) );
  INVX1 U2177 ( .A(n3686), .Y(n3679) );
  INVX1 U2178 ( .A(n3687), .Y(n3678) );
  INVX1 U2179 ( .A(n3647), .Y(n3638) );
  MUX4X1 U2180 ( .D0(n3275), .D1(n3276), .D2(n3277), .D3(n3278), .S0(n3635), 
        .S1(n3656), .Y(n3264) );
  NOR3XL U2181 ( .A(n3682), .B(n3708), .C(A[343]), .Y(n3277) );
  NOR3XL U2182 ( .A(n3680), .B(n3707), .C(A[351]), .Y(n3278) );
  NOR21XL U2183 ( .B(n3280), .A(n3694), .Y(n3275) );
  MUX4X1 U2184 ( .D0(n3267), .D1(n3268), .D2(n3269), .D3(n3270), .S0(n3652), 
        .S1(n3637), .Y(n3266) );
  NOR3XL U2185 ( .A(n3683), .B(n3708), .C(A[367]), .Y(n3269) );
  NOR3XL U2186 ( .A(n3682), .B(n3708), .C(A[359]), .Y(n3267) );
  NOR3XL U2187 ( .A(n3681), .B(n3707), .C(A[375]), .Y(n3268) );
  MUX4X1 U2188 ( .D0(n3517), .D1(n3518), .D2(n3519), .D3(n3520), .S0(n3635), 
        .S1(n3655), .Y(n3506) );
  NOR3XL U2189 ( .A(n3678), .B(n3699), .C(A[338]), .Y(n3519) );
  NOR3XL U2190 ( .A(n3678), .B(n3699), .C(A[346]), .Y(n3520) );
  NOR21XL U2191 ( .B(n3522), .A(n3716), .Y(n3517) );
  MUX4X1 U2192 ( .D0(n3569), .D1(n3570), .D2(n3571), .D3(n3572), .S0(n3636), 
        .S1(n3656), .Y(n3558) );
  NOR3XL U2193 ( .A(n3682), .B(n3700), .C(A[337]), .Y(n3571) );
  NOR3XL U2194 ( .A(n3690), .B(n3700), .C(A[345]), .Y(n3572) );
  NOR21XL U2195 ( .B(n3574), .A(n3716), .Y(n3569) );
  MUX4X1 U2196 ( .D0(n3419), .D1(n3420), .D2(n3421), .D3(n3422), .S0(n3636), 
        .S1(n3655), .Y(n3408) );
  NOR3XL U2197 ( .A(n3690), .B(n3704), .C(A[340]), .Y(n3421) );
  NOR3XL U2198 ( .A(n3684), .B(n3704), .C(A[348]), .Y(n3422) );
  NOR21XL U2199 ( .B(n3424), .A(SH[9]), .Y(n3419) );
  MUX4X1 U2200 ( .D0(n3370), .D1(n3371), .D2(n3372), .D3(n3373), .S0(n3636), 
        .S1(n3656), .Y(n3359) );
  NOR3XL U2201 ( .A(n3679), .B(n3705), .C(A[341]), .Y(n3372) );
  NOR3XL U2202 ( .A(n3691), .B(n3715), .C(A[349]), .Y(n3373) );
  NOR21XL U2203 ( .B(n3375), .A(SH[9]), .Y(n3370) );
  MUX4X1 U2204 ( .D0(n3468), .D1(n3469), .D2(n3470), .D3(n3471), .S0(n3636), 
        .S1(n3655), .Y(n3457) );
  NOR3XL U2205 ( .A(n3679), .B(n3697), .C(A[339]), .Y(n3470) );
  NOR3XL U2206 ( .A(n3690), .B(n3697), .C(A[347]), .Y(n3471) );
  NOR21XL U2207 ( .B(n3473), .A(n3694), .Y(n3468) );
  MUX4X1 U2208 ( .D0(n3561), .D1(n3562), .D2(n3563), .D3(n3564), .S0(n3653), 
        .S1(n3638), .Y(n3560) );
  NOR3XL U2209 ( .A(n3690), .B(n3700), .C(A[361]), .Y(n3563) );
  NOR3XL U2210 ( .A(n3684), .B(n3700), .C(A[353]), .Y(n3561) );
  NOR3XL U2211 ( .A(n3690), .B(n3700), .C(A[369]), .Y(n3562) );
  MUX4X1 U2212 ( .D0(n3411), .D1(n3412), .D2(n3413), .D3(n3414), .S0(n3654), 
        .S1(n3637), .Y(n3410) );
  NOR3XL U2213 ( .A(n3690), .B(n3704), .C(A[364]), .Y(n3413) );
  NOR3XL U2214 ( .A(n3681), .B(n3704), .C(A[356]), .Y(n3411) );
  NOR3XL U2215 ( .A(n3680), .B(n3704), .C(A[372]), .Y(n3412) );
  MUX4X1 U2216 ( .D0(n3362), .D1(n3363), .D2(n3364), .D3(n3365), .S0(n3653), 
        .S1(n3641), .Y(n3361) );
  NOR3XL U2217 ( .A(n3680), .B(n3716), .C(A[365]), .Y(n3364) );
  NOR3XL U2218 ( .A(n3679), .B(n3716), .C(A[357]), .Y(n3362) );
  NOR3XL U2219 ( .A(n3679), .B(n3716), .C(A[373]), .Y(n3363) );
  MUX4X1 U2220 ( .D0(n3460), .D1(n3461), .D2(n3462), .D3(n3463), .S0(n3657), 
        .S1(n3638), .Y(n3459) );
  NOR3XL U2221 ( .A(n3681), .B(n3702), .C(A[363]), .Y(n3462) );
  NOR3XL U2222 ( .A(n3679), .B(n3698), .C(A[355]), .Y(n3460) );
  NOR3XL U2223 ( .A(n3691), .B(n3702), .C(A[371]), .Y(n3461) );
  MUX4X1 U2224 ( .D0(n3509), .D1(n3510), .D2(n3511), .D3(n3512), .S0(n3654), 
        .S1(n3638), .Y(n3508) );
  NOR3XL U2225 ( .A(n3678), .B(n3698), .C(A[362]), .Y(n3511) );
  NOR3XL U2226 ( .A(n3678), .B(n3698), .C(A[354]), .Y(n3509) );
  NOR3XL U2227 ( .A(n3678), .B(n3698), .C(A[370]), .Y(n3510) );
  MUX4X1 U2228 ( .D0(n3621), .D1(n3622), .D2(n3623), .D3(n3624), .S0(n3636), 
        .S1(n3656), .Y(n3610) );
  NOR3XL U2229 ( .A(n3690), .B(n3702), .C(A[336]), .Y(n3623) );
  NOR3XL U2230 ( .A(n3679), .B(n3702), .C(A[344]), .Y(n3624) );
  NOR21XL U2231 ( .B(n3626), .A(n3692), .Y(n3621) );
  MUX4X1 U2232 ( .D0(n3322), .D1(n3323), .D2(n3324), .D3(n3325), .S0(n3636), 
        .S1(n3655), .Y(n3311) );
  NOR3XL U2233 ( .A(n3691), .B(n3706), .C(A[342]), .Y(n3324) );
  NOR3XL U2234 ( .A(n3681), .B(n3706), .C(A[350]), .Y(n3325) );
  NOR21XL U2235 ( .B(n3327), .A(n3694), .Y(n3322) );
  MUX4X1 U2236 ( .D0(n3613), .D1(n3614), .D2(n3615), .D3(n3616), .S0(n3652), 
        .S1(n3639), .Y(n3612) );
  NOR3XL U2237 ( .A(n3682), .B(n3701), .C(A[360]), .Y(n3615) );
  NOR3XL U2238 ( .A(n3690), .B(n3702), .C(A[352]), .Y(n3613) );
  NOR3XL U2239 ( .A(n3682), .B(n3702), .C(A[368]), .Y(n3614) );
  MUX4X1 U2240 ( .D0(n3314), .D1(n3315), .D2(n3316), .D3(n3317), .S0(n3653), 
        .S1(n3638), .Y(n3313) );
  NOR3XL U2241 ( .A(n3682), .B(n3707), .C(A[366]), .Y(n3316) );
  NOR3XL U2242 ( .A(n3681), .B(n3707), .C(A[358]), .Y(n3314) );
  NOR3XL U2243 ( .A(n3680), .B(n3706), .C(A[374]), .Y(n3315) );
  NOR3XL U2244 ( .A(A[175]), .B(n3706), .C(n3673), .Y(n3254) );
  INVX1 U2245 ( .A(n3685), .Y(n3683) );
  INVX1 U2246 ( .A(n3689), .Y(n3687) );
  INVX1 U2247 ( .A(n3711), .Y(n3715) );
  INVX1 U2248 ( .A(n3689), .Y(n3688) );
  INVX1 U2249 ( .A(n3711), .Y(n3716) );
  INVX1 U2250 ( .A(n3685), .Y(n3684) );
  INVX1 U2251 ( .A(n3658), .Y(n3656) );
  BUFX3 U2252 ( .A(n3651), .Y(n3642) );
  BUFX3 U2253 ( .A(n3651), .Y(n3646) );
  BUFX3 U2254 ( .A(n3651), .Y(n3644) );
  BUFX3 U2255 ( .A(n3651), .Y(n3648) );
  BUFX3 U2256 ( .A(n3649), .Y(n3643) );
  BUFX3 U2257 ( .A(n3651), .Y(n3649) );
  INVX1 U2258 ( .A(n3685), .Y(n3682) );
  INVX1 U2259 ( .A(n3718), .Y(n3717) );
  INVX1 U2260 ( .A(n3690), .Y(n3686) );
  INVX1 U2261 ( .A(n3658), .Y(n3655) );
  INVX1 U2262 ( .A(n3658), .Y(n3657) );
  INVX1 U2263 ( .A(n3658), .Y(n3653) );
  INVX1 U2264 ( .A(n3658), .Y(n3654) );
  BUFX3 U2265 ( .A(n3650), .Y(n3645) );
  BUFX3 U2266 ( .A(n3650), .Y(n3647) );
  BUFX3 U2267 ( .A(n3651), .Y(n3650) );
  MUX2IX1 U2268 ( .D0(n3239), .D1(n3240), .S(SH[7]), .Y(B[7]) );
  MUX4X1 U2269 ( .D0(n3241), .D1(n3242), .D2(n3243), .D3(n3244), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3240) );
  MUX4X1 U2270 ( .D0(n3263), .D1(n3264), .D2(n3265), .D3(n3266), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3239) );
  MUX3X1 U2271 ( .D0(n3253), .D1(n3254), .D2(n3255), .S0(n3640), .S1(n3657), 
        .Y(n3242) );
  MUX2IX1 U2272 ( .D0(A[71]), .D1(A[327]), .S(n3665), .Y(n3280) );
  NOR21XL U2273 ( .B(n3271), .A(n3692), .Y(n3270) );
  MUX2IX1 U2274 ( .D0(A[127]), .D1(A[383]), .S(n3665), .Y(n3271) );
  NOR21XL U2275 ( .B(n3279), .A(n3693), .Y(n3276) );
  MUX2IX1 U2276 ( .D0(A[79]), .D1(A[335]), .S(n3665), .Y(n3279) );
  MUX2IX1 U2277 ( .D0(A[15]), .D1(A[271]), .S(n3664), .Y(n3285) );
  MUX2X1 U2278 ( .D0(n3281), .D1(n3282), .S(n3655), .Y(n3263) );
  NOR4XL U2279 ( .A(n3695), .B(n3667), .C(n3636), .D(A[23]), .Y(n3282) );
  MUX2IX1 U2280 ( .D0(n3283), .D1(n3284), .S(n3635), .Y(n3281) );
  NAND2X1 U2281 ( .A(n3285), .B(n3711), .Y(n3284) );
  NAND2X1 U2282 ( .A(n3286), .B(n3711), .Y(n3283) );
  MUX2IX1 U2283 ( .D0(A[7]), .D1(A[263]), .S(n3665), .Y(n3286) );
  MUX2IX1 U2284 ( .D0(A[9]), .D1(A[265]), .S(n3663), .Y(n3579) );
  MUX2IX1 U2285 ( .D0(A[10]), .D1(A[266]), .S(n3660), .Y(n3527) );
  MUX2IX1 U2286 ( .D0(n3529), .D1(n3530), .S(SH[7]), .Y(B[1]) );
  MUX4X1 U2287 ( .D0(n3531), .D1(n3532), .D2(n3533), .D3(n3534), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3530) );
  MUX4X1 U2288 ( .D0(n3557), .D1(n3558), .D2(n3559), .D3(n3560), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3529) );
  MUX4X1 U2289 ( .D0(n3535), .D1(n3536), .D2(n3537), .D3(n3538), .S0(n3654), 
        .S1(n3639), .Y(n3534) );
  MUX2IX1 U2290 ( .D0(n3382), .D1(n3383), .S(SH[7]), .Y(B[4]) );
  MUX4X1 U2291 ( .D0(n3384), .D1(n3385), .D2(n3386), .D3(n3387), .S0(SH[5]), 
        .S1(n3634), .Y(n3383) );
  MUX4X1 U2292 ( .D0(n3407), .D1(n3408), .D2(n3409), .D3(n3410), .S0(SH[6]), 
        .S1(n3633), .Y(n3382) );
  MUX4X1 U2293 ( .D0(n3392), .D1(n3393), .D2(n3394), .D3(n3395), .S0(n3654), 
        .S1(n3637), .Y(n3386) );
  MUX2IX1 U2294 ( .D0(n3334), .D1(n3335), .S(SH[7]), .Y(B[5]) );
  MUX4X1 U2295 ( .D0(n3336), .D1(n3337), .D2(n3338), .D3(n3339), .S0(n3633), 
        .S1(n3634), .Y(n3335) );
  MUX4X1 U2296 ( .D0(n3358), .D1(n3359), .D2(n3360), .D3(n3361), .S0(n3634), 
        .S1(n3633), .Y(n3334) );
  MUX3X1 U2297 ( .D0(n3340), .D1(n3341), .D2(n3342), .S0(n3640), .S1(n3657), 
        .Y(n3339) );
  MUX2IX1 U2298 ( .D0(n3431), .D1(n3432), .S(SH[7]), .Y(B[3]) );
  MUX4X1 U2299 ( .D0(n3433), .D1(n3434), .D2(n3435), .D3(n3436), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3432) );
  MUX4X1 U2300 ( .D0(n3456), .D1(n3457), .D2(n3458), .D3(n3459), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3431) );
  MUX4X1 U2301 ( .D0(n3441), .D1(n3442), .D2(n3443), .D3(n3444), .S0(n3657), 
        .S1(n3637), .Y(n3435) );
  MUX2IX1 U2302 ( .D0(n3480), .D1(n3481), .S(SH[7]), .Y(B[2]) );
  MUX4X1 U2303 ( .D0(n3482), .D1(n3483), .D2(n3484), .D3(n3485), .S0(SH[5]), 
        .S1(n3634), .Y(n3481) );
  MUX4X1 U2304 ( .D0(n3505), .D1(n3506), .D2(n3507), .D3(n3508), .S0(SH[6]), 
        .S1(n3633), .Y(n3480) );
  MUX4X1 U2305 ( .D0(n3490), .D1(n3491), .D2(n3492), .D3(n3493), .S0(SH[4]), 
        .S1(n3638), .Y(n3484) );
  MUX2IX1 U2306 ( .D0(A[65]), .D1(A[321]), .S(n3663), .Y(n3574) );
  NOR21XL U2307 ( .B(n3565), .A(n3715), .Y(n3564) );
  MUX2IX1 U2308 ( .D0(A[121]), .D1(A[377]), .S(n3662), .Y(n3565) );
  MUX2IX1 U2309 ( .D0(A[68]), .D1(A[324]), .S(n3661), .Y(n3424) );
  MUX2IX1 U2310 ( .D0(A[69]), .D1(A[325]), .S(n3662), .Y(n3375) );
  NOR21XL U2311 ( .B(n3415), .A(n3694), .Y(n3414) );
  MUX2IX1 U2312 ( .D0(A[124]), .D1(A[380]), .S(n3661), .Y(n3415) );
  MUX2IX1 U2313 ( .D0(A[67]), .D1(A[323]), .S(n3659), .Y(n3473) );
  NOR21XL U2314 ( .B(n3366), .A(n3716), .Y(n3365) );
  MUX2IX1 U2315 ( .D0(A[125]), .D1(A[381]), .S(n3662), .Y(n3366) );
  MUX2IX1 U2316 ( .D0(A[66]), .D1(A[322]), .S(n3660), .Y(n3522) );
  NOR21XL U2317 ( .B(n3464), .A(n3692), .Y(n3463) );
  MUX2IX1 U2318 ( .D0(A[123]), .D1(A[379]), .S(n3660), .Y(n3464) );
  NOR21XL U2319 ( .B(n3513), .A(n3695), .Y(n3512) );
  MUX2IX1 U2320 ( .D0(A[122]), .D1(A[378]), .S(n3659), .Y(n3513) );
  NOR21XL U2321 ( .B(n3573), .A(n3694), .Y(n3570) );
  MUX2IX1 U2322 ( .D0(A[73]), .D1(A[329]), .S(n3662), .Y(n3573) );
  NOR21XL U2323 ( .B(n3423), .A(SH[9]), .Y(n3420) );
  MUX2IX1 U2324 ( .D0(A[76]), .D1(A[332]), .S(n3661), .Y(n3423) );
  NOR21XL U2325 ( .B(n3374), .A(n3695), .Y(n3371) );
  MUX2IX1 U2326 ( .D0(A[77]), .D1(A[333]), .S(n3662), .Y(n3374) );
  NOR21XL U2327 ( .B(n3472), .A(n3693), .Y(n3469) );
  MUX2IX1 U2328 ( .D0(A[75]), .D1(A[331]), .S(n3659), .Y(n3472) );
  NOR21XL U2329 ( .B(n3521), .A(n3695), .Y(n3518) );
  MUX2IX1 U2330 ( .D0(A[74]), .D1(A[330]), .S(n3659), .Y(n3521) );
  MUX2X1 U2331 ( .D0(n3575), .D1(n3576), .S(SH[4]), .Y(n3557) );
  NOR4XL U2332 ( .A(n3696), .B(n3666), .C(n3636), .D(A[17]), .Y(n3576) );
  MUX2IX1 U2333 ( .D0(n3577), .D1(n3578), .S(n3635), .Y(n3575) );
  NAND2X1 U2334 ( .A(n3579), .B(n3712), .Y(n3578) );
  MUX2X1 U2335 ( .D0(n3523), .D1(n3524), .S(SH[4]), .Y(n3505) );
  NOR4XL U2336 ( .A(n3696), .B(n3666), .C(n3641), .D(A[18]), .Y(n3524) );
  MUX2IX1 U2337 ( .D0(n3525), .D1(n3526), .S(n3635), .Y(n3523) );
  NAND2X1 U2338 ( .A(n3527), .B(n3718), .Y(n3526) );
  NAND2X1 U2339 ( .A(n3580), .B(n3713), .Y(n3577) );
  MUX2IX1 U2340 ( .D0(A[1]), .D1(A[257]), .S(n3663), .Y(n3580) );
  NAND2X1 U2341 ( .A(n3528), .B(n3718), .Y(n3525) );
  MUX2IX1 U2342 ( .D0(A[2]), .D1(A[258]), .S(n3660), .Y(n3528) );
  MUX2IX1 U2343 ( .D0(n3287), .D1(n3288), .S(SH[7]), .Y(B[6]) );
  MUX4X1 U2344 ( .D0(n3289), .D1(n3290), .D2(n3291), .D3(n3292), .S0(n3633), 
        .S1(n3634), .Y(n3288) );
  MUX4X1 U2345 ( .D0(n3310), .D1(n3311), .D2(n3312), .D3(n3313), .S0(n3634), 
        .S1(n3633), .Y(n3287) );
  MUX2X1 U2346 ( .D0(n3301), .D1(n3302), .S(n3655), .Y(n3290) );
  MUX2IX1 U2347 ( .D0(A[12]), .D1(A[268]), .S(n3660), .Y(n3429) );
  MUX2IX1 U2348 ( .D0(A[5]), .D1(A[261]), .S(n3662), .Y(n3381) );
  MUX2IX1 U2349 ( .D0(A[11]), .D1(A[267]), .S(n3659), .Y(n3478) );
  NAND2X1 U2350 ( .A(n3380), .B(n3713), .Y(n3379) );
  MUX2IX1 U2351 ( .D0(A[13]), .D1(A[269]), .S(n3662), .Y(n3380) );
  MUX2IX1 U2352 ( .D0(A[6]), .D1(A[262]), .S(n3663), .Y(n3333) );
  NAND2X1 U2353 ( .A(n3332), .B(n3711), .Y(n3331) );
  MUX2IX1 U2354 ( .D0(A[14]), .D1(A[270]), .S(n3663), .Y(n3332) );
  MUX2IX1 U2355 ( .D0(n3581), .D1(n3582), .S(SH[7]), .Y(B[0]) );
  MUX4X1 U2356 ( .D0(n3583), .D1(n3584), .D2(n3585), .D3(n3586), .S0(SH[5]), 
        .S1(n3634), .Y(n3582) );
  MUX4X1 U2357 ( .D0(n3609), .D1(n3610), .D2(n3611), .D3(n3612), .S0(SH[6]), 
        .S1(n3633), .Y(n3581) );
  MUX4X1 U2358 ( .D0(n3587), .D1(n3588), .D2(n3589), .D3(n3590), .S0(n3653), 
        .S1(n3639), .Y(n3586) );
  MUX2IX1 U2359 ( .D0(A[64]), .D1(A[320]), .S(n3665), .Y(n3626) );
  MUX2IX1 U2360 ( .D0(A[70]), .D1(A[326]), .S(n3663), .Y(n3327) );
  NOR21XL U2361 ( .B(n3625), .A(n3692), .Y(n3622) );
  MUX2IX1 U2362 ( .D0(A[72]), .D1(A[328]), .S(n3665), .Y(n3625) );
  NOR21XL U2363 ( .B(n3326), .A(SH[9]), .Y(n3323) );
  MUX2IX1 U2364 ( .D0(A[78]), .D1(A[334]), .S(n3663), .Y(n3326) );
  NOR21XL U2365 ( .B(n3617), .A(n3692), .Y(n3616) );
  MUX2IX1 U2366 ( .D0(A[120]), .D1(A[376]), .S(n3664), .Y(n3617) );
  NOR21XL U2367 ( .B(n3318), .A(SH[9]), .Y(n3317) );
  MUX2IX1 U2368 ( .D0(A[126]), .D1(A[382]), .S(n3664), .Y(n3318) );
  MUX2X1 U2369 ( .D0(n3425), .D1(n3426), .S(n3655), .Y(n3407) );
  NOR4XL U2370 ( .A(n3695), .B(n3666), .C(n3641), .D(A[20]), .Y(n3426) );
  MUX2IX1 U2371 ( .D0(n3427), .D1(n3428), .S(n3635), .Y(n3425) );
  NAND2X1 U2372 ( .A(n3429), .B(n3718), .Y(n3428) );
  MUX2X1 U2373 ( .D0(n3376), .D1(n3377), .S(n3655), .Y(n3358) );
  NOR4XL U2374 ( .A(n3696), .B(n3666), .C(n3636), .D(A[21]), .Y(n3377) );
  MUX2IX1 U2375 ( .D0(n3378), .D1(n3379), .S(n3635), .Y(n3376) );
  NAND2X1 U2376 ( .A(n3381), .B(n3712), .Y(n3378) );
  MUX2X1 U2377 ( .D0(n3474), .D1(n3475), .S(n3655), .Y(n3456) );
  NOR4XL U2378 ( .A(n3695), .B(n3666), .C(n3641), .D(A[19]), .Y(n3475) );
  MUX2IX1 U2379 ( .D0(n3476), .D1(n3477), .S(n3635), .Y(n3474) );
  NAND2X1 U2380 ( .A(n3478), .B(n3718), .Y(n3477) );
  MUX2X1 U2381 ( .D0(n3627), .D1(n3628), .S(SH[4]), .Y(n3609) );
  NOR4XL U2382 ( .A(n3696), .B(n3667), .C(n3641), .D(A[16]), .Y(n3628) );
  MUX2IX1 U2383 ( .D0(n3629), .D1(n3630), .S(n3635), .Y(n3627) );
  NAND2X1 U2384 ( .A(n3631), .B(n3714), .Y(n3630) );
  MUX2X1 U2385 ( .D0(n3328), .D1(n3329), .S(n3655), .Y(n3310) );
  NOR4XL U2386 ( .A(n3696), .B(n3666), .C(n3636), .D(A[22]), .Y(n3329) );
  MUX2IX1 U2387 ( .D0(n3330), .D1(n3331), .S(n3635), .Y(n3328) );
  NAND2X1 U2388 ( .A(n3333), .B(n3718), .Y(n3330) );
  MUX2IX1 U2389 ( .D0(A[8]), .D1(A[264]), .S(n3665), .Y(n3631) );
  NAND2X1 U2390 ( .A(n3632), .B(n3711), .Y(n3629) );
  MUX2IX1 U2391 ( .D0(A[0]), .D1(A[256]), .S(n3659), .Y(n3632) );
  NAND2X1 U2392 ( .A(n3430), .B(n3718), .Y(n3427) );
  MUX2IX1 U2393 ( .D0(A[4]), .D1(A[260]), .S(n3660), .Y(n3430) );
  NAND2X1 U2394 ( .A(n3479), .B(n3718), .Y(n3476) );
  MUX2IX1 U2395 ( .D0(A[3]), .D1(A[259]), .S(n3659), .Y(n3479) );
  MUX2IX1 U2396 ( .D0(A[135]), .D1(A[391]), .S(n3664), .Y(n3262) );
  MUX2IX1 U2397 ( .D0(A[143]), .D1(A[399]), .S(n3664), .Y(n3260) );
  MUX4X1 U2398 ( .D0(n3249), .D1(n3250), .D2(n3251), .D3(n3252), .S0(n3652), 
        .S1(n3639), .Y(n3243) );
  AOI21X1 U2399 ( .B(A[207]), .C(n3684), .A(n3710), .Y(n3251) );
  AOI21X1 U2400 ( .B(A[199]), .C(n3683), .A(n3710), .Y(n3249) );
  AOI21X1 U2401 ( .B(A[215]), .C(n3684), .A(n3710), .Y(n3250) );
  MUX4X1 U2402 ( .D0(n3602), .D1(n3603), .D2(n3604), .D3(n3605), .S0(n3652), 
        .S1(n3639), .Y(n3583) );
  NOR3XL U2403 ( .A(A[152]), .B(n3701), .C(n3687), .Y(n3605) );
  NOR21XL U2404 ( .B(n3606), .A(n3693), .Y(n3604) );
  NOR21XL U2405 ( .B(n3607), .A(n3692), .Y(n3603) );
  MUX4X1 U2406 ( .D0(n3256), .D1(n3257), .D2(n3258), .D3(n3259), .S0(n3652), 
        .S1(n3637), .Y(n3241) );
  NOR3XL U2407 ( .A(A[159]), .B(n3708), .C(n3672), .Y(n3259) );
  NOR21XL U2408 ( .B(n3260), .A(n3692), .Y(n3258) );
  NOR21XL U2409 ( .B(n3262), .A(n3693), .Y(n3256) );
  MUX4X1 U2410 ( .D0(n3245), .D1(n3246), .D2(n3247), .D3(n3248), .S0(n3652), 
        .S1(n3639), .Y(n3244) );
  NOR3XL U2411 ( .A(A[239]), .B(n3703), .C(n3668), .Y(n3247) );
  NOR3XL U2412 ( .A(A[255]), .B(n3697), .C(n3668), .Y(n3248) );
  NOR3XL U2413 ( .A(A[231]), .B(n3708), .C(n3673), .Y(n3245) );
  MUX3X1 U2414 ( .D0(n3272), .D1(n3273), .D2(n3274), .S0(n3640), .S1(n3657), 
        .Y(n3265) );
  NOR4XL U2415 ( .A(n3696), .B(n3667), .C(A[63]), .D(n3649), .Y(n3274) );
  NOR3XL U2416 ( .A(A[47]), .B(n3708), .C(n3672), .Y(n3273) );
  NOR3XL U2417 ( .A(A[39]), .B(n3707), .C(n3672), .Y(n3272) );
  NOR21XL U2418 ( .B(n3608), .A(n3693), .Y(n3602) );
  MUX2IX1 U2419 ( .D0(A[128]), .D1(A[384]), .S(n3665), .Y(n3608) );
  NOR21XL U2420 ( .B(n3261), .A(n3693), .Y(n3257) );
  MUX2IX1 U2421 ( .D0(A[151]), .D1(A[407]), .S(n3665), .Y(n3261) );
  NOR3XL U2422 ( .A(A[167]), .B(n3707), .C(n3672), .Y(n3253) );
  NOR3XL U2423 ( .A(A[247]), .B(n3708), .C(n3673), .Y(n3246) );
  NOR3XL U2424 ( .A(A[223]), .B(n3707), .C(n3673), .Y(n3252) );
  INVX1 U2425 ( .A(n3691), .Y(n3685) );
  INVX1 U2426 ( .A(SH[8]), .Y(n3691) );
  INVX1 U2427 ( .A(SH[8]), .Y(n3689) );
  INVX1 U2428 ( .A(n3658), .Y(n3652) );
  INVX1 U2429 ( .A(SH[4]), .Y(n3658) );
  INVX1 U2430 ( .A(SH[3]), .Y(n3651) );
  AOI211X1 U2431 ( .C(n3641), .D(A[191]), .A(n3709), .B(n3673), .Y(n3255) );
  INVX1 U2432 ( .A(SH[8]), .Y(n3690) );
  INVX1 U2433 ( .A(SH[9]), .Y(n3718) );
  MUX2IX1 U2434 ( .D0(A[129]), .D1(A[385]), .S(n3661), .Y(n3556) );
  MUX2IX1 U2435 ( .D0(A[137]), .D1(A[393]), .S(n3661), .Y(n3554) );
  MUX2IX1 U2436 ( .D0(A[193]), .D1(A[449]), .S(n3661), .Y(n3545) );
  MUX2IX1 U2437 ( .D0(A[201]), .D1(A[457]), .S(n3663), .Y(n3543) );
  MUX2IX1 U2438 ( .D0(A[132]), .D1(A[388]), .S(n3661), .Y(n3406) );
  MUX2IX1 U2439 ( .D0(A[140]), .D1(A[396]), .S(n3661), .Y(n3404) );
  MUX2IX1 U2440 ( .D0(A[133]), .D1(A[389]), .S(n3662), .Y(n3357) );
  MUX2IX1 U2441 ( .D0(A[141]), .D1(A[397]), .S(n3662), .Y(n3355) );
  MUX2IX1 U2442 ( .D0(A[131]), .D1(A[387]), .S(n3660), .Y(n3455) );
  MUX2IX1 U2443 ( .D0(A[139]), .D1(A[395]), .S(n3660), .Y(n3453) );
  MUX2IX1 U2444 ( .D0(A[144]), .D1(A[400]), .S(n3665), .Y(n3607) );
  MUX2IX1 U2445 ( .D0(A[136]), .D1(A[392]), .S(n3664), .Y(n3606) );
  MUX2IX1 U2446 ( .D0(A[192]), .D1(A[448]), .S(n3664), .Y(n3597) );
  MUX2IX1 U2447 ( .D0(A[200]), .D1(A[456]), .S(n3663), .Y(n3595) );
  MUX2IX1 U2448 ( .D0(A[130]), .D1(A[386]), .S(n3659), .Y(n3504) );
  MUX2IX1 U2449 ( .D0(A[138]), .D1(A[394]), .S(n3659), .Y(n3502) );
  MUX2IX1 U2450 ( .D0(A[134]), .D1(A[390]), .S(n3664), .Y(n3309) );
  MUX2IX1 U2451 ( .D0(A[142]), .D1(A[398]), .S(n3664), .Y(n3307) );
  NOR21XL U2452 ( .B(n3308), .A(n3693), .Y(n3304) );
  MUX2IX1 U2453 ( .D0(A[150]), .D1(A[406]), .S(n3663), .Y(n3308) );
  MUX4X1 U2454 ( .D0(n3539), .D1(n3540), .D2(n3541), .D3(n3542), .S0(n3654), 
        .S1(n3639), .Y(n3533) );
  NOR3XL U2455 ( .A(A[217]), .B(n3699), .C(SH[8]), .Y(n3542) );
  NOR21XL U2456 ( .B(n3543), .A(n3693), .Y(n3541) );
  NOR21XL U2457 ( .B(n3545), .A(n3717), .Y(n3539) );
  MUX4X1 U2458 ( .D0(n3343), .D1(n3344), .D2(n3345), .D3(n3346), .S0(n3653), 
        .S1(n3637), .Y(n3338) );
  AOI21X1 U2459 ( .B(A[205]), .C(n3678), .A(n3710), .Y(n3345) );
  AOI21X1 U2460 ( .B(A[197]), .C(n3678), .A(n3710), .Y(n3343) );
  AOI21X1 U2461 ( .B(A[213]), .C(n3690), .A(n3709), .Y(n3344) );
  MUX4X1 U2462 ( .D0(n3591), .D1(n3592), .D2(n3593), .D3(n3594), .S0(n3652), 
        .S1(n3640), .Y(n3585) );
  NOR3XL U2463 ( .A(A[216]), .B(n3701), .C(n3687), .Y(n3594) );
  NOR21XL U2464 ( .B(n3595), .A(n3693), .Y(n3593) );
  NOR21XL U2465 ( .B(n3597), .A(n3694), .Y(n3591) );
  MUX4X1 U2466 ( .D0(n3546), .D1(n3547), .D2(n3548), .D3(n3549), .S0(n3653), 
        .S1(n3639), .Y(n3532) );
  NOR3XL U2467 ( .A(A[169]), .B(n3699), .C(n3688), .Y(n3548) );
  NOR3XL U2468 ( .A(A[185]), .B(n3699), .C(n3688), .Y(n3549) );
  NOR3XL U2469 ( .A(A[161]), .B(n3700), .C(n3685), .Y(n3546) );
  MUX4X1 U2470 ( .D0(n3396), .D1(n3397), .D2(n3398), .D3(n3399), .S0(n3654), 
        .S1(n3637), .Y(n3385) );
  NOR3XL U2471 ( .A(A[172]), .B(n3705), .C(n3671), .Y(n3398) );
  NOR3XL U2472 ( .A(A[188]), .B(n3705), .C(n3671), .Y(n3399) );
  NOR3XL U2473 ( .A(A[164]), .B(n3704), .C(n3670), .Y(n3396) );
  MUX4X1 U2474 ( .D0(n3347), .D1(n3348), .D2(n3349), .D3(n3350), .S0(n3653), 
        .S1(n3641), .Y(n3337) );
  NOR3XL U2475 ( .A(A[173]), .B(n3706), .C(n3685), .Y(n3349) );
  NOR3XL U2476 ( .A(A[189]), .B(n3706), .C(n3686), .Y(n3350) );
  NOR3XL U2477 ( .A(A[165]), .B(n3715), .C(n3685), .Y(n3347) );
  MUX4X1 U2478 ( .D0(n3445), .D1(n3446), .D2(n3447), .D3(n3448), .S0(n3657), 
        .S1(n3638), .Y(n3434) );
  NOR3XL U2479 ( .A(A[171]), .B(n3703), .C(n3669), .Y(n3447) );
  NOR3XL U2480 ( .A(A[187]), .B(n3703), .C(n3670), .Y(n3448) );
  NOR3XL U2481 ( .A(A[163]), .B(n3703), .C(n3669), .Y(n3445) );
  MUX4X1 U2482 ( .D0(n3598), .D1(n3599), .D2(n3600), .D3(n3601), .S0(n3652), 
        .S1(n3639), .Y(n3584) );
  NOR3XL U2483 ( .A(A[168]), .B(n3701), .C(n3688), .Y(n3600) );
  NOR3XL U2484 ( .A(A[184]), .B(n3701), .C(SH[8]), .Y(n3601) );
  NOR3XL U2485 ( .A(A[160]), .B(n3701), .C(n3688), .Y(n3598) );
  MUX4X1 U2486 ( .D0(n3494), .D1(n3495), .D2(n3496), .D3(n3497), .S0(n3657), 
        .S1(n3638), .Y(n3483) );
  NOR3XL U2487 ( .A(A[170]), .B(n3697), .C(n3668), .Y(n3496) );
  NOR3XL U2488 ( .A(A[186]), .B(n3697), .C(n3668), .Y(n3497) );
  NOR3XL U2489 ( .A(A[162]), .B(n3698), .C(n3668), .Y(n3494) );
  MUX4X1 U2490 ( .D0(n3550), .D1(n3551), .D2(n3552), .D3(n3553), .S0(n3653), 
        .S1(n3639), .Y(n3531) );
  NOR3XL U2491 ( .A(A[153]), .B(n3700), .C(SH[8]), .Y(n3553) );
  NOR21XL U2492 ( .B(n3554), .A(n3717), .Y(n3552) );
  NOR21XL U2493 ( .B(n3556), .A(n3717), .Y(n3550) );
  MUX4X1 U2494 ( .D0(n3400), .D1(n3401), .D2(n3402), .D3(n3403), .S0(n3654), 
        .S1(n3637), .Y(n3384) );
  NOR3XL U2495 ( .A(A[156]), .B(n3704), .C(n3670), .Y(n3403) );
  NOR21XL U2496 ( .B(n3404), .A(n3717), .Y(n3402) );
  NOR21XL U2497 ( .B(n3406), .A(n3717), .Y(n3400) );
  MUX4X1 U2498 ( .D0(n3351), .D1(n3352), .D2(n3353), .D3(n3354), .S0(n3653), 
        .S1(n3641), .Y(n3336) );
  NOR3XL U2499 ( .A(A[157]), .B(n3715), .C(n3686), .Y(n3354) );
  NOR21XL U2500 ( .B(n3355), .A(n3716), .Y(n3353) );
  NOR21XL U2501 ( .B(n3357), .A(n3716), .Y(n3351) );
  MUX4X1 U2502 ( .D0(n3449), .D1(n3450), .D2(n3451), .D3(n3452), .S0(n3657), 
        .S1(n3638), .Y(n3433) );
  NOR3XL U2503 ( .A(A[155]), .B(n3702), .C(n3669), .Y(n3452) );
  NOR21XL U2504 ( .B(n3453), .A(n3692), .Y(n3451) );
  NOR21XL U2505 ( .B(n3455), .A(n3692), .Y(n3449) );
  MUX4X1 U2506 ( .D0(n3498), .D1(n3499), .D2(n3500), .D3(n3501), .S0(n3654), 
        .S1(n3638), .Y(n3482) );
  NOR3XL U2507 ( .A(A[154]), .B(n3698), .C(n3673), .Y(n3501) );
  NOR21XL U2508 ( .B(n3502), .A(n3717), .Y(n3500) );
  NOR21XL U2509 ( .B(n3504), .A(n3695), .Y(n3498) );
  MUX4X1 U2510 ( .D0(n3303), .D1(n3304), .D2(n3305), .D3(n3306), .S0(n3653), 
        .S1(SH[3]), .Y(n3289) );
  NOR3XL U2511 ( .A(A[158]), .B(n3707), .C(n3672), .Y(n3306) );
  NOR21XL U2512 ( .B(n3307), .A(n3693), .Y(n3305) );
  NOR21XL U2513 ( .B(n3309), .A(SH[9]), .Y(n3303) );
  MUX4X1 U2514 ( .D0(n3388), .D1(n3389), .D2(n3390), .D3(n3391), .S0(n3654), 
        .S1(n3637), .Y(n3387) );
  NOR3XL U2515 ( .A(A[236]), .B(n3705), .C(n3671), .Y(n3390) );
  NOR3XL U2516 ( .A(A[252]), .B(n3705), .C(n3671), .Y(n3391) );
  NOR3XL U2517 ( .A(A[228]), .B(n3705), .C(n3671), .Y(n3388) );
  MUX4X1 U2518 ( .D0(n3437), .D1(n3438), .D2(n3439), .D3(n3440), .S0(n3654), 
        .S1(n3638), .Y(n3436) );
  NOR3XL U2519 ( .A(A[235]), .B(n3703), .C(n3670), .Y(n3439) );
  NOR3XL U2520 ( .A(A[251]), .B(n3703), .C(n3670), .Y(n3440) );
  NOR3XL U2521 ( .A(A[227]), .B(n3703), .C(n3670), .Y(n3437) );
  MUX4X1 U2522 ( .D0(n3486), .D1(n3487), .D2(n3488), .D3(n3489), .S0(n3657), 
        .S1(n3637), .Y(n3485) );
  NOR3XL U2523 ( .A(A[234]), .B(n3697), .C(n3669), .Y(n3488) );
  NOR3XL U2524 ( .A(A[250]), .B(n3698), .C(n3669), .Y(n3489) );
  NOR3XL U2525 ( .A(A[226]), .B(n3697), .C(n3669), .Y(n3486) );
  MUX3X1 U2526 ( .D0(n3566), .D1(n3567), .D2(n3568), .S0(n3640), .S1(n3656), 
        .Y(n3559) );
  NOR4XL U2527 ( .A(n3695), .B(n3666), .C(A[57]), .D(n3642), .Y(n3568) );
  NOR3XL U2528 ( .A(A[41]), .B(n3700), .C(n3667), .Y(n3567) );
  NOR3XL U2529 ( .A(A[33]), .B(n3700), .C(n3667), .Y(n3566) );
  MUX3X1 U2530 ( .D0(n3416), .D1(n3417), .D2(n3418), .S0(n3640), .S1(n3656), 
        .Y(n3409) );
  NOR4XL U2531 ( .A(n3696), .B(n3666), .C(A[60]), .D(n3645), .Y(n3418) );
  NOR3XL U2532 ( .A(A[44]), .B(n3704), .C(n3670), .Y(n3417) );
  NOR3XL U2533 ( .A(A[36]), .B(n3704), .C(n3670), .Y(n3416) );
  MUX3X1 U2534 ( .D0(n3367), .D1(n3368), .D2(n3369), .S0(n3640), .S1(n3656), 
        .Y(n3360) );
  NOR4XL U2535 ( .A(n3696), .B(n3666), .C(A[61]), .D(n3646), .Y(n3369) );
  NOR3XL U2536 ( .A(A[45]), .B(n3705), .C(n3671), .Y(n3368) );
  NOR3XL U2537 ( .A(A[37]), .B(n3717), .C(n3671), .Y(n3367) );
  MUX3X1 U2538 ( .D0(n3465), .D1(n3466), .D2(n3467), .S0(n3641), .S1(n3656), 
        .Y(n3458) );
  NOR4XL U2539 ( .A(n3695), .B(n3667), .C(A[59]), .D(n3644), .Y(n3467) );
  NOR3XL U2540 ( .A(A[43]), .B(n3698), .C(n3669), .Y(n3466) );
  NOR3XL U2541 ( .A(A[35]), .B(n3697), .C(n3669), .Y(n3465) );
  MUX3X1 U2542 ( .D0(n3618), .D1(n3619), .D2(n3620), .S0(n3640), .S1(n3657), 
        .Y(n3611) );
  NOR4XL U2543 ( .A(n3695), .B(n3667), .C(A[56]), .D(n3648), .Y(n3620) );
  NOR3XL U2544 ( .A(A[40]), .B(n3702), .C(n3688), .Y(n3619) );
  NOR3XL U2545 ( .A(A[32]), .B(n3702), .C(n3668), .Y(n3618) );
  MUX3X1 U2546 ( .D0(n3514), .D1(n3515), .D2(n3516), .S0(n3640), .S1(n3656), 
        .Y(n3507) );
  NOR4XL U2547 ( .A(n3696), .B(n3667), .C(A[58]), .D(n3643), .Y(n3516) );
  NOR3XL U2548 ( .A(A[42]), .B(n3698), .C(n3668), .Y(n3515) );
  NOR3XL U2549 ( .A(A[34]), .B(n3699), .C(n3688), .Y(n3514) );
  NOR21XL U2550 ( .B(n3555), .A(n3694), .Y(n3551) );
  MUX2IX1 U2551 ( .D0(A[145]), .D1(A[401]), .S(n3661), .Y(n3555) );
  NOR21XL U2552 ( .B(n3544), .A(n3694), .Y(n3540) );
  MUX2IX1 U2553 ( .D0(A[209]), .D1(A[465]), .S(n3660), .Y(n3544) );
  NOR21XL U2554 ( .B(n3405), .A(SH[9]), .Y(n3401) );
  MUX2IX1 U2555 ( .D0(A[148]), .D1(A[404]), .S(n3661), .Y(n3405) );
  NOR21XL U2556 ( .B(n3356), .A(n3694), .Y(n3352) );
  MUX2IX1 U2557 ( .D0(A[149]), .D1(A[405]), .S(n3662), .Y(n3356) );
  NOR21XL U2558 ( .B(n3454), .A(n3692), .Y(n3450) );
  MUX2IX1 U2559 ( .D0(A[147]), .D1(A[403]), .S(n3660), .Y(n3454) );
  NOR21XL U2560 ( .B(n3596), .A(n3694), .Y(n3592) );
  MUX2IX1 U2561 ( .D0(A[208]), .D1(A[464]), .S(n3664), .Y(n3596) );
  NOR21XL U2562 ( .B(n3503), .A(n3717), .Y(n3499) );
  MUX2IX1 U2563 ( .D0(A[146]), .D1(A[402]), .S(n3659), .Y(n3503) );
  AOI211X1 U2564 ( .C(A[245]), .D(n3650), .A(n3708), .B(n3673), .Y(n3342) );
  NOR3XL U2565 ( .A(A[237]), .B(n3706), .C(n3685), .Y(n3341) );
  AOI21X1 U2566 ( .B(A[204]), .C(n3680), .A(n3710), .Y(n3394) );
  AOI21X1 U2567 ( .B(A[203]), .C(n3683), .A(n3709), .Y(n3443) );
  AOI21X1 U2568 ( .B(A[202]), .C(n3680), .A(n3710), .Y(n3492) );
  AOI21X1 U2569 ( .B(A[212]), .C(n3682), .A(n3709), .Y(n3393) );
  AOI21X1 U2570 ( .B(A[211]), .C(n3683), .A(n3710), .Y(n3442) );
  AOI21X1 U2571 ( .B(A[210]), .C(n3679), .A(n3709), .Y(n3491) );
  AOI21X1 U2572 ( .B(A[196]), .C(n3691), .A(n3709), .Y(n3392) );
  AOI21X1 U2573 ( .B(A[195]), .C(n3682), .A(n3709), .Y(n3441) );
  AOI21X1 U2574 ( .B(A[194]), .C(n3684), .A(n3710), .Y(n3490) );
  NOR3XL U2575 ( .A(A[229]), .B(n3705), .C(n3686), .Y(n3340) );
  NOR3XL U2576 ( .A(A[221]), .B(n3715), .C(n3685), .Y(n3346) );
  NOR3XL U2577 ( .A(A[244]), .B(n3704), .C(n3671), .Y(n3389) );
  NOR3XL U2578 ( .A(A[233]), .B(n3702), .C(n3668), .Y(n3537) );
  NOR3XL U2579 ( .A(A[232]), .B(n3701), .C(n3667), .Y(n3589) );
  NOR3XL U2580 ( .A(A[243]), .B(n3703), .C(n3670), .Y(n3438) );
  NOR3XL U2581 ( .A(A[242]), .B(n3698), .C(n3669), .Y(n3487) );
  NOR3XL U2582 ( .A(A[241]), .B(n3699), .C(SH[8]), .Y(n3536) );
  NOR3XL U2583 ( .A(A[240]), .B(n3701), .C(n3667), .Y(n3588) );
  NOR3XL U2584 ( .A(A[177]), .B(n3699), .C(n3673), .Y(n3547) );
  NOR3XL U2585 ( .A(A[180]), .B(n3705), .C(n3671), .Y(n3397) );
  NOR3XL U2586 ( .A(A[181]), .B(n3715), .C(n3685), .Y(n3348) );
  NOR3XL U2587 ( .A(A[179]), .B(n3703), .C(n3669), .Y(n3446) );
  NOR3XL U2588 ( .A(A[176]), .B(n3701), .C(SH[8]), .Y(n3599) );
  NOR3XL U2589 ( .A(A[178]), .B(n3697), .C(n3668), .Y(n3495) );
  NOR3XL U2590 ( .A(A[224]), .B(n3701), .C(n3688), .Y(n3587) );
  NOR3XL U2591 ( .A(A[249]), .B(n3699), .C(SH[8]), .Y(n3538) );
  NOR3XL U2592 ( .A(A[219]), .B(n3703), .C(n3670), .Y(n3444) );
  NOR3XL U2593 ( .A(A[248]), .B(n3700), .C(n3687), .Y(n3590) );
  NOR3XL U2594 ( .A(A[225]), .B(n3699), .C(n3688), .Y(n3535) );
  NOR3XL U2595 ( .A(A[220]), .B(n3705), .C(n3671), .Y(n3395) );
  NOR3XL U2596 ( .A(A[218]), .B(n3697), .C(n3668), .Y(n3493) );
  MUX4X1 U2597 ( .D0(n3297), .D1(n3298), .D2(n3299), .D3(n3300), .S0(n3652), 
        .S1(SH[3]), .Y(n3291) );
  AOI21X1 U2598 ( .B(A[206]), .C(n3683), .A(n3709), .Y(n3299) );
  AOI21X1 U2599 ( .B(A[198]), .C(n3682), .A(n3709), .Y(n3297) );
  AOI21X1 U2600 ( .B(A[214]), .C(n3681), .A(n3710), .Y(n3298) );
  MUX4X1 U2601 ( .D0(n3293), .D1(n3294), .D2(n3295), .D3(n3296), .S0(n3652), 
        .S1(SH[3]), .Y(n3292) );
  NOR3XL U2602 ( .A(A[238]), .B(n3706), .C(n3672), .Y(n3295) );
  NOR3XL U2603 ( .A(A[254]), .B(n3707), .C(n3672), .Y(n3296) );
  NOR3XL U2604 ( .A(A[230]), .B(n3706), .C(n3672), .Y(n3293) );
  AOI211X1 U2605 ( .C(A[166]), .D(n3650), .A(n3709), .B(n3673), .Y(n3301) );
  AOI211X1 U2606 ( .C(n3641), .D(A[190]), .A(n3708), .B(n3673), .Y(n3302) );
  MUX3X1 U2607 ( .D0(n3319), .D1(n3320), .D2(n3321), .S0(n3640), .S1(n3656), 
        .Y(n3312) );
  NOR4XL U2608 ( .A(n3696), .B(n3666), .C(A[62]), .D(n3647), .Y(n3321) );
  NOR3XL U2609 ( .A(A[38]), .B(n3715), .C(n3686), .Y(n3319) );
  NOR3XL U2610 ( .A(A[46]), .B(n3706), .C(n3685), .Y(n3320) );
  NOR3XL U2611 ( .A(A[246]), .B(n3708), .C(n3672), .Y(n3294) );
  NOR3XL U2612 ( .A(A[222]), .B(n3707), .C(n3672), .Y(n3300) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regx_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N16, N17, N18, N19, N20,
         net8993, n12, n3, n4, n5, n6, n7, n8, n9, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net8993), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N20), .SIN(db_cnt_2_), .SMC(test_se), .C(net8993), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N18), .SIN(db_cnt_0_), .SMC(test_se), .C(net8993), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N17), .SIN(o_dbc), .SMC(test_se), .C(net8993), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N19), .SIN(db_cnt_1_), .SMC(test_se), .C(net8993), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n12), .SIN(d_org_0_), .SMC(test_se), .C(net8993), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n6), .Y(n1) );
  NOR21XL U4 ( .B(n3), .A(n4), .Y(n6) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  OAI22X1 U6 ( .A(db_cnt_2_), .B(n5), .C(n7), .D(n2), .Y(N19) );
  AOI21BBXL U7 ( .B(n1), .C(db_cnt_1_), .A(N17), .Y(n7) );
  AO22AXL U8 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR2X1 U9 ( .A(n3), .B(n4), .Y(o_chg) );
  NOR2X1 U10 ( .A(n1), .B(db_cnt_0_), .Y(N17) );
  NAND4X1 U11 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(db_cnt_0_), .Y(
        n3) );
  NAND3X1 U12 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(n6), .Y(n5) );
  ENOX1 U13 ( .A(n2), .B(n5), .C(test_so), .D(n6), .Y(N20) );
  NOR2X1 U14 ( .A(n8), .B(n1), .Y(N18) );
  XNOR2XL U15 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n8) );
  NAND31X1 U16 ( .C(db_cnt_0_), .A(n4), .B(n9), .Y(N16) );
  NOR3XL U17 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n9) );
  INVX1 U18 ( .A(db_cnt_2_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N16, N17, N18, N19, N20,
         net9011, n12, n3, n4, n5, n6, n7, n8, n9, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9011), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N20), .SIN(db_cnt_2_), .SMC(test_se), .C(net9011), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N18), .SIN(db_cnt_0_), .SMC(test_se), .C(net9011), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N17), .SIN(o_dbc), .SMC(test_se), .C(net9011), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N19), .SIN(db_cnt_1_), .SMC(test_se), .C(net9011), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n12), .SIN(d_org_0_), .SMC(test_se), .C(net9011), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n6), .Y(n1) );
  NOR21XL U4 ( .B(n3), .A(n4), .Y(n6) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  OAI22X1 U6 ( .A(db_cnt_2_), .B(n5), .C(n7), .D(n2), .Y(N19) );
  AOI21BBXL U7 ( .B(n1), .C(db_cnt_1_), .A(N17), .Y(n7) );
  AO22AXL U8 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR2X1 U9 ( .A(n3), .B(n4), .Y(o_chg) );
  NOR2X1 U10 ( .A(n1), .B(db_cnt_0_), .Y(N17) );
  NAND4X1 U11 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(db_cnt_0_), .Y(
        n3) );
  NAND3X1 U12 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(n6), .Y(n5) );
  ENOX1 U13 ( .A(n2), .B(n5), .C(test_so), .D(n6), .Y(N20) );
  NOR2X1 U14 ( .A(n8), .B(n1), .Y(N18) );
  XNOR2XL U15 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n8) );
  NAND31X1 U16 ( .C(db_cnt_0_), .A(n4), .B(n9), .Y(N16) );
  NOR3XL U17 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n9) );
  INVX1 U18 ( .A(db_cnt_2_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_4 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_5 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_6 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module glreg_a0_7 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9029;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_7 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9029), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9029), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9029), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9029), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9029), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9029), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9029), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9029), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9029), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_8 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9047;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_8 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9047), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9047), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9047), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9047), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9047), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9047), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9047), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9047), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9047), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_9 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9065;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_9 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9065), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9065), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9065), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9065), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9065), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9065), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9065), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9065), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9065), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH7_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9083;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9083), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9083), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9083), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9083), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9083), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9083), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9083), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9083), 
        .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_7 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module glreg_a0_10 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9101;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_10 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9101), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9101), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9101), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9101), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9101), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9101), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9101), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9101), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9101), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_11 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9119;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_11 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9119), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9119), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9119), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9119), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9119), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9119), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9119), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9119), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9119), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_12 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9137;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_12 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9137), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9137), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9137), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9137), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9137), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9137), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9137), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9137), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9137), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_13 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9155;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_13 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9155), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9155), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9155), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9155), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9155), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9155), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9155), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9155), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9155), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_14 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9173;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_14 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9173), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9173), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9173), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9173), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9173), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9173), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9173), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9173), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9173), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9191;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9191), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9191), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9191), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9191), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9191), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9191), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9191), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9209;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9209), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9209), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9209), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9209), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9209), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9209), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9209), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_15 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9227;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_15 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9227), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9227), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9227), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9227), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9227), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9227), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9227), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9227), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9227), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_6_00000002 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9245;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9245), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9245), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9245), 
        .XS(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9245), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9245), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9245), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9245), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_a0_16 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9263;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_16 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9263), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9263), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9263), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9263), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9263), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9263), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9263), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9263), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9263), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_17 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9281;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_17 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9281), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9281), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9281), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9281), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9281), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9281), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9281), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9281), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9281), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_18 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9299;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_18 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9299), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9299), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9299), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9299), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9299), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9299), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9299), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9299), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9299), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module cvctl_a0 ( r_cvcwr, wdat, r_sdischg, r_vcomp, r_idacsh, r_cvofsx, 
        r_cvofs, sdischg_duty, r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, 
        r_fw_pwrv, r_dac0, r_dac3, clk_100k, clk, srstz, test_si, test_se );
  input [5:0] r_cvcwr;
  input [7:0] wdat;
  output [7:0] r_sdischg;
  output [7:0] r_vcomp;
  output [7:0] r_idacsh;
  output [7:0] r_cvofsx;
  output [15:0] r_cvofs;
  input [11:0] r_fw_pwrv;
  output [10:0] r_dac0;
  output [5:0] r_dac3;
  input r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, clk_100k, clk, srstz,
         test_si, test_se;
  output sdischg_duty;
  wire   clk_5k, N29, N34, N35, N36, N38, N39, N40, N41, N42, N47, N84, N94,
         N95, N96, N97, N98, N99, N106, N107, N108, N109, N115, N121, N122,
         N123, N126, N127, N128, N129, N130, net9317, n81, N68, N67, N66, N65,
         N64, N63, N62, N61, N60, n2, n4, n5, n6, n7, n8, n9, N83, N82, N81,
         N80, N79, N78, N77, N76, N75, N74, N73, N72, N59, N58, N57, N56, N55,
         N54, N53, N52, N51, N50, N49, N48, n34, n35, n36, n37, n38, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, add_62_carry_1_, add_62_carry_2_, add_62_carry_3_,
         add_62_carry_4_, add_62_carry_5_, n3, n12, n17, n18, n19, n20, n21,
         n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33;
  wire   [4:0] div20_cnt;
  wire   [10:1] cv_code;
  wire   [4:0] sdischg_cnt;
  wire   [4:2] add_81_carry;
  wire   [4:2] add_41_carry;
  wire   [2:1] add_3_root_sub_0_root_add_46_3_carry;

  HAD1X1 add_81_U1_1_1 ( .A(sdischg_cnt[1]), .B(sdischg_cnt[0]), .CO(
        add_81_carry[2]), .SO(N121) );
  HAD1X1 add_81_U1_1_2 ( .A(sdischg_cnt[2]), .B(add_81_carry[2]), .CO(
        add_81_carry[3]), .SO(N122) );
  HAD1X1 add_81_U1_1_3 ( .A(sdischg_cnt[3]), .B(add_81_carry[3]), .CO(
        add_81_carry[4]), .SO(N123) );
  HAD1X1 add_41_U1_1_1 ( .A(div20_cnt[1]), .B(div20_cnt[0]), .CO(
        add_41_carry[2]), .SO(N34) );
  HAD1X1 add_41_U1_1_2 ( .A(div20_cnt[2]), .B(add_41_carry[2]), .CO(
        add_41_carry[3]), .SO(N35) );
  HAD1X1 add_41_U1_1_3 ( .A(div20_cnt[3]), .B(add_41_carry[3]), .CO(
        add_41_carry[4]), .SO(N36) );
  FAD1X1 add_3_root_sub_0_root_add_46_3_U1_1 ( .A(N47), .B(r_vcomp[1]), .CI(
        add_3_root_sub_0_root_add_46_3_carry[1]), .CO(
        add_3_root_sub_0_root_add_46_3_carry[2]), .SO(N61) );
  INVX1 U4 ( .A(n9), .Y(n8) );
  INVX1 U5 ( .A(n9), .Y(n4) );
  INVX1 U6 ( .A(n9), .Y(n5) );
  INVX1 U7 ( .A(n9), .Y(n6) );
  INVX1 U8 ( .A(n9), .Y(n7) );
  INVX1 U9 ( .A(n9), .Y(n2) );
  INVX1 U10 ( .A(srstz), .Y(n9) );
  glreg_a0_24 u0_v_comp ( .clk(clk), .arstz(n8), .we(r_cvcwr[3]), .wdat(wdat), 
        .rdat(r_vcomp), .test_si(r_sdischg[7]), .test_se(test_se) );
  glreg_a0_23 u0_idac_shift ( .clk(clk), .arstz(n7), .we(r_cvcwr[4]), .wdat(
        wdat), .rdat(r_idacsh), .test_si(r_cvofs[15]), .test_se(test_se) );
  glreg_a0_22 u0_cv_ofsx ( .clk(clk), .arstz(n6), .we(r_cvcwr[5]), .wdat(wdat), 
        .rdat(r_cvofsx), .test_si(sdischg_duty), .test_se(test_se) );
  glreg_a0_21 u0_cvofs01 ( .clk(clk), .arstz(n5), .we(r_cvcwr[0]), .wdat(wdat), 
        .rdat(r_cvofs[7:0]), .test_si(r_cvofsx[7]), .test_se(test_se) );
  glreg_a0_20 u0_cvofs23 ( .clk(clk), .arstz(n4), .we(r_cvcwr[1]), .wdat(wdat), 
        .rdat(r_cvofs[15:8]), .test_si(r_cvofs[7]), .test_se(test_se) );
  glreg_a0_19 u0_sdischg ( .clk(clk), .arstz(n2), .we(r_cvcwr[2]), .wdat(wdat), 
        .rdat(r_sdischg), .test_si(r_idacsh[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_cvctl_a0 clk_gate_sdischg_cnt_reg ( .CLK(clk_100k), 
        .EN(N115), .ENCLK(net9317), .TE(test_se) );
  cvctl_a0_DW01_sub_1 sub_2_root_sub_0_root_add_46_3 ( .A(r_fw_pwrv), .B({1'b0, 
        1'b0, 1'b0, 1'b0, r_idacsh}), .CI(1'b0), .DIFF({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .CO() );
  cvctl_a0_DW01_add_2 add_1_root_sub_0_root_add_46_3 ( .A({r_cvofsx[7], 
        r_cvofsx[7], r_cvofsx[7], r_cvofsx[7], r_cvofsx}), .B({1'b0, 1'b0, 
        1'b0, N68, N67, N66, N65, N64, N63, N62, N61, N60}), .CI(1'b0), .SUM({
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}), .CO() );
  cvctl_a0_DW01_add_1 add_0_root_sub_0_root_add_46_3 ( .A({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .B({N83, N82, N81, N80, N79, 
        N78, N77, N76, N75, N74, N73, N72}), .CI(1'b0), .SUM({N84, cv_code, 
        r_dac0[0]}), .CO() );
  FAD1X1 add_62_U1_1 ( .A(N95), .B(N107), .CI(add_62_carry_1_), .CO(
        add_62_carry_2_), .SO(r_dac3[1]) );
  FAD1X1 add_62_U1_2 ( .A(N96), .B(N108), .CI(add_62_carry_2_), .CO(
        add_62_carry_3_), .SO(r_dac3[2]) );
  FAD1X1 add_62_U1_3 ( .A(N97), .B(N109), .CI(add_62_carry_3_), .CO(
        add_62_carry_4_), .SO(r_dac3[3]) );
  SDFFRQX1 sdischg_cnt_reg_0_ ( .D(N126), .SIN(div20_cnt[4]), .SMC(test_se), 
        .C(net9317), .XR(srstz), .Q(sdischg_cnt[0]) );
  SDFFRQX1 sdischg_cnt_reg_4_ ( .D(N130), .SIN(sdischg_cnt[3]), .SMC(test_se), 
        .C(net9317), .XR(n6), .Q(sdischg_cnt[4]) );
  SDFFRQX1 sdischg_cnt_reg_1_ ( .D(N127), .SIN(sdischg_cnt[0]), .SMC(test_se), 
        .C(net9317), .XR(srstz), .Q(sdischg_cnt[1]) );
  SDFFRQX1 sdischg_cnt_reg_2_ ( .D(N128), .SIN(sdischg_cnt[1]), .SMC(test_se), 
        .C(net9317), .XR(n4), .Q(sdischg_cnt[2]) );
  SDFFRQX1 div20_cnt_reg_2_ ( .D(N40), .SIN(div20_cnt[1]), .SMC(test_se), .C(
        clk_100k), .XR(n2), .Q(div20_cnt[2]) );
  SDFFRQX1 div20_cnt_reg_1_ ( .D(N39), .SIN(div20_cnt[0]), .SMC(test_se), .C(
        clk_100k), .XR(n5), .Q(div20_cnt[1]) );
  SDFFRQX1 div20_cnt_reg_3_ ( .D(N41), .SIN(div20_cnt[2]), .SMC(test_se), .C(
        clk_100k), .XR(n4), .Q(div20_cnt[3]) );
  SDFFRQX1 div20_cnt_reg_0_ ( .D(N38), .SIN(clk_5k), .SMC(test_se), .C(
        clk_100k), .XR(n8), .Q(div20_cnt[0]) );
  SDFFRQX1 div20_cnt_reg_4_ ( .D(N42), .SIN(div20_cnt[3]), .SMC(test_se), .C(
        clk_100k), .XR(n8), .Q(div20_cnt[4]) );
  SDFFRQX1 sdischg_cnt_reg_3_ ( .D(N129), .SIN(sdischg_cnt[2]), .SMC(test_se), 
        .C(net9317), .XR(n7), .Q(sdischg_cnt[3]) );
  SDFFRQX1 sdischg_reg ( .D(n81), .SIN(sdischg_cnt[4]), .SMC(test_se), .C(
        net9317), .XR(n6), .Q(sdischg_duty) );
  SDFFRQX1 clk_5k_reg ( .D(N29), .SIN(test_si), .SMC(test_se), .C(clk_100k), 
        .XR(n5), .Q(clk_5k) );
  INVX1 U11 ( .A(N84), .Y(n3) );
  INVX1 U14 ( .A(N98), .Y(n12) );
  NOR2X1 U19 ( .A(n26), .B(n52), .Y(n50) );
  NOR2X1 U20 ( .A(n72), .B(r_dac0[10]), .Y(n75) );
  NOR2X1 U21 ( .A(n76), .B(r_dac0[9]), .Y(n73) );
  INVX1 U22 ( .A(n76), .Y(r_dac0[10]) );
  NOR2X1 U23 ( .A(n23), .B(cv_code[1]), .Y(N94) );
  NOR2X1 U24 ( .A(n51), .B(n23), .Y(N98) );
  XNOR2XL U25 ( .A(cv_code[5]), .B(n50), .Y(n51) );
  NAND2X1 U26 ( .A(n28), .B(n23), .Y(r_dac0[1]) );
  NAND2X1 U27 ( .A(n27), .B(n23), .Y(r_dac0[2]) );
  NAND2X1 U28 ( .A(n25), .B(n3), .Y(r_dac0[6]) );
  NAND2X1 U29 ( .A(n26), .B(n3), .Y(r_dac0[4]) );
  INVX1 U30 ( .A(cv_code[2]), .Y(n27) );
  INVX1 U31 ( .A(cv_code[4]), .Y(n26) );
  XNOR2XL U32 ( .A(cv_code[2]), .B(cv_code[1]), .Y(n55) );
  INVX1 U33 ( .A(cv_code[6]), .Y(n25) );
  NAND2X1 U34 ( .A(cv_code[5]), .B(n50), .Y(n49) );
  INVX1 U35 ( .A(cv_code[1]), .Y(n28) );
  NAND3X1 U36 ( .A(cv_code[2]), .B(cv_code[1]), .C(cv_code[3]), .Y(n52) );
  NOR2X1 U37 ( .A(N84), .B(cv_code[10]), .Y(n76) );
  XOR2X1 U38 ( .A(add_62_carry_4_), .B(N98), .Y(r_dac3[4]) );
  XOR2X1 U39 ( .A(N99), .B(add_62_carry_5_), .Y(r_dac3[5]) );
  NOR2X1 U40 ( .A(n48), .B(n23), .Y(N99) );
  NOR21XL U41 ( .B(add_62_carry_4_), .A(n12), .Y(add_62_carry_5_) );
  XNOR2XL U42 ( .A(n49), .B(n25), .Y(n48) );
  INVX1 U43 ( .A(N106), .Y(n17) );
  NOR2X1 U44 ( .A(r_dac0[10]), .B(cv_code[9]), .Y(n72) );
  INVX1 U45 ( .A(N84), .Y(n23) );
  NAND21X1 U46 ( .B(cv_code[9]), .A(n23), .Y(r_dac0[9]) );
  OAI21BBX1 U47 ( .A(cv_code[10]), .B(cv_code[9]), .C(n23), .Y(n74) );
  XOR2X1 U48 ( .A(N94), .B(N106), .Y(r_dac3[0]) );
  NOR3XL U49 ( .A(n29), .B(n58), .C(n30), .Y(n56) );
  OR2X1 U50 ( .A(cv_code[7]), .B(N84), .Y(r_dac0[7]) );
  OR2X1 U51 ( .A(cv_code[8]), .B(N84), .Y(r_dac0[8]) );
  OR2X1 U52 ( .A(cv_code[3]), .B(N84), .Y(r_dac0[3]) );
  OR2X1 U53 ( .A(cv_code[5]), .B(N84), .Y(r_dac0[5]) );
  NOR21XL U54 ( .B(N35), .A(n62), .Y(N40) );
  NOR21XL U55 ( .B(N36), .A(n62), .Y(N41) );
  NOR21XL U56 ( .B(N34), .A(n62), .Y(N39) );
  INVX1 U57 ( .A(n37), .Y(n19) );
  NOR21XL U58 ( .B(N123), .A(n37), .Y(N129) );
  NOR21XL U59 ( .B(N122), .A(n37), .Y(N128) );
  NOR21XL U60 ( .B(N121), .A(n37), .Y(N127) );
  NOR2X1 U61 ( .A(n53), .B(n23), .Y(N97) );
  AO2222XL U62 ( .A(r_cvofs[7]), .B(n72), .C(r_cvofs[15]), .D(n73), .E(
        r_cvofs[14]), .F(n74), .G(r_cvofs[6]), .H(n75), .Y(N109) );
  XNOR2XL U63 ( .A(n52), .B(n26), .Y(n53) );
  XOR2X1 U64 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .Y(N62) );
  XNOR2XL U65 ( .A(r_vcomp[3]), .B(n60), .Y(N63) );
  NAND2X1 U66 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .Y(n60) );
  XNOR2XL U67 ( .A(r_vcomp[4]), .B(n58), .Y(N64) );
  XNOR2XL U68 ( .A(n59), .B(n30), .Y(N65) );
  NOR2X1 U69 ( .A(n58), .B(n29), .Y(n59) );
  XOR2X1 U70 ( .A(n56), .B(r_vcomp[6]), .Y(N66) );
  XNOR2XL U71 ( .A(r_vcomp[7]), .B(n57), .Y(N67) );
  NAND2X1 U72 ( .A(r_vcomp[6]), .B(n56), .Y(n57) );
  GEN2XL U73 ( .D(N84), .E(n27), .C(N94), .B(cv_code[3]), .A(n54), .Y(N96) );
  AO2222XL U74 ( .A(r_cvofs[2]), .B(n72), .C(r_cvofs[10]), .D(n73), .E(
        r_cvofs[13]), .F(n74), .G(r_cvofs[5]), .H(n75), .Y(N108) );
  NOR4XL U75 ( .A(cv_code[3]), .B(n28), .C(n27), .D(n23), .Y(n54) );
  NOR32XL U76 ( .B(r_hlsb_en), .C(clk_5k), .A(r_hlsb_sel), .Y(N47) );
  NOR21XL U77 ( .B(r_vcomp[0]), .A(n47), .Y(
        add_3_root_sub_0_root_add_46_3_carry[1]) );
  AND3X1 U78 ( .A(r_vcomp[7]), .B(n56), .C(r_vcomp[6]), .Y(N68) );
  AO2222XL U79 ( .A(r_cvofs[0]), .B(n72), .C(r_cvofs[8]), .D(n73), .E(
        r_cvofs[11]), .F(n74), .G(r_cvofs[3]), .H(n75), .Y(N106) );
  NOR2X1 U80 ( .A(n55), .B(n23), .Y(N95) );
  AO2222XL U81 ( .A(r_cvofs[1]), .B(n72), .C(r_cvofs[9]), .D(n73), .E(
        r_cvofs[12]), .F(n74), .G(r_cvofs[4]), .H(n75), .Y(N107) );
  NOR21XL U82 ( .B(N94), .A(n17), .Y(add_62_carry_1_) );
  XNOR2XL U83 ( .A(r_vcomp[0]), .B(n47), .Y(N60) );
  NAND3X1 U84 ( .A(r_hlsb_en), .B(clk_5k), .C(r_hlsb_sel), .Y(n47) );
  NAND3X1 U85 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .C(r_vcomp[3]), .Y(n58) );
  INVX1 U86 ( .A(r_vcomp[4]), .Y(n29) );
  INVX1 U87 ( .A(r_vcomp[5]), .Y(n30) );
  NOR21XL U88 ( .B(sdischg_cnt[3]), .A(r_sdischg[3]), .Y(n46) );
  OAI32X1 U89 ( .A(n22), .B(sdischg_cnt[2]), .C(n46), .D(sdischg_cnt[3]), .E(
        n21), .Y(n44) );
  INVX1 U90 ( .A(r_sdischg[3]), .Y(n21) );
  AO222X1 U91 ( .A(n34), .B(n19), .C(n35), .D(n36), .E(sdischg_duty), .F(n37), 
        .Y(n81) );
  AOI22BXL U92 ( .B(N126), .A(n38), .D(r_sdischg[1]), .C(sdischg_cnt[1]), .Y(
        n35) );
  OAI22AX1 U93 ( .D(n36), .C(n43), .A(sdischg_cnt[4]), .B(n20), .Y(n34) );
  EORX1 U94 ( .A(n20), .B(sdischg_cnt[4]), .C(n45), .D(n44), .Y(n36) );
  AOI21X1 U95 ( .B(sdischg_cnt[2]), .C(n22), .A(n46), .Y(n45) );
  AOI21BX1 U96 ( .C(sdischg_cnt[1]), .B(r_sdischg[1]), .A(n44), .Y(n43) );
  OAI221X1 U97 ( .A(n63), .B(n18), .C(n64), .D(n33), .E(r_hlsb_en), .Y(n62) );
  INVX1 U98 ( .A(r_hlsb_freq), .Y(n18) );
  AOI211X1 U99 ( .C(div20_cnt[1]), .D(div20_cnt[0]), .A(div20_cnt[3]), .B(
        div20_cnt[2]), .Y(n64) );
  AOI21X1 U100 ( .B(div20_cnt[0]), .C(div20_cnt[3]), .A(n65), .Y(n63) );
  NOR2X1 U101 ( .A(r_sdischg[6]), .B(r_sdischg[5]), .Y(n37) );
  NAND2X1 U102 ( .A(n33), .B(n68), .Y(n65) );
  OAI21X1 U103 ( .B(div20_cnt[1]), .C(div20_cnt[2]), .A(div20_cnt[3]), .Y(n68)
         );
  INVX1 U104 ( .A(div20_cnt[4]), .Y(n33) );
  INVX1 U105 ( .A(r_sdischg[4]), .Y(n20) );
  NOR2X1 U106 ( .A(n37), .B(sdischg_cnt[0]), .Y(N126) );
  INVX1 U107 ( .A(r_sdischg[2]), .Y(n22) );
  NAND2X1 U108 ( .A(r_sdischg[0]), .B(n19), .Y(n38) );
  NOR2X1 U109 ( .A(n61), .B(n62), .Y(N42) );
  XNOR2XL U110 ( .A(div20_cnt[4]), .B(add_41_carry[4]), .Y(n61) );
  NOR2X1 U111 ( .A(div20_cnt[0]), .B(n62), .Y(N38) );
  NOR2X1 U112 ( .A(n37), .B(n70), .Y(N130) );
  XNOR2XL U113 ( .A(sdischg_cnt[4]), .B(add_81_carry[4]), .Y(n70) );
  OAI21BX1 U114 ( .C(n69), .B(div20_cnt[3]), .A(r_hlsb_freq), .Y(n66) );
  OAI31XL U115 ( .A(div20_cnt[1]), .B(r_hlsb_duty), .C(div20_cnt[0]), .D(
        div20_cnt[2]), .Y(n69) );
  AOI31X1 U116 ( .A(n66), .B(n67), .C(n32), .D(n31), .Y(N29) );
  INVX1 U117 ( .A(r_hlsb_en), .Y(n31) );
  NAND3X1 U118 ( .A(div20_cnt[0]), .B(div20_cnt[3]), .C(r_hlsb_duty), .Y(n67)
         );
  INVX1 U119 ( .A(n65), .Y(n32) );
  NAND42X1 U120 ( .C(sdischg_cnt[0]), .D(sdischg_cnt[1]), .A(n37), .B(n71), 
        .Y(N115) );
  NOR3XL U121 ( .A(sdischg_cnt[2]), .B(sdischg_cnt[4]), .C(sdischg_cnt[3]), 
        .Y(n71) );
endmodule


module cvctl_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module cvctl_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  XOR2X1 U2 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U4 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  XOR2X1 U5 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U6 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  AND2X1 U7 ( .A(carry[10]), .B(A[10]), .Y(carry[11]) );
endmodule


module cvctl_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n11, n12, n13, n14, n15, n16, n17, n18, n19;
  wire   [10:1] carry;

  FAD1X1 U2_7 ( .A(A[7]), .B(n18), .CI(carry[7]), .CO(carry[8]), .SO(DIFF[7])
         );
  FAD1X1 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n14), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n15), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n12), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n16), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n17), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR2X1 U1 ( .A(n1), .B(A[11]), .Y(DIFF[11]) );
  NOR2X1 U2 ( .A(A[10]), .B(carry[10]), .Y(n1) );
  XNOR2XL U3 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2XL U4 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2XL U5 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  INVX1 U6 ( .A(B[2]), .Y(n16) );
  INVX1 U7 ( .A(B[3]), .Y(n12) );
  INVX1 U8 ( .A(B[4]), .Y(n15) );
  INVX1 U9 ( .A(B[5]), .Y(n14) );
  INVX1 U10 ( .A(B[6]), .Y(n11) );
  INVX1 U11 ( .A(B[1]), .Y(n17) );
  NAND21X1 U12 ( .B(n13), .A(n19), .Y(carry[1]) );
  INVX1 U13 ( .A(A[0]), .Y(n19) );
  INVX1 U14 ( .A(B[7]), .Y(n18) );
  INVX1 U15 ( .A(B[0]), .Y(n13) );
  XNOR2XL U16 ( .A(n13), .B(A[0]), .Y(DIFF[0]) );
  OR2X1 U17 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  OR2X1 U18 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_cvctl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_19 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9335;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_19 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9335), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9335), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9335), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9335), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9335), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9335), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9335), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9335), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9335), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_20 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9353;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_20 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9353), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9353), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9353), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9353), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9353), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9353), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9353), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9353), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9353), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_21 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9371;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_21 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9371), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9371), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9371), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9371), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9371), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9371), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9371), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9371), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9371), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_22 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9389;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_22 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9389), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9389), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9389), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9389), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9389), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9389), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9389), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9389), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9389), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_23 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9407;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_23 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9407), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9407), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9407), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9407), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9407), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9407), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9407), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9407), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9407), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_24 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9425;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_24 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9425), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9425), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9425), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9425), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9425), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9425), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9425), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9425), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9425), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcp_a0 ( dp_comp, dm_comp, id_comp, intr, tx_en, tx_dat, r_dat, r_sta, 
        r_ctl, r_msk, r_crc, r_acc, r_dpdmsta, r_wdat, r_wr, r_re, clk, srstz, 
        r_tui, test_si, test_so, test_se );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  output [7:0] r_crc;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input [7:0] r_wdat;
  input [6:0] r_wr;
  output [7:0] r_tui;
  input dp_comp, dm_comp, id_comp, r_re, clk, srstz, test_si, test_se;
  output intr, tx_en, tx_dat, test_so;
  wire   r_dm, r_dmchg, r_acc_int, r_wr_last, r_wr_other, n3, n4, n1;

  INVX1 U3 ( .A(n4), .Y(n3) );
  INVX1 U4 ( .A(srstz), .Y(n4) );
  dpdmacc_a0 u0_dpdmacc ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(
        id_comp), .r_re_0(r_re), .r_wr_1(r_wr[6]), .r_wdat(r_wdat), .r_acc(
        r_acc), .r_dpdmsta(r_dpdmsta), .r_dm(r_dm), .r_dmchg(r_dmchg), .r_int(
        r_acc_int), .clk(clk), .rstz(srstz), .test_si(test_si), .test_se(
        test_se) );
  fcpegn_a0 u0_fcpegn ( .intr(intr), .tx_en(tx_en), .tx_dat(tx_dat), .r_dat(
        r_dat), .r_sta(r_sta), .r_ctl(r_ctl), .r_msk(r_msk), .r_wr(r_wr[4:0]), 
        .r_wdat(r_wdat), .ff_idn(r_dm), .ff_chg(n1), .r_acc_int(r_acc_int), 
        .clk(clk), .srstz(n3), .r_tui(r_tui), .test_si(r_crc[7]), .test_so(
        test_so), .test_se(test_se) );
  fcpcrc_a0 u0_fcpcrc ( .tx_crc(r_crc), .crc_din(r_wdat), .crc_en(r_ctl[2]), 
        .crc_shfi(r_wr_other), .crc_shfl(r_wr_last), .clk(clk), .srstz(n3), 
        .test_si(r_dpdmsta[5]), .test_se(test_se) );
  BUFX3 U1 ( .A(r_dmchg), .Y(n1) );
  AND2X1 U2 ( .A(r_wr[5]), .B(r_ctl[3]), .Y(r_wr_last) );
  NOR21XL U5 ( .B(r_wr[5]), .A(r_ctl[3]), .Y(r_wr_other) );
endmodule


module fcpcrc_a0 ( tx_crc, crc_din, crc_en, crc_shfi, crc_shfl, clk, srstz, 
        test_si, test_se );
  output [7:0] tx_crc;
  input [7:0] crc_din;
  input crc_en, crc_shfi, crc_shfl, clk, srstz, test_si, test_se;
  wire   N81, N82, N83, N84, N85, N86, N87, N88, N89, net9443, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n1;

  SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 clk_gate_crc8_r_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net9443), .TE(test_se) );
  SDFFRQX1 crc8_r_reg_0_ ( .D(N82), .SIN(test_si), .SMC(test_se), .C(net9443), 
        .XR(srstz), .Q(tx_crc[0]) );
  SDFFRQX1 crc8_r_reg_2_ ( .D(N84), .SIN(tx_crc[1]), .SMC(test_se), .C(net9443), .XR(srstz), .Q(tx_crc[2]) );
  SDFFRQX1 crc8_r_reg_4_ ( .D(N86), .SIN(tx_crc[3]), .SMC(test_se), .C(net9443), .XR(srstz), .Q(tx_crc[4]) );
  SDFFRQX1 crc8_r_reg_3_ ( .D(N85), .SIN(tx_crc[2]), .SMC(test_se), .C(net9443), .XR(srstz), .Q(tx_crc[3]) );
  SDFFRQX1 crc8_r_reg_1_ ( .D(N83), .SIN(tx_crc[0]), .SMC(test_se), .C(net9443), .XR(srstz), .Q(tx_crc[1]) );
  SDFFRQX1 crc8_r_reg_6_ ( .D(N88), .SIN(tx_crc[5]), .SMC(test_se), .C(net9443), .XR(srstz), .Q(tx_crc[6]) );
  SDFFRQX1 crc8_r_reg_7_ ( .D(N89), .SIN(tx_crc[6]), .SMC(test_se), .C(net9443), .XR(srstz), .Q(tx_crc[7]) );
  SDFFRQX1 crc8_r_reg_5_ ( .D(N87), .SIN(tx_crc[4]), .SMC(test_se), .C(net9443), .XR(srstz), .Q(tx_crc[5]) );
  XNOR2XL U3 ( .A(n36), .B(n37), .Y(n15) );
  XNOR2XL U4 ( .A(n35), .B(n34), .Y(n19) );
  XNOR2XL U5 ( .A(n8), .B(n1), .Y(n35) );
  XNOR2XL U6 ( .A(n28), .B(n24), .Y(n13) );
  XNOR2XL U7 ( .A(n13), .B(n23), .Y(n8) );
  XNOR2XL U8 ( .A(n2), .B(n9), .Y(n28) );
  OAI22X1 U9 ( .A(n15), .B(n3), .C(n16), .D(n5), .Y(N87) );
  XNOR2XL U10 ( .A(n17), .B(n18), .Y(n16) );
  XNOR2XL U11 ( .A(n6), .B(n15), .Y(n18) );
  XNOR2XL U12 ( .A(n19), .B(n14), .Y(n17) );
  XOR2X1 U13 ( .A(n20), .B(n2), .Y(n23) );
  XNOR2XL U14 ( .A(n27), .B(n26), .Y(n6) );
  XNOR2XL U15 ( .A(n15), .B(n28), .Y(n27) );
  XNOR2XL U16 ( .A(n38), .B(n39), .Y(n20) );
  XNOR2XL U17 ( .A(crc_din[4]), .B(n40), .Y(n39) );
  OAI22X1 U18 ( .A(n20), .B(n3), .C(n21), .D(n5), .Y(N86) );
  XOR2X1 U19 ( .A(n19), .B(n22), .Y(n21) );
  XNOR2XL U20 ( .A(n14), .B(n23), .Y(n22) );
  OAI22X1 U21 ( .A(n2), .B(n3), .C(n4), .D(n5), .Y(N89) );
  XOR2X1 U22 ( .A(n6), .B(n7), .Y(n4) );
  XNOR2XL U23 ( .A(n8), .B(n2), .Y(n7) );
  OAI22X1 U24 ( .A(n9), .B(n3), .C(n10), .D(n5), .Y(N88) );
  XNOR2XL U25 ( .A(n11), .B(n12), .Y(n10) );
  XNOR2XL U26 ( .A(n13), .B(n9), .Y(n12) );
  XNOR2XL U27 ( .A(n14), .B(n6), .Y(n11) );
  OAI22X1 U28 ( .A(n24), .B(n3), .C(n25), .D(n5), .Y(N85) );
  XNOR2XL U29 ( .A(n19), .B(n13), .Y(n25) );
  OAI22X1 U30 ( .A(n34), .B(n3), .C(n19), .D(n5), .Y(N82) );
  XNOR2XL U31 ( .A(n31), .B(n32), .Y(n14) );
  XNOR2XL U32 ( .A(n1), .B(n30), .Y(n32) );
  XNOR2XL U33 ( .A(n23), .B(n9), .Y(n31) );
  XNOR2XL U34 ( .A(n41), .B(n42), .Y(n24) );
  XNOR2XL U35 ( .A(crc_din[3]), .B(n43), .Y(n42) );
  INVX1 U36 ( .A(n15), .Y(n1) );
  XNOR2XL U37 ( .A(crc_din[1]), .B(n33), .Y(n30) );
  OAI22X1 U38 ( .A(n30), .B(n3), .C(n14), .D(n5), .Y(N83) );
  OAI22X1 U39 ( .A(n26), .B(n3), .C(n6), .D(n5), .Y(N84) );
  XNOR2XL U40 ( .A(crc_din[2]), .B(n29), .Y(n26) );
  XNOR2XL U41 ( .A(crc_din[0]), .B(n41), .Y(n34) );
  XOR2X1 U42 ( .A(n41), .B(n33), .Y(n38) );
  XNOR2XL U43 ( .A(n43), .B(n40), .Y(n51) );
  XNOR2XL U44 ( .A(n44), .B(n45), .Y(n9) );
  XNOR2XL U45 ( .A(n33), .B(n43), .Y(n45) );
  XNOR2XL U46 ( .A(n29), .B(n48), .Y(n44) );
  XNOR2XL U47 ( .A(tx_crc[6]), .B(crc_din[6]), .Y(n48) );
  XNOR2XL U48 ( .A(n49), .B(n50), .Y(n2) );
  XOR2X1 U49 ( .A(n51), .B(n29), .Y(n49) );
  XNOR2XL U50 ( .A(tx_crc[7]), .B(crc_din[7]), .Y(n50) );
  XNOR2XL U51 ( .A(n38), .B(n29), .Y(n36) );
  XNOR2XL U52 ( .A(tx_crc[5]), .B(crc_din[5]), .Y(n37) );
  NAND21X1 U53 ( .B(crc_shfl), .A(crc_en), .Y(n3) );
  NAND2X1 U54 ( .A(crc_shfl), .B(crc_en), .Y(n5) );
  OR2X1 U55 ( .A(crc_shfi), .B(n3), .Y(N81) );
  XOR2X1 U56 ( .A(n46), .B(n47), .Y(n33) );
  XOR2X1 U57 ( .A(tx_crc[5]), .B(tx_crc[6]), .Y(n46) );
  XNOR2XL U58 ( .A(tx_crc[1]), .B(n40), .Y(n47) );
  XNOR2XL U59 ( .A(tx_crc[3]), .B(n53), .Y(n43) );
  XNOR2XL U60 ( .A(tx_crc[7]), .B(tx_crc[4]), .Y(n40) );
  XNOR2XL U61 ( .A(n51), .B(n54), .Y(n41) );
  XOR2X1 U62 ( .A(tx_crc[0]), .B(tx_crc[5]), .Y(n54) );
  XOR2X1 U63 ( .A(tx_crc[7]), .B(tx_crc[6]), .Y(n53) );
  XNOR2XL U64 ( .A(n52), .B(n53), .Y(n29) );
  XNOR2XL U65 ( .A(tx_crc[5]), .B(tx_crc[2]), .Y(n52) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcpegn_a0 ( intr, tx_en, tx_dat, r_dat, r_sta, r_ctl, r_msk, r_wr, 
        r_wdat, ff_idn, ff_chg, r_acc_int, clk, srstz, r_tui, test_si, test_so, 
        test_se );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  input [4:0] r_wr;
  input [7:0] r_wdat;
  output [7:0] r_tui;
  input ff_idn, ff_chg, r_acc_int, clk, srstz, test_si, test_se;
  output intr, tx_en, tx_dat, test_so;
  wire   N22, upd_dbuf_en, us_cnt_2_, us_cnt_1_, us_cnt_0_, N85, N87, N88,
         N141, N142, N144, N145, N172, N173, adp_tx_ui_7_, adp_tx_ui_6_, N205,
         N221, N222, N223, N224, N225, N226, N227, N228, N260, N261, N348,
         N349, N356, N362, N363, N444, rx_trans_8_chg, N1005, N1006, N1007,
         N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1043,
         net9465, net9469, net9472, net9473, net9474, net9475, net9476,
         net9477, net9480, net9483, net9488, net9493, net9498, n26, n27, n28,
         n29, n30, n31, n32, n516, n525, n526, N1259, N1258, N1257, N1256,
         N1255, N1254, N1253, N1252, N161, N160, N159, N108, N107, n41, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n461, n464, n4, n83, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n463, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n517, n518, n519, n520, n521, n522,
         n523, n524, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n20, n21, n22, n23, n24, n25, n33, n34, n35, n36, n37, n38, n39,
         n40, n42, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3;
  wire   [6:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;
  wire   [7:0] upd_dbuf;
  wire   [10:0] rxtx_buf;
  wire   [4:1] rx_ui_3_8;
  wire   [4:1] rx_ui_5_8;
  wire   [5:0] catch_sync;
  wire   [7:0] ui_intv_cnt;
  wire   [6:2] symb_cnt;
  wire   [6:0] adp_tx_1_4;
  wire   [7:0] tui_wdat;
  wire   [11:0] trans_buf;
  wire   [1:0] new_rx_sync_cnt;
  wire   [3:0] fcp_state;
  wire   [5:1] add_264_carry;
  wire   [5:1] add_263_carry;
  wire   [8:6] add_274_2_carry;
  wire   [8:6] add_274_carry;

  FAD1X1 add_264_U1_1 ( .A(n69), .B(n73), .CI(add_264_carry[1]), .CO(
        add_264_carry[2]), .SO(rx_ui_5_8[1]) );
  FAD1X1 add_264_U1_2 ( .A(n71), .B(n72), .CI(add_264_carry[2]), .CO(
        add_264_carry[3]), .SO(rx_ui_5_8[2]) );
  FAD1X1 add_264_U1_3 ( .A(n73), .B(n67), .CI(add_264_carry[3]), .CO(
        add_264_carry[4]), .SO(rx_ui_5_8[3]) );
  FAD1X1 add_264_U1_4 ( .A(n72), .B(n68), .CI(add_264_carry[4]), .CO(
        add_264_carry[5]), .SO(rx_ui_5_8[4]) );
  FAD1X1 add_263_U1_1 ( .A(n71), .B(n73), .CI(add_263_carry[1]), .CO(
        add_263_carry[2]), .SO(rx_ui_3_8[1]) );
  FAD1X1 add_263_U1_2 ( .A(n73), .B(n72), .CI(add_263_carry[2]), .CO(
        add_263_carry[3]), .SO(rx_ui_3_8[2]) );
  FAD1X1 add_263_U1_3 ( .A(n72), .B(n67), .CI(add_263_carry[3]), .CO(
        add_263_carry[4]), .SO(rx_ui_3_8[3]) );
  FAD1X1 add_263_U1_4 ( .A(n67), .B(n5), .CI(add_263_carry[4]), .CO(
        add_263_carry[5]), .SO(rx_ui_3_8[4]) );
  FAD1X1 add_274_2_U1_6 ( .A(N160), .B(ui_intv_cnt[6]), .CI(add_274_2_carry[6]), .CO(add_274_2_carry[7]), .SO(N172) );
  FAD1X1 add_274_2_U1_7 ( .A(N161), .B(ui_intv_cnt[7]), .CI(add_274_2_carry[7]), .CO(add_274_2_carry[8]), .SO(N173) );
  FAD1X1 add_274_U1_6 ( .A(N107), .B(ui_intv_cnt[6]), .CI(add_274_carry[6]), 
        .CO(add_274_carry[7]), .SO(N144) );
  FAD1X1 add_274_U1_7 ( .A(N108), .B(ui_intv_cnt[7]), .CI(add_274_carry[7]), 
        .CO(add_274_carry[8]), .SO(N145) );
  INVX1 U23 ( .A(n51), .Y(n46) );
  INVX1 U24 ( .A(n51), .Y(n47) );
  INVX1 U25 ( .A(n51), .Y(n48) );
  INVX1 U26 ( .A(n51), .Y(n49) );
  INVX1 U27 ( .A(n51), .Y(n50) );
  INVX1 U28 ( .A(n51), .Y(n45) );
  INVX1 U29 ( .A(n51), .Y(n43) );
  INVX1 U30 ( .A(n51), .Y(n44) );
  INVX1 U31 ( .A(n51), .Y(n41) );
  INVX1 U32 ( .A(srstz), .Y(n51) );
  MAJ3X1 U619 ( .A(rx_ui_3_8[1]), .B(n447), .C(n117), .Y(n446) );
  glreg_8_00000000 u0_fcpctl ( .clk(clk), .arstz(n46), .we(r_wr[0]), .wdat({
        r_wdat[7:3], n23, r_wdat[1:0]}), .rdat({n464, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, r_ctl[4:0]}), .test_si(r_ctl[7]), .test_se(
        test_se) );
  glsta_a0_0 u0_fcpsta ( .clk(clk), .arstz(n45), .rst0(1'b0), .set2({r_acc_int, 
        setsta[6:5], n536, setsta[3], n525, n4, setsta[0]}), .clr1(clrsta), 
        .rdat(r_sta), .irq(r_irq), .test_si(r_msk[7]), .test_se(test_se) );
  glreg_a0_4 u0_fcpmsk ( .clk(clk), .arstz(n44), .we(r_wr[2]), .wdat({
        r_wdat[7:3], n23, r_wdat[1:0]}), .rdat(r_msk), .test_si(r_dat[7]), 
        .test_se(test_se) );
  glreg_a0_3 u0_fcpdat ( .clk(clk), .arstz(n43), .we(upd_dbuf_en), .wdat(
        upd_dbuf), .rdat(r_dat), .test_si(n464), .test_se(test_se) );
  glreg_a0_2 u0_fcptui ( .clk(clk), .arstz(n41), .we(n83), .wdat(tui_wdat), 
        .rdat(r_tui), .test_si(r_sta[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 clk_gate_catch_sync_reg ( .CLK(clk), .EN(
        n526), .ENCLK(net9465), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 clk_gate_ui_intv_cnt_reg ( .CLK(clk), .EN(
        N205), .ENCLK(net9483), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 clk_gate_rxtx_buf_reg ( .CLK(clk), .EN(N22), 
        .ENCLK(net9488), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 clk_gate_fcp_state_reg ( .CLK(clk), .EN(
        N1005), .ENCLK(net9493), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 clk_gate_symb_cnt_reg ( .CLK(clk), .EN(
        N1043), .ENCLK(net9498), .TE(test_se) );
  fcpegn_a0_DW01_inc_0 r611 ( .A({symb_cnt[6:4], n14, n12, n7, n16}), .SUM({
        n26, n27, n28, n29, n30, n31, n32}) );
  fcpegn_a0_DW01_inc_1 add_283_round ( .A({1'b0, adp_tx_ui_7_, adp_tx_ui_6_, 
        n75, r_tui[4:1]}), .SUM({adp_tx_1_4, SYNOPSYS_UNCONNECTED_3}) );
  fcpegn_a0_DW01_inc_2 add_316_aco ( .A({N1259, N1258, N1257, N1256, N1255, 
        N1254, N1253, N1252}), .SUM({N228, N227, N226, N225, N224, N223, N222, 
        N221}) );
  SDFFRQX1 rxtx_buf_reg_8_ ( .D(trans_buf[8]), .SIN(rxtx_buf[7]), .SMC(test_se), .C(net9488), .XR(n47), .Q(rxtx_buf[8]) );
  SDFFRQX1 rxtx_buf_reg_10_ ( .D(trans_buf[10]), .SIN(rxtx_buf[9]), .SMC(
        test_se), .C(net9488), .XR(n47), .Q(rxtx_buf[10]) );
  SDFFRQX1 rxtx_buf_reg_9_ ( .D(trans_buf[9]), .SIN(rxtx_buf[8]), .SMC(test_se), .C(net9488), .XR(n47), .Q(rxtx_buf[9]) );
  SDFFRQX1 rxtx_buf_reg_0_ ( .D(trans_buf[0]), .SIN(rx_trans_8_chg), .SMC(
        test_se), .C(net9488), .XR(n48), .Q(rxtx_buf[0]) );
  SDFFRQX1 rxtx_buf_reg_4_ ( .D(trans_buf[4]), .SIN(rxtx_buf[3]), .SMC(test_se), .C(net9488), .XR(n47), .Q(rxtx_buf[4]) );
  SDFFRQX1 rxtx_buf_reg_6_ ( .D(trans_buf[6]), .SIN(rxtx_buf[5]), .SMC(test_se), .C(net9488), .XR(n47), .Q(rxtx_buf[6]) );
  SDFFRQX1 rxtx_buf_reg_7_ ( .D(trans_buf[7]), .SIN(rxtx_buf[6]), .SMC(test_se), .C(net9488), .XR(n47), .Q(rxtx_buf[7]) );
  SDFFRQX1 rxtx_buf_reg_3_ ( .D(trans_buf[3]), .SIN(rxtx_buf[2]), .SMC(test_se), .C(net9488), .XR(n48), .Q(rxtx_buf[3]) );
  SDFFRQX1 rxtx_buf_reg_5_ ( .D(trans_buf[5]), .SIN(rxtx_buf[4]), .SMC(test_se), .C(net9488), .XR(n47), .Q(rxtx_buf[5]) );
  SDFFRQX1 rxtx_buf_reg_1_ ( .D(trans_buf[1]), .SIN(rxtx_buf[0]), .SMC(test_se), .C(net9488), .XR(n49), .Q(rxtx_buf[1]) );
  SDFFRQX1 rx_byte_pchk_reg ( .D(N356), .SIN(new_rx_sync_cnt[1]), .SMC(test_se), .C(clk), .XR(n50), .Q(setsta[5]) );
  SDFFRQX1 rxtx_buf_reg_2_ ( .D(trans_buf[2]), .SIN(rxtx_buf[1]), .SMC(test_se), .C(net9488), .XR(n47), .Q(rxtx_buf[2]) );
  SDFFRQX1 new_rx_sync_cnt_reg_1_ ( .D(N349), .SIN(new_rx_sync_cnt[0]), .SMC(
        test_se), .C(clk), .XR(n44), .Q(new_rx_sync_cnt[1]) );
  SDFFRQX1 new_rx_sync_cnt_reg_0_ ( .D(N348), .SIN(fcp_state[3]), .SMC(test_se), .C(clk), .XR(n41), .Q(new_rx_sync_cnt[0]) );
  SDFFQX1 rx_trans_8_chg_reg ( .D(n516), .SIN(setsta[5]), .SMC(test_se), .C(
        clk), .Q(rx_trans_8_chg) );
  SDFFRQX1 us_cnt_reg_3_ ( .D(N88), .SIN(us_cnt_2_), .SMC(test_se), .C(clk), 
        .XR(n43), .Q(test_so) );
  SDFFRQX1 us_cnt_reg_2_ ( .D(N87), .SIN(us_cnt_1_), .SMC(test_se), .C(clk), 
        .XR(n45), .Q(us_cnt_2_) );
  SDFFRQX1 us_cnt_reg_1_ ( .D(n461), .SIN(us_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(srstz), .Q(us_cnt_1_) );
  SDFFRQX1 us_cnt_reg_0_ ( .D(N85), .SIN(ui_intv_cnt[7]), .SMC(test_se), .C(
        clk), .XR(n47), .Q(us_cnt_0_) );
  SDFFRQX1 ui_intv_cnt_reg_6_ ( .D(net9472), .SIN(n11), .SMC(test_se), .C(
        net9483), .XR(n49), .Q(ui_intv_cnt[6]) );
  SDFFRQX1 ui_intv_cnt_reg_7_ ( .D(net9469), .SIN(ui_intv_cnt[6]), .SMC(
        test_se), .C(net9483), .XR(n49), .Q(ui_intv_cnt[7]) );
  SDFFRQX1 ui_intv_cnt_reg_4_ ( .D(net9474), .SIN(N141), .SMC(test_se), .C(
        net9483), .XR(n49), .Q(N142) );
  SDFFRQX1 ui_intv_cnt_reg_1_ ( .D(net9477), .SIN(ui_intv_cnt[0]), .SMC(
        test_se), .C(net9483), .XR(n48), .Q(ui_intv_cnt[1]) );
  SDFFRQX1 ui_intv_cnt_reg_3_ ( .D(net9475), .SIN(ui_intv_cnt[2]), .SMC(
        test_se), .C(net9483), .XR(n48), .Q(N141) );
  SDFFRQX1 ui_intv_cnt_reg_0_ ( .D(net9480), .SIN(r_tui[7]), .SMC(test_se), 
        .C(net9483), .XR(n48), .Q(ui_intv_cnt[0]) );
  SDFFRQX1 ui_intv_cnt_reg_2_ ( .D(net9476), .SIN(ui_intv_cnt[1]), .SMC(
        test_se), .C(net9483), .XR(n48), .Q(ui_intv_cnt[2]) );
  SDFFRQX1 ui_intv_cnt_reg_5_ ( .D(net9473), .SIN(n3), .SMC(test_se), .C(
        net9483), .XR(n49), .Q(ui_intv_cnt[5]) );
  SDFFSQX1 catch_sync_reg_5_ ( .D(n11), .SIN(catch_sync[4]), .SMC(test_se), 
        .C(net9465), .XS(n46), .Q(catch_sync[5]) );
  SDFFRQX1 catch_sync_reg_4_ ( .D(n3), .SIN(catch_sync[3]), .SMC(test_se), .C(
        net9465), .XR(n48), .Q(catch_sync[4]) );
  SDFFRQX1 sync_length_reg_1_ ( .D(N261), .SIN(N362), .SMC(test_se), .C(
        net9483), .XR(n49), .Q(N363) );
  SDFFRQX1 symb_cnt_reg_4_ ( .D(N1014), .SIN(n14), .SMC(test_se), .C(net9498), 
        .XR(n50), .Q(symb_cnt[4]) );
  SDFFRQX1 symb_cnt_reg_5_ ( .D(N1015), .SIN(symb_cnt[4]), .SMC(test_se), .C(
        net9498), .XR(n50), .Q(symb_cnt[5]) );
  SDFFRQX1 symb_cnt_reg_6_ ( .D(N1016), .SIN(symb_cnt[5]), .SMC(test_se), .C(
        net9498), .XR(n49), .Q(symb_cnt[6]) );
  SDFFRQX1 sync_length_reg_0_ ( .D(N260), .SIN(symb_cnt[6]), .SMC(test_se), 
        .C(net9483), .XR(n49), .Q(N362) );
  SDFFRQX1 symb_cnt_reg_3_ ( .D(N1013), .SIN(n12), .SMC(test_se), .C(net9498), 
        .XR(n50), .Q(symb_cnt[3]) );
  SDFFSQX1 catch_sync_reg_3_ ( .D(N141), .SIN(catch_sync[2]), .SMC(test_se), 
        .C(net9465), .XS(n46), .Q(catch_sync[3]) );
  SDFFRQX1 symb_cnt_reg_1_ ( .D(N1011), .SIN(n16), .SMC(test_se), .C(net9498), 
        .XR(n50), .Q(N160) );
  SDFFRQX1 symb_cnt_reg_2_ ( .D(N1012), .SIN(n7), .SMC(test_se), .C(net9498), 
        .XR(n50), .Q(symb_cnt[2]) );
  SDFFRQX1 symb_cnt_reg_0_ ( .D(N1010), .SIN(tx_dat), .SMC(test_se), .C(
        net9498), .XR(n50), .Q(N159) );
  SDFFRQX1 catch_sync_reg_1_ ( .D(ui_intv_cnt[1]), .SIN(catch_sync[0]), .SMC(
        test_se), .C(net9465), .XR(n48), .Q(catch_sync[1]) );
  SDFFRQX1 catch_sync_reg_2_ ( .D(ui_intv_cnt[2]), .SIN(catch_sync[1]), .SMC(
        test_se), .C(net9465), .XR(n48), .Q(catch_sync[2]) );
  SDFFRQX1 catch_sync_reg_0_ ( .D(ui_intv_cnt[0]), .SIN(test_si), .SMC(test_se), .C(net9465), .XR(n48), .Q(catch_sync[0]) );
  SDFFRQX1 rxtx_buf_reg_11_ ( .D(trans_buf[11]), .SIN(rxtx_buf[10]), .SMC(
        test_se), .C(net9488), .XR(n49), .Q(tx_dat) );
  SDFFSQX1 tx_dbuf_keep_empty_reg ( .D(N444), .SIN(N363), .SMC(test_se), .C(
        clk), .XS(n47), .Q(r_ctl[7]) );
  SDFFRQX1 fcp_state_reg_3_ ( .D(N1009), .SIN(fcp_state[2]), .SMC(test_se), 
        .C(net9493), .XR(n49), .Q(fcp_state[3]) );
  SDFFRQX1 fcp_state_reg_0_ ( .D(N1006), .SIN(catch_sync[5]), .SMC(test_se), 
        .C(net9493), .XR(n50), .Q(fcp_state[0]) );
  SDFFRQX1 fcp_state_reg_1_ ( .D(N1007), .SIN(fcp_state[0]), .SMC(test_se), 
        .C(net9493), .XR(n50), .Q(fcp_state[1]) );
  SDFFRQX1 fcp_state_reg_2_ ( .D(N1008), .SIN(fcp_state[1]), .SMC(test_se), 
        .C(net9493), .XR(n50), .Q(fcp_state[2]) );
  BUFX3 U4 ( .A(n270), .Y(n2) );
  BUFX3 U5 ( .A(N142), .Y(n3) );
  INVX1 U6 ( .A(n333), .Y(n5) );
  INVX1 U7 ( .A(n122), .Y(n6) );
  INVX1 U8 ( .A(n131), .Y(n7) );
  INVX1 U9 ( .A(ff_idn), .Y(n8) );
  INVX1 U10 ( .A(n100), .Y(n9) );
  INVX1 U11 ( .A(n58), .Y(n10) );
  INVX1 U12 ( .A(n123), .Y(n11) );
  INVX1 U13 ( .A(n128), .Y(n12) );
  INVX1 U14 ( .A(r_ctl[0]), .Y(n13) );
  INVX1 U15 ( .A(n126), .Y(n14) );
  INVX1 U16 ( .A(r_wr[3]), .Y(n15) );
  BUFX3 U17 ( .A(N159), .Y(n16) );
  INVX1 U18 ( .A(N141), .Y(n17) );
  XNOR2XL U19 ( .A(n186), .B(n187), .Y(n157) );
  XNOR2XL U20 ( .A(n184), .B(n185), .Y(n159) );
  INVX1 U21 ( .A(n24), .Y(n23) );
  INVX1 U22 ( .A(n295), .Y(n542) );
  INVX1 U33 ( .A(r_wr[3]), .Y(n80) );
  INVX1 U34 ( .A(r_wr[4]), .Y(n81) );
  NOR2X1 U35 ( .A(n34), .B(n78), .Y(clrsta[5]) );
  NOR2X1 U36 ( .A(n22), .B(n78), .Y(clrsta[1]) );
  NOR2X1 U37 ( .A(n33), .B(n78), .Y(clrsta[4]) );
  NOR2X1 U38 ( .A(n21), .B(n78), .Y(clrsta[0]) );
  INVX1 U39 ( .A(r_wdat[7]), .Y(n36) );
  INVX1 U40 ( .A(r_wdat[6]), .Y(n35) );
  INVX1 U41 ( .A(r_wdat[4]), .Y(n33) );
  INVX1 U42 ( .A(r_wdat[3]), .Y(n25) );
  INVX1 U43 ( .A(r_wdat[5]), .Y(n34) );
  NOR2X1 U44 ( .A(n35), .B(n78), .Y(clrsta[6]) );
  NOR2X1 U45 ( .A(n24), .B(n78), .Y(clrsta[2]) );
  NOR2X1 U46 ( .A(n36), .B(n78), .Y(clrsta[7]) );
  NOR2X1 U47 ( .A(n25), .B(n78), .Y(clrsta[3]) );
  INVX1 U48 ( .A(r_wdat[2]), .Y(n24) );
  INVX1 U49 ( .A(r_wdat[1]), .Y(n22) );
  INVX1 U50 ( .A(r_wdat[0]), .Y(n21) );
  NOR2X1 U51 ( .A(n542), .B(n541), .Y(n264) );
  NOR2X1 U52 ( .A(n549), .B(n543), .Y(n295) );
  INVX1 U53 ( .A(n269), .Y(n79) );
  INVX1 U54 ( .A(n257), .Y(n42) );
  INVX1 U55 ( .A(r_wr[1]), .Y(n78) );
  OAI221X1 U56 ( .A(n155), .B(n104), .C(n33), .D(n81), .E(n158), .Y(
        tui_wdat[4]) );
  OAI221X1 U57 ( .A(n103), .B(n155), .C(n34), .D(n81), .E(n158), .Y(
        tui_wdat[5]) );
  OAI221X1 U58 ( .A(n105), .B(n155), .C(n25), .D(n81), .E(n158), .Y(
        tui_wdat[3]) );
  INVX1 U59 ( .A(n159), .Y(n105) );
  INVX1 U60 ( .A(n167), .Y(n101) );
  INVX1 U61 ( .A(n157), .Y(n103) );
  INVX1 U62 ( .A(n173), .Y(n104) );
  INVX1 U63 ( .A(n316), .Y(n66) );
  NAND2X1 U64 ( .A(n159), .B(n160), .Y(n179) );
  INVX1 U65 ( .A(n505), .Y(n113) );
  INVX1 U66 ( .A(n348), .Y(n549) );
  INVX1 U67 ( .A(n377), .Y(n543) );
  INVX1 U68 ( .A(n420), .Y(n541) );
  NOR2X1 U69 ( .A(n293), .B(n80), .Y(n269) );
  INVX1 U70 ( .A(n256), .Y(n52) );
  NAND2X1 U71 ( .A(n253), .B(n58), .Y(n257) );
  INVX1 U72 ( .A(n249), .Y(n58) );
  NAND31X1 U73 ( .C(n162), .A(n81), .B(n154), .Y(n155) );
  OAI222XL U74 ( .A(r_wr[4]), .B(n154), .C(n155), .D(n156), .E(n35), .F(n81), 
        .Y(tui_wdat[6]) );
  XNOR2XL U75 ( .A(n101), .B(n157), .Y(n156) );
  OAI2B11X1 U76 ( .D(N221), .C(n90), .A(n278), .B(n38), .Y(net9480) );
  NAND2X1 U77 ( .A(n162), .B(n81), .Y(n158) );
  OAI2B11X1 U78 ( .D(n160), .C(n155), .A(n158), .B(n161), .Y(tui_wdat[2]) );
  EORX1 U79 ( .A(r_wr[4]), .B(n23), .C(n154), .D(r_wr[4]), .Y(n161) );
  ENOX1 U80 ( .A(n280), .B(n278), .C(N225), .D(n279), .Y(net9474) );
  ENOX1 U81 ( .A(n280), .B(n278), .C(N227), .D(n279), .Y(net9472) );
  INVX1 U82 ( .A(n280), .Y(n38) );
  XNOR2XL U83 ( .A(n36), .B(n54), .Y(n342) );
  AND2X1 U84 ( .A(N224), .B(n279), .Y(net9475) );
  AND2X1 U85 ( .A(N226), .B(n279), .Y(net9473) );
  AND2X1 U86 ( .A(N223), .B(n279), .Y(net9476) );
  AND2X1 U87 ( .A(N222), .B(n279), .Y(net9477) );
  NAND3X1 U88 ( .A(n278), .B(n90), .C(n38), .Y(N205) );
  XNOR2XL U89 ( .A(n68), .B(add_263_carry[5]), .Y(n449) );
  XNOR2XL U90 ( .A(n177), .B(n176), .Y(n167) );
  AOI21X1 U91 ( .B(n176), .C(n177), .A(n175), .Y(n169) );
  OAI21BBX1 U92 ( .A(n216), .B(n233), .C(n239), .Y(n231) );
  OAI21X1 U93 ( .B(n216), .C(n233), .A(n235), .Y(n239) );
  NOR32XL U94 ( .B(n186), .C(n181), .A(n180), .Y(n177) );
  NOR21XL U95 ( .B(n181), .A(n180), .Y(n187) );
  XNOR2XL U96 ( .A(n180), .B(n181), .Y(n173) );
  XNOR2XL U97 ( .A(n233), .B(n234), .Y(n196) );
  XOR2X1 U98 ( .A(n235), .B(n216), .Y(n234) );
  NOR2X1 U99 ( .A(n132), .B(n114), .Y(n505) );
  AOI211X1 U100 ( .C(n111), .D(n309), .A(n245), .B(n307), .Y(n308) );
  NAND2X1 U101 ( .A(n132), .B(n130), .Y(N107) );
  INVX1 U102 ( .A(n418), .Y(n130) );
  INVX1 U103 ( .A(n339), .Y(n70) );
  NOR21XL U104 ( .B(n183), .A(n182), .Y(n185) );
  NAND32X1 U105 ( .B(n184), .C(n182), .A(n183), .Y(n180) );
  XNOR2XL U106 ( .A(n341), .B(n68), .Y(n316) );
  NAND2X1 U107 ( .A(n72), .B(n67), .Y(n341) );
  XNOR2XL U108 ( .A(n72), .B(n67), .Y(n318) );
  NOR2X1 U109 ( .A(n545), .B(n245), .Y(n393) );
  INVX1 U110 ( .A(n307), .Y(n37) );
  XNOR2XL U111 ( .A(n182), .B(n183), .Y(n160) );
  OAI21X1 U112 ( .B(n72), .C(n67), .A(n68), .Y(n321) );
  NOR2X1 U113 ( .A(n491), .B(n54), .Y(n427) );
  AOI32X1 U114 ( .A(n545), .B(n112), .C(n492), .D(n283), .E(n548), .Y(n491) );
  NAND2X1 U115 ( .A(n67), .B(add_264_carry[5]), .Y(n142) );
  INVX1 U116 ( .A(n309), .Y(n109) );
  INVX1 U117 ( .A(n509), .Y(n55) );
  INVX1 U118 ( .A(n492), .Y(n111) );
  INVX1 U119 ( .A(n486), .Y(n57) );
  NOR4XL U120 ( .A(n283), .B(n284), .C(n40), .D(n54), .Y(n525) );
  NAND2X1 U121 ( .A(n285), .B(n548), .Y(n284) );
  OAI211X1 U122 ( .C(n549), .D(n113), .A(n110), .B(n542), .Y(N1043) );
  INVX1 U123 ( .A(n293), .Y(n546) );
  BUFX3 U124 ( .A(ff_idn), .Y(r_ctl[5]) );
  NAND2X1 U125 ( .A(n493), .B(n544), .Y(n377) );
  NOR2X1 U126 ( .A(n550), .B(n352), .Y(n420) );
  NAND2X1 U127 ( .A(n535), .B(n551), .Y(n348) );
  NOR2X1 U128 ( .A(n533), .B(n551), .Y(n493) );
  INVX1 U129 ( .A(n376), .Y(n550) );
  XNOR2XL U130 ( .A(n265), .B(n266), .Y(n261) );
  XNOR2XL U131 ( .A(n271), .B(n272), .Y(n265) );
  XNOR2XL U132 ( .A(n267), .B(n268), .Y(n266) );
  XNOR2XL U133 ( .A(n252), .B(n251), .Y(n271) );
  XNOR2XL U134 ( .A(n263), .B(n255), .Y(n267) );
  XNOR2XL U135 ( .A(n250), .B(n248), .Y(n272) );
  XNOR2XL U136 ( .A(n258), .B(n254), .Y(n268) );
  OAI21X1 U137 ( .B(n85), .C(n58), .A(n259), .Y(trans_buf[1]) );
  AOI32X1 U138 ( .A(n42), .B(n260), .C(n261), .D(n52), .E(n61), .Y(n259) );
  OAI211X1 U139 ( .C(n2), .D(n342), .A(n58), .B(n343), .Y(n256) );
  AOI21X1 U140 ( .B(n344), .C(n79), .A(n77), .Y(n343) );
  NOR2X1 U141 ( .A(n269), .B(n270), .Y(n249) );
  AO33X1 U142 ( .A(n249), .B(n264), .C(ff_idn), .D(n261), .E(n260), .F(n52), 
        .Y(trans_buf[0]) );
  AOI22X1 U143 ( .A(n52), .B(n263), .C(n59), .D(n253), .Y(n247) );
  NOR2X1 U144 ( .A(n77), .B(n52), .Y(n253) );
  OAI222XL U145 ( .A(n255), .B(n256), .C(n254), .D(n257), .E(n86), .F(n58), 
        .Y(trans_buf[3]) );
  OAI222XL U146 ( .A(n254), .B(n256), .C(n258), .D(n257), .E(n82), .F(n58), 
        .Y(trans_buf[2]) );
  INVX1 U147 ( .A(n495), .Y(n39) );
  NOR32XL U148 ( .B(n281), .C(n278), .A(n280), .Y(n279) );
  OAI2B11X1 U149 ( .D(n264), .C(n40), .A(n79), .B(n346), .Y(n280) );
  INVX1 U150 ( .A(n243), .Y(n83) );
  AOI31X1 U151 ( .A(ff_chg), .B(n244), .C(n245), .D(r_wr[4]), .Y(n243) );
  OAI22X1 U152 ( .A(n36), .B(n81), .C(r_wr[4]), .D(n74), .Y(tui_wdat[7]) );
  OAI22X1 U153 ( .A(n21), .B(n81), .C(n166), .D(n155), .Y(tui_wdat[0]) );
  XNOR2XL U154 ( .A(n125), .B(n17), .Y(n166) );
  OAI22X1 U155 ( .A(n100), .B(n58), .C(n345), .D(n13), .Y(N260) );
  EORX1 U156 ( .A(n2), .B(n344), .C(n342), .D(n79), .Y(n345) );
  INVX1 U157 ( .A(n263), .Y(n59) );
  INVX1 U158 ( .A(n258), .Y(n61) );
  INVX1 U159 ( .A(n255), .Y(n60) );
  OAI22X1 U160 ( .A(r_wr[3]), .B(n85), .C(n80), .D(n21), .Y(upd_dbuf[0]) );
  OAI22X1 U161 ( .A(r_wr[3]), .B(n82), .C(n80), .D(n22), .Y(upd_dbuf[1]) );
  OAI22X1 U162 ( .A(r_wr[3]), .B(n86), .C(n80), .D(n24), .Y(upd_dbuf[2]) );
  AND2X1 U163 ( .A(N228), .B(n279), .Y(net9469) );
  NOR2X1 U164 ( .A(n383), .B(n121), .Y(N1259) );
  OAI211X1 U165 ( .C(n110), .D(n305), .A(n10), .B(n346), .Y(N22) );
  OAI21X1 U166 ( .B(n133), .C(n134), .A(n15), .Y(upd_dbuf_en) );
  NAND4X1 U167 ( .A(n146), .B(n147), .C(n148), .D(n149), .Y(n133) );
  NAND4X1 U168 ( .A(n135), .B(n136), .C(n137), .D(n138), .Y(n134) );
  NOR3XL U169 ( .A(n150), .B(n151), .C(n90), .Y(n149) );
  AOI21X1 U170 ( .B(n538), .C(n277), .A(r_wr[3]), .Y(N444) );
  INVX1 U171 ( .A(n334), .Y(n72) );
  INVX1 U172 ( .A(n153), .Y(n67) );
  AOI31X1 U173 ( .A(n543), .B(n126), .C(n276), .D(n408), .Y(n406) );
  INVX1 U174 ( .A(n330), .Y(n73) );
  INVX1 U175 ( .A(n291), .Y(n71) );
  OAI221X1 U176 ( .A(n56), .B(n423), .C(n424), .D(n54), .E(n425), .Y(n408) );
  AOI221XL U177 ( .A(n415), .B(n541), .C(n543), .D(n405), .E(n549), .Y(n423)
         );
  AOI221XL U178 ( .A(n473), .B(n474), .C(n421), .D(n419), .E(n475), .Y(n424)
         );
  AOI31X1 U179 ( .A(n296), .B(n541), .C(n98), .D(n426), .Y(n425) );
  OAI31XL U180 ( .A(n151), .B(n422), .C(n409), .D(n53), .Y(n426) );
  INVX1 U181 ( .A(n427), .Y(n53) );
  NOR2X1 U182 ( .A(n340), .B(n291), .Y(add_263_carry[1]) );
  AOI22X1 U183 ( .A(rx_ui_3_8[3]), .B(n124), .C(rx_ui_3_8[2]), .D(n122), .Y(
        n443) );
  ENOX1 U184 ( .A(n406), .B(n119), .C(n27), .D(n407), .Y(N1015) );
  ENOX1 U185 ( .A(n406), .B(n116), .C(n28), .D(n407), .Y(N1014) );
  ENOX1 U186 ( .A(n406), .B(n128), .C(n30), .D(n407), .Y(N1012) );
  ENOX1 U187 ( .A(n406), .B(n131), .C(n31), .D(n407), .Y(N1011) );
  INVX1 U188 ( .A(n445), .Y(n63) );
  NOR32XL U189 ( .B(n204), .C(n205), .A(n208), .Y(n213) );
  NAND31X1 U190 ( .C(n172), .A(n171), .B(n174), .Y(n162) );
  AOI33X1 U191 ( .A(n175), .B(n176), .C(n177), .D(n101), .E(n102), .F(n178), 
        .Y(n174) );
  AOI22X1 U192 ( .A(n157), .B(n179), .C(n104), .D(n157), .Y(n178) );
  INVX1 U193 ( .A(n169), .Y(n102) );
  XNOR2XL U194 ( .A(n218), .B(n238), .Y(n204) );
  XNOR2XL U195 ( .A(n231), .B(n232), .Y(n238) );
  OAI22X1 U196 ( .A(n206), .B(n20), .C(n106), .D(n207), .Y(n175) );
  AOI21X1 U197 ( .B(n203), .C(n202), .A(n210), .Y(n206) );
  XNOR2XL U198 ( .A(n208), .B(n209), .Y(n207) );
  NAND2X1 U199 ( .A(n205), .B(n204), .Y(n209) );
  OAI211X1 U200 ( .C(n409), .D(n305), .A(n410), .B(n411), .Y(n407) );
  AOI31X1 U201 ( .A(ff_idn), .B(n419), .C(n89), .D(n363), .Y(n410) );
  AOI22AXL U202 ( .A(n412), .B(n413), .D(n414), .C(n56), .Y(n411) );
  INVX1 U203 ( .A(n421), .Y(n89) );
  OAI211X1 U204 ( .C(n167), .D(n168), .A(n169), .B(n170), .Y(n154) );
  OAI31XL U205 ( .A(n173), .B(n159), .C(n160), .D(n103), .Y(n168) );
  NOR21XL U206 ( .B(n171), .A(n172), .Y(n170) );
  OAI21X1 U207 ( .B(n232), .C(n237), .A(n240), .Y(n233) );
  OAI21BBX1 U208 ( .A(n237), .B(n232), .C(N107), .Y(n240) );
  OAI22X1 U209 ( .A(n106), .B(n200), .C(n20), .D(n201), .Y(n176) );
  XNOR2XL U210 ( .A(n202), .B(n203), .Y(n201) );
  XNOR2XL U211 ( .A(n204), .B(n205), .Y(n200) );
  NAND2X1 U212 ( .A(n129), .B(n404), .Y(n235) );
  INVX1 U213 ( .A(n375), .Y(n132) );
  NAND2X1 U214 ( .A(n235), .B(n537), .Y(n237) );
  INVX1 U215 ( .A(n405), .Y(n129) );
  NOR32XL U216 ( .B(add_274_carry[8]), .C(n193), .A(n196), .Y(n205) );
  NOR21XL U217 ( .B(n231), .A(n232), .Y(n215) );
  XNOR2XL U218 ( .A(N107), .B(n236), .Y(n193) );
  XNOR2XL U219 ( .A(n232), .B(n237), .Y(n236) );
  OAI21X1 U220 ( .B(n241), .C(n116), .A(n230), .Y(n216) );
  INVX1 U221 ( .A(n333), .Y(n68) );
  NOR2X1 U222 ( .A(n504), .B(n505), .Y(n492) );
  NOR2X1 U223 ( .A(n131), .B(n537), .Y(n418) );
  OAI22X1 U224 ( .A(n106), .B(n190), .C(n20), .D(n191), .Y(n181) );
  XNOR2XL U225 ( .A(add_274_2_carry[8]), .B(n192), .Y(n191) );
  XNOR2XL U226 ( .A(add_274_carry[8]), .B(n193), .Y(n190) );
  NOR2X1 U227 ( .A(n107), .B(n71), .Y(n339) );
  OAI22X1 U228 ( .A(n20), .B(n194), .C(n106), .D(n195), .Y(n186) );
  XNOR2XL U229 ( .A(n198), .B(n199), .Y(n194) );
  XNOR2XL U230 ( .A(n196), .B(n197), .Y(n195) );
  NAND2X1 U231 ( .A(add_274_2_carry[8]), .B(n192), .Y(n199) );
  NAND2X1 U232 ( .A(n382), .B(n100), .Y(n372) );
  OAI21X1 U233 ( .B(n126), .C(n372), .A(n380), .Y(n369) );
  AOI21X1 U234 ( .B(n117), .C(n69), .A(add_263_carry[1]), .Y(n327) );
  INVX1 U235 ( .A(n340), .Y(n69) );
  INVX1 U236 ( .A(n380), .Y(n115) );
  NAND2X1 U237 ( .A(n241), .B(n116), .Y(n230) );
  NAND2X1 U238 ( .A(n119), .B(n116), .Y(n274) );
  OAI221X1 U239 ( .A(n275), .B(n112), .C(n40), .D(n293), .E(n310), .Y(n307) );
  NAND4X1 U240 ( .A(n311), .B(n121), .C(n312), .D(n313), .Y(n310) );
  AOI32X1 U241 ( .A(n319), .B(n120), .C(n320), .D(n151), .E(n282), .Y(n312) );
  NOR3XL U242 ( .A(n309), .B(n314), .C(n40), .Y(n313) );
  INVX1 U243 ( .A(n518), .Y(n114) );
  NAND2X1 U244 ( .A(add_274_carry[8]), .B(n193), .Y(n197) );
  NAND2X1 U245 ( .A(n382), .B(n130), .Y(n373) );
  NOR2X1 U246 ( .A(n115), .B(n360), .Y(n351) );
  INVX1 U247 ( .A(n347), .Y(n95) );
  OAI31XL U248 ( .A(n348), .B(n96), .C(n349), .D(n350), .Y(n347) );
  AOI33X1 U249 ( .A(n351), .B(n352), .C(n353), .D(n354), .E(n355), .F(n99), 
        .Y(n350) );
  INVX1 U250 ( .A(n356), .Y(n99) );
  NOR32XL U251 ( .B(n494), .C(n552), .A(n551), .Y(n245) );
  NOR32XL U252 ( .B(add_274_2_carry[8]), .C(n192), .A(n198), .Y(n203) );
  XNOR2XL U253 ( .A(n225), .B(n126), .Y(n202) );
  XNOR2XL U254 ( .A(n20), .B(n189), .Y(n164) );
  AOI21X1 U255 ( .B(n537), .C(n123), .A(add_274_2_carry[6]), .Y(n189) );
  XNOR2XL U256 ( .A(adp_tx_1_4[5]), .B(n123), .Y(n469) );
  NOR2X1 U257 ( .A(n383), .B(n122), .Y(N1254) );
  NOR2X1 U258 ( .A(n383), .B(n17), .Y(N1255) );
  NOR2X1 U259 ( .A(n383), .B(n125), .Y(N1256) );
  NOR2X1 U260 ( .A(n383), .B(n123), .Y(N1257) );
  NOR2X1 U261 ( .A(n383), .B(n117), .Y(N1253) );
  XNOR2XL U262 ( .A(adp_tx_1_4[6]), .B(n120), .Y(n470) );
  XNOR2XL U263 ( .A(adp_tx_1_4[4]), .B(n125), .Y(n468) );
  XNOR2XL U264 ( .A(adp_tx_1_4[3]), .B(n124), .Y(n467) );
  AOI22X1 U265 ( .A(N172), .B(n106), .C(N144), .D(n20), .Y(n182) );
  NOR2X1 U266 ( .A(n383), .B(n120), .Y(N1258) );
  XNOR2XL U267 ( .A(n120), .B(adp_tx_ui_6_), .Y(n528) );
  NOR3XL U268 ( .A(n538), .B(n95), .C(n276), .Y(setsta[0]) );
  NAND3X1 U269 ( .A(n552), .B(n551), .C(n494), .Y(n293) );
  INVX1 U270 ( .A(n151), .Y(n545) );
  NOR2X1 U271 ( .A(n383), .B(n107), .Y(N1252) );
  NOR3XL U272 ( .A(n124), .B(n125), .C(n164), .Y(n183) );
  AND2X1 U273 ( .A(n230), .B(n119), .Y(n218) );
  AOI22X1 U274 ( .A(N173), .B(n106), .C(N145), .D(n20), .Y(n184) );
  INVX1 U275 ( .A(n277), .Y(n4) );
  AOI221XL U276 ( .A(n72), .B(n545), .C(n393), .D(n75), .E(n245), .Y(n396) );
  NOR31X1 U277 ( .C(n357), .A(n358), .B(n359), .Y(n353) );
  INVX1 U278 ( .A(n504), .Y(n110) );
  NOR2X1 U279 ( .A(n537), .B(n123), .Y(add_274_2_carry[6]) );
  NOR2X1 U280 ( .A(n100), .B(n537), .Y(n358) );
  NAND2X1 U281 ( .A(n376), .B(n377), .Y(n354) );
  NOR2X1 U282 ( .A(n291), .B(n144), .Y(add_264_carry[1]) );
  XNOR2XL U283 ( .A(n220), .B(n127), .Y(n198) );
  XNOR2XL U284 ( .A(n116), .B(n128), .Y(n220) );
  NOR21XL U285 ( .B(n459), .A(n460), .Y(n454) );
  XNOR2XL U286 ( .A(n124), .B(n73), .Y(n460) );
  XNOR2XL U287 ( .A(n120), .B(n68), .Y(n141) );
  XNOR2XL U288 ( .A(n145), .B(n121), .Y(n135) );
  NAND21X1 U289 ( .B(n142), .A(n68), .Y(n145) );
  XNOR2XL U290 ( .A(n125), .B(n72), .Y(n458) );
  XNOR2XL U291 ( .A(adp_tx_1_4[1]), .B(n117), .Y(n471) );
  XNOR2XL U292 ( .A(adp_tx_ui_7_), .B(n121), .Y(n530) );
  XNOR2XL U293 ( .A(n123), .B(n75), .Y(n529) );
  NOR2X1 U294 ( .A(n305), .B(n150), .Y(n536) );
  NAND2X1 U295 ( .A(n366), .B(n131), .Y(n309) );
  NAND4X1 U296 ( .A(n122), .B(n123), .C(n17), .D(n480), .Y(n421) );
  NOR2X1 U297 ( .A(n120), .B(n478), .Y(n480) );
  NAND2X1 U298 ( .A(n56), .B(n349), .Y(n509) );
  NOR3XL U299 ( .A(n333), .B(n153), .C(n334), .Y(n315) );
  ENOX1 U300 ( .A(n153), .B(n151), .C(adp_tx_ui_6_), .D(n393), .Y(n401) );
  NOR3XL U301 ( .A(n415), .B(n420), .C(n296), .Y(n363) );
  INVX1 U302 ( .A(n20), .Y(n106) );
  INVX1 U303 ( .A(n276), .Y(n56) );
  NOR3XL U304 ( .A(n282), .B(n476), .C(n413), .Y(n475) );
  NAND2X1 U305 ( .A(n422), .B(n545), .Y(n305) );
  NOR2X1 U306 ( .A(n355), .B(n276), .Y(n487) );
  NAND2X1 U307 ( .A(n334), .B(n17), .Y(n328) );
  NOR2X1 U308 ( .A(n139), .B(n140), .Y(n137) );
  XNOR2XL U309 ( .A(rx_ui_5_8[3]), .B(n17), .Y(n139) );
  XNOR2XL U310 ( .A(n141), .B(n142), .Y(n140) );
  INVX1 U311 ( .A(n281), .Y(n90) );
  NAND2X1 U312 ( .A(n116), .B(n217), .Y(n210) );
  INVX1 U313 ( .A(n227), .Y(n127) );
  INVX1 U314 ( .A(n428), .Y(n112) );
  INVX1 U315 ( .A(n415), .Y(n98) );
  INVX1 U316 ( .A(ff_chg), .Y(n40) );
  XNOR2XL U317 ( .A(adp_tx_1_4[0]), .B(n107), .Y(n472) );
  XNOR2XL U318 ( .A(n117), .B(n69), .Y(n456) );
  NOR4XL U319 ( .A(n130), .B(n110), .C(n276), .D(n128), .Y(n486) );
  AND2X1 U320 ( .A(n534), .B(n115), .Y(n283) );
  NAND4X1 U321 ( .A(n404), .B(n126), .C(n119), .D(n118), .Y(n534) );
  OAI22X1 U322 ( .A(n479), .B(n283), .C(n473), .D(n539), .Y(n419) );
  INVX1 U323 ( .A(n479), .Y(n548) );
  INVX1 U324 ( .A(n217), .Y(n108) );
  NOR21XL U325 ( .B(n496), .A(n497), .Y(n488) );
  OAI21X1 U326 ( .B(n126), .C(n128), .A(n380), .Y(n285) );
  INVX1 U327 ( .A(ff_idn), .Y(n54) );
  NOR2X1 U328 ( .A(n377), .B(n150), .Y(n497) );
  OAI211X1 U329 ( .C(n55), .D(n376), .A(n502), .B(n503), .Y(n484) );
  NAND4X1 U330 ( .A(ff_idn), .B(n492), .C(n545), .D(n112), .Y(n503) );
  OAI31XL U331 ( .A(n276), .B(n504), .C(n113), .D(n543), .Y(n502) );
  NOR3XL U332 ( .A(n54), .B(n476), .C(n282), .Y(n412) );
  NAND2X1 U333 ( .A(ff_chg), .B(n545), .Y(n275) );
  OAI21BBX1 U334 ( .A(n56), .B(n497), .C(n496), .Y(n513) );
  INVX1 U335 ( .A(n474), .Y(n539) );
  NAND21X1 U336 ( .B(n285), .A(n222), .Y(n244) );
  NAND3X1 U337 ( .A(n545), .B(n244), .C(ff_idn), .Y(n278) );
  INVX1 U338 ( .A(n282), .Y(n547) );
  OAI21X1 U339 ( .B(n94), .C(n93), .A(n293), .Y(n286) );
  INVX1 U340 ( .A(n352), .Y(n540) );
  AOI21X1 U341 ( .B(n93), .C(n94), .A(n286), .Y(n461) );
  NOR2X1 U342 ( .A(n40), .B(n282), .Y(n526) );
  NOR32XL U343 ( .B(fcp_state[0]), .C(fcp_state[3]), .A(fcp_state[2]), .Y(n535) );
  NOR3XL U344 ( .A(n533), .B(fcp_state[1]), .C(n544), .Y(n352) );
  NAND2X1 U345 ( .A(n535), .B(fcp_state[1]), .Y(n376) );
  INVX1 U346 ( .A(fcp_state[1]), .Y(n551) );
  INVX1 U347 ( .A(fcp_state[2]), .Y(n544) );
  INVX1 U348 ( .A(fcp_state[0]), .Y(n552) );
  NAND2X1 U349 ( .A(fcp_state[3]), .B(n552), .Y(n533) );
  AOI22X1 U350 ( .A(r_wdat[1]), .B(n269), .C(r_dat[1]), .D(n270), .Y(n254) );
  AOI22X1 U351 ( .A(r_wdat[7]), .B(n269), .C(n270), .D(r_dat[7]), .Y(n263) );
  AOI22X1 U352 ( .A(r_wdat[0]), .B(n269), .C(r_dat[0]), .D(n270), .Y(n258) );
  AOI22X1 U353 ( .A(n23), .B(n269), .C(r_dat[2]), .D(n270), .Y(n255) );
  ENOX1 U354 ( .A(n35), .B(n79), .C(r_dat[6]), .D(n270), .Y(n251) );
  ENOX1 U355 ( .A(n33), .B(n79), .C(r_dat[4]), .D(n270), .Y(n250) );
  ENOX1 U356 ( .A(n25), .B(n79), .C(r_dat[3]), .D(n270), .Y(n252) );
  ENOX1 U357 ( .A(n34), .B(n79), .C(r_dat[5]), .D(n270), .Y(n248) );
  OAI32X1 U358 ( .A(n76), .B(n512), .C(n79), .D(r_ctl[7]), .E(n514), .Y(n495)
         );
  INVX1 U359 ( .A(r_ctl[4]), .Y(n76) );
  AOI22X1 U360 ( .A(n487), .B(n352), .C(n55), .D(n550), .Y(n514) );
  AO2222XL U361 ( .A(n249), .B(rxtx_buf[7]), .C(n250), .D(n77), .E(n52), .F(
        n59), .G(n42), .H(n251), .Y(trans_buf[8]) );
  AO2222XL U362 ( .A(rxtx_buf[9]), .B(n249), .C(n251), .D(n77), .E(n52), .F(
        n59), .G(n42), .H(n263), .Y(trans_buf[10]) );
  NAND32X1 U363 ( .B(n498), .C(n484), .A(n499), .Y(N1007) );
  AOI32X1 U364 ( .A(n547), .B(ff_idn), .C(n476), .D(n500), .E(n501), .Y(n499)
         );
  OAI21BBX1 U365 ( .A(n77), .B(r_ctl[1]), .C(n260), .Y(n501) );
  GEN2XL U366 ( .D(n486), .E(n549), .C(n497), .B(n538), .A(n495), .Y(n500) );
  NAND4X1 U367 ( .A(n287), .B(n288), .C(n289), .D(n290), .Y(intr) );
  AOI22X1 U368 ( .A(r_msk[2]), .B(r_irq[2]), .C(r_msk[3]), .D(r_irq[3]), .Y(
        n289) );
  AOI22X1 U369 ( .A(r_msk[4]), .B(r_irq[4]), .C(r_msk[5]), .D(r_irq[5]), .Y(
        n288) );
  AOI22X1 U370 ( .A(r_msk[6]), .B(r_irq[6]), .C(r_msk[7]), .D(r_irq[7]), .Y(
        n287) );
  OAI221X1 U371 ( .A(n487), .B(n540), .C(n54), .D(n539), .E(n489), .Y(N1008)
         );
  AOI31X1 U372 ( .A(r_ctl[0]), .B(n490), .C(r_ctl[1]), .D(n427), .Y(n489) );
  OAI31XL U373 ( .A(n276), .B(r_ctl[7]), .C(n488), .D(n39), .Y(n490) );
  NAND2X1 U374 ( .A(n262), .B(n247), .Y(trans_buf[11]) );
  AOI22X1 U375 ( .A(n59), .B(n13), .C(rxtx_buf[10]), .D(n249), .Y(n262) );
  NAND2X1 U376 ( .A(n246), .B(n247), .Y(trans_buf[9]) );
  AOI22X1 U377 ( .A(n248), .B(n13), .C(rxtx_buf[8]), .D(n249), .Y(n246) );
  AO2222XL U378 ( .A(n249), .B(rxtx_buf[5]), .C(n52), .D(n248), .E(n60), .F(
        n77), .G(n253), .H(n250), .Y(trans_buf[6]) );
  AO2222XL U379 ( .A(n249), .B(rxtx_buf[4]), .C(n52), .D(n250), .E(n62), .F(
        n77), .G(n253), .H(n252), .Y(trans_buf[5]) );
  INVX1 U380 ( .A(n254), .Y(n62) );
  AO2222XL U381 ( .A(n249), .B(rxtx_buf[6]), .C(n252), .D(n77), .E(n52), .F(
        n251), .G(n253), .H(n248), .Y(trans_buf[7]) );
  AO2222XL U382 ( .A(n249), .B(rxtx_buf[3]), .C(n52), .D(n252), .E(n61), .F(
        n77), .G(n253), .H(n60), .Y(trans_buf[4]) );
  OAI22X1 U383 ( .A(n22), .B(n81), .C(n155), .D(n163), .Y(tui_wdat[1]) );
  XNOR2XL U384 ( .A(n164), .B(n165), .Y(n163) );
  NAND2X1 U385 ( .A(N141), .B(N142), .Y(n165) );
  OAI211X1 U386 ( .C(r_ctl[1]), .D(n506), .A(n507), .B(n508), .Y(N1006) );
  AOI31X1 U387 ( .A(r_ctl[4]), .B(n546), .C(n512), .D(n412), .Y(n507) );
  AOI221XL U388 ( .A(n549), .B(n57), .C(n550), .D(n509), .E(n498), .Y(n508) );
  AOI21X1 U389 ( .B(n513), .C(n538), .A(n495), .Y(n506) );
  OAI21BBX1 U390 ( .A(N363), .B(n10), .C(n256), .Y(N261) );
  NAND31X1 U391 ( .C(n484), .A(n39), .B(n485), .Y(N1009) );
  OA222X1 U392 ( .A(n348), .B(n486), .C(n540), .D(n487), .E(n488), .F(r_ctl[7]), .Y(n485) );
  ENOX1 U393 ( .A(n15), .B(n33), .C(n80), .D(rxtx_buf[4]), .Y(upd_dbuf[4]) );
  ENOX1 U394 ( .A(n15), .B(n25), .C(n80), .D(rxtx_buf[3]), .Y(upd_dbuf[3]) );
  ENOX1 U395 ( .A(n15), .B(n34), .C(n80), .D(rxtx_buf[5]), .Y(upd_dbuf[5]) );
  ENOX1 U396 ( .A(n15), .B(n35), .C(n80), .D(rxtx_buf[6]), .Y(upd_dbuf[6]) );
  ENOX1 U397 ( .A(n36), .B(n80), .C(n80), .D(rxtx_buf[7]), .Y(upd_dbuf[7]) );
  OAI22X1 U398 ( .A(r_tui[7]), .B(n75), .C(catch_sync[3]), .D(n74), .Y(n334)
         );
  OAI22X1 U399 ( .A(r_tui[7]), .B(r_tui[3]), .C(catch_sync[1]), .D(n74), .Y(
        n291) );
  OAI22X1 U400 ( .A(catch_sync[4]), .B(n74), .C(r_tui[7]), .D(adp_tx_ui_6_), 
        .Y(n153) );
  OAI22X1 U401 ( .A(r_tui[7]), .B(r_tui[4]), .C(catch_sync[2]), .D(n74), .Y(
        n330) );
  OAI22X1 U402 ( .A(r_tui[7]), .B(r_tui[2]), .C(catch_sync[0]), .D(n74), .Y(
        n340) );
  OAI21X1 U403 ( .B(r_tui[6]), .C(n75), .A(adp_tx_ui_7_), .Y(adp_tx_ui_6_) );
  AO22X1 U404 ( .A(n408), .B(n14), .C(n29), .D(n407), .Y(N1013) );
  INVX1 U405 ( .A(r_tui[7]), .Y(n74) );
  INVX1 U406 ( .A(r_tui[5]), .Y(n75) );
  NAND2X1 U407 ( .A(n449), .B(ui_intv_cnt[5]), .Y(n445) );
  NAND2X1 U408 ( .A(r_tui[6]), .B(n75), .Y(adp_tx_ui_7_) );
  OAI221X1 U409 ( .A(rx_ui_3_8[3]), .B(n124), .C(rx_ui_3_8[2]), .D(n122), .E(
        n446), .Y(n444) );
  NOR2X1 U410 ( .A(ui_intv_cnt[0]), .B(n448), .Y(n447) );
  XNOR2XL U411 ( .A(n69), .B(n71), .Y(n448) );
  AOI32X1 U412 ( .A(n428), .B(n88), .C(n87), .D(n111), .E(n429), .Y(n409) );
  OR4X1 U413 ( .A(n430), .B(n431), .C(n40), .D(n84), .Y(n429) );
  OAI31XL U414 ( .A(n432), .B(ui_intv_cnt[6]), .C(ui_intv_cnt[5]), .D(n110), 
        .Y(n431) );
  AOI21BX1 U415 ( .C(n439), .B(n440), .A(n441), .Y(n430) );
  OAI21X1 U416 ( .B(ui_intv_cnt[5]), .C(n449), .A(n450), .Y(n440) );
  AOI33X1 U417 ( .A(n445), .B(n125), .C(rx_ui_3_8[4]), .D(n68), .E(n120), .F(
        add_263_carry[5]), .Y(n450) );
  AOI211X1 U418 ( .C(N142), .D(n64), .A(n442), .B(n439), .Y(n441) );
  INVX1 U419 ( .A(rx_ui_3_8[4]), .Y(n64) );
  GEN2XL U420 ( .D(N141), .E(n65), .C(n443), .B(n444), .A(n63), .Y(n442) );
  INVX1 U421 ( .A(rx_ui_3_8[3]), .Y(n65) );
  ENOX1 U422 ( .A(n406), .B(n118), .C(n26), .D(n407), .Y(N1016) );
  ENOX1 U423 ( .A(n406), .B(n537), .C(n32), .D(n407), .Y(N1010) );
  NOR21XL U424 ( .B(n211), .A(n212), .Y(n171) );
  OAI31XL U425 ( .A(n213), .B(n106), .C(n214), .D(n118), .Y(n212) );
  AOI33X1 U426 ( .A(n106), .B(n108), .C(symb_cnt[4]), .D(n214), .E(n20), .F(
        n213), .Y(n211) );
  NAND2X1 U427 ( .A(n215), .B(n216), .Y(n214) );
  AOI21X1 U428 ( .B(n129), .C(symb_cnt[3]), .A(n241), .Y(n232) );
  NOR2X1 U429 ( .A(n132), .B(symb_cnt[2]), .Y(n405) );
  NOR2X1 U430 ( .A(N159), .B(N160), .Y(n375) );
  NAND2X1 U431 ( .A(n121), .B(n451), .Y(n439) );
  OAI21BBX1 U432 ( .A(n68), .B(add_263_carry[5]), .C(ui_intv_cnt[6]), .Y(n451)
         );
  NOR2X1 U433 ( .A(n129), .B(symb_cnt[3]), .Y(n241) );
  NAND2X1 U434 ( .A(symb_cnt[2]), .B(n132), .Y(n404) );
  XNOR2XL U435 ( .A(N159), .B(n235), .Y(N108) );
  GEN2XL U436 ( .D(n515), .E(n373), .C(symb_cnt[2]), .B(symb_cnt[3]), .A(n369), 
        .Y(n349) );
  NAND21X1 U437 ( .B(n358), .A(n131), .Y(n515) );
  XNOR2XL U438 ( .A(N363), .B(n9), .Y(n382) );
  OAI22X1 U439 ( .A(catch_sync[5]), .B(n74), .C(r_tui[7]), .D(adp_tx_ui_7_), 
        .Y(n333) );
  XOR2X1 U440 ( .A(n215), .B(n229), .Y(n208) );
  OAI21X1 U441 ( .B(n230), .C(symb_cnt[5]), .A(n216), .Y(n229) );
  INVX1 U442 ( .A(N159), .Y(n537) );
  AOI21BBXL U443 ( .B(n337), .C(n73), .A(n338), .Y(n336) );
  AOI21X1 U444 ( .B(n73), .C(n337), .A(n122), .Y(n338) );
  OAI221X1 U445 ( .A(ui_intv_cnt[1]), .B(n339), .C(ui_intv_cnt[0]), .D(n291), 
        .E(n327), .Y(n337) );
  INVX1 U446 ( .A(N160), .Y(n131) );
  OAI32X1 U447 ( .A(n218), .B(n106), .C(n213), .D(n219), .E(n20), .Y(n172) );
  AOI31X1 U448 ( .A(n202), .B(n210), .C(n203), .D(symb_cnt[5]), .Y(n219) );
  NOR3XL U449 ( .A(n95), .B(r_ctl[7]), .C(n276), .Y(n270) );
  INVX1 U450 ( .A(n367), .Y(n96) );
  GEN2XL U451 ( .D(n97), .E(symb_cnt[2]), .C(symb_cnt[3]), .B(n368), .A(n369), 
        .Y(n367) );
  INVX1 U452 ( .A(n372), .Y(n97) );
  NAND2X1 U453 ( .A(n370), .B(n371), .Y(n368) );
  NOR2X1 U454 ( .A(n274), .B(symb_cnt[6]), .Y(n380) );
  NOR2X1 U455 ( .A(n115), .B(symb_cnt[2]), .Y(n518) );
  INVX1 U456 ( .A(symb_cnt[4]), .Y(n116) );
  OAI211X1 U457 ( .C(n517), .D(n114), .A(n378), .B(n492), .Y(n355) );
  AOI22X1 U458 ( .A(N363), .B(n130), .C(N362), .D(n131), .Y(n517) );
  OAI21X1 U459 ( .B(N160), .C(symb_cnt[2]), .A(n372), .Y(n371) );
  OAI21X1 U460 ( .B(N362), .C(N159), .A(n373), .Y(n370) );
  INVX1 U461 ( .A(symb_cnt[5]), .Y(n119) );
  OAI32X1 U462 ( .A(n87), .B(new_rx_sync_cnt[1]), .C(n37), .D(n306), .E(n88), 
        .Y(N349) );
  AOI21X1 U463 ( .B(n307), .C(n87), .A(n308), .Y(n306) );
  OAI22X1 U464 ( .A(N141), .B(n153), .C(ui_intv_cnt[2]), .D(n334), .Y(n437) );
  OAI21BBX1 U465 ( .A(n331), .B(n315), .C(n332), .Y(n311) );
  OAI21X1 U466 ( .B(n315), .C(n331), .A(n120), .Y(n332) );
  OAI221X1 U467 ( .A(N142), .B(n318), .C(ui_intv_cnt[5]), .D(n66), .E(n335), 
        .Y(n331) );
  OAI22AX1 U468 ( .D(n328), .C(n336), .A(n17), .B(n334), .Y(n335) );
  OAI21X1 U469 ( .B(n68), .C(n125), .A(n433), .Y(n432) );
  OAI22X1 U470 ( .A(N142), .B(n333), .C(n434), .D(n435), .Y(n433) );
  AOI21X1 U471 ( .B(n67), .C(n124), .A(n436), .Y(n435) );
  AOI211X1 U472 ( .C(n73), .D(n70), .A(n437), .B(n438), .Y(n434) );
  NAND3X1 U473 ( .A(n110), .B(n378), .C(n379), .Y(n360) );
  NAND41X1 U474 ( .D(n359), .A(n380), .B(n381), .C(n357), .Y(n379) );
  OAI22X1 U475 ( .A(N362), .B(N159), .C(N160), .D(n382), .Y(n381) );
  AOI22X1 U476 ( .A(N141), .B(n153), .C(ui_intv_cnt[2]), .D(n334), .Y(n436) );
  AOI21X1 U477 ( .B(n339), .C(n330), .A(ui_intv_cnt[1]), .Y(n438) );
  NAND3X1 U478 ( .A(N362), .B(n518), .C(N363), .Y(n378) );
  NAND2X1 U479 ( .A(n382), .B(N160), .Y(n357) );
  XNOR2XL U480 ( .A(n537), .B(symb_cnt[2]), .Y(N161) );
  NOR2X1 U481 ( .A(N159), .B(n123), .Y(add_274_carry[6]) );
  AND4X1 U482 ( .A(n384), .B(n385), .C(n386), .D(n387), .Y(n383) );
  XNOR2XL U483 ( .A(n402), .B(n107), .Y(n384) );
  XNOR2XL U484 ( .A(ui_intv_cnt[6]), .B(n401), .Y(n385) );
  NOR2X1 U485 ( .A(n397), .B(n398), .Y(n386) );
  OAI21X1 U486 ( .B(n228), .C(n221), .A(n222), .Y(n227) );
  NOR2X1 U487 ( .A(N160), .B(symb_cnt[3]), .Y(n228) );
  OAI31XL U488 ( .A(n114), .B(n365), .C(n374), .D(n110), .Y(n356) );
  AOI21X1 U489 ( .B(N362), .C(n537), .A(n131), .Y(n374) );
  OAI211X1 U490 ( .C(n56), .D(n541), .A(n109), .B(n294), .Y(n277) );
  AOI211X1 U491 ( .C(n295), .D(n296), .A(n16), .B(n264), .Y(n294) );
  INVX1 U492 ( .A(N141), .Y(n124) );
  NAND3X1 U493 ( .A(fcp_state[0]), .B(n494), .C(fcp_state[1]), .Y(n151) );
  INVX1 U494 ( .A(ui_intv_cnt[5]), .Y(n123) );
  XNOR2XL U495 ( .A(n392), .B(n122), .Y(n391) );
  ENOX1 U496 ( .A(n151), .B(n340), .C(r_tui[2]), .D(n393), .Y(n392) );
  NOR3XL U497 ( .A(n292), .B(us_cnt_2_), .C(n91), .Y(n281) );
  NAND4X1 U498 ( .A(n519), .B(n281), .C(n520), .D(n521), .Y(n276) );
  XNOR2XL U499 ( .A(n6), .B(r_tui[2]), .Y(n519) );
  NOR4XL U500 ( .A(n522), .B(n523), .C(n524), .D(n527), .Y(n521) );
  NOR3XL U501 ( .A(n528), .B(n529), .C(n530), .Y(n520) );
  OAI21X1 U502 ( .B(n221), .C(n222), .A(n223), .Y(n192) );
  AOI32X1 U503 ( .A(n221), .B(n131), .C(symb_cnt[3]), .D(n224), .E(n126), .Y(
        n223) );
  XNOR2XL U504 ( .A(N160), .B(n221), .Y(n224) );
  NOR2X1 U505 ( .A(n115), .B(symb_cnt[3]), .Y(n504) );
  INVX1 U506 ( .A(symb_cnt[2]), .Y(n128) );
  INVX1 U507 ( .A(ui_intv_cnt[1]), .Y(n117) );
  BUFX3 U508 ( .A(n188), .Y(n20) );
  GEN2XL U509 ( .D(N142), .E(n242), .C(ui_intv_cnt[5]), .B(ui_intv_cnt[6]), 
        .A(ui_intv_cnt[7]), .Y(n188) );
  NAND4X1 U510 ( .A(n124), .B(n107), .C(n117), .D(n122), .Y(n242) );
  INVX1 U511 ( .A(ui_intv_cnt[2]), .Y(n122) );
  OAI22X1 U512 ( .A(n127), .B(n128), .C(n226), .D(n116), .Y(n225) );
  NOR2X1 U513 ( .A(symb_cnt[2]), .B(n227), .Y(n226) );
  INVX1 U514 ( .A(ui_intv_cnt[0]), .Y(n107) );
  INVX1 U515 ( .A(N362), .Y(n100) );
  AOI21X1 U516 ( .B(N362), .C(N363), .A(n128), .Y(n359) );
  AOI21X1 U517 ( .B(n375), .C(N362), .A(N363), .Y(n365) );
  ENOX1 U518 ( .A(n144), .B(n151), .C(r_tui[1]), .D(n393), .Y(n395) );
  ENOX1 U519 ( .A(n291), .B(n151), .C(r_tui[3]), .D(n393), .Y(n394) );
  NOR2X1 U520 ( .A(fcp_state[2]), .B(fcp_state[3]), .Y(n494) );
  NOR4XL U521 ( .A(n388), .B(n389), .C(n390), .D(n391), .Y(n387) );
  XNOR2XL U522 ( .A(ui_intv_cnt[5]), .B(n396), .Y(n388) );
  XNOR2XL U523 ( .A(n395), .B(n117), .Y(n389) );
  XNOR2XL U524 ( .A(n394), .B(n124), .Y(n390) );
  NAND2X1 U525 ( .A(symb_cnt[2]), .B(N159), .Y(n221) );
  NAND4X1 U526 ( .A(n463), .B(n459), .C(n465), .D(n466), .Y(n296) );
  XNOR2XL U527 ( .A(ui_intv_cnt[2]), .B(adp_tx_1_4[2]), .Y(n463) );
  NOR2X1 U528 ( .A(n471), .B(n472), .Y(n465) );
  NOR4XL U529 ( .A(n467), .B(n468), .C(n469), .D(n470), .Y(n466) );
  AOI221XL U530 ( .A(n315), .B(n120), .C(n316), .D(n123), .E(n317), .Y(n314)
         );
  AOI22X1 U531 ( .A(n66), .B(ui_intv_cnt[5]), .C(n318), .D(N142), .Y(n317) );
  ENOX1 U532 ( .A(new_rx_sync_cnt[0]), .B(n37), .C(new_rx_sync_cnt[0]), .D(
        n308), .Y(N348) );
  NAND3X1 U533 ( .A(us_cnt_0_), .B(n293), .C(us_cnt_1_), .Y(n292) );
  AOI22X1 U534 ( .A(r_msk[0]), .B(r_irq[0]), .C(r_msk[1]), .D(r_irq[1]), .Y(
        n290) );
  NOR43XL U535 ( .B(n477), .C(n120), .D(ui_intv_cnt[2]), .A(n478), .Y(n413) );
  XNOR2XL U536 ( .A(n123), .B(n124), .Y(n477) );
  AOI22AXL U537 ( .A(n482), .B(n109), .D(n483), .C(N363), .Y(n415) );
  AOI21X1 U538 ( .B(n366), .C(n482), .A(n109), .Y(n483) );
  NAND2X1 U539 ( .A(N159), .B(n100), .Y(n482) );
  XNOR2XL U540 ( .A(n152), .B(n153), .Y(n148) );
  XNOR2XL U541 ( .A(n11), .B(add_264_carry[5]), .Y(n152) );
  AND4X1 U542 ( .A(n452), .B(n453), .C(n454), .D(n455), .Y(n422) );
  XNOR2XL U543 ( .A(n71), .B(ui_intv_cnt[2]), .Y(n453) );
  XNOR2XL U544 ( .A(n67), .B(ui_intv_cnt[5]), .Y(n452) );
  NOR4XL U545 ( .A(n456), .B(n457), .C(n458), .D(n141), .Y(n455) );
  XNOR2XL U546 ( .A(n117), .B(r_tui[1]), .Y(n524) );
  XNOR2XL U547 ( .A(ui_intv_cnt[7]), .B(n399), .Y(n398) );
  AOI221XL U548 ( .A(n545), .B(n68), .C(n393), .D(adp_tx_ui_7_), .E(n245), .Y(
        n399) );
  XNOR2XL U549 ( .A(n125), .B(r_tui[4]), .Y(n527) );
  XNOR2XL U550 ( .A(n400), .B(n125), .Y(n397) );
  ENOX1 U551 ( .A(n151), .B(n330), .C(r_tui[4]), .D(n393), .Y(n400) );
  XNOR2XL U552 ( .A(n107), .B(r_tui[0]), .Y(n523) );
  XNOR2XL U553 ( .A(n124), .B(r_tui[3]), .Y(n522) );
  INVX1 U554 ( .A(symb_cnt[3]), .Y(n126) );
  NOR4XL U555 ( .A(n537), .B(n126), .C(n114), .D(N160), .Y(n428) );
  INVX1 U556 ( .A(N142), .Y(n125) );
  NAND21X1 U557 ( .B(n403), .A(r_tui[0]), .Y(n402) );
  AOI21X1 U558 ( .B(n74), .C(n545), .A(n393), .Y(n403) );
  INVX1 U559 ( .A(ui_intv_cnt[6]), .Y(n120) );
  INVX1 U560 ( .A(ui_intv_cnt[7]), .Y(n121) );
  NAND2X1 U561 ( .A(symb_cnt[3]), .B(n225), .Y(n217) );
  NOR2X1 U562 ( .A(n110), .B(n12), .Y(n366) );
  NOR2X1 U563 ( .A(n90), .B(ui_intv_cnt[7]), .Y(n459) );
  NAND4X1 U564 ( .A(n459), .B(N142), .C(n107), .D(n117), .Y(n478) );
  OAI22X1 U565 ( .A(n322), .B(n323), .C(ui_intv_cnt[5]), .D(n321), .Y(n319) );
  NOR2X1 U566 ( .A(n324), .B(n318), .Y(n323) );
  AOI21X1 U567 ( .B(n324), .C(n318), .A(n125), .Y(n322) );
  AND2X1 U568 ( .A(n325), .B(n326), .Y(n324) );
  NAND2X1 U569 ( .A(r_tui[1]), .B(n74), .Y(n144) );
  AOI31X1 U570 ( .A(n56), .B(n361), .C(n362), .D(n363), .Y(n346) );
  AO21X1 U571 ( .B(n309), .C(n364), .A(n365), .Y(n362) );
  AO222X1 U572 ( .A(n352), .B(n360), .C(n354), .D(n356), .E(n96), .F(n549), 
        .Y(n361) );
  NAND3X1 U573 ( .A(N362), .B(n537), .C(n366), .Y(n364) );
  AOI32X1 U574 ( .A(n330), .B(n328), .C(ui_intv_cnt[2]), .D(n72), .E(N141), 
        .Y(n325) );
  NAND2X1 U575 ( .A(N160), .B(symb_cnt[3]), .Y(n222) );
  OAI211X1 U576 ( .C(ui_intv_cnt[0]), .D(n327), .A(n328), .B(n329), .Y(n326)
         );
  AOI22X1 U577 ( .A(n73), .B(n122), .C(n71), .D(n117), .Y(n329) );
  AOI221XL U578 ( .A(n543), .B(n126), .C(n415), .D(n416), .E(n417), .Y(n414)
         );
  AOI21X1 U579 ( .B(n418), .C(n12), .A(n348), .Y(n417) );
  ENOX1 U580 ( .A(n349), .B(n376), .C(n355), .D(n352), .Y(n416) );
  NAND2X1 U581 ( .A(n11), .B(n321), .Y(n320) );
  NOR32XL U582 ( .B(n7), .C(n366), .A(N159), .Y(n476) );
  AOI21X1 U583 ( .B(n493), .C(fcp_state[2]), .A(n245), .Y(n479) );
  XNOR2XL U584 ( .A(rx_ui_5_8[4]), .B(N142), .Y(n146) );
  XNOR2XL U585 ( .A(n144), .B(ui_intv_cnt[0]), .Y(n457) );
  NOR3XL U586 ( .A(n40), .B(n16), .C(n309), .Y(n512) );
  INVX1 U587 ( .A(test_so), .Y(n91) );
  NOR21XL U588 ( .B(n536), .A(n297), .Y(N356) );
  XNOR2XL U589 ( .A(rxtx_buf[0]), .B(n298), .Y(n297) );
  XNOR2XL U590 ( .A(n299), .B(n300), .Y(n298) );
  XNOR2XL U591 ( .A(n301), .B(n302), .Y(n300) );
  XNOR2XL U592 ( .A(ui_intv_cnt[2]), .B(rx_ui_5_8[2]), .Y(n147) );
  XNOR2XL U593 ( .A(r_dat[7]), .B(n8), .Y(n344) );
  NOR4XL U594 ( .A(n544), .B(fcp_state[0]), .C(fcp_state[1]), .D(fcp_state[3]), 
        .Y(n474) );
  NAND3X1 U595 ( .A(n494), .B(n551), .C(fcp_state[0]), .Y(n282) );
  NOR3XL U596 ( .A(n88), .B(new_rx_sync_cnt[0]), .C(n275), .Y(setsta[3]) );
  AND3X1 U597 ( .A(symb_cnt[5]), .B(n481), .C(symb_cnt[6]), .Y(n473) );
  NAND3X1 U598 ( .A(n126), .B(n116), .C(n128), .Y(n481) );
  NAND2X1 U599 ( .A(n14), .B(n505), .Y(n150) );
  INVX1 U600 ( .A(symb_cnt[6]), .Y(n118) );
  NAND4X1 U601 ( .A(n418), .B(n504), .C(n549), .D(n12), .Y(n496) );
  NAND2X1 U602 ( .A(n510), .B(n511), .Y(n498) );
  NAND4X1 U603 ( .A(n547), .B(n109), .C(n16), .D(n54), .Y(n511) );
  OAI21X1 U604 ( .B(n428), .C(n111), .A(n545), .Y(n510) );
  INVX1 U605 ( .A(rx_trans_8_chg), .Y(n84) );
  NOR3XL U606 ( .A(n273), .B(n54), .C(n539), .Y(setsta[6]) );
  NAND3X1 U607 ( .A(symb_cnt[6]), .B(n274), .C(ff_chg), .Y(n273) );
  XNOR2XL U608 ( .A(ui_intv_cnt[1]), .B(rx_ui_5_8[1]), .Y(n138) );
  XNOR2XL U609 ( .A(n143), .B(n144), .Y(n136) );
  XNOR2XL U610 ( .A(n71), .B(ui_intv_cnt[0]), .Y(n143) );
  XNOR2XL U611 ( .A(n303), .B(n304), .Y(n299) );
  XNOR2XL U612 ( .A(rxtx_buf[3]), .B(rxtx_buf[2]), .Y(n304) );
  XNOR2XL U613 ( .A(n82), .B(n54), .Y(n303) );
  INVX1 U614 ( .A(r_ctl[0]), .Y(n77) );
  OAI32X1 U615 ( .A(n292), .B(us_cnt_2_), .C(n281), .D(n286), .E(n92), .Y(N87)
         );
  INVX1 U616 ( .A(r_ctl[7]), .Y(n538) );
  INVX1 U617 ( .A(new_rx_sync_cnt[0]), .Y(n87) );
  INVX1 U618 ( .A(new_rx_sync_cnt[1]), .Y(n88) );
  XNOR2XL U620 ( .A(rxtx_buf[5]), .B(rxtx_buf[4]), .Y(n301) );
  XNOR2XL U621 ( .A(rxtx_buf[7]), .B(rxtx_buf[6]), .Y(n302) );
  OAI32X1 U622 ( .A(n275), .B(rx_trans_8_chg), .C(n150), .D(ff_chg), .E(n84), 
        .Y(n516) );
  OAI32X1 U623 ( .A(n92), .B(test_so), .C(n292), .D(n91), .E(n286), .Y(N88) );
  OR2X1 U624 ( .A(r_ctl[1]), .B(n77), .Y(n260) );
  INVX1 U625 ( .A(rxtx_buf[1]), .Y(n82) );
  NAND4X1 U626 ( .A(n151), .B(n264), .C(n531), .D(n532), .Y(N1005) );
  AOI211X1 U627 ( .C(ff_chg), .D(n285), .A(n54), .B(n551), .Y(n532) );
  AOI21X1 U628 ( .B(fcp_state[2]), .C(n533), .A(n283), .Y(n531) );
  INVX1 U629 ( .A(us_cnt_0_), .Y(n94) );
  INVX1 U630 ( .A(rxtx_buf[2]), .Y(n86) );
  INVX1 U631 ( .A(us_cnt_1_), .Y(n93) );
  NOR2X1 U632 ( .A(us_cnt_0_), .B(n546), .Y(N85) );
  INVX1 U633 ( .A(us_cnt_2_), .Y(n92) );
  INVX1 U634 ( .A(rxtx_buf[0]), .Y(n85) );
  BUFX3 U635 ( .A(r_ctl[6]), .Y(tx_en) );
  INVX1 U636 ( .A(n264), .Y(r_ctl[6]) );
endmodule


module fcpegn_a0_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module fcpegn_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(SUM[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
endmodule


module fcpegn_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9515;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9515), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9515), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9515), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9515), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9515), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9515), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9515), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9515), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9515), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9533;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9533), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9533), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9533), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9533), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9533), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9533), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9533), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9533), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9533), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9551;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9551), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9551), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9551), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9551), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9551), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9551), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9551), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9551), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9551), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_0 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_0 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[2]), .Y(n2) );
  INVX1 U3 ( .A(set2[0]), .Y(n14) );
  INVX1 U4 ( .A(set2[1]), .Y(n13) );
  INVX1 U5 ( .A(set2[4]), .Y(n15) );
  NOR3XL U6 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NAND3X1 U7 ( .A(n4), .B(n1), .C(n16), .Y(n21) );
  INVX1 U8 ( .A(set2[3]), .Y(n3) );
  INVX1 U9 ( .A(set2[7]), .Y(n1) );
  NOR2X1 U10 ( .A(rdat[6]), .B(n4), .Y(irq[6]) );
  NOR2X1 U11 ( .A(rdat[7]), .B(n1), .Y(irq[7]) );
  NAND4X1 U12 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U13 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR4XL U14 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U15 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  AOI211X1 U16 ( .C(n14), .D(n12), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U17 ( .A(rdat[0]), .Y(n12) );
  AOI211X1 U18 ( .C(n13), .D(n11), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U19 ( .A(rdat[1]), .Y(n11) );
  AOI211X1 U20 ( .C(n2), .D(n10), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U21 ( .A(rdat[2]), .Y(n10) );
  AOI211X1 U22 ( .C(n3), .D(n9), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U23 ( .A(rdat[3]), .Y(n9) );
  AOI211X1 U24 ( .C(n16), .D(n8), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U25 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U26 ( .C(n4), .D(n7), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U27 ( .A(rdat[6]), .Y(n7) );
  AOI211X1 U28 ( .C(n1), .D(n6), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U29 ( .A(rdat[7]), .Y(n6) );
  AOI211X1 U30 ( .C(n15), .D(n5), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U31 ( .A(rdat[4]), .Y(n5) );
  NOR2X1 U32 ( .A(rdat[0]), .B(n14), .Y(irq[0]) );
  NOR2X1 U33 ( .A(rdat[1]), .B(n13), .Y(irq[1]) );
  NOR2X1 U34 ( .A(rdat[4]), .B(n15), .Y(irq[4]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n2), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[3]), .B(n3), .Y(irq[3]) );
  INVX1 U37 ( .A(set2[6]), .Y(n4) );
  INVX1 U38 ( .A(set2[5]), .Y(n16) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9569;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9569), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9569), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9569), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9569), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9569), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9569), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9569), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9569), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9569), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000000 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9587;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9587), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9587), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9587), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9587), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9587), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9587), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9587), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9587), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9587), 
        .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dpdmacc_a0 ( dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, r_wdat, r_acc, 
        r_dpdmsta, r_dm, r_dmchg, r_int, clk, rstz, test_si, test_se );
  input [7:0] r_wdat;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, clk, rstz, test_si, test_se;
  output r_dm, r_dmchg, r_int;
  wire   dp_chg, dp_rise, dm_fall, dp_active_acc, dp_inacti_acc, dm_active_acc,
         dm_inacti_acc, upd00, n3, n4, n5, n6, n27, n28, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n2, n7, n8, n9, n10, n11, n38;
  wire   [7:0] wd00;

  INVX1 U5 ( .A(n6), .Y(n4) );
  INVX1 U6 ( .A(n6), .Y(n3) );
  INVX1 U7 ( .A(n6), .Y(n5) );
  INVX1 U8 ( .A(rstz), .Y(n6) );
  ff_sync_2 u0_dpsync ( .i_org(dp_comp), .o_dbc(r_dpdmsta[6]), .o_chg(dp_chg), 
        .clk(clk), .rstz(n4), .test_si(n27), .test_se(test_se) );
  ff_sync_1 u0_dmsync ( .i_org(dm_comp), .o_dbc(r_dpdmsta[7]), .o_chg(r_dmchg), 
        .clk(clk), .rstz(n4), .test_si(n28), .test_se(test_se) );
  ff_sync_0 u0_idsync ( .i_org(id_comp), .o_dbc(r_dpdmsta[5]), .o_chg(), .clk(
        clk), .rstz(n5), .test_si(r_dpdmsta[6]), .test_se(test_se) );
  filter150us_a0_1 u0_dpfltr ( .active_hit(dp_active_acc), .inacti_hit(
        dp_inacti_acc), .start_edge(dp_rise), .any_edge(dp_chg), .clk(clk), 
        .rstz(n5), .test_si(r_dpdmsta[4]), .test_so(n27), .test_se(test_se) );
  filter150us_a0_0 u0_dmfltr ( .active_hit(dm_active_acc), .inacti_hit(
        dm_inacti_acc), .start_edge(dm_fall), .any_edge(r_dmchg), .clk(clk), 
        .rstz(n5), .test_si(r_acc[7]), .test_so(n28), .test_se(test_se) );
  glreg_a0_5 u0_accmltr ( .clk(clk), .arstz(n3), .we(upd00), .wdat(wd00), 
        .rdat(r_acc), .test_si(test_si), .test_se(test_se) );
  glreg_WIDTH5_0 u0_dpdmsta ( .clk(clk), .arstz(n4), .we(r_wr_1), .wdat(
        r_wdat[4:0]), .rdat(r_dpdmsta[4:0]), .test_si(r_dpdmsta[7]), .test_se(
        test_se) );
  NAND2X1 U3 ( .A(n32), .B(n38), .Y(upd00) );
  INVX1 U4 ( .A(r_re_0), .Y(n38) );
  NOR2X1 U9 ( .A(n2), .B(n7), .Y(n32) );
  OAI22X1 U10 ( .A(n38), .B(n29), .C(r_re_0), .D(n30), .Y(wd00[0]) );
  XNOR2XL U11 ( .A(n26), .B(n11), .Y(n30) );
  OAI22X1 U12 ( .A(n18), .B(n38), .C(r_re_0), .D(n19), .Y(wd00[4]) );
  XNOR2XL U13 ( .A(n17), .B(n10), .Y(n19) );
  INVX1 U14 ( .A(n29), .Y(n7) );
  INVX1 U15 ( .A(n18), .Y(n2) );
  NOR2X1 U16 ( .A(n17), .B(n10), .Y(n15) );
  NOR2X1 U17 ( .A(n26), .B(n11), .Y(n24) );
  BUFX3 U18 ( .A(r_dpdmsta[7]), .Y(r_dm) );
  OAI21X1 U19 ( .B(n32), .C(n38), .A(n33), .Y(r_int) );
  AOI33X1 U20 ( .A(n7), .B(n11), .C(n34), .D(n2), .E(n10), .F(n35), .Y(n33) );
  NOR3XL U21 ( .A(r_acc[5]), .B(r_acc[7]), .C(r_acc[6]), .Y(n35) );
  AOI21BX1 U22 ( .C(r_acc[7]), .B(n12), .A(r_re_0), .Y(wd00[7]) );
  NAND21X1 U23 ( .B(n13), .A(r_acc[6]), .Y(n12) );
  AOI21BX1 U24 ( .C(r_acc[3]), .B(n21), .A(r_re_0), .Y(wd00[3]) );
  NAND21X1 U25 ( .B(n22), .A(r_acc[2]), .Y(n21) );
  NOR2X1 U26 ( .A(r_re_0), .B(n25), .Y(wd00[1]) );
  XNOR2XL U27 ( .A(r_acc[1]), .B(n24), .Y(n25) );
  NOR2X1 U28 ( .A(r_re_0), .B(n16), .Y(wd00[5]) );
  XNOR2XL U29 ( .A(r_acc[5]), .B(n15), .Y(n16) );
  NOR2X1 U30 ( .A(r_re_0), .B(n23), .Y(wd00[2]) );
  XOR2X1 U31 ( .A(n22), .B(r_acc[2]), .Y(n23) );
  NOR2X1 U32 ( .A(r_re_0), .B(n14), .Y(wd00[6]) );
  XOR2X1 U33 ( .A(n13), .B(r_acc[6]), .Y(n14) );
  OAI21X1 U34 ( .B(dm_inacti_acc), .C(n9), .A(n37), .Y(n18) );
  OAI21BX1 U35 ( .C(dm_active_acc), .B(r_dpdmsta[7]), .A(n9), .Y(n37) );
  INVX1 U36 ( .A(r_dpdmsta[1]), .Y(n9) );
  OAI21X1 U37 ( .B(dp_inacti_acc), .C(n8), .A(n36), .Y(n29) );
  OAI21BBX1 U38 ( .A(r_dpdmsta[6]), .B(dp_active_acc), .C(n8), .Y(n36) );
  INVX1 U39 ( .A(r_dpdmsta[0]), .Y(n8) );
  NOR21XL U40 ( .B(dp_chg), .A(r_dpdmsta[6]), .Y(dp_rise) );
  AND2X1 U41 ( .A(r_dpdmsta[7]), .B(r_dmchg), .Y(dm_fall) );
  NAND2X1 U42 ( .A(n2), .B(n20), .Y(n17) );
  NAND4X1 U43 ( .A(r_acc[6]), .B(r_acc[5]), .C(r_acc[4]), .D(r_acc[7]), .Y(n20) );
  NAND2X1 U44 ( .A(n15), .B(r_acc[5]), .Y(n13) );
  INVX1 U45 ( .A(r_acc[0]), .Y(n11) );
  NOR3XL U46 ( .A(r_acc[1]), .B(r_acc[3]), .C(r_acc[2]), .Y(n34) );
  NAND2X1 U47 ( .A(n7), .B(n31), .Y(n26) );
  NAND4X1 U48 ( .A(r_acc[2]), .B(r_acc[1]), .C(r_acc[0]), .D(r_acc[3]), .Y(n31) );
  NAND2X1 U49 ( .A(n24), .B(r_acc[1]), .Y(n22) );
  INVX1 U50 ( .A(r_acc[4]), .Y(n10) );
endmodule


module glreg_WIDTH5_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9605;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9605), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9605), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9605), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9605), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9605), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9605), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9623;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9623), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9623), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9623), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9623), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9623), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9623), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9623), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9623), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9623), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_0 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz, test_si, test_so, test_se );
  input start_edge, any_edge, clk, rstz, test_si, test_se;
  output active_hit, inacti_hit, test_so;
  wire   dbcnt_10_, dbcnt_9_, dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_,
         dbcnt_3_, dbcnt_2_, dbcnt_1_, dbcnt_0_, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, net9641, n2, n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n4, n14;

  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9641), .TE(test_se) );
  filter150us_a0_0_DW01_inc_0 add_76 ( .A({test_so, dbcnt_10_, dbcnt_9_, 
        dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_, dbcnt_3_, dbcnt_2_, 
        dbcnt_1_, dbcnt_0_}), .SUM({N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12}) );
  SDFFRQX1 dbcnt_reg_4_ ( .D(N29), .SIN(dbcnt_3_), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_4_) );
  SDFFRQX1 dbcnt_reg_3_ ( .D(N28), .SIN(dbcnt_2_), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_3_) );
  SDFFRQX1 dbcnt_reg_11_ ( .D(N36), .SIN(dbcnt_10_), .SMC(test_se), .C(net9641), .XR(n2), .Q(test_so) );
  SDFFRQX1 dbcnt_reg_2_ ( .D(N27), .SIN(dbcnt_1_), .SMC(test_se), .C(net9641), 
        .XR(rstz), .Q(dbcnt_2_) );
  SDFFRQX1 dbcnt_reg_1_ ( .D(N26), .SIN(dbcnt_0_), .SMC(test_se), .C(net9641), 
        .XR(rstz), .Q(dbcnt_1_) );
  SDFFRQX1 dbcnt_reg_0_ ( .D(N25), .SIN(test_si), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_0_) );
  SDFFRQX1 dbcnt_reg_7_ ( .D(N32), .SIN(dbcnt_6_), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_7_) );
  SDFFRQX1 dbcnt_reg_5_ ( .D(N30), .SIN(dbcnt_4_), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_5_) );
  SDFFRQX1 dbcnt_reg_6_ ( .D(N31), .SIN(dbcnt_5_), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_6_) );
  SDFFRQX1 dbcnt_reg_9_ ( .D(N34), .SIN(dbcnt_8_), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_9_) );
  SDFFRQX1 dbcnt_reg_8_ ( .D(N33), .SIN(dbcnt_7_), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_8_) );
  SDFFRQX1 dbcnt_reg_10_ ( .D(N35), .SIN(dbcnt_9_), .SMC(test_se), .C(net9641), 
        .XR(n2), .Q(dbcnt_10_) );
  BUFX3 U3 ( .A(n9), .Y(n1) );
  INVX1 U6 ( .A(any_edge), .Y(n4) );
  AND2X1 U7 ( .A(N22), .B(n9), .Y(N35) );
  AND2X1 U8 ( .A(N20), .B(n9), .Y(N33) );
  AND2X1 U9 ( .A(N21), .B(n9), .Y(N34) );
  NOR3XL U10 ( .A(n11), .B(any_edge), .C(n14), .Y(n9) );
  AND2X1 U11 ( .A(N16), .B(n9), .Y(N29) );
  AND2X1 U12 ( .A(N15), .B(n9), .Y(N28) );
  AND2X1 U13 ( .A(N19), .B(n9), .Y(N32) );
  AND2X1 U14 ( .A(N17), .B(n9), .Y(N30) );
  AND2X1 U15 ( .A(N18), .B(n9), .Y(N31) );
  AND2X1 U16 ( .A(N14), .B(n1), .Y(N27) );
  AND2X1 U17 ( .A(N13), .B(n1), .Y(N26) );
  INVX1 U18 ( .A(n5), .Y(n14) );
  OR2X1 U19 ( .A(n1), .B(any_edge), .Y(N24) );
  AOI211X1 U20 ( .C(n5), .D(n6), .A(n4), .B(start_edge), .Y(inacti_hit) );
  AOI21X1 U21 ( .B(n7), .C(n8), .A(test_so), .Y(n5) );
  NAND32X1 U22 ( .B(dbcnt_4_), .C(dbcnt_3_), .A(n13), .Y(n7) );
  NOR3XL U23 ( .A(dbcnt_5_), .B(dbcnt_7_), .C(dbcnt_6_), .Y(n13) );
  AND3X1 U24 ( .A(dbcnt_8_), .B(dbcnt_10_), .C(dbcnt_9_), .Y(n8) );
  NOR3XL U25 ( .A(n6), .B(test_so), .C(n7), .Y(active_hit) );
  NAND4X1 U26 ( .A(dbcnt_2_), .B(dbcnt_1_), .C(dbcnt_0_), .D(n8), .Y(n6) );
  AND2X1 U27 ( .A(N23), .B(n1), .Y(N36) );
  NOR4XL U28 ( .A(dbcnt_0_), .B(dbcnt_10_), .C(n7), .D(n12), .Y(n11) );
  OR4X1 U29 ( .A(dbcnt_9_), .B(dbcnt_8_), .C(dbcnt_2_), .D(dbcnt_1_), .Y(n12)
         );
  OAI21BBX1 U30 ( .A(N12), .B(n9), .C(n10), .Y(N25) );
  OAI21X1 U31 ( .B(n11), .C(n14), .A(any_edge), .Y(n10) );
endmodule


module filter150us_a0_0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_1 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz, test_si, test_so, test_se );
  input start_edge, any_edge, clk, rstz, test_si, test_se;
  output active_hit, inacti_hit, test_so;
  wire   dbcnt_10_, dbcnt_9_, dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_,
         dbcnt_3_, dbcnt_2_, dbcnt_1_, dbcnt_0_, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, net9659, n2, n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n4, n14;

  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9659), .TE(test_se) );
  filter150us_a0_1_DW01_inc_0 add_76 ( .A({test_so, dbcnt_10_, dbcnt_9_, 
        dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_, dbcnt_3_, dbcnt_2_, 
        dbcnt_1_, dbcnt_0_}), .SUM({N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12}) );
  SDFFRQX1 dbcnt_reg_4_ ( .D(N29), .SIN(dbcnt_3_), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_4_) );
  SDFFRQX1 dbcnt_reg_3_ ( .D(N28), .SIN(dbcnt_2_), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_3_) );
  SDFFRQX1 dbcnt_reg_11_ ( .D(N36), .SIN(dbcnt_10_), .SMC(test_se), .C(net9659), .XR(n2), .Q(test_so) );
  SDFFRQX1 dbcnt_reg_2_ ( .D(N27), .SIN(dbcnt_1_), .SMC(test_se), .C(net9659), 
        .XR(rstz), .Q(dbcnt_2_) );
  SDFFRQX1 dbcnt_reg_1_ ( .D(N26), .SIN(dbcnt_0_), .SMC(test_se), .C(net9659), 
        .XR(rstz), .Q(dbcnt_1_) );
  SDFFRQX1 dbcnt_reg_0_ ( .D(N25), .SIN(test_si), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_0_) );
  SDFFRQX1 dbcnt_reg_7_ ( .D(N32), .SIN(dbcnt_6_), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_7_) );
  SDFFRQX1 dbcnt_reg_5_ ( .D(N30), .SIN(dbcnt_4_), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_5_) );
  SDFFRQX1 dbcnt_reg_6_ ( .D(N31), .SIN(dbcnt_5_), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_6_) );
  SDFFRQX1 dbcnt_reg_9_ ( .D(N34), .SIN(dbcnt_8_), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_9_) );
  SDFFRQX1 dbcnt_reg_8_ ( .D(N33), .SIN(dbcnt_7_), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_8_) );
  SDFFRQX1 dbcnt_reg_10_ ( .D(N35), .SIN(dbcnt_9_), .SMC(test_se), .C(net9659), 
        .XR(n2), .Q(dbcnt_10_) );
  BUFX3 U3 ( .A(n9), .Y(n1) );
  INVX1 U6 ( .A(any_edge), .Y(n14) );
  AND2X1 U7 ( .A(N22), .B(n9), .Y(N35) );
  AND2X1 U8 ( .A(N20), .B(n9), .Y(N33) );
  AND2X1 U9 ( .A(N21), .B(n9), .Y(N34) );
  NOR3XL U10 ( .A(n11), .B(any_edge), .C(n4), .Y(n9) );
  AND2X1 U11 ( .A(N15), .B(n9), .Y(N28) );
  AND2X1 U12 ( .A(N19), .B(n9), .Y(N32) );
  AND2X1 U13 ( .A(N17), .B(n9), .Y(N30) );
  AND2X1 U14 ( .A(N18), .B(n9), .Y(N31) );
  AND2X1 U15 ( .A(N14), .B(n9), .Y(N27) );
  AND2X1 U16 ( .A(N13), .B(n1), .Y(N26) );
  AND2X1 U17 ( .A(N16), .B(n1), .Y(N29) );
  INVX1 U18 ( .A(n5), .Y(n4) );
  OR2X1 U19 ( .A(n1), .B(any_edge), .Y(N24) );
  AOI211X1 U20 ( .C(n5), .D(n6), .A(n14), .B(start_edge), .Y(inacti_hit) );
  AOI21X1 U21 ( .B(n7), .C(n8), .A(test_so), .Y(n5) );
  NAND32X1 U22 ( .B(dbcnt_4_), .C(dbcnt_3_), .A(n13), .Y(n7) );
  NOR3XL U23 ( .A(dbcnt_5_), .B(dbcnt_7_), .C(dbcnt_6_), .Y(n13) );
  AND3X1 U24 ( .A(dbcnt_8_), .B(dbcnt_10_), .C(dbcnt_9_), .Y(n8) );
  NOR3XL U25 ( .A(n6), .B(test_so), .C(n7), .Y(active_hit) );
  NAND4X1 U26 ( .A(dbcnt_2_), .B(dbcnt_1_), .C(dbcnt_0_), .D(n8), .Y(n6) );
  AND2X1 U27 ( .A(N23), .B(n1), .Y(N36) );
  NOR4XL U28 ( .A(dbcnt_0_), .B(dbcnt_10_), .C(n7), .D(n12), .Y(n11) );
  OR4X1 U29 ( .A(dbcnt_9_), .B(dbcnt_8_), .C(dbcnt_2_), .D(dbcnt_1_), .Y(n12)
         );
  OAI21BBX1 U30 ( .A(N12), .B(n9), .C(n10), .Y(N25) );
  OAI21X1 U31 ( .B(n11), .C(n4), .A(any_edge), .Y(n10) );
endmodule


module filter150us_a0_1_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ff_sync_0 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg;
  wire   d_org_0_;

  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_1 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg;
  wire   d_org_0_;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_2 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg;
  wire   d_org_0_;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module dacmux_a0 ( clk, srstz, i_comp, r_comp_opt, r_wdat, r_adofs, r_isofs, 
        r_wr, dacv_wr, o_dacv, o_shrst, o_hold, o_dac1, o_daci_sel, o_dat, 
        r_dac_en, r_sar_en, o_dactl, o_cmpsta, x_daclsb, o_intr, o_smpl, 
        test_si2, test_si1, test_so1, test_se );
  input [2:0] r_comp_opt;
  input [7:0] r_wdat;
  output [7:0] r_adofs;
  output [7:0] r_isofs;
  input [10:0] r_wr;
  input [17:0] dacv_wr;
  output [143:0] o_dacv;
  output [9:0] o_dac1;
  output [17:0] o_daci_sel;
  output [17:0] o_dat;
  output [17:0] r_dac_en;
  output [17:0] r_sar_en;
  output [7:0] o_dactl;
  output [7:0] o_cmpsta;
  output [5:0] x_daclsb;
  output [4:0] o_smpl;
  input clk, srstz, i_comp, test_si2, test_si1, test_se;
  output o_shrst, o_hold, o_intr, test_so1;
  wire   dacyc_done, updcmp, semi_start, sacyc_done, sar_ini, sar_nxt,
         sampl_begn, sampl_done, ps_md4ch, ps_sample, updlsb, wda_6_, N1239,
         N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1250, N1251,
         N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1261, N1262, N1263,
         N1264, N1265, N1266, N1267, N1268, N1269, N1272, N1273, N1274, N1275,
         N1276, N1277, N1278, N1279, N1280, N1283, N1284, N1285, N1286, N1287,
         N1288, N1289, N1290, N1291, N1294, N1295, N1296, N1297, N1298, N1299,
         N1300, N1301, N1302, N1305, N1306, N1307, N1308, N1309, N1310, N1311,
         N1312, N1313, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323,
         N1324, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335,
         N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1349,
         N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1360, N1361,
         N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1371, N1372, N1373,
         N1374, N1375, N1376, N1377, N1378, N1379, N1382, N1383, N1384, N1385,
         N1386, N1387, N1388, N1389, N1390, N1393, N1394, N1395, N1396, N1397,
         N1398, N1399, N1400, N1401, N1404, N1405, N1406, N1407, N1408, N1409,
         N1410, N1411, N1412, N1415, N1416, N1417, N1418, N1419, N1420, N1421,
         N1422, N1423, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433,
         N1434, n544, n536, n538, n537, n540, n541, n539, n85, n87, n535, n141,
         n142, n143, n144, n145, n146, n147, n148, n151, n153, n154, n155,
         n156, n157, n158, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n542, n543, n65, n88, n89,
         n90, n130, n131, n132, n133, n134, n136, n139, n140, n149, n150, n152,
         n159, n160, n176, n177, n178, n179, n181, n182, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n210, n211, n212,
         n214, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n301, n302, n303, n305, n306, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n327, n330, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n411, n412, n413, n414, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n86, n92, n94, n96, n98, n100, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n113, n114, n115, n116, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n135, n137, n138, n180, n183, n197, n198, n199, n209, n213, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n300, n304, n307, n308,
         n309, n310, n311, n312, n326, n328, n329, n331, n410, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n435, n436,
         n437, n438, n439, n440, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534;
  wire   [1:0] syn_comp;
  wire   [4:0] cs_ptr;
  wire   [17:0] datcmp;
  wire   [4:0] ps_ptr;
  wire   [9:0] r_dac1v;
  wire   [9:0] r_rpt_v;
  wire   [17:0] app_dacis;
  wire   [17:0] pos_dacis;
  wire   [5:0] wdlsb;
  wire   [17:0] upd;
  wire   [143:0] r_dacvs;
  wire   [7:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;

  INVX1 U126 ( .A(n173), .Y(n172) );
  INVX1 U127 ( .A(n173), .Y(n166) );
  INVX1 U128 ( .A(n173), .Y(n165) );
  INVX1 U129 ( .A(n174), .Y(n164) );
  INVX1 U130 ( .A(n175), .Y(n163) );
  INVX1 U131 ( .A(n175), .Y(n162) );
  INVX1 U132 ( .A(n174), .Y(n161) );
  INVX1 U133 ( .A(n173), .Y(n158) );
  INVX1 U134 ( .A(n174), .Y(n156) );
  INVX1 U135 ( .A(n174), .Y(n155) );
  INVX1 U136 ( .A(n175), .Y(n154) );
  INVX1 U137 ( .A(n173), .Y(n153) );
  INVX1 U138 ( .A(n174), .Y(n151) );
  INVX1 U139 ( .A(n175), .Y(n148) );
  INVX1 U140 ( .A(n174), .Y(n147) );
  INVX1 U141 ( .A(n174), .Y(n146) );
  INVX1 U142 ( .A(n175), .Y(n145) );
  INVX1 U143 ( .A(n175), .Y(n144) );
  INVX1 U144 ( .A(n175), .Y(n157) );
  INVX1 U145 ( .A(n175), .Y(n143) );
  INVX1 U146 ( .A(n174), .Y(n170) );
  INVX1 U147 ( .A(n174), .Y(n169) );
  INVX1 U148 ( .A(n174), .Y(n168) );
  INVX1 U149 ( .A(n173), .Y(n167) );
  INVX1 U150 ( .A(n175), .Y(n142) );
  INVX1 U151 ( .A(n173), .Y(n171) );
  INVX1 U154 ( .A(srstz), .Y(n173) );
  INVX1 U178 ( .A(n175), .Y(n141) );
  INVX1 U179 ( .A(srstz), .Y(n175) );
  INVX1 U180 ( .A(srstz), .Y(n174) );
  glreg_00000012 u0_compi ( .clk(clk), .arstz(n163), .we(updcmp), .wdat(datcmp), .rdat(o_dat), .test_si(o_cmpsta[7]), .test_se(test_se) );
  dac2sar_a0 u0_dac2sar ( .r_dac_t(o_dactl[3:2]), .r_dacyc(o_dactl[7]), 
        .r_sar10(n65), .sar_ini(sar_ini), .sar_nxt(sar_nxt), .semi_nxt(n88), 
        .auto_sar(n456), .busy(o_dactl[0]), .stop(n71), .sync_i(syn_comp[1]), 
        .sampl_begn(sampl_begn), .sampl_done(sampl_done), .sh_rst(o_shrst), 
        .dacyc_done(dacyc_done), .sacyc_done(sacyc_done), .dac_v(r_dac1v), 
        .rpt_v(r_rpt_v), .clk(clk), .srstz(srstz), .test_si2(o_dat[17]), 
        .test_si1(test_si1), .test_so1(n543), .test_se(test_se) );
  shmux_00000005_00000012_00000012 u0_shmux ( .ps_sample(ps_sample), 
        .ps_md4ch(ps_md4ch), .r_comp_swtch(r_comp_opt[2]), .r_semi(n90), 
        .r_loop(o_dactl[1]), .r_dac_en(r_dac_en), .wr_dacv(dacv_wr), .busy(
        o_dactl[0]), .sh_hold(o_hold), .stop(n71), .semi_start(semi_start), 
        .auto_start(n457), .mxcyc_done(n87), .sampl_begn(sampl_begn), 
        .sampl_done(sampl_done), .app_dacis(app_dacis), .pos_dacis(pos_dacis), 
        .cs_ptr(cs_ptr), .ps_ptr(ps_ptr), .clk(clk), .srstz(n171), .test_si2(
        r_sar_en[7]), .test_si1(o_shrst), .test_so1(test_so1), .test_se(
        test_se) );
  glreg_WIDTH7_1 u0_dactl ( .clk(clk), .arstz(n171), .we(n89), .wdat({
        r_wdat[7], n8, n10, n6, r_wdat[3], n4, n60}), .rdat(o_dactl[7:1]), 
        .test_si(x_daclsb[5]), .test_se(test_se) );
  glreg_a0_48 u0_dacen ( .clk(clk), .arstz(n141), .we(r_wr[1]), .wdat({
        r_wdat[7], n8, r_wdat[5], n6, r_wdat[3], n4, n60, n78}), .rdat(
        r_dac_en[7:0]), .test_si(n543), .test_se(test_se) );
  glreg_a0_47 u0_saren ( .clk(clk), .arstz(n142), .we(r_wr[2]), .wdat({
        r_wdat[7], n8, n10, n6, r_wdat[3], n4, r_wdat[1], n78}), .rdat(
        r_sar_en[7:0]), .test_si(r_isofs[7]), .test_se(test_se) );
  glreg_WIDTH6_2 u0_daclsb ( .clk(clk), .arstz(n172), .we(updlsb), .wdat(wdlsb), .rdat(x_daclsb), .test_si(r_dac_en[7]), .test_se(test_se) );
  glreg_a0_46 dacvs_0__u0 ( .clk(clk), .arstz(n143), .we(upd[0]), .wdat({n59, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[7:0]), .test_si(
        test_si2), .test_se(test_se) );
  glreg_a0_45 dacvs_1__u0 ( .clk(clk), .arstz(n157), .we(upd[1]), .wdat({n58, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[15:8]), .test_si(
        r_dacvs[7]), .test_se(test_se) );
  glreg_a0_44 dacvs_2__u0 ( .clk(clk), .arstz(n144), .we(upd[2]), .wdat({n59, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[23:16]), .test_si(
        r_dacvs[15]), .test_se(test_se) );
  glreg_a0_43 dacvs_3__u0 ( .clk(clk), .arstz(n145), .we(upd[3]), .wdat({n59, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[31:24]), .test_si(
        r_dacvs[23]), .test_se(test_se) );
  glreg_a0_42 dacvs_4__u0 ( .clk(clk), .arstz(n146), .we(upd[4]), .wdat({n58, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[39:32]), .test_si(
        r_dacvs[31]), .test_se(test_se) );
  glreg_a0_41 dacvs_5__u0 ( .clk(clk), .arstz(n147), .we(upd[5]), .wdat({n58, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[47:40]), .test_si(
        r_dacvs[39]), .test_se(test_se) );
  glreg_a0_40 dacvs_6__u0 ( .clk(clk), .arstz(n148), .we(upd[6]), .wdat({n59, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[55:48]), .test_si(
        r_dacvs[47]), .test_se(test_se) );
  glreg_a0_39 dacvs_7__u0 ( .clk(clk), .arstz(n151), .we(upd[7]), .wdat({n58, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[63:56]), .test_si(
        r_dacvs[55]), .test_se(test_se) );
  glreg_a0_38 dacvs_8__u0 ( .clk(clk), .arstz(n153), .we(upd[8]), .wdat({n58, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[71:64]), .test_si(
        r_dacvs[63]), .test_se(test_se) );
  glreg_a0_37 dacvs_9__u0 ( .clk(clk), .arstz(n154), .we(upd[9]), .wdat({n59, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[79:72]), .test_si(
        r_dacvs[71]), .test_se(test_se) );
  glreg_a0_36 dacvs_10__u0 ( .clk(clk), .arstz(n155), .we(upd[10]), .wdat({n59, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[87:80]), .test_si(
        r_dacvs[79]), .test_se(test_se) );
  glreg_a0_35 dacvs_11__u0 ( .clk(clk), .arstz(n156), .we(upd[11]), .wdat({n58, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[95:88]), .test_si(
        r_dacvs[87]), .test_se(test_se) );
  glreg_a0_34 dacvs_12__u0 ( .clk(clk), .arstz(n158), .we(upd[12]), .wdat({n59, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[103:96]), .test_si(
        r_dacvs[95]), .test_se(test_se) );
  glreg_a0_33 dacvs_13__u0 ( .clk(clk), .arstz(n161), .we(upd[13]), .wdat({n59, 
        n16, n18, n38, n41, n48, n52, n44}), .rdat(r_dacvs[111:104]), 
        .test_si(r_dacvs[103]), .test_se(test_se) );
  glreg_a0_32 dacvs_14__u0 ( .clk(clk), .arstz(n162), .we(upd[14]), .wdat({n58, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[119:112]), 
        .test_si(r_dacvs[111]), .test_se(test_se) );
  glreg_a0_31 dacvs_15__u0 ( .clk(clk), .arstz(n163), .we(upd[15]), .wdat({n59, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[127:120]), 
        .test_si(r_dacvs[119]), .test_se(test_se) );
  glreg_a0_30 dacvs_16__u0 ( .clk(clk), .arstz(n164), .we(upd[16]), .wdat({n58, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[135:128]), 
        .test_si(r_dacvs[127]), .test_se(test_se) );
  glreg_a0_29 dacvs_17__u0 ( .clk(clk), .arstz(n165), .we(upd[17]), .wdat({n58, 
        n15, n17, n19, n40, n47, n51, n43}), .rdat(r_dacvs[143:136]), 
        .test_si(r_dacvs[135]), .test_se(test_se) );
  glsta_a0_1 u0_cmpsta ( .clk(clk), .arstz(n166), .rst0(1'b0), .set2(setsta), 
        .clr1(clrsta), .rdat(o_cmpsta), .irq(r_irq), .test_si(r_adofs[7]), 
        .test_se(test_se) );
  glreg_a0_28 u0_adofs ( .clk(clk), .arstz(n167), .we(r_wr[5]), .wdat({
        r_wdat[7], n8, n10, n6, r_wdat[3], n4, n60, n14}), .rdat({n535, n536, 
        n537, n538, n539, n540, n541, n544}), .test_si(syn_comp[1]), .test_se(
        test_se) );
  glreg_a0_27 u0_isofs ( .clk(clk), .arstz(n168), .we(r_wr[6]), .wdat({
        r_wdat[7], n8, n10, n6, r_wdat[3], n4, n60, n78}), .rdat(r_isofs), 
        .test_si(o_dactl[7]), .test_se(test_se) );
  glreg_a0_26 u1_dacen ( .clk(clk), .arstz(n169), .we(r_wr[7]), .wdat({
        r_wdat[7], n8, n10, n6, r_wdat[3], n4, n60, n78}), .rdat(
        r_dac_en[15:8]), .test_si(pos_dacis[17]), .test_se(test_se) );
  glreg_a0_25 u1_saren ( .clk(clk), .arstz(n170), .we(r_wr[8]), .wdat({
        r_wdat[7], n8, n10, n6, r_wdat[3], n4, r_wdat[1], n78}), .rdat(
        r_sar_en[15:8]), .test_si(r_dac_en[15]), .test_se(test_se) );
  glreg_WIDTH2_1 u2_dacen ( .clk(clk), .arstz(n172), .we(r_wr[9]), .wdat({n60, 
        n14}), .rdat(r_dac_en[17:16]), .test_si(r_sar_en[15]), .test_so(n542), 
        .test_se(test_se) );
  glreg_WIDTH2_0 u2_saren ( .clk(clk), .arstz(n172), .we(r_wr[10]), .wdat({n60, 
        n78}), .rdat(r_sar_en[17:16]), .test_si(n542), .test_se(test_se) );
  dacmux_a0_DW01_add_0 add_230_I18 ( .A({1'b0, r_dacvs[143:136]}), .B({
        r_adofs[7], n114, n100, n98, n96, n94, n92, n86, r_adofs[0]}), .CI(
        1'b0), .SUM({N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, 
        N1426}), .CO() );
  dacmux_a0_DW01_add_1 add_230_I17 ( .A({1'b0, r_dacvs[135:128]}), .B({
        r_adofs[7], n114, r_adofs[6:0]}), .CI(1'b0), .SUM({N1423, N1422, N1421, 
        N1420, N1419, N1418, N1417, N1416, N1415}), .CO() );
  dacmux_a0_DW01_add_2 add_230_I16 ( .A({1'b0, r_dacvs[127:120]}), .B({n116, 
        n114, n100, n98, n96, n94, n92, n86, n111}), .CI(1'b0), .SUM({N1412, 
        N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404}), .CO() );
  dacmux_a0_DW01_add_3 add_230_I15 ( .A({1'b0, r_dacvs[119:112]}), .B({n116, 
        n114, r_adofs[6:1], n111}), .CI(1'b0), .SUM({N1401, N1400, N1399, 
        N1398, N1397, N1396, N1395, N1394, N1393}), .CO() );
  dacmux_a0_DW01_add_4 add_230_I14 ( .A({1'b0, r_dacvs[111:104]}), .B({n116, 
        n114, n100, n98, n96, n94, n92, n86, n111}), .CI(1'b0), .SUM({N1390, 
        N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382}), .CO() );
  dacmux_a0_DW01_add_5 add_230_I13 ( .A({1'b0, r_dacvs[103:96]}), .B({n116, 
        n114, r_adofs[6:1], n111}), .CI(1'b0), .SUM({N1379, N1378, N1377, 
        N1376, N1375, N1374, N1373, N1372, N1371}), .CO() );
  dacmux_a0_DW01_add_6 add_230_I12 ( .A({1'b0, r_dacvs[95:88]}), .B({n116, 
        n114, n100, n98, n96, n94, n92, n86, n111}), .CI(1'b0), .SUM({N1368, 
        N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360}), .CO() );
  dacmux_a0_DW01_add_7 add_230_I11 ( .A({1'b0, r_dacvs[87:80]}), .B({n116, 
        n114, r_adofs[6:1], n110}), .CI(1'b0), .SUM({N1357, N1356, N1355, 
        N1354, N1353, N1352, N1351, N1350, N1349}), .CO() );
  dacmux_a0_DW01_add_8 add_230_I10 ( .A({1'b0, r_dacvs[79:72]}), .B({n115, 
        n114, n100, n98, n96, n94, n92, n86, n110}), .CI(1'b0), .SUM({N1346, 
        N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338}), .CO() );
  dacmux_a0_DW01_add_9 add_230_I9 ( .A({1'b0, r_dacvs[71:64]}), .B({n115, n114, 
        r_adofs[6:1], n110}), .CI(1'b0), .SUM({N1335, N1334, N1333, N1332, 
        N1331, N1330, N1329, N1328, N1327}), .CO() );
  dacmux_a0_DW01_add_10 add_230_I8 ( .A({1'b0, r_dacvs[63:56]}), .B({n115, 
        n115, n100, n98, n96, n94, n92, n86, n110}), .CI(1'b0), .SUM({N1324, 
        N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316}), .CO() );
  dacmux_a0_DW01_add_11 add_230_I7 ( .A({1'b0, r_dacvs[55:48]}), .B({n116, 
        n115, r_adofs[6:1], n110}), .CI(1'b0), .SUM({N1313, N1312, N1311, 
        N1310, N1309, N1308, N1307, N1306, N1305}), .CO() );
  dacmux_a0_DW01_add_12 add_230_I6 ( .A({1'b0, r_dacvs[47:40]}), .B({n116, 
        n115, n100, n98, n96, n94, n92, n86, r_adofs[0]}), .CI(1'b0), .SUM({
        N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294}), .CO()
         );
  dacmux_a0_DW01_add_13 add_230_I5 ( .A({1'b0, r_dacvs[39:32]}), .B({n116, 
        n115, r_adofs[6:0]}), .CI(1'b0), .SUM({N1291, N1290, N1289, N1288, 
        N1287, N1286, N1285, N1284, N1283}), .CO() );
  dacmux_a0_DW01_add_14 add_230_I4 ( .A({1'b0, r_dacvs[31:24]}), .B({
        r_adofs[7], n115, n100, n98, n96, n94, n92, n86, n544}), .CI(1'b0), 
        .SUM({N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272}), 
        .CO() );
  dacmux_a0_DW01_add_15 add_230_I3 ( .A({1'b0, r_dacvs[23:16]}), .B({
        r_isofs[7], r_isofs}), .CI(1'b0), .SUM({N1269, N1268, N1267, N1266, 
        N1265, N1264, N1263, N1262, N1261}), .CO() );
  dacmux_a0_DW01_add_16 add_230_I2 ( .A({1'b0, r_dacvs[15:8]}), .B({n116, n115, 
        r_adofs[6:1], n544}), .CI(1'b0), .SUM({N1258, N1257, N1256, N1255, 
        N1254, N1253, N1252, N1251, N1250}), .CO() );
  dacmux_a0_DW01_add_17 add_230 ( .A({1'b0, r_dacvs[7:0]}), .B({r_adofs[7], 
        n115, n100, n98, n96, n94, n92, n86, n544}), .CI(1'b0), .SUM({N1247, 
        N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239}), .CO() );
  SDFFQX1 syn_comp_reg_1_ ( .D(syn_comp[0]), .SIN(syn_comp[0]), .SMC(test_se), 
        .C(clk), .Q(syn_comp[1]) );
  SDFFQX1 syn_comp_reg_0_ ( .D(i_comp), .SIN(r_dacvs[143]), .SMC(test_se), .C(
        clk), .Q(syn_comp[0]) );
  NAND32X2 U21 ( .B(n90), .C(n71), .A(n89), .Y(n135) );
  AO21X4 U22 ( .B(r_wr[0]), .C(n220), .A(n71), .Y(n89) );
  NAND21XL U23 ( .B(ps_ptr[1]), .A(ps_ptr[2]), .Y(n230) );
  BUFX6 U24 ( .A(n72), .Y(n1) );
  NOR2XL U25 ( .A(n227), .B(n73), .Y(n72) );
  NAND21X1 U26 ( .B(ps_ptr[2]), .A(n227), .Y(n228) );
  INVX1 U27 ( .A(n228), .Y(n241) );
  INVX2 U28 ( .A(n229), .Y(n240) );
  INVX1 U29 ( .A(n230), .Y(n242) );
  INVX2 U30 ( .A(n135), .Y(n457) );
  BUFX3 U31 ( .A(r_wdat[1]), .Y(n60) );
  AND3X1 U32 ( .A(n497), .B(n498), .C(n503), .Y(n2) );
  INVXL U33 ( .A(r_wdat[2]), .Y(n3) );
  INVXL U34 ( .A(n3), .Y(n4) );
  INVXL U35 ( .A(r_wdat[4]), .Y(n5) );
  INVXL U36 ( .A(n5), .Y(n6) );
  INVXL U37 ( .A(r_wdat[6]), .Y(n7) );
  INVXL U38 ( .A(n7), .Y(n8) );
  INVXL U39 ( .A(r_wdat[5]), .Y(n9) );
  INVXL U40 ( .A(n9), .Y(n10) );
  INVXL U41 ( .A(n409), .Y(n11) );
  INVXL U42 ( .A(n409), .Y(n12) );
  INVXL U43 ( .A(n78), .Y(n13) );
  INVXL U44 ( .A(n13), .Y(n14) );
  BUFX3 U45 ( .A(n312), .Y(wda_6_) );
  INVX1 U46 ( .A(wda_6_), .Y(n15) );
  INVX1 U47 ( .A(wda_6_), .Y(n16) );
  BUFX3 U48 ( .A(n326), .Y(n455) );
  INVX1 U49 ( .A(n455), .Y(n17) );
  INVX1 U50 ( .A(n455), .Y(n18) );
  BUFX3 U51 ( .A(n328), .Y(n454) );
  INVX1 U52 ( .A(n454), .Y(n19) );
  INVX1 U53 ( .A(n454), .Y(n38) );
  INVX1 U54 ( .A(n491), .Y(n39) );
  BUFX3 U55 ( .A(n331), .Y(n453) );
  INVX1 U56 ( .A(n453), .Y(n40) );
  INVX1 U57 ( .A(n453), .Y(n41) );
  NOR2X1 U58 ( .A(n179), .B(n106), .Y(n42) );
  BUFX3 U59 ( .A(n417), .Y(n451) );
  INVX1 U60 ( .A(n451), .Y(n43) );
  INVX1 U61 ( .A(n451), .Y(n44) );
  INVX1 U62 ( .A(n460), .Y(n45) );
  NOR2X1 U63 ( .A(n108), .B(n179), .Y(n46) );
  BUFX3 U64 ( .A(n410), .Y(n452) );
  INVX1 U65 ( .A(n452), .Y(n47) );
  INVX1 U66 ( .A(n452), .Y(n48) );
  BUFX3 U67 ( .A(n334), .Y(n49) );
  NOR2X1 U68 ( .A(n108), .B(n136), .Y(n50) );
  BUFX3 U69 ( .A(n416), .Y(n85) );
  INVX1 U70 ( .A(n85), .Y(n51) );
  INVX1 U71 ( .A(n85), .Y(n52) );
  INVX1 U72 ( .A(n490), .Y(n53) );
  AO21X4 U73 ( .B(n308), .C(n309), .A(n307), .Y(sar_ini) );
  BUFX3 U74 ( .A(n332), .Y(n54) );
  NOR2X1 U75 ( .A(o_dactl[0]), .B(semi_start), .Y(n462) );
  INVX1 U76 ( .A(n462), .Y(n55) );
  INVX1 U77 ( .A(n462), .Y(n56) );
  NOR2X1 U78 ( .A(n108), .B(n159), .Y(n57) );
  MUX2IX1 U79 ( .D0(r_rpt_v[9]), .D1(r_wdat[7]), .S(n130), .Y(n68) );
  INVX1 U80 ( .A(n68), .Y(n58) );
  INVX1 U81 ( .A(n68), .Y(n59) );
  NAND3X1 U82 ( .A(cs_ptr[4]), .B(n107), .C(n492), .Y(n333) );
  INVX1 U83 ( .A(n333), .Y(n61) );
  INVX1 U84 ( .A(n333), .Y(n62) );
  NOR2X1 U85 ( .A(n136), .B(n106), .Y(n63) );
  NOR2X1 U86 ( .A(n108), .B(n149), .Y(n64) );
  INVX1 U87 ( .A(n424), .Y(n66) );
  INVX1 U88 ( .A(r_wr[0]), .Y(n67) );
  INVXL U89 ( .A(dacv_wr[13]), .Y(n423) );
  INVXL U90 ( .A(dacv_wr[14]), .Y(n422) );
  INVXL U91 ( .A(dacv_wr[9]), .Y(n437) );
  INVXL U92 ( .A(dacv_wr[17]), .Y(n311) );
  INVXL U93 ( .A(dacv_wr[10]), .Y(n436) );
  INVXL U94 ( .A(ps_ptr[2]), .Y(n73) );
  NOR2X2 U95 ( .A(r_wdat[0]), .B(n67), .Y(n71) );
  NAND21XL U96 ( .B(n307), .A(n225), .Y(semi_start) );
  AND2XL U97 ( .A(r_wr[4]), .B(r_wdat[7]), .Y(clrsta[7]) );
  INVXL U98 ( .A(n221), .Y(n223) );
  OAI222XL U99 ( .A(n202), .B(n495), .C(n203), .D(n496), .E(cs_ptr[4]), .F(
        n426), .Y(n133) );
  INVX1 U100 ( .A(n520), .Y(n491) );
  INVX1 U101 ( .A(dacv_wr[5]), .Y(n458) );
  INVX1 U102 ( .A(dacv_wr[4]), .Y(n459) );
  INVX1 U103 ( .A(dacv_wr[7]), .Y(n439) );
  INVX1 U104 ( .A(dacv_wr[6]), .Y(n440) );
  NAND21X1 U105 ( .B(n106), .A(n104), .Y(n520) );
  NAND2X1 U106 ( .A(n106), .B(n104), .Y(n184) );
  INVX1 U107 ( .A(n519), .Y(n490) );
  NAND21X1 U108 ( .B(n104), .A(n70), .Y(n152) );
  NAND21X1 U109 ( .B(n104), .A(n69), .Y(n182) );
  INVX1 U110 ( .A(ps_ptr[1]), .Y(n227) );
  INVX1 U111 ( .A(dacv_wr[16]), .Y(n419) );
  INVXL U112 ( .A(dacv_wr[8]), .Y(n438) );
  INVX1 U113 ( .A(dacv_wr[15]), .Y(n421) );
  INVXL U114 ( .A(dacv_wr[11]), .Y(n435) );
  INVXL U115 ( .A(dacv_wr[12]), .Y(n425) );
  AND2X1 U116 ( .A(r_wr[4]), .B(n14), .Y(clrsta[0]) );
  NAND21X1 U117 ( .B(n104), .A(n107), .Y(n519) );
  INVX1 U118 ( .A(n105), .Y(n104) );
  INVX1 U119 ( .A(n107), .Y(n106) );
  NAND2X1 U120 ( .A(n106), .B(n105), .Y(n186) );
  NOR2X1 U121 ( .A(n105), .B(n12), .Y(n318) );
  NOR2X1 U122 ( .A(n11), .B(n104), .Y(n320) );
  NOR2X1 U123 ( .A(n108), .B(n136), .Y(n69) );
  NOR2X1 U124 ( .A(n108), .B(n159), .Y(n70) );
  NOR2X1 U125 ( .A(n159), .B(n106), .Y(n334) );
  NOR2X1 U152 ( .A(n136), .B(n106), .Y(n330) );
  NAND21X1 U153 ( .B(n105), .A(n57), .Y(n150) );
  NAND21X1 U155 ( .B(n105), .A(n75), .Y(n139) );
  NAND21X1 U156 ( .B(n104), .A(n64), .Y(n140) );
  NAND21X1 U157 ( .B(n105), .A(n74), .Y(n177) );
  NAND21X1 U158 ( .B(n105), .A(n50), .Y(n181) );
  NAND21X1 U159 ( .B(n104), .A(n46), .Y(n178) );
  NAND21XL U160 ( .B(ps_ptr[2]), .A(ps_ptr[1]), .Y(n229) );
  INVX1 U161 ( .A(n60), .Y(n415) );
  INVX1 U162 ( .A(r_wdat[3]), .Y(n329) );
  INVX1 U163 ( .A(n226), .Y(n87) );
  INVX1 U164 ( .A(N1346), .Y(n505) );
  INVX1 U165 ( .A(N1335), .Y(n504) );
  OAI22AX1 U166 ( .D(dacv_wr[1]), .C(n56), .A(n159), .B(n461), .Y(upd[1]) );
  OAI22AX1 U167 ( .D(dacv_wr[0]), .C(n56), .A(n159), .B(n463), .Y(upd[0]) );
  OAI22X1 U168 ( .A(n149), .B(n461), .C(n458), .D(n55), .Y(upd[5]) );
  OAI22X1 U169 ( .A(n149), .B(n463), .C(n459), .D(n55), .Y(upd[4]) );
  OAI22X1 U170 ( .A(n136), .B(n463), .C(n438), .D(n55), .Y(upd[8]) );
  OAI22X1 U171 ( .A(n179), .B(n461), .C(n423), .D(n55), .Y(upd[13]) );
  OAI22X1 U172 ( .A(n179), .B(n463), .C(n425), .D(n55), .Y(upd[12]) );
  OAI22X1 U173 ( .A(n136), .B(n461), .C(n437), .D(n55), .Y(upd[9]) );
  OAI22X1 U174 ( .A(n311), .B(n55), .C(n160), .D(n130), .Y(upd[17]) );
  OAI22X1 U175 ( .A(n419), .B(n55), .C(n176), .D(n130), .Y(upd[16]) );
  OAI22X1 U176 ( .A(n421), .B(n56), .C(n177), .D(n66), .Y(upd[15]) );
  OAI22X1 U177 ( .A(n422), .B(n56), .C(n178), .D(n66), .Y(upd[14]) );
  OAI22X1 U181 ( .A(n435), .B(n56), .C(n181), .D(n66), .Y(upd[11]) );
  OAI22X1 U182 ( .A(n436), .B(n56), .C(n182), .D(n66), .Y(upd[10]) );
  OAI22X1 U183 ( .A(n439), .B(n56), .C(n139), .D(n66), .Y(upd[7]) );
  OAI22X1 U184 ( .A(n440), .B(n56), .C(n140), .D(n66), .Y(upd[6]) );
  OAI22AX1 U185 ( .D(dacv_wr[3]), .C(n56), .A(n150), .B(n66), .Y(upd[3]) );
  OAI22AX1 U186 ( .D(dacv_wr[2]), .C(n56), .A(n152), .B(n66), .Y(upd[2]) );
  INVX1 U187 ( .A(n225), .Y(n88) );
  INVX1 U188 ( .A(N1423), .Y(n512) );
  INVX1 U189 ( .A(N1434), .Y(n513) );
  INVX1 U190 ( .A(N1379), .Y(n508) );
  INVX1 U191 ( .A(N1412), .Y(n511) );
  INVX1 U192 ( .A(N1368), .Y(n507) );
  INVX1 U193 ( .A(N1357), .Y(n506) );
  INVX1 U194 ( .A(N1401), .Y(n510) );
  INVX1 U195 ( .A(N1390), .Y(n509) );
  INVX1 U196 ( .A(N1280), .Y(n475) );
  INVX1 U197 ( .A(N1247), .Y(n466) );
  INVX1 U198 ( .A(N1324), .Y(n487) );
  INVX1 U199 ( .A(N1291), .Y(n478) );
  INVX1 U200 ( .A(N1302), .Y(n481) );
  INVX1 U201 ( .A(N1258), .Y(n469) );
  INVX1 U202 ( .A(N1313), .Y(n484) );
  INVX1 U203 ( .A(n473), .Y(n474) );
  NAND21X1 U204 ( .B(n535), .A(N1280), .Y(n473) );
  INVX1 U205 ( .A(n464), .Y(n465) );
  NAND21X1 U206 ( .B(n535), .A(N1247), .Y(n464) );
  INVX1 U207 ( .A(n485), .Y(n486) );
  NAND21X1 U208 ( .B(r_adofs[7]), .A(N1324), .Y(n485) );
  INVX1 U209 ( .A(n476), .Y(n477) );
  NAND21X1 U210 ( .B(r_adofs[7]), .A(N1291), .Y(n476) );
  INVX1 U211 ( .A(n479), .Y(n480) );
  NAND21X1 U212 ( .B(r_adofs[7]), .A(N1302), .Y(n479) );
  INVX1 U213 ( .A(n467), .Y(n468) );
  NAND21X1 U214 ( .B(n535), .A(N1258), .Y(n467) );
  AND2X1 U215 ( .A(r_wr[4]), .B(n10), .Y(clrsta[5]) );
  AND2X1 U216 ( .A(r_wr[4]), .B(n4), .Y(clrsta[2]) );
  AND2X1 U217 ( .A(n60), .B(r_wr[4]), .Y(clrsta[1]) );
  AND2X1 U218 ( .A(r_wr[4]), .B(n8), .Y(clrsta[6]) );
  AND2X1 U219 ( .A(n6), .B(r_wr[4]), .Y(clrsta[4]) );
  AND2X1 U220 ( .A(r_wr[4]), .B(r_wdat[3]), .Y(clrsta[3]) );
  INVX1 U221 ( .A(cs_ptr[1]), .Y(n107) );
  INVX1 U222 ( .A(cs_ptr[0]), .Y(n105) );
  INVX1 U223 ( .A(dacyc_done), .Y(n518) );
  NOR2X1 U224 ( .A(n520), .B(n185), .Y(setsta[5]) );
  NOR2X1 U225 ( .A(n520), .B(n188), .Y(setsta[1]) );
  NOR2X1 U226 ( .A(n186), .B(n185), .Y(setsta[6]) );
  NOR2X1 U227 ( .A(n519), .B(n188), .Y(setsta[0]) );
  NOR2X1 U228 ( .A(n186), .B(n188), .Y(setsta[2]) );
  NAND2X1 U229 ( .A(cs_ptr[4]), .B(n105), .Y(n203) );
  NAND2X1 U230 ( .A(cs_ptr[4]), .B(n104), .Y(n202) );
  NOR2X1 U231 ( .A(n519), .B(n185), .Y(setsta[4]) );
  NAND21X1 U232 ( .B(cs_ptr[4]), .A(n488), .Y(n136) );
  NOR2X1 U233 ( .A(n179), .B(n106), .Y(n327) );
  NOR2X1 U234 ( .A(n184), .B(n185), .Y(setsta[7]) );
  NOR2X1 U235 ( .A(n184), .B(n188), .Y(setsta[3]) );
  NAND21X1 U236 ( .B(cs_ptr[4]), .A(n492), .Y(n159) );
  INVX1 U237 ( .A(n424), .Y(n130) );
  NAND21X1 U238 ( .B(n520), .A(n424), .Y(n461) );
  NAND21X1 U239 ( .B(n519), .A(n424), .Y(n463) );
  NOR2X1 U240 ( .A(n108), .B(n179), .Y(n74) );
  NOR2X1 U241 ( .A(n108), .B(n149), .Y(n75) );
  NOR2X1 U242 ( .A(n149), .B(n106), .Y(n332) );
  INVX1 U243 ( .A(cs_ptr[1]), .Y(n108) );
  NAND21X1 U244 ( .B(n520), .A(n418), .Y(n160) );
  NAND21X1 U245 ( .B(n519), .A(n418), .Y(n176) );
  AO21X1 U246 ( .B(N1265), .C(n472), .A(n471), .Y(o_dacv[20]) );
  AO21X1 U247 ( .B(N1251), .C(n469), .A(n468), .Y(o_dacv[9]) );
  AO21X1 U248 ( .B(N1263), .C(n472), .A(n471), .Y(o_dacv[18]) );
  AO21X1 U249 ( .B(N1243), .C(n466), .A(n465), .Y(o_dacv[4]) );
  AO21X1 U250 ( .B(N1242), .C(n466), .A(n465), .Y(o_dacv[3]) );
  AO21X1 U251 ( .B(N1245), .C(n466), .A(n465), .Y(o_dacv[6]) );
  AO21X1 U252 ( .B(N1246), .C(n466), .A(n465), .Y(o_dacv[7]) );
  AO21X1 U253 ( .B(N1244), .C(n466), .A(n465), .Y(o_dacv[5]) );
  AO21X1 U254 ( .B(N1240), .C(n466), .A(n465), .Y(o_dacv[1]) );
  AO21X1 U255 ( .B(N1241), .C(n466), .A(n465), .Y(o_dacv[2]) );
  AO21X1 U256 ( .B(N1266), .C(n472), .A(n471), .Y(o_dacv[21]) );
  AO21X1 U257 ( .B(N1262), .C(n472), .A(n471), .Y(o_dacv[17]) );
  AO21X1 U258 ( .B(N1264), .C(n472), .A(n471), .Y(o_dacv[19]) );
  AO21X1 U259 ( .B(N1261), .C(n472), .A(n471), .Y(o_dacv[16]) );
  AO21X1 U260 ( .B(N1267), .C(n472), .A(n471), .Y(o_dacv[22]) );
  AO21X1 U261 ( .B(N1268), .C(n472), .A(n471), .Y(o_dacv[23]) );
  INVX1 U262 ( .A(n222), .Y(n307) );
  NAND6XL U263 ( .A(r_wdat[6]), .B(n14), .C(n223), .D(n3), .E(n329), .F(n9), 
        .Y(n222) );
  NAND6XL U264 ( .A(n10), .B(r_wdat[3]), .C(n4), .D(n223), .E(n13), .F(n7), 
        .Y(n225) );
  INVX1 U265 ( .A(n113), .Y(n110) );
  INVX1 U266 ( .A(n113), .Y(n111) );
  NAND2X1 U267 ( .A(N1346), .B(n118), .Y(n305) );
  NAND2X1 U268 ( .A(N1335), .B(n118), .Y(n306) );
  NAND2X1 U269 ( .A(N1412), .B(n118), .Y(n315) );
  AO21X1 U270 ( .B(N1275), .C(n475), .A(n474), .Y(o_dacv[27]) );
  AO21X1 U271 ( .B(N1299), .C(n481), .A(n480), .Y(o_dacv[45]) );
  AO21X1 U272 ( .B(N1278), .C(n475), .A(n474), .Y(o_dacv[30]) );
  AO21X1 U273 ( .B(N1300), .C(n481), .A(n480), .Y(o_dacv[46]) );
  AO21X1 U274 ( .B(N1279), .C(n475), .A(n474), .Y(o_dacv[31]) );
  AO21X1 U275 ( .B(N1253), .C(n469), .A(n468), .Y(o_dacv[11]) );
  AO21X1 U276 ( .B(N1257), .C(n469), .A(n468), .Y(o_dacv[15]) );
  AO21X1 U277 ( .B(N1322), .C(n487), .A(n486), .Y(o_dacv[62]) );
  AO21X1 U278 ( .B(N1323), .C(n487), .A(n486), .Y(o_dacv[63]) );
  AO21X1 U279 ( .B(N1285), .C(n478), .A(n477), .Y(o_dacv[34]) );
  INVX1 U280 ( .A(n482), .Y(n483) );
  NAND21X1 U281 ( .B(r_adofs[7]), .A(N1313), .Y(n482) );
  NAND2X1 U282 ( .A(N1423), .B(n118), .Y(n314) );
  NAND2X1 U283 ( .A(N1434), .B(n118), .Y(n313) );
  NAND2X1 U284 ( .A(N1379), .B(n118), .Y(n301) );
  NAND2X1 U285 ( .A(N1368), .B(n118), .Y(n302) );
  NAND2X1 U286 ( .A(N1357), .B(n118), .Y(n303) );
  NAND2X1 U287 ( .A(N1401), .B(n118), .Y(n316) );
  NAND2X1 U288 ( .A(N1390), .B(n119), .Y(n317) );
  INVX1 U289 ( .A(n113), .Y(r_adofs[0]) );
  OAI21BBX1 U290 ( .A(N1367), .B(n507), .C(n302), .Y(o_dacv[95]) );
  OAI21BBX1 U291 ( .A(N1356), .B(n506), .C(n303), .Y(o_dacv[87]) );
  OAI21BBX1 U292 ( .A(N1400), .B(n510), .C(n316), .Y(o_dacv[119]) );
  OAI21BBX1 U293 ( .A(N1378), .B(n508), .C(n301), .Y(o_dacv[103]) );
  OAI21BBX1 U294 ( .A(N1389), .B(n509), .C(n317), .Y(o_dacv[111]) );
  AO21X1 U295 ( .B(N1295), .C(n481), .A(n480), .Y(o_dacv[41]) );
  AO21X1 U296 ( .B(N1273), .C(n475), .A(n474), .Y(o_dacv[25]) );
  INVX1 U297 ( .A(N1269), .Y(n472) );
  OAI21BBX1 U298 ( .A(N1361), .B(n507), .C(n302), .Y(o_dacv[89]) );
  OAI21BBX1 U299 ( .A(N1350), .B(n506), .C(n303), .Y(o_dacv[81]) );
  OAI21BBX1 U300 ( .A(N1394), .B(n510), .C(n316), .Y(o_dacv[113]) );
  OAI21BBX1 U301 ( .A(N1372), .B(n508), .C(n301), .Y(o_dacv[97]) );
  OAI21BBX1 U302 ( .A(N1383), .B(n509), .C(n317), .Y(o_dacv[105]) );
  OAI21BBX1 U303 ( .A(N1364), .B(n507), .C(n302), .Y(o_dacv[92]) );
  OAI21BBX1 U304 ( .A(N1353), .B(n506), .C(n303), .Y(o_dacv[84]) );
  OAI21BBX1 U305 ( .A(N1397), .B(n510), .C(n316), .Y(o_dacv[116]) );
  OAI21BBX1 U306 ( .A(N1375), .B(n508), .C(n301), .Y(o_dacv[100]) );
  OAI21BBX1 U307 ( .A(N1386), .B(n509), .C(n317), .Y(o_dacv[108]) );
  OAI21BBX1 U308 ( .A(N1365), .B(n507), .C(n302), .Y(o_dacv[93]) );
  OAI21BBX1 U309 ( .A(N1354), .B(n506), .C(n303), .Y(o_dacv[85]) );
  OAI21BBX1 U310 ( .A(N1398), .B(n510), .C(n316), .Y(o_dacv[117]) );
  OAI21BBX1 U311 ( .A(N1376), .B(n508), .C(n301), .Y(o_dacv[101]) );
  OAI21BBX1 U312 ( .A(N1387), .B(n509), .C(n317), .Y(o_dacv[109]) );
  OAI21BBX1 U313 ( .A(N1362), .B(n507), .C(n302), .Y(o_dacv[90]) );
  OAI21BBX1 U314 ( .A(N1351), .B(n506), .C(n303), .Y(o_dacv[82]) );
  OAI21BBX1 U315 ( .A(N1395), .B(n510), .C(n316), .Y(o_dacv[114]) );
  OAI21BBX1 U316 ( .A(N1373), .B(n508), .C(n301), .Y(o_dacv[98]) );
  OAI21BBX1 U317 ( .A(N1384), .B(n509), .C(n317), .Y(o_dacv[106]) );
  OAI21BBX1 U318 ( .A(N1363), .B(n507), .C(n302), .Y(o_dacv[91]) );
  OAI21BBX1 U319 ( .A(N1352), .B(n506), .C(n303), .Y(o_dacv[83]) );
  OAI21BBX1 U320 ( .A(N1396), .B(n510), .C(n316), .Y(o_dacv[115]) );
  OAI21BBX1 U321 ( .A(N1374), .B(n508), .C(n301), .Y(o_dacv[99]) );
  OAI21BBX1 U322 ( .A(N1385), .B(n509), .C(n317), .Y(o_dacv[107]) );
  OAI21BBX1 U323 ( .A(N1366), .B(n507), .C(n302), .Y(o_dacv[94]) );
  OAI21BBX1 U324 ( .A(N1355), .B(n506), .C(n303), .Y(o_dacv[86]) );
  OAI21BBX1 U325 ( .A(N1399), .B(n510), .C(n316), .Y(o_dacv[118]) );
  OAI21BBX1 U326 ( .A(N1377), .B(n508), .C(n301), .Y(o_dacv[102]) );
  OAI21BBX1 U327 ( .A(N1388), .B(n509), .C(n317), .Y(o_dacv[110]) );
  GEN2XL U328 ( .D(n288), .E(n289), .C(n290), .B(n528), .A(n291), .Y(n284) );
  AOI21X1 U329 ( .B(n287), .C(n289), .A(n528), .Y(n291) );
  NOR21XL U330 ( .B(n285), .A(n271), .Y(n287) );
  AOI21X1 U331 ( .B(n527), .C(n284), .A(n286), .Y(n273) );
  AOI31X1 U332 ( .A(n287), .B(n528), .C(n279), .D(n527), .Y(n286) );
  INVX1 U333 ( .A(n119), .Y(n114) );
  INVX1 U334 ( .A(n119), .Y(n115) );
  OR3XL U335 ( .A(n255), .B(n246), .C(n250), .Y(n254) );
  OAI21X1 U336 ( .B(n273), .C(n274), .A(n275), .Y(n264) );
  OAI211X1 U337 ( .C(n527), .D(n284), .A(n528), .B(n285), .Y(n283) );
  INVX1 U338 ( .A(n119), .Y(n116) );
  INVX1 U339 ( .A(n293), .Y(n532) );
  NAND2X1 U340 ( .A(n272), .B(n264), .Y(n267) );
  INVX1 U341 ( .A(n289), .Y(n529) );
  AOI21BBXL U342 ( .B(n266), .C(n525), .A(n265), .Y(n252) );
  AOI211X1 U343 ( .C(n268), .D(n269), .A(n524), .B(n270), .Y(n266) );
  NAND3X1 U344 ( .A(n528), .B(n527), .C(n271), .Y(n269) );
  NAND32X1 U345 ( .B(n273), .C(n276), .A(n268), .Y(n277) );
  AOI21BX1 U346 ( .C(n283), .B(n268), .A(n281), .Y(n276) );
  OAI21X1 U347 ( .B(n252), .C(n523), .A(n247), .Y(o_smpl[1]) );
  NAND3X1 U348 ( .A(n529), .B(n528), .C(n288), .Y(n279) );
  OAI21X1 U349 ( .B(n523), .C(n255), .A(n254), .Y(o_smpl[0]) );
  NAND2X1 U350 ( .A(n280), .B(n268), .Y(n274) );
  INVX1 U351 ( .A(n280), .Y(n524) );
  INVX1 U352 ( .A(n263), .Y(n525) );
  OAI21AX1 U353 ( .B(n66), .C(n131), .A(r_wr[3]), .Y(updlsb) );
  INVX1 U354 ( .A(n245), .Y(n523) );
  INVX1 U355 ( .A(n200), .Y(n90) );
  AND3X1 U356 ( .A(n501), .B(n502), .C(n517), .Y(n76) );
  MUX2BXL U357 ( .D0(n518), .D1(sacyc_done), .S(n456), .Y(n226) );
  INVX1 U358 ( .A(n129), .Y(n456) );
  NAND21X1 U359 ( .B(n90), .A(n133), .Y(n129) );
  INVX1 U360 ( .A(n522), .Y(n488) );
  INVX1 U361 ( .A(o_dactl[0]), .Y(n220) );
  INVX1 U362 ( .A(n460), .Y(n492) );
  OAI22X1 U363 ( .A(n522), .B(n500), .C(n521), .D(n515), .Y(n434) );
  INVX1 U364 ( .A(n196), .Y(n521) );
  INVX1 U365 ( .A(n131), .Y(n65) );
  NAND21X1 U366 ( .B(n149), .A(n187), .Y(n185) );
  NAND21X1 U367 ( .B(n159), .A(n187), .Y(n188) );
  NAND2X1 U368 ( .A(o_dactl[0]), .B(n133), .Y(n409) );
  NAND2X1 U369 ( .A(n298), .B(n299), .Y(o_intr) );
  NOR4XL U370 ( .A(r_irq[3]), .B(r_irq[2]), .C(r_irq[1]), .D(r_irq[0]), .Y(
        n298) );
  NOR4XL U371 ( .A(r_irq[7]), .B(r_irq[6]), .C(r_irq[5]), .D(r_irq[4]), .Y(
        n299) );
  NAND21X1 U372 ( .B(n494), .A(n77), .Y(n149) );
  NAND21X1 U373 ( .B(cs_ptr[4]), .A(n489), .Y(n179) );
  AO21X1 U374 ( .B(n90), .C(dacyc_done), .A(sacyc_done), .Y(n424) );
  AOI21X1 U375 ( .B(n200), .C(n201), .A(n518), .Y(sar_nxt) );
  NAND2X1 U376 ( .A(n134), .B(n133), .Y(n201) );
  NOR2X1 U377 ( .A(n132), .B(n518), .Y(updcmp) );
  XNOR2XL U378 ( .A(n133), .B(n134), .Y(n132) );
  OAI22X1 U379 ( .A(n159), .B(n441), .C(n447), .D(n534), .Y(datcmp[1]) );
  NOR2X1 U380 ( .A(n520), .B(n159), .Y(n447) );
  OAI22X1 U381 ( .A(n149), .B(n441), .C(n445), .D(n533), .Y(datcmp[5]) );
  NOR2X1 U382 ( .A(n520), .B(n149), .Y(n445) );
  INVX1 U383 ( .A(n310), .Y(n418) );
  NAND21X1 U384 ( .B(n460), .A(cs_ptr[4]), .Y(n310) );
  NAND2X1 U385 ( .A(n245), .B(n246), .Y(o_smpl[4]) );
  AO21X1 U386 ( .B(N1321), .C(n487), .A(n486), .Y(o_dacv[61]) );
  AO21X1 U387 ( .B(N1309), .C(n484), .A(n483), .Y(o_dacv[52]) );
  AO21X1 U388 ( .B(N1316), .C(n487), .A(n486), .Y(o_dacv[56]) );
  AO21X1 U389 ( .B(N1305), .C(n484), .A(n483), .Y(o_dacv[48]) );
  AO21X1 U390 ( .B(N1306), .C(n484), .A(n483), .Y(o_dacv[49]) );
  AO21X1 U391 ( .B(N1311), .C(n484), .A(n483), .Y(o_dacv[54]) );
  AO21X1 U392 ( .B(N1312), .C(n484), .A(n483), .Y(o_dacv[55]) );
  AO21X1 U393 ( .B(N1319), .C(n487), .A(n486), .Y(o_dacv[59]) );
  AO21X1 U394 ( .B(N1317), .C(n487), .A(n486), .Y(o_dacv[57]) );
  AO21X1 U395 ( .B(N1288), .C(n478), .A(n477), .Y(o_dacv[37]) );
  AO21X1 U396 ( .B(N1286), .C(n478), .A(n477), .Y(o_dacv[35]) );
  AO21X1 U397 ( .B(N1297), .C(n481), .A(n480), .Y(o_dacv[43]) );
  AO21X1 U398 ( .B(N1298), .C(n481), .A(n480), .Y(o_dacv[44]) );
  AO21X1 U399 ( .B(N1284), .C(n478), .A(n477), .Y(o_dacv[33]) );
  AO21X1 U400 ( .B(N1289), .C(n478), .A(n477), .Y(o_dacv[38]) );
  AO21X1 U401 ( .B(N1255), .C(n469), .A(n468), .Y(o_dacv[13]) );
  AO21X1 U402 ( .B(N1256), .C(n469), .A(n468), .Y(o_dacv[14]) );
  AO21X1 U403 ( .B(N1250), .C(n469), .A(n468), .Y(o_dacv[8]) );
  AO21X1 U404 ( .B(N1301), .C(n481), .A(n480), .Y(o_dacv[47]) );
  AO21X1 U405 ( .B(N1276), .C(n475), .A(n474), .Y(o_dacv[28]) );
  AO21X1 U406 ( .B(N1296), .C(n481), .A(n480), .Y(o_dacv[42]) );
  AO21X1 U407 ( .B(N1277), .C(n475), .A(n474), .Y(o_dacv[29]) );
  AO21X1 U408 ( .B(N1287), .C(n478), .A(n477), .Y(o_dacv[36]) );
  AO21X1 U409 ( .B(N1290), .C(n478), .A(n477), .Y(o_dacv[39]) );
  AO21X1 U410 ( .B(N1254), .C(n469), .A(n468), .Y(o_dacv[12]) );
  AO21X1 U411 ( .B(N1283), .C(n478), .A(n477), .Y(o_dacv[32]) );
  AO21X1 U412 ( .B(N1318), .C(n487), .A(n486), .Y(o_dacv[58]) );
  AO21X1 U413 ( .B(N1274), .C(n475), .A(n474), .Y(o_dacv[26]) );
  AO21X1 U414 ( .B(N1307), .C(n484), .A(n483), .Y(o_dacv[50]) );
  AO21X1 U415 ( .B(N1308), .C(n484), .A(n483), .Y(o_dacv[51]) );
  AO21X1 U416 ( .B(N1239), .C(n466), .A(n465), .Y(o_dacv[0]) );
  AO21X1 U417 ( .B(N1252), .C(n469), .A(n468), .Y(o_dacv[10]) );
  AO21X1 U418 ( .B(N1310), .C(n484), .A(n483), .Y(o_dacv[53]) );
  AO21X1 U419 ( .B(N1320), .C(n487), .A(n486), .Y(o_dacv[60]) );
  MUX2X1 U420 ( .D0(n10), .D1(o_dactl[5]), .S(n224), .Y(ps_md4ch) );
  OAI221X1 U421 ( .A(n458), .B(n180), .C(n514), .D(n459), .E(n138), .Y(n217)
         );
  INVX1 U422 ( .A(r_sar_en[5]), .Y(n180) );
  OA222X1 U423 ( .A(n515), .B(n440), .C(n438), .D(n137), .E(n516), .F(n439), 
        .Y(n138) );
  INVX1 U424 ( .A(r_sar_en[8]), .Y(n137) );
  OAI221X1 U425 ( .A(n422), .B(n199), .C(n423), .D(n198), .E(n197), .Y(n216)
         );
  INVX1 U426 ( .A(r_sar_en[14]), .Y(n199) );
  INVX1 U427 ( .A(r_sar_en[13]), .Y(n198) );
  OA222X1 U428 ( .A(n421), .B(n183), .C(n496), .D(n419), .E(n495), .F(n311), 
        .Y(n197) );
  NAND6XL U429 ( .A(r_wdat[7]), .B(n90), .C(n220), .D(n219), .E(n415), .F(n5), 
        .Y(n221) );
  NAND43X1 U430 ( .B(n218), .C(n217), .D(n216), .A(n215), .Y(n219) );
  AO2222XL U431 ( .A(r_sar_en[2]), .B(dacv_wr[2]), .C(r_sar_en[3]), .D(
        dacv_wr[3]), .E(r_sar_en[0]), .F(dacv_wr[0]), .G(r_sar_en[1]), .H(
        dacv_wr[1]), .Y(n218) );
  MUX2X1 U432 ( .D0(n6), .D1(o_dactl[4]), .S(n224), .Y(ps_sample) );
  OA2222XL U433 ( .A(n500), .B(n436), .C(n499), .D(n437), .E(n425), .F(n213), 
        .G(n435), .H(n209), .Y(n215) );
  INVX1 U434 ( .A(r_sar_en[12]), .Y(n213) );
  INVX1 U435 ( .A(r_sar_en[11]), .Y(n209) );
  OAI21BBX1 U436 ( .A(N1334), .B(n504), .C(n306), .Y(o_dacv[71]) );
  OAI21BBX1 U437 ( .A(N1411), .B(n511), .C(n315), .Y(o_dacv[127]) );
  OAI21BBX1 U438 ( .A(N1345), .B(n505), .C(n305), .Y(o_dacv[79]) );
  INVX1 U439 ( .A(n544), .Y(n113) );
  OAI21BBX1 U440 ( .A(N1433), .B(n513), .C(n313), .Y(o_dacv[143]) );
  AO21X1 U441 ( .B(N1294), .C(n481), .A(n480), .Y(o_dacv[40]) );
  AO21X1 U442 ( .B(N1272), .C(n475), .A(n474), .Y(o_dacv[24]) );
  BUFX3 U443 ( .A(n541), .Y(n86) );
  BUFX3 U444 ( .A(n541), .Y(r_adofs[1]) );
  OAI21BBX1 U445 ( .A(N1422), .B(n512), .C(n314), .Y(o_dacv[135]) );
  OAI21BBX1 U446 ( .A(N1427), .B(n513), .C(n313), .Y(o_dacv[137]) );
  OAI21BBX1 U447 ( .A(N1428), .B(n513), .C(n313), .Y(o_dacv[138]) );
  OAI21BBX1 U448 ( .A(N1328), .B(n504), .C(n306), .Y(o_dacv[65]) );
  OAI21BBX1 U449 ( .A(N1405), .B(n511), .C(n315), .Y(o_dacv[121]) );
  OAI21BBX1 U450 ( .A(N1331), .B(n504), .C(n306), .Y(o_dacv[68]) );
  OAI21BBX1 U451 ( .A(N1332), .B(n504), .C(n306), .Y(o_dacv[69]) );
  OAI21BBX1 U452 ( .A(N1408), .B(n511), .C(n315), .Y(o_dacv[124]) );
  OAI21BBX1 U453 ( .A(N1330), .B(n504), .C(n306), .Y(o_dacv[67]) );
  OAI21BBX1 U454 ( .A(N1409), .B(n511), .C(n315), .Y(o_dacv[125]) );
  OAI21BBX1 U455 ( .A(N1329), .B(n504), .C(n306), .Y(o_dacv[66]) );
  OAI21BBX1 U456 ( .A(N1407), .B(n511), .C(n315), .Y(o_dacv[123]) );
  OAI21BBX1 U457 ( .A(N1406), .B(n511), .C(n315), .Y(o_dacv[122]) );
  MUX2AXL U458 ( .D0(r_rpt_v[7]), .D1(n9), .S(n130), .Y(n326) );
  MUX2AXL U459 ( .D0(r_rpt_v[5]), .D1(n329), .S(n130), .Y(n331) );
  OAI21BBX1 U460 ( .A(N1339), .B(n505), .C(n305), .Y(o_dacv[73]) );
  OAI21BBX1 U461 ( .A(N1342), .B(n505), .C(n305), .Y(o_dacv[76]) );
  OAI21BBX1 U462 ( .A(N1343), .B(n505), .C(n305), .Y(o_dacv[77]) );
  OAI21BBX1 U463 ( .A(N1341), .B(n505), .C(n305), .Y(o_dacv[75]) );
  OAI21BBX1 U464 ( .A(N1340), .B(n505), .C(n305), .Y(o_dacv[74]) );
  BUFX3 U465 ( .A(n540), .Y(n92) );
  BUFX3 U466 ( .A(n539), .Y(n94) );
  MUX2X1 U467 ( .D0(r_rpt_v[0]), .D1(n78), .S(r_wr[3]), .Y(wdlsb[0]) );
  BUFX3 U468 ( .A(n539), .Y(r_adofs[3]) );
  BUFX3 U469 ( .A(n540), .Y(r_adofs[2]) );
  MUX2X1 U470 ( .D0(x_daclsb[4]), .D1(n10), .S(r_wr[3]), .Y(wdlsb[4]) );
  MUX2X1 U471 ( .D0(r_rpt_v[1]), .D1(n60), .S(r_wr[3]), .Y(wdlsb[1]) );
  MUX2X1 U472 ( .D0(x_daclsb[5]), .D1(n8), .S(r_wr[3]), .Y(wdlsb[5]) );
  MUX2X1 U473 ( .D0(x_daclsb[2]), .D1(n4), .S(r_wr[3]), .Y(wdlsb[2]) );
  MUX2X1 U474 ( .D0(x_daclsb[3]), .D1(n6), .S(r_wr[3]), .Y(wdlsb[3]) );
  MUX2AXL U475 ( .D0(r_rpt_v[3]), .D1(n415), .S(n130), .Y(n416) );
  MUX2AXL U476 ( .D0(r_rpt_v[4]), .D1(n3), .S(n130), .Y(n410) );
  MUX2AXL U477 ( .D0(r_rpt_v[2]), .D1(n13), .S(n130), .Y(n417) );
  MUX2AXL U478 ( .D0(r_rpt_v[6]), .D1(n5), .S(n130), .Y(n328) );
  MUX2AXL U479 ( .D0(r_rpt_v[8]), .D1(n7), .S(n130), .Y(n312) );
  INVX1 U480 ( .A(n470), .Y(n471) );
  NAND21X1 U481 ( .B(r_isofs[7]), .A(N1269), .Y(n470) );
  OAI21BBX1 U482 ( .A(N1416), .B(n512), .C(n314), .Y(o_dacv[129]) );
  OAI21BBX1 U483 ( .A(N1417), .B(n512), .C(n314), .Y(o_dacv[130]) );
  OAI21BBX1 U484 ( .A(N1430), .B(n513), .C(n313), .Y(o_dacv[140]) );
  OAI21BBX1 U485 ( .A(N1420), .B(n512), .C(n314), .Y(o_dacv[133]) );
  OAI21BBX1 U486 ( .A(N1429), .B(n513), .C(n313), .Y(o_dacv[139]) );
  OAI21BBX1 U487 ( .A(N1431), .B(n513), .C(n313), .Y(o_dacv[141]) );
  OAI21BBX1 U488 ( .A(N1421), .B(n512), .C(n314), .Y(o_dacv[134]) );
  OAI21BBX1 U489 ( .A(N1432), .B(n513), .C(n313), .Y(o_dacv[142]) );
  OAI21BBX1 U490 ( .A(N1327), .B(n504), .C(n306), .Y(o_dacv[64]) );
  OAI21BBX1 U491 ( .A(N1333), .B(n504), .C(n306), .Y(o_dacv[70]) );
  OAI21BBX1 U492 ( .A(N1338), .B(n505), .C(n305), .Y(o_dacv[72]) );
  OAI21BBX1 U493 ( .A(N1344), .B(n505), .C(n305), .Y(o_dacv[78]) );
  OAI21BBX1 U494 ( .A(N1404), .B(n511), .C(n315), .Y(o_dacv[120]) );
  OAI21BBX1 U495 ( .A(N1410), .B(n511), .C(n315), .Y(o_dacv[126]) );
  BUFX3 U496 ( .A(n538), .Y(n96) );
  BUFX3 U497 ( .A(n538), .Y(r_adofs[4]) );
  OAI21BBX1 U498 ( .A(N1426), .B(n513), .C(n313), .Y(o_dacv[136]) );
  OAI21BBX1 U499 ( .A(N1415), .B(n512), .C(n314), .Y(o_dacv[128]) );
  OAI21BBX1 U500 ( .A(N1419), .B(n512), .C(n314), .Y(o_dacv[132]) );
  OAI21BBX1 U501 ( .A(N1418), .B(n512), .C(n314), .Y(o_dacv[131]) );
  OAI21BBX1 U502 ( .A(N1360), .B(n507), .C(n302), .Y(o_dacv[88]) );
  OAI21BBX1 U503 ( .A(N1349), .B(n506), .C(n303), .Y(o_dacv[80]) );
  OAI21BBX1 U504 ( .A(N1393), .B(n510), .C(n316), .Y(o_dacv[112]) );
  OAI21BBX1 U505 ( .A(N1371), .B(n508), .C(n301), .Y(o_dacv[96]) );
  OAI21BBX1 U506 ( .A(N1382), .B(n509), .C(n317), .Y(o_dacv[104]) );
  BUFX3 U507 ( .A(n537), .Y(n98) );
  BUFX3 U508 ( .A(n536), .Y(n100) );
  BUFX3 U509 ( .A(n537), .Y(r_adofs[5]) );
  BUFX3 U510 ( .A(n536), .Y(r_adofs[6]) );
  XNOR2XL U511 ( .A(pos_dacis[1]), .B(pos_dacis[0]), .Y(n293) );
  OAI22AX1 U512 ( .D(pos_dacis[3]), .C(n296), .A(pos_dacis[3]), .B(n297), .Y(
        n289) );
  NOR3XL U513 ( .A(n297), .B(pos_dacis[0]), .C(n532), .Y(n296) );
  OAI32X1 U514 ( .A(n530), .B(pos_dacis[0]), .C(n532), .D(pos_dacis[2]), .E(
        n293), .Y(n297) );
  INVX1 U515 ( .A(pos_dacis[2]), .Y(n530) );
  AO22X1 U516 ( .A(pos_dacis[12]), .B(pos_dacis[13]), .C(n525), .D(n267), .Y(
        n265) );
  OA21X1 U517 ( .B(n256), .C(pos_dacis[16]), .A(n253), .Y(n250) );
  NOR4XL U518 ( .A(pos_dacis[15]), .B(pos_dacis[14]), .C(n525), .D(n257), .Y(
        n256) );
  OAI21X1 U519 ( .B(pos_dacis[15]), .C(n258), .A(n259), .Y(n246) );
  NAND4X1 U520 ( .A(pos_dacis[15]), .B(n258), .C(n260), .D(n526), .Y(n259) );
  OAI22BX1 U521 ( .B(pos_dacis[9]), .A(n281), .D(pos_dacis[8]), .C(n282), .Y(
        n270) );
  NOR2X1 U522 ( .A(n273), .B(n283), .Y(n282) );
  OAI22X1 U523 ( .A(n261), .B(n526), .C(pos_dacis[14]), .D(n262), .Y(n258) );
  NOR43XL U524 ( .B(n257), .C(n249), .D(n260), .A(n252), .Y(n261) );
  AOI21X1 U525 ( .B(n263), .C(n264), .A(n265), .Y(n262) );
  NOR42XL U526 ( .C(n251), .D(n253), .A(pos_dacis[14]), .B(pos_dacis[15]), .Y(
        n247) );
  AOI221XL U527 ( .A(n277), .B(n524), .C(pos_dacis[10]), .D(pos_dacis[11]), 
        .E(n270), .Y(n275) );
  OAI21X1 U528 ( .B(n255), .C(n246), .A(pos_dacis[16]), .Y(n253) );
  AOI211X1 U529 ( .C(n529), .D(pos_dacis[5]), .A(pos_dacis[4]), .B(n531), .Y(
        n285) );
  INVX1 U530 ( .A(n294), .Y(n531) );
  NOR3XL U531 ( .A(n273), .B(pos_dacis[8]), .C(n283), .Y(n281) );
  INVX1 U532 ( .A(n535), .Y(n119) );
  NAND2X1 U533 ( .A(pos_dacis[17]), .B(n254), .Y(n251) );
  NAND2X1 U534 ( .A(n247), .B(n248), .Y(o_smpl[3]) );
  OAI21X1 U535 ( .B(pos_dacis[13]), .C(n249), .A(n245), .Y(n248) );
  NOR21XL U536 ( .B(n292), .A(n290), .Y(n271) );
  OAI31XL U537 ( .A(n293), .B(pos_dacis[3]), .C(pos_dacis[2]), .D(n288), .Y(
        n292) );
  OAI21X1 U538 ( .B(pos_dacis[17]), .C(n250), .A(n251), .Y(o_smpl[2]) );
  ENOX1 U539 ( .A(pos_dacis[12]), .B(n267), .C(n272), .D(n263), .Y(n260) );
  OAI2B11X1 U540 ( .D(pos_dacis[15]), .C(n258), .A(n260), .B(n526), .Y(n255)
         );
  AOI31X1 U541 ( .A(n294), .B(n289), .C(n295), .D(n288), .Y(n290) );
  NAND2X1 U542 ( .A(pos_dacis[4]), .B(pos_dacis[5]), .Y(n295) );
  OAI22X1 U543 ( .A(n276), .B(n524), .C(pos_dacis[10]), .D(n277), .Y(n272) );
  INVX1 U544 ( .A(n118), .Y(r_adofs[7]) );
  AOI211X1 U545 ( .C(n532), .D(pos_dacis[3]), .A(pos_dacis[0]), .B(
        pos_dacis[2]), .Y(n294) );
  INVX1 U546 ( .A(n535), .Y(n118) );
  NAND2X1 U547 ( .A(n275), .B(n278), .Y(n257) );
  OAI21AX1 U548 ( .B(pos_dacis[7]), .C(n279), .A(n274), .Y(n278) );
  NOR2X1 U549 ( .A(pos_dacis[4]), .B(pos_dacis[5]), .Y(n288) );
  NAND32X1 U550 ( .B(pos_dacis[12]), .C(n274), .A(n273), .Y(n249) );
  INVX1 U551 ( .A(pos_dacis[6]), .Y(n528) );
  INVX1 U552 ( .A(pos_dacis[7]), .Y(n527) );
  NOR21XL U553 ( .B(app_dacis[9]), .A(n103), .Y(o_daci_sel[9]) );
  NOR21XL U554 ( .B(app_dacis[8]), .A(n102), .Y(o_daci_sel[8]) );
  NOR21XL U555 ( .B(app_dacis[2]), .A(n102), .Y(o_daci_sel[2]) );
  NOR21XL U556 ( .B(app_dacis[3]), .A(n103), .Y(o_daci_sel[3]) );
  NOR21XL U557 ( .B(app_dacis[10]), .A(n103), .Y(o_daci_sel[10]) );
  NOR21XL U558 ( .B(app_dacis[7]), .A(n103), .Y(o_daci_sel[7]) );
  NOR21XL U559 ( .B(app_dacis[5]), .A(n103), .Y(o_daci_sel[5]) );
  NOR21XL U560 ( .B(app_dacis[13]), .A(n102), .Y(o_daci_sel[13]) );
  NOR21XL U561 ( .B(app_dacis[15]), .A(n102), .Y(o_daci_sel[15]) );
  NOR21XL U562 ( .B(app_dacis[6]), .A(n102), .Y(o_daci_sel[6]) );
  NOR21XL U563 ( .B(app_dacis[0]), .A(n102), .Y(o_daci_sel[0]) );
  NOR21XL U564 ( .B(app_dacis[1]), .A(n103), .Y(o_daci_sel[1]) );
  NOR21XL U565 ( .B(app_dacis[17]), .A(n102), .Y(o_daci_sel[17]) );
  NOR21XL U566 ( .B(app_dacis[11]), .A(n102), .Y(o_daci_sel[11]) );
  NOR21XL U567 ( .B(app_dacis[12]), .A(n103), .Y(o_daci_sel[12]) );
  NOR21XL U568 ( .B(app_dacis[14]), .A(n103), .Y(o_daci_sel[14]) );
  NOR21XL U569 ( .B(app_dacis[4]), .A(n102), .Y(o_daci_sel[4]) );
  NOR21XL U570 ( .B(app_dacis[16]), .A(n103), .Y(o_daci_sel[16]) );
  NOR2X1 U571 ( .A(pos_dacis[8]), .B(pos_dacis[9]), .Y(n268) );
  NOR2X1 U572 ( .A(pos_dacis[11]), .B(pos_dacis[10]), .Y(n280) );
  NOR2X1 U573 ( .A(pos_dacis[12]), .B(pos_dacis[13]), .Y(n263) );
  INVX1 U574 ( .A(pos_dacis[14]), .Y(n526) );
  NOR2X1 U575 ( .A(pos_dacis[16]), .B(pos_dacis[17]), .Y(n245) );
  NAND42X1 U576 ( .C(r_dac_en[3]), .D(n128), .A(n127), .B(n126), .Y(n200) );
  NOR43XL U577 ( .B(n125), .C(n124), .D(n123), .A(n122), .Y(n126) );
  NAND21X1 U578 ( .B(r_dac_en[1]), .A(n120), .Y(n128) );
  NOR32XL U579 ( .B(n493), .C(n76), .A(n121), .Y(n127) );
  INVX1 U580 ( .A(r_dac_en[7]), .Y(n517) );
  OR4X1 U581 ( .A(r_dac_en[4]), .B(r_dac_en[5]), .C(r_dac_en[11]), .D(
        r_dac_en[10]), .Y(n122) );
  NAND21X1 U582 ( .B(r_dac_en[0]), .A(n2), .Y(n121) );
  INVX1 U583 ( .A(r_dac_en[15]), .Y(n503) );
  INVX1 U584 ( .A(r_dac_en[17]), .Y(n498) );
  INVX1 U585 ( .A(r_dac_en[8]), .Y(n501) );
  INVX1 U586 ( .A(r_dac_en[2]), .Y(n120) );
  INVX1 U587 ( .A(r_dac_en[16]), .Y(n497) );
  INVX1 U588 ( .A(r_dac_en[6]), .Y(n493) );
  INVX1 U589 ( .A(r_dac_en[13]), .Y(n125) );
  INVX1 U590 ( .A(r_dac_en[9]), .Y(n502) );
  INVX1 U591 ( .A(r_dac_en[14]), .Y(n123) );
  INVX1 U592 ( .A(r_dac_en[12]), .Y(n124) );
  NAND21X1 U593 ( .B(cs_ptr[2]), .A(cs_ptr[3]), .Y(n522) );
  OA2222XL U594 ( .A(n427), .B(n186), .C(n428), .D(n184), .E(n429), .F(n39), 
        .G(n430), .H(n53), .Y(n426) );
  AOI221XL U595 ( .A(r_sar_en[2]), .B(n492), .C(r_sar_en[14]), .D(n489), .E(
        n434), .Y(n427) );
  AOI221XL U596 ( .A(r_sar_en[1]), .B(n492), .C(r_sar_en[13]), .D(n489), .E(
        n432), .Y(n429) );
  NOR2X1 U597 ( .A(n494), .B(cs_ptr[3]), .Y(n196) );
  AOI221XL U598 ( .A(r_sar_en[0]), .B(n492), .C(r_sar_en[12]), .D(n489), .E(
        n431), .Y(n430) );
  ENOX1 U599 ( .A(n521), .B(n514), .C(n488), .D(r_sar_en[8]), .Y(n431) );
  AOI221XL U600 ( .A(r_sar_en[3]), .B(n492), .C(r_sar_en[15]), .D(n489), .E(
        n433), .Y(n428) );
  ENOX1 U601 ( .A(n521), .B(n516), .C(n488), .D(r_sar_en[11]), .Y(n433) );
  ENOX1 U602 ( .A(n522), .B(n499), .C(n196), .D(r_sar_en[5]), .Y(n432) );
  NAND21X1 U603 ( .B(cs_ptr[3]), .A(n494), .Y(n460) );
  XNOR2XL U604 ( .A(n107), .B(x_daclsb[4]), .Y(n414) );
  INVX1 U605 ( .A(n420), .Y(n489) );
  NAND21X1 U606 ( .B(n494), .A(cs_ptr[3]), .Y(n420) );
  INVX1 U607 ( .A(cs_ptr[2]), .Y(n494) );
  NAND4X1 U608 ( .A(o_dactl[6]), .B(n77), .C(n411), .D(n412), .Y(n131) );
  NOR2X1 U609 ( .A(n413), .B(n414), .Y(n412) );
  XNOR2XL U610 ( .A(x_daclsb[3]), .B(n104), .Y(n411) );
  XNOR2XL U611 ( .A(n494), .B(x_daclsb[5]), .Y(n413) );
  INVX1 U612 ( .A(r_sar_en[9]), .Y(n499) );
  INVX1 U613 ( .A(r_sar_en[7]), .Y(n516) );
  INVX1 U614 ( .A(r_sar_en[6]), .Y(n515) );
  INVX1 U615 ( .A(r_sar_en[4]), .Y(n514) );
  INVX1 U616 ( .A(r_sar_en[10]), .Y(n500) );
  NOR43XL U617 ( .B(n189), .C(o_dactl[1]), .D(dacyc_done), .A(n133), .Y(n187)
         );
  XNOR2XL U618 ( .A(syn_comp[1]), .B(n190), .Y(n189) );
  AOI221XL U619 ( .A(n491), .B(n191), .C(n490), .D(n192), .E(n193), .Y(n190)
         );
  OAI22X1 U620 ( .A(n460), .B(n534), .C(n521), .D(n533), .Y(n191) );
  AO222X1 U621 ( .A(n318), .B(n369), .C(n320), .D(n370), .E(r_dac1v[5]), .F(
        n11), .Y(o_dac1[5]) );
  NAND4X1 U622 ( .A(n375), .B(n376), .C(n377), .D(n378), .Y(n369) );
  NAND4X1 U623 ( .A(n371), .B(n372), .C(n373), .D(n374), .Y(n370) );
  AOI22X1 U624 ( .A(r_dacvs[139]), .B(n61), .C(r_dacvs[11]), .D(n334), .Y(n375) );
  AO222X1 U625 ( .A(n318), .B(n319), .C(n320), .D(n321), .E(r_dac1v[9]), .F(
        n12), .Y(o_dac1[9]) );
  NAND4X1 U626 ( .A(n335), .B(n336), .C(n337), .D(n338), .Y(n319) );
  NAND4X1 U627 ( .A(n322), .B(n323), .C(n324), .D(n325), .Y(n321) );
  AOI22X1 U628 ( .A(r_dacvs[143]), .B(n61), .C(r_dacvs[15]), .D(n334), .Y(n335) );
  AO222X1 U629 ( .A(n318), .B(n399), .C(n320), .D(n400), .E(r_dac1v[2]), .F(
        n12), .Y(o_dac1[2]) );
  NAND4X1 U630 ( .A(n405), .B(n406), .C(n407), .D(n408), .Y(n399) );
  NAND4X1 U631 ( .A(n401), .B(n402), .C(n403), .D(n404), .Y(n400) );
  AOI22X1 U632 ( .A(r_dacvs[136]), .B(n62), .C(r_dacvs[8]), .D(n49), .Y(n405)
         );
  AO222X1 U633 ( .A(n318), .B(n389), .C(n320), .D(n390), .E(r_dac1v[3]), .F(
        n11), .Y(o_dac1[3]) );
  NAND4X1 U634 ( .A(n395), .B(n396), .C(n397), .D(n398), .Y(n389) );
  NAND4X1 U635 ( .A(n391), .B(n392), .C(n393), .D(n394), .Y(n390) );
  AOI22X1 U636 ( .A(r_dacvs[137]), .B(n62), .C(r_dacvs[9]), .D(n49), .Y(n395)
         );
  AO222X1 U637 ( .A(n318), .B(n379), .C(n320), .D(n380), .E(r_dac1v[4]), .F(
        n12), .Y(o_dac1[4]) );
  NAND4X1 U638 ( .A(n385), .B(n386), .C(n387), .D(n388), .Y(n379) );
  NAND4X1 U639 ( .A(n381), .B(n382), .C(n383), .D(n384), .Y(n380) );
  AOI22X1 U640 ( .A(r_dacvs[138]), .B(n62), .C(r_dacvs[10]), .D(n49), .Y(n385)
         );
  AO222X1 U641 ( .A(n318), .B(n339), .C(n320), .D(n340), .E(r_dac1v[8]), .F(
        n11), .Y(o_dac1[8]) );
  NAND4X1 U642 ( .A(n345), .B(n346), .C(n347), .D(n348), .Y(n339) );
  NAND4X1 U643 ( .A(n341), .B(n342), .C(n343), .D(n344), .Y(n340) );
  AOI22X1 U644 ( .A(r_dacvs[142]), .B(n62), .C(r_dacvs[14]), .D(n49), .Y(n345)
         );
  AO222X1 U645 ( .A(n318), .B(n359), .C(n320), .D(n360), .E(r_dac1v[6]), .F(
        n11), .Y(o_dac1[6]) );
  NAND4X1 U646 ( .A(n365), .B(n366), .C(n367), .D(n368), .Y(n359) );
  NAND4X1 U647 ( .A(n361), .B(n362), .C(n363), .D(n364), .Y(n360) );
  AOI22X1 U648 ( .A(r_dacvs[140]), .B(n62), .C(r_dacvs[12]), .D(n334), .Y(n365) );
  NOR2X1 U649 ( .A(cs_ptr[4]), .B(cs_ptr[3]), .Y(n77) );
  OAI22X1 U650 ( .A(n194), .B(n184), .C(n195), .D(n186), .Y(n193) );
  AOI22X1 U651 ( .A(o_dat[7]), .B(n196), .C(o_dat[3]), .D(n492), .Y(n194) );
  AOI22X1 U652 ( .A(o_dat[6]), .B(n196), .C(o_dat[2]), .D(n492), .Y(n195) );
  INVX1 U653 ( .A(r_sar_en[17]), .Y(n495) );
  INVX1 U654 ( .A(r_sar_en[16]), .Y(n496) );
  INVX1 U655 ( .A(r_sar_en[15]), .Y(n183) );
  AO222X1 U656 ( .A(n318), .B(n349), .C(n320), .D(n350), .E(r_dac1v[7]), .F(
        n11), .Y(o_dac1[7]) );
  NAND4X1 U657 ( .A(n355), .B(n356), .C(n357), .D(n358), .Y(n349) );
  NAND4X1 U658 ( .A(n351), .B(n352), .C(n353), .D(n354), .Y(n350) );
  AOI22X1 U659 ( .A(r_dacvs[141]), .B(n62), .C(r_dacvs[13]), .D(n49), .Y(n355)
         );
  AO22X1 U660 ( .A(x_daclsb[0]), .B(n409), .C(r_dac1v[0]), .D(n12), .Y(
        o_dac1[0]) );
  AO22X1 U661 ( .A(x_daclsb[1]), .B(n409), .C(r_dac1v[1]), .D(n12), .Y(
        o_dac1[1]) );
  AO22X1 U662 ( .A(n492), .B(o_dat[0]), .C(n196), .D(o_dat[4]), .Y(n192) );
  AOI222XL U663 ( .A(r_dacvs[115]), .B(n74), .C(r_dacvs[99]), .D(n327), .E(
        r_dacvs[83]), .F(n69), .Y(n374) );
  AOI222XL U664 ( .A(r_dacvs[116]), .B(n74), .C(r_dacvs[100]), .D(n327), .E(
        r_dacvs[84]), .F(n69), .Y(n364) );
  AOI222XL U665 ( .A(r_dacvs[119]), .B(n46), .C(r_dacvs[103]), .D(n42), .E(
        r_dacvs[87]), .F(n50), .Y(n325) );
  AOI222XL U666 ( .A(r_dacvs[112]), .B(n46), .C(r_dacvs[96]), .D(n42), .E(
        r_dacvs[80]), .F(n50), .Y(n404) );
  AOI222XL U667 ( .A(r_dacvs[120]), .B(n74), .C(r_dacvs[104]), .D(n327), .E(
        r_dacvs[88]), .F(n69), .Y(n408) );
  AOI222XL U668 ( .A(r_dacvs[113]), .B(n74), .C(r_dacvs[97]), .D(n327), .E(
        r_dacvs[81]), .F(n69), .Y(n394) );
  AOI222XL U669 ( .A(r_dacvs[121]), .B(n46), .C(r_dacvs[105]), .D(n42), .E(
        r_dacvs[89]), .F(n50), .Y(n398) );
  AOI222XL U670 ( .A(r_dacvs[114]), .B(n46), .C(r_dacvs[98]), .D(n42), .E(
        r_dacvs[82]), .F(n50), .Y(n384) );
  AOI222XL U671 ( .A(r_dacvs[122]), .B(n74), .C(r_dacvs[106]), .D(n327), .E(
        r_dacvs[90]), .F(n69), .Y(n388) );
  AOI222XL U672 ( .A(r_dacvs[123]), .B(n46), .C(r_dacvs[107]), .D(n42), .E(
        r_dacvs[91]), .F(n50), .Y(n378) );
  AOI222XL U673 ( .A(r_dacvs[124]), .B(n74), .C(r_dacvs[108]), .D(n327), .E(
        r_dacvs[92]), .F(n69), .Y(n368) );
  AOI222XL U674 ( .A(r_dacvs[117]), .B(n46), .C(r_dacvs[101]), .D(n42), .E(
        r_dacvs[85]), .F(n50), .Y(n354) );
  AOI222XL U675 ( .A(r_dacvs[125]), .B(n46), .C(r_dacvs[109]), .D(n42), .E(
        r_dacvs[93]), .F(n50), .Y(n358) );
  AOI222XL U676 ( .A(r_dacvs[118]), .B(n46), .C(r_dacvs[102]), .D(n42), .E(
        r_dacvs[86]), .F(n50), .Y(n344) );
  AOI222XL U677 ( .A(r_dacvs[126]), .B(n74), .C(r_dacvs[110]), .D(n327), .E(
        r_dacvs[94]), .F(n69), .Y(n348) );
  AOI222XL U678 ( .A(r_dacvs[127]), .B(n74), .C(r_dacvs[111]), .D(n327), .E(
        r_dacvs[95]), .F(n69), .Y(n338) );
  AOI22X1 U679 ( .A(r_dacvs[16]), .B(n57), .C(r_dacvs[64]), .D(n63), .Y(n403)
         );
  AOI22X1 U680 ( .A(r_dacvs[24]), .B(n70), .C(r_dacvs[72]), .D(n330), .Y(n407)
         );
  AOI22X1 U681 ( .A(r_dacvs[17]), .B(n70), .C(r_dacvs[65]), .D(n330), .Y(n393)
         );
  AOI22X1 U682 ( .A(r_dacvs[25]), .B(n57), .C(r_dacvs[73]), .D(n63), .Y(n397)
         );
  AOI22X1 U683 ( .A(r_dacvs[18]), .B(n57), .C(r_dacvs[66]), .D(n63), .Y(n383)
         );
  AOI22X1 U684 ( .A(r_dacvs[26]), .B(n70), .C(r_dacvs[74]), .D(n330), .Y(n387)
         );
  AOI22X1 U685 ( .A(r_dacvs[19]), .B(n70), .C(r_dacvs[67]), .D(n330), .Y(n373)
         );
  AOI22X1 U686 ( .A(r_dacvs[27]), .B(n57), .C(r_dacvs[75]), .D(n63), .Y(n377)
         );
  AOI22X1 U687 ( .A(r_dacvs[20]), .B(n70), .C(r_dacvs[68]), .D(n330), .Y(n363)
         );
  AOI22X1 U688 ( .A(r_dacvs[28]), .B(n70), .C(r_dacvs[76]), .D(n330), .Y(n367)
         );
  AOI22X1 U689 ( .A(r_dacvs[21]), .B(n57), .C(r_dacvs[69]), .D(n63), .Y(n353)
         );
  AOI22X1 U690 ( .A(r_dacvs[29]), .B(n57), .C(r_dacvs[77]), .D(n63), .Y(n357)
         );
  AOI22X1 U691 ( .A(r_dacvs[22]), .B(n57), .C(r_dacvs[70]), .D(n63), .Y(n343)
         );
  AOI22X1 U692 ( .A(r_dacvs[30]), .B(n70), .C(r_dacvs[78]), .D(n330), .Y(n347)
         );
  AOI22X1 U693 ( .A(r_dacvs[23]), .B(n57), .C(r_dacvs[71]), .D(n63), .Y(n324)
         );
  AOI22X1 U694 ( .A(r_dacvs[31]), .B(n70), .C(r_dacvs[79]), .D(n330), .Y(n337)
         );
  AOI22X1 U695 ( .A(r_dacvs[48]), .B(n64), .C(r_dacvs[32]), .D(n332), .Y(n402)
         );
  AOI22X1 U696 ( .A(r_dacvs[56]), .B(n75), .C(r_dacvs[40]), .D(n54), .Y(n406)
         );
  AOI22X1 U697 ( .A(r_dacvs[49]), .B(n75), .C(r_dacvs[33]), .D(n332), .Y(n392)
         );
  AOI22X1 U698 ( .A(r_dacvs[57]), .B(n64), .C(r_dacvs[41]), .D(n54), .Y(n396)
         );
  AOI22X1 U699 ( .A(r_dacvs[50]), .B(n64), .C(r_dacvs[34]), .D(n332), .Y(n382)
         );
  AOI22X1 U700 ( .A(r_dacvs[58]), .B(n75), .C(r_dacvs[42]), .D(n54), .Y(n386)
         );
  AOI22X1 U701 ( .A(r_dacvs[51]), .B(n75), .C(r_dacvs[35]), .D(n332), .Y(n372)
         );
  AOI22X1 U702 ( .A(r_dacvs[59]), .B(n64), .C(r_dacvs[43]), .D(n332), .Y(n376)
         );
  AOI22X1 U703 ( .A(r_dacvs[52]), .B(n75), .C(r_dacvs[36]), .D(n332), .Y(n362)
         );
  AOI22X1 U704 ( .A(r_dacvs[60]), .B(n75), .C(r_dacvs[44]), .D(n332), .Y(n366)
         );
  AOI22X1 U705 ( .A(r_dacvs[53]), .B(n64), .C(r_dacvs[37]), .D(n54), .Y(n352)
         );
  AOI22X1 U706 ( .A(r_dacvs[61]), .B(n64), .C(r_dacvs[45]), .D(n54), .Y(n356)
         );
  AOI22X1 U707 ( .A(r_dacvs[54]), .B(n64), .C(r_dacvs[38]), .D(n54), .Y(n342)
         );
  AOI22X1 U708 ( .A(r_dacvs[62]), .B(n75), .C(r_dacvs[46]), .D(n54), .Y(n346)
         );
  AOI22X1 U709 ( .A(r_dacvs[55]), .B(n64), .C(r_dacvs[39]), .D(n332), .Y(n323)
         );
  AOI22X1 U710 ( .A(r_dacvs[63]), .B(n75), .C(r_dacvs[47]), .D(n332), .Y(n336)
         );
  AOI22X1 U711 ( .A(r_dacvs[128]), .B(n61), .C(r_dacvs[0]), .D(n334), .Y(n401)
         );
  AOI22X1 U712 ( .A(r_dacvs[129]), .B(n62), .C(r_dacvs[1]), .D(n334), .Y(n391)
         );
  AOI22X1 U713 ( .A(r_dacvs[130]), .B(n62), .C(r_dacvs[2]), .D(n334), .Y(n381)
         );
  AOI22X1 U714 ( .A(r_dacvs[131]), .B(n61), .C(r_dacvs[3]), .D(n334), .Y(n371)
         );
  AOI22X1 U715 ( .A(r_dacvs[132]), .B(n61), .C(r_dacvs[4]), .D(n334), .Y(n361)
         );
  AOI22X1 U716 ( .A(r_dacvs[133]), .B(n62), .C(r_dacvs[5]), .D(n49), .Y(n351)
         );
  AOI22X1 U717 ( .A(r_dacvs[134]), .B(n62), .C(r_dacvs[6]), .D(n49), .Y(n341)
         );
  AOI22X1 U718 ( .A(r_dacvs[135]), .B(n61), .C(r_dacvs[7]), .D(n334), .Y(n322)
         );
  INVX1 U719 ( .A(o_dat[5]), .Y(n533) );
  INVX1 U720 ( .A(o_dat[1]), .Y(n534) );
  OAI222XL U721 ( .A(n202), .B(n498), .C(n203), .D(n497), .E(cs_ptr[4]), .F(
        n204), .Y(n134) );
  OA2222XL U722 ( .A(n205), .B(n186), .C(n206), .D(n184), .E(n207), .F(n520), 
        .G(n208), .H(n519), .Y(n204) );
  AOI221XL U723 ( .A(r_dac_en[2]), .B(n45), .C(r_dac_en[14]), .D(n489), .E(
        n214), .Y(n205) );
  AOI221XL U724 ( .A(r_dac_en[1]), .B(n45), .C(r_dac_en[13]), .D(n489), .E(
        n211), .Y(n207) );
  AOI221XL U725 ( .A(r_dac_en[0]), .B(n45), .C(r_dac_en[12]), .D(n489), .E(
        n210), .Y(n208) );
  ENOX1 U726 ( .A(n522), .B(n501), .C(n196), .D(r_dac_en[4]), .Y(n210) );
  AOI221XL U727 ( .A(r_dac_en[3]), .B(n45), .C(r_dac_en[15]), .D(n489), .E(
        n212), .Y(n206) );
  ENOX1 U728 ( .A(n521), .B(n517), .C(n488), .D(r_dac_en[11]), .Y(n212) );
  ENOX1 U729 ( .A(n522), .B(n502), .C(n196), .D(r_dac_en[5]), .Y(n211) );
  ENOX1 U730 ( .A(n521), .B(n493), .C(n488), .D(r_dac_en[10]), .Y(n214) );
  NAND2X1 U731 ( .A(syn_comp[1]), .B(n491), .Y(n441) );
  BUFX3 U732 ( .A(r_comp_opt[0]), .Y(n102) );
  BUFX3 U733 ( .A(r_comp_opt[0]), .Y(n103) );
  OAI21X1 U734 ( .B(n149), .C(n443), .A(n446), .Y(datcmp[4]) );
  OAI21X1 U735 ( .B(n519), .C(n149), .A(o_dat[4]), .Y(n446) );
  OAI21X1 U736 ( .B(n136), .C(n443), .A(n444), .Y(datcmp[8]) );
  OAI21X1 U737 ( .B(n519), .C(n136), .A(o_dat[8]), .Y(n444) );
  OAI21X1 U738 ( .B(n179), .C(n443), .A(n449), .Y(datcmp[12]) );
  OAI21X1 U739 ( .B(n519), .C(n179), .A(o_dat[12]), .Y(n449) );
  OAI21X1 U740 ( .B(n159), .C(n443), .A(n450), .Y(datcmp[0]) );
  OAI21X1 U741 ( .B(n519), .C(n159), .A(o_dat[0]), .Y(n450) );
  OAI21X1 U742 ( .B(n136), .C(n441), .A(n442), .Y(datcmp[9]) );
  OAI21X1 U743 ( .B(n520), .C(n136), .A(o_dat[9]), .Y(n442) );
  OAI21X1 U744 ( .B(n179), .C(n441), .A(n448), .Y(datcmp[13]) );
  OAI21X1 U745 ( .B(n520), .C(n179), .A(o_dat[13]), .Y(n448) );
  ENOX1 U746 ( .A(n150), .B(n109), .C(n150), .D(o_dat[3]), .Y(datcmp[3]) );
  ENOX1 U747 ( .A(n139), .B(n109), .C(n139), .D(o_dat[7]), .Y(datcmp[7]) );
  ENOX1 U748 ( .A(n152), .B(n109), .C(n152), .D(o_dat[2]), .Y(datcmp[2]) );
  ENOX1 U749 ( .A(n140), .B(n109), .C(n140), .D(o_dat[6]), .Y(datcmp[6]) );
  ENOX1 U750 ( .A(n177), .B(n109), .C(o_dat[15]), .D(n177), .Y(datcmp[15]) );
  ENOX1 U751 ( .A(n176), .B(n109), .C(o_dat[16]), .D(n176), .Y(datcmp[16]) );
  ENOX1 U752 ( .A(n182), .B(n109), .C(o_dat[10]), .D(n182), .Y(datcmp[10]) );
  ENOX1 U753 ( .A(n160), .B(n109), .C(o_dat[17]), .D(n160), .Y(datcmp[17]) );
  ENOX1 U754 ( .A(n181), .B(n109), .C(o_dat[11]), .D(n181), .Y(datcmp[11]) );
  ENOX1 U755 ( .A(n178), .B(n109), .C(o_dat[14]), .D(n178), .Y(datcmp[14]) );
  NAND2X1 U756 ( .A(syn_comp[1]), .B(n490), .Y(n443) );
  INVX1 U757 ( .A(syn_comp[1]), .Y(n109) );
  NOR2X2 U758 ( .A(ps_ptr[4]), .B(n228), .Y(n84) );
  BUFXL U759 ( .A(r_wdat[0]), .Y(n78) );
  INVXL U760 ( .A(n89), .Y(n224) );
  NOR2X1 U761 ( .A(n80), .B(n81), .Y(n304) );
  MUX2X2 U762 ( .D0(n304), .D1(n300), .S(ps_ptr[0]), .Y(n308) );
  AOI21AX1 U763 ( .B(ps_ptr[4]), .C(r_dac_en[17]), .A(n79), .Y(n83) );
  MUX2IX1 U764 ( .D0(n244), .D1(n243), .S(ps_ptr[3]), .Y(n79) );
  AOI21XL U765 ( .B(ps_ptr[4]), .C(r_dac_en[16]), .A(n233), .Y(n80) );
  AOI21XL U766 ( .B(ps_ptr[4]), .C(r_sar_en[16]), .A(n236), .Y(n81) );
  NOR2XL U767 ( .A(n82), .B(n83), .Y(n300) );
  AOI21XL U768 ( .B(ps_ptr[4]), .C(r_sar_en[17]), .A(n239), .Y(n82) );
  MUX2X1 U769 ( .D0(n235), .D1(n234), .S(ps_ptr[3]), .Y(n236) );
  MUX2X1 U770 ( .D0(n232), .D1(n231), .S(ps_ptr[3]), .Y(n233) );
  MUX2X1 U771 ( .D0(n238), .D1(n237), .S(ps_ptr[3]), .Y(n239) );
  AO2222X1 U772 ( .A(n1), .B(r_sar_en[6]), .C(n84), .D(r_sar_en[0]), .E(n240), 
        .F(r_sar_en[2]), .G(n242), .H(r_sar_en[4]), .Y(n235) );
  AO2222X1 U773 ( .A(n1), .B(r_sar_en[7]), .C(n84), .D(r_sar_en[1]), .E(n240), 
        .F(r_sar_en[3]), .G(n242), .H(r_sar_en[5]), .Y(n238) );
  AO2222X1 U774 ( .A(n1), .B(r_dac_en[7]), .C(r_dac_en[1]), .D(n84), .E(
        r_dac_en[3]), .F(n240), .G(r_dac_en[5]), .H(n242), .Y(n244) );
  AO2222X1 U775 ( .A(n242), .B(r_sar_en[12]), .C(n1), .D(r_sar_en[14]), .E(
        n241), .F(r_sar_en[8]), .G(n240), .H(r_sar_en[10]), .Y(n234) );
  AO2222X1 U776 ( .A(r_dac_en[13]), .B(n242), .C(n1), .D(r_dac_en[15]), .E(
        r_dac_en[9]), .F(n241), .G(r_dac_en[11]), .H(n240), .Y(n243) );
  AO2222X1 U777 ( .A(n1), .B(r_dac_en[6]), .C(r_dac_en[0]), .D(n84), .E(
        r_dac_en[2]), .F(n240), .G(r_dac_en[4]), .H(n242), .Y(n232) );
  AO2222X1 U778 ( .A(r_dac_en[12]), .B(n242), .C(r_dac_en[14]), .D(n1), .E(
        r_dac_en[8]), .F(n241), .G(r_dac_en[10]), .H(n240), .Y(n231) );
  AO2222X1 U779 ( .A(n242), .B(r_sar_en[13]), .C(n1), .D(r_sar_en[15]), .E(
        n241), .F(r_sar_en[9]), .G(n240), .H(r_sar_en[11]), .Y(n237) );
  NAND21XL U780 ( .B(n457), .A(n226), .Y(n309) );
endmodule


module dacmux_a0_DW01_add_17 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_16 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_15 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_14 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_13 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_12 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_11 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_10 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_9 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_6 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_5 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module glreg_WIDTH2_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n4, n5;

  SDFFRQX1 mem_reg_1_ ( .D(n4), .SIN(rdat[0]), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(n5), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  MUX2XL U2 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n5) );
  MUX2XL U3 ( .D0(rdat[1]), .D1(wdat[1]), .S(we), .Y(n4) );
endmodule


module glreg_WIDTH2_1 ( clk, arstz, we, wdat, rdat, test_si, test_so, test_se
 );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  output test_so;
  wire   n6, n7, n1;

  SDFFRQX1 mem_reg_0_ ( .D(n7), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(n6), .SIN(n1), .SMC(test_se), .C(clk), .XR(arstz), 
        .Q(rdat[1]) );
  BUFX3 U2 ( .A(rdat[0]), .Y(n1) );
  MUX2XL U3 ( .D0(n1), .D1(wdat[0]), .S(we), .Y(n7) );
  MUX2XL U4 ( .D0(rdat[1]), .D1(wdat[1]), .S(we), .Y(n6) );
  BUFX3 U5 ( .A(rdat[1]), .Y(test_so) );
endmodule


module glreg_a0_25 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9677;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_25 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9677), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9677), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9677), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9677), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9677), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9677), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9677), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9677), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9677), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_26 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n3, net9695, n1;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_26 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9695), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(n3), .SMC(test_se), .C(net9695), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9695), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9695), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9695), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9695), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9695), 
        .XR(arstz), .Q(n3) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9695), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9695), 
        .XR(arstz), .Q(rdat[7]) );
  INVXL U2 ( .A(n3), .Y(n1) );
  INVXL U3 ( .A(n1), .Y(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_27 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9713;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_27 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9713), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9713), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9713), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9713), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9713), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9713), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9713), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9713), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9713), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_28 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9731;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_28 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9731), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9731), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9731), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9731), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9731), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9731), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9731), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9731), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9731), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_1 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21;
  wire   [7:0] wd_r;

  glreg_WIDTH8_1 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[5]), .Y(n16) );
  INVX1 U3 ( .A(set2[1]), .Y(n20) );
  NAND21X1 U4 ( .B(set2[5]), .A(n15), .Y(n1) );
  INVX1 U5 ( .A(set2[6]), .Y(n15) );
  INVX1 U6 ( .A(set2[0]), .Y(n21) );
  INVX1 U7 ( .A(set2[2]), .Y(n19) );
  INVX1 U8 ( .A(set2[4]), .Y(n17) );
  INVX1 U9 ( .A(set2[7]), .Y(n14) );
  INVX1 U10 ( .A(set2[3]), .Y(n18) );
  NAND42X1 U11 ( .C(n5), .D(n4), .A(n3), .B(n2), .Y(upd_r) );
  NOR43XL U12 ( .B(n14), .C(n18), .D(n17), .A(n1), .Y(n2) );
  NAND21X1 U13 ( .B(set2[1]), .A(n19), .Y(n4) );
  NAND21X1 U14 ( .B(clr1[0]), .A(n21), .Y(n5) );
  NOR8XL U15 ( .A(clr1[4]), .B(clr1[5]), .C(clr1[6]), .D(clr1[7]), .E(rst0), 
        .F(clr1[1]), .G(clr1[2]), .H(clr1[3]), .Y(n3) );
  AOI211X1 U16 ( .C(n19), .D(n11), .A(clr1[2]), .B(rst0), .Y(wd_r[2]) );
  INVX1 U17 ( .A(rdat[2]), .Y(n11) );
  AOI211X1 U18 ( .C(n17), .D(n9), .A(clr1[4]), .B(rst0), .Y(wd_r[4]) );
  INVX1 U19 ( .A(rdat[4]), .Y(n9) );
  AOI211X1 U20 ( .C(n21), .D(n13), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U21 ( .A(rdat[0]), .Y(n13) );
  AOI211X1 U22 ( .C(n20), .D(n12), .A(clr1[1]), .B(rst0), .Y(wd_r[1]) );
  INVX1 U23 ( .A(rdat[1]), .Y(n12) );
  AOI211X1 U24 ( .C(n18), .D(n10), .A(clr1[3]), .B(rst0), .Y(wd_r[3]) );
  INVX1 U25 ( .A(rdat[3]), .Y(n10) );
  AOI211X1 U26 ( .C(n16), .D(n8), .A(clr1[5]), .B(rst0), .Y(wd_r[5]) );
  INVX1 U27 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U28 ( .C(n15), .D(n7), .A(clr1[6]), .B(rst0), .Y(wd_r[6]) );
  INVX1 U29 ( .A(rdat[6]), .Y(n7) );
  AOI211X1 U30 ( .C(n14), .D(n6), .A(clr1[7]), .B(rst0), .Y(wd_r[7]) );
  INVX1 U31 ( .A(rdat[7]), .Y(n6) );
  NOR2X1 U32 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
  NOR2X1 U33 ( .A(rdat[1]), .B(n20), .Y(irq[1]) );
  NOR2X1 U34 ( .A(rdat[0]), .B(n21), .Y(irq[0]) );
  NOR2X1 U35 ( .A(rdat[4]), .B(n17), .Y(irq[4]) );
  NOR2X1 U36 ( .A(rdat[6]), .B(n15), .Y(irq[6]) );
  NOR2X1 U37 ( .A(rdat[2]), .B(n19), .Y(irq[2]) );
  NOR2X1 U38 ( .A(rdat[7]), .B(n14), .Y(irq[7]) );
  NOR2X1 U39 ( .A(rdat[3]), .B(n18), .Y(irq[3]) );
endmodule


module glreg_WIDTH8_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9749;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9749), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9749), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9749), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9749), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9749), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9749), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9749), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9749), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9749), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_29 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9767;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_29 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9767), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9767), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9767), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9767), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9767), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9767), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9767), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9767), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9767), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_30 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9785;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_30 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9785), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9785), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9785), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9785), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9785), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9785), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9785), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9785), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9785), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_31 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9803;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_31 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9803), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9803), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9803), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9803), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9803), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9803), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9803), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9803), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9803), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_32 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9821;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_32 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9821), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9821), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9821), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9821), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9821), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9821), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9821), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9821), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9821), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_33 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9839;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_33 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9839), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9839), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9839), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9839), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9839), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9839), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9839), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9839), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9839), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_34 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9857;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_34 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9857), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9857), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9857), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9857), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9857), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9857), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9857), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9857), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9857), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_35 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9875;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_35 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9875), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9875), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9875), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9875), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9875), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9875), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9875), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9875), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9875), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_36 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9893;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_36 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9893), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9893), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9893), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9893), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9893), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9893), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9893), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9893), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9893), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_37 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9911;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_37 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9911), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9911), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9911), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9911), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9911), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9911), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9911), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9911), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9911), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_38 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9929;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_38 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9929), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9929), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9929), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9929), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9929), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9929), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9929), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9929), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9929), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_39 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9947;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_39 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9947), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9947), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9947), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9947), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9947), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9947), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9947), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9947), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9947), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_40 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9965;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_40 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9965), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9965), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9965), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9965), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9965), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9965), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9965), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9965), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9965), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_41 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9983;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_41 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9983), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9983), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9983), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9983), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9983), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9983), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9983), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9983), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9983), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_42 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10001;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_42 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10001), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10001), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10001), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10001), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10001), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10001), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10001), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10001), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10001), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_43 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10019;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_43 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10019), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10019), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10019), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10019), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10019), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10019), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10019), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10019), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10019), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_44 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10037;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_44 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10037), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10037), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10037), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10037), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10037), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10037), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10037), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10037), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10037), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_45 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10055;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_45 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10055), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10055), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10055), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10055), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10055), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10055), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10055), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10055), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10055), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_46 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10073;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_46 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10073), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10073), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10073), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10073), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10073), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10073), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10073), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10073), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10073), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10091;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10091), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10091), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10091), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10091), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10091), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10091), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10091), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_47 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10109;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_47 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10109), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10109), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10109), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10109), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10109), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10109), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10109), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10109), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10109), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_48 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n11, n12, n13, n14, n15, net10127, n1, n3, n5, n7, n9;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_48 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10127), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(n14), .SMC(test_se), .C(net10127), 
        .XR(arstz), .Q(n13) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(n13), .SMC(test_se), .C(net10127), 
        .XR(arstz), .Q(n12) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(n12), .SMC(test_se), .C(net10127), 
        .XR(arstz), .Q(n11) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(n11), .SMC(test_se), .C(net10127), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10127), .XR(arstz), .Q(n14) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(n15), .SMC(test_se), .C(net10127), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10127), .XR(arstz), .Q(n15) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10127), .XR(arstz), .Q(rdat[7]) );
  INVXL U2 ( .A(n14), .Y(n1) );
  INVXL U3 ( .A(n1), .Y(rdat[2]) );
  INVXL U4 ( .A(n11), .Y(n3) );
  INVXL U5 ( .A(n3), .Y(rdat[5]) );
  INVXL U6 ( .A(n12), .Y(n5) );
  INVXL U7 ( .A(n5), .Y(rdat[4]) );
  INVXL U8 ( .A(n13), .Y(n7) );
  INVXL U9 ( .A(n7), .Y(rdat[3]) );
  INVX1 U10 ( .A(n15), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH7_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10145;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10145), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10145), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10145), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10145), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10145), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10145), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10145), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10145), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module shmux_00000005_00000012_00000012 ( ps_sample, ps_md4ch, r_comp_swtch, 
        r_semi, r_loop, r_dac_en, wr_dacv, busy, sh_hold, stop, semi_start, 
        auto_start, mxcyc_done, sampl_begn, sampl_done, app_dacis, pos_dacis, 
        cs_ptr, ps_ptr, clk, srstz, test_si2, test_si1, test_so1, test_se );
  input [17:0] r_dac_en;
  input [17:0] wr_dacv;
  output [17:0] app_dacis;
  output [17:0] pos_dacis;
  output [4:0] cs_ptr;
  output [4:0] ps_ptr;
  input ps_sample, ps_md4ch, r_comp_swtch, r_semi, r_loop, stop, semi_start,
         auto_start, mxcyc_done, sampl_begn, sampl_done, clk, srstz, test_si2,
         test_si1, test_se;
  output busy, sh_hold, test_so1;
  wire   cs_mux_5_, neg_dacis_16_, neg_dacis_15_, neg_dacis_14_, neg_dacis_13_,
         neg_dacis_12_, neg_dacis_11_, neg_dacis_10_, neg_dacis_9_,
         neg_dacis_8_, neg_dacis_7_, neg_dacis_6_, neg_dacis_5_, neg_dacis_4_,
         neg_dacis_3_, neg_dacis_2_, neg_dacis_1_, neg_dacis_0_, N956, N957,
         N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, N973, N1002, N1003, N1004, N1005, N1006,
         N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016,
         N1017, N1018, N1019, N1020, N1030, N1031, N1032, N1033, N1034, N1035,
         N1175, N1184, N1225, N1257, N1266, N1298, N1307, N1339, N1348, N1380,
         N1389, N1421, N1430, N1585, N1594, N1708, N1717, net10163, net10169,
         n660, sub_395_S2_I14_aco_carry_4_, n52, n53, n54, n55, n56, n66, n67,
         n68, n71, n729, n728, n727, n726, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n197, n202, n203, n204, n205, n207, n209,
         n210, n211, n213, n215, n217, n218, n219, n220, n221, n222, n223,
         n270, n271, n276, n291, n306, n307, n311, n327, n328, n330, n331,
         n338, n344, n345, n354, n355, n356, n367, n403, n404, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n474, n476, n477, n478, n479, n480, n481, n482,
         n483, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n522, n523, n527, n528, n529, n530, n531, n555, n563, n569, n570,
         n571, n572, n573, n575, n576, n577, n583, n584, n586, n588, n590,
         n591, n592, n593, n594, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n644, n646, n647, n648, n649, n652,
         n653, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n42, n43, n44,
         n46, n47, n49, n50, n51, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n69, n70, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n198, n199, n200, n201, n206, n208, n212, n214, n216, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n272, n273, n274, n275, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n308,
         n309, n310, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n329, n332, n333, n334, n335,
         n336, n337, n339, n340, n341, n342, n343, n346, n347, n348, n349,
         n350, n351, n352, n353, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n405, n420, n421, n422, n423, n424,
         n471, n472, n473, n475, n484, n517, n518, n519, n520, n521, n524,
         n525, n526, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n556, n557, n558, n559, n560, n561, n562, n564,
         n565, n566, n567, n568, n574, n578, n579, n580, n581, n582, n585,
         n587, n589, n595, n596, n642, n643, n645, n650, n651, n654, n655,
         n656, n657, n658, n659, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725;
  wire   [5:4] sub_395_S2_aco_carry;
  wire   [5:4] sub_395_S2_I2_aco_carry;
  wire   [5:4] sub_395_S2_I3_aco_carry;
  wire   [5:4] sub_395_S2_I4_aco_carry;
  wire   [5:4] sub_395_S2_I5_aco_carry;
  wire   [5:4] sub_395_S2_I6_aco_carry;
  wire   [5:4] sub_395_S2_I7_aco_carry;
  wire   [5:4] sub_395_S2_I11_aco_carry;

  FAD1X1 sub_395_S2_aco_U2_4 ( .A(N1175), .B(n55), .CI(sub_395_S2_aco_carry[4]), .CO(sub_395_S2_aco_carry[5]), .SO(N1184) );
  FAD1X1 sub_395_S2_I2_aco_U2_4 ( .A(n51), .B(n71), .CI(
        sub_395_S2_I2_aco_carry[4]), .CO(sub_395_S2_I2_aco_carry[5]), .SO(
        N1225) );
  FAD1X1 sub_395_S2_I3_aco_U2_4 ( .A(N1257), .B(n56), .CI(
        sub_395_S2_I3_aco_carry[4]), .CO(sub_395_S2_I3_aco_carry[5]), .SO(
        N1266) );
  FAD1X1 sub_395_S2_I4_aco_U2_4 ( .A(N1298), .B(n67), .CI(
        sub_395_S2_I4_aco_carry[4]), .CO(sub_395_S2_I4_aco_carry[5]), .SO(
        N1307) );
  FAD1X1 sub_395_S2_I5_aco_U2_4 ( .A(N1339), .B(n54), .CI(
        sub_395_S2_I5_aco_carry[4]), .CO(sub_395_S2_I5_aco_carry[5]), .SO(
        N1348) );
  FAD1X1 sub_395_S2_I6_aco_U2_4 ( .A(N1380), .B(n68), .CI(
        sub_395_S2_I6_aco_carry[4]), .CO(sub_395_S2_I6_aco_carry[5]), .SO(
        N1389) );
  FAD1X1 sub_395_S2_I7_aco_U2_4 ( .A(N1421), .B(n52), .CI(
        sub_395_S2_I7_aco_carry[4]), .CO(sub_395_S2_I7_aco_carry[5]), .SO(
        N1430) );
  FAD1X1 sub_395_S2_I11_aco_U2_4 ( .A(N1585), .B(n53), .CI(
        sub_395_S2_I11_aco_carry[4]), .CO(sub_395_S2_I11_aco_carry[5]), .SO(
        N1594) );
  INVX8 U741 ( .A(srstz), .Y(n177) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 clk_gate_r_dacis_reg ( 
        .CLK(clk), .EN(N1002), .ENCLK(net10163), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 clk_gate_cs_mux_reg ( 
        .CLK(clk), .EN(N1030), .ENCLK(net10169), .TE(test_se) );
  SDFFQX1 cs_mux_reg_4_ ( .D(N1035), .SIN(cs_ptr[3]), .SMC(test_se), .C(
        net10169), .Q(n726) );
  SDFFQX1 cs_mux_reg_0_ ( .D(N1031), .SIN(test_si2), .SMC(test_se), .C(
        net10169), .Q(n729) );
  SDFFQX1 cs_mux_reg_2_ ( .D(N1033), .SIN(n728), .SMC(test_se), .C(net10169), 
        .Q(cs_ptr[2]) );
  SDFFQX1 cs_mux_reg_3_ ( .D(N1034), .SIN(n11), .SMC(test_se), .C(net10169), 
        .Q(n727) );
  SDFFQX1 cs_mux_reg_1_ ( .D(N1032), .SIN(n42), .SMC(test_se), .C(net10169), 
        .Q(n728) );
  SDFFQX1 r_dacis_reg_16_ ( .D(N1019), .SIN(pos_dacis[15]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[16]) );
  SDFFQX1 r_dacis_reg_17_ ( .D(N1020), .SIN(pos_dacis[16]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[17]) );
  SDFFQX1 r_dacis_reg_11_ ( .D(N1014), .SIN(pos_dacis[10]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[11]) );
  SDFFQX1 r_dacis_reg_10_ ( .D(N1013), .SIN(pos_dacis[9]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[10]) );
  SDFFQX1 r_dacis_reg_13_ ( .D(N1016), .SIN(pos_dacis[12]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[13]) );
  SDFFQX1 r_dacis_reg_12_ ( .D(N1015), .SIN(pos_dacis[11]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[12]) );
  SDFFQX1 r_dacis_reg_15_ ( .D(N1018), .SIN(pos_dacis[14]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[15]) );
  SDFFQX1 r_dacis_reg_14_ ( .D(N1017), .SIN(pos_dacis[13]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[14]) );
  SDFFQX1 r_dacis_reg_9_ ( .D(N1012), .SIN(pos_dacis[8]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[9]) );
  SDFFQX1 r_dacis_reg_8_ ( .D(N1011), .SIN(pos_dacis[7]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[8]) );
  SDFFNQX1 neg_dacis_reg_0_ ( .D(N956), .SIN(test_si1), .SMC(test_se), .XC(clk), .Q(neg_dacis_0_) );
  SDFFNQX1 neg_dacis_reg_1_ ( .D(N957), .SIN(neg_dacis_0_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_1_) );
  SDFFNQX1 neg_dacis_reg_2_ ( .D(N958), .SIN(neg_dacis_1_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_2_) );
  SDFFNQX1 neg_dacis_reg_3_ ( .D(N959), .SIN(neg_dacis_2_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_3_) );
  SDFFNQX1 neg_dacis_reg_4_ ( .D(N960), .SIN(neg_dacis_3_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_4_) );
  SDFFNQX1 neg_dacis_reg_5_ ( .D(N961), .SIN(neg_dacis_4_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_5_) );
  SDFFNQX1 neg_dacis_reg_6_ ( .D(N962), .SIN(neg_dacis_5_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_6_) );
  SDFFNQX1 neg_dacis_reg_7_ ( .D(N963), .SIN(neg_dacis_6_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_7_) );
  SDFFNQX1 neg_dacis_reg_8_ ( .D(N964), .SIN(neg_dacis_7_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_8_) );
  SDFFNQX1 neg_dacis_reg_9_ ( .D(N965), .SIN(neg_dacis_8_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_9_) );
  SDFFNQX1 neg_dacis_reg_10_ ( .D(N966), .SIN(neg_dacis_9_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_10_) );
  SDFFNQX1 neg_dacis_reg_11_ ( .D(N967), .SIN(neg_dacis_10_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_11_) );
  SDFFNQX1 neg_dacis_reg_12_ ( .D(N968), .SIN(neg_dacis_11_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_12_) );
  SDFFNQX1 neg_dacis_reg_13_ ( .D(N969), .SIN(neg_dacis_12_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_13_) );
  SDFFNQX1 neg_dacis_reg_14_ ( .D(N970), .SIN(neg_dacis_13_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_14_) );
  SDFFNQX1 neg_dacis_reg_15_ ( .D(N971), .SIN(neg_dacis_14_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_15_) );
  SDFFNQX1 neg_dacis_reg_16_ ( .D(N972), .SIN(neg_dacis_15_), .SMC(test_se), 
        .XC(clk), .Q(neg_dacis_16_) );
  SDFFNQX1 neg_dacis_reg_17_ ( .D(N973), .SIN(neg_dacis_16_), .SMC(test_se), 
        .XC(clk), .Q(test_so1) );
  SDFFQX1 r_dacis_reg_6_ ( .D(N1009), .SIN(pos_dacis[5]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[6]) );
  SDFFQX1 r_dacis_reg_7_ ( .D(N1010), .SIN(pos_dacis[6]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[7]) );
  SDFFQX1 r_dacis_reg_4_ ( .D(N1007), .SIN(pos_dacis[3]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[4]) );
  SDFFQX1 r_dacis_reg_5_ ( .D(N1008), .SIN(pos_dacis[4]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[5]) );
  SDFFQX1 cs_mux_reg_5_ ( .D(n660), .SIN(n50), .SMC(test_se), .C(clk), .Q(
        cs_mux_5_) );
  SDFFQX1 r_dacis_reg_3_ ( .D(N1006), .SIN(pos_dacis[2]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[3]) );
  SDFFQX1 r_dacis_reg_1_ ( .D(N1004), .SIN(pos_dacis[0]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[1]) );
  SDFFQX1 r_dacis_reg_2_ ( .D(N1005), .SIN(pos_dacis[1]), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[2]) );
  SDFFQX1 r_dacis_reg_0_ ( .D(N1003), .SIN(cs_mux_5_), .SMC(test_se), .C(
        net10163), .Q(pos_dacis[0]) );
  INVX3 U3 ( .A(n153), .Y(n201) );
  NAND21X1 U4 ( .B(r_semi), .A(n152), .Y(n153) );
  GEN2XL U5 ( .D(n594), .E(n664), .C(n669), .B(n28), .A(n597), .Y(n590) );
  OA222X1 U6 ( .A(n387), .B(n334), .C(n528), .D(n129), .E(n655), .F(n386), .Y(
        n130) );
  GEN2XL U7 ( .D(n241), .E(n728), .C(n159), .B(n158), .A(n238), .Y(n160) );
  INVX1 U8 ( .A(auto_start), .Y(n152) );
  INVX1 U9 ( .A(n361), .Y(n195) );
  NOR2X1 U10 ( .A(n363), .B(n163), .Y(n17) );
  GEN3XL U11 ( .F(n326), .G(n325), .E(n324), .D(n323), .C(n322), .B(n321), .A(
        n320), .Y(n329) );
  OAI211X1 U12 ( .C(n301), .D(n361), .A(n300), .B(n299), .Y(ps_ptr[3]) );
  OA222X1 U13 ( .A(n27), .B(n348), .C(n574), .D(n353), .E(n298), .F(n347), .Y(
        n299) );
  OA222X1 U14 ( .A(n272), .B(n348), .C(n269), .D(n353), .E(n268), .F(n347), 
        .Y(n273) );
  NAND32X1 U15 ( .B(n177), .C(stop), .A(n537), .Y(n660) );
  AND2X1 U16 ( .A(n414), .B(n581), .Y(n1) );
  OAI21X1 U17 ( .B(n608), .C(n609), .A(n610), .Y(n2) );
  AOI21X1 U18 ( .B(n658), .C(n80), .A(n79), .Y(n3) );
  AND4X1 U19 ( .A(n512), .B(n419), .C(n511), .D(n632), .Y(n4) );
  AOI21X1 U20 ( .B(n580), .C(n282), .A(n281), .Y(n5) );
  OA21X1 U21 ( .B(n494), .C(n495), .A(n78), .Y(n6) );
  AOI21X1 U22 ( .B(n230), .C(n509), .A(n685), .Y(n7) );
  BUFXL U23 ( .A(r_dac_en[11]), .Y(n8) );
  INVXL U24 ( .A(n312), .Y(n9) );
  INVX1 U25 ( .A(cs_ptr[3]), .Y(n10) );
  INVX1 U26 ( .A(n12), .Y(n11) );
  GEN2XL U27 ( .D(n241), .E(n11), .C(n256), .B(n33), .A(n240), .Y(n249) );
  OR3X1 U28 ( .A(wr_dacv[0]), .B(n201), .C(r_dac_en[0]), .Y(n363) );
  BUFX3 U29 ( .A(n587), .Y(n12) );
  BUFX3 U30 ( .A(n727), .Y(cs_ptr[3]) );
  NAND2X1 U31 ( .A(sampl_done), .B(srstz), .Y(n14) );
  INVX1 U32 ( .A(n36), .Y(n15) );
  NAND42X1 U33 ( .C(n275), .D(n21), .A(n274), .B(n273), .Y(ps_ptr[4]) );
  INVXL U34 ( .A(n534), .Y(n341) );
  INVX1 U35 ( .A(n262), .Y(n16) );
  NAND32X1 U36 ( .B(n224), .C(n216), .A(n214), .Y(n347) );
  INVXL U37 ( .A(ps_ptr[3]), .Y(n388) );
  AOI21BXL U38 ( .C(n16), .B(n261), .A(n534), .Y(n21) );
  AOI32XL U39 ( .A(n297), .B(n323), .C(n296), .D(n341), .E(n295), .Y(n300) );
  INVXL U40 ( .A(ps_ptr[0]), .Y(n395) );
  INVXL U41 ( .A(n256), .Y(n285) );
  AOI211XL U42 ( .C(n395), .D(n41), .A(n374), .B(n373), .Y(n375) );
  XNOR2XL U43 ( .A(n466), .B(cs_ptr[1]), .Y(n327) );
  INVXL U44 ( .A(n237), .Y(n158) );
  NAND32XL U45 ( .B(n332), .C(n257), .A(n17), .Y(n258) );
  INVXL U46 ( .A(n286), .Y(n241) );
  INVXL U47 ( .A(n363), .Y(n198) );
  MUX2IXL U48 ( .D0(n43), .D1(n395), .S(ps_sample), .Y(n35) );
  OAI211XL U49 ( .C(n589), .D(n286), .A(n33), .B(n285), .Y(n296) );
  AND4XL U50 ( .A(ps_sample), .B(n376), .C(n420), .D(n375), .Y(n384) );
  AND2XL U51 ( .A(n558), .B(ps_ptr[0]), .Y(N1031) );
  AND2XL U52 ( .A(n558), .B(ps_ptr[3]), .Y(N1034) );
  XNOR2XL U53 ( .A(n587), .B(n589), .Y(n180) );
  OAI222XL U54 ( .A(n270), .B(n625), .C(n626), .D(n695), .E(n431), .F(n696), 
        .Y(n584) );
  XNOR2XL U55 ( .A(n589), .B(n710), .Y(n501) );
  NOR21XL U56 ( .B(n655), .A(wr_dacv[10]), .Y(n317) );
  AOI31XL U57 ( .A(n309), .B(n308), .C(n305), .D(n304), .Y(n314) );
  NAND32XL U58 ( .B(wr_dacv[3]), .C(r_dac_en[3]), .A(n329), .Y(n333) );
  INVXL U59 ( .A(n302), .Y(n326) );
  XNOR2XL U60 ( .A(n516), .B(n727), .Y(n514) );
  AND2X1 U61 ( .A(n389), .B(n388), .Y(n390) );
  AND2X1 U62 ( .A(n543), .B(n402), .Y(N1005) );
  INVX1 U63 ( .A(n549), .Y(n556) );
  INVX1 U64 ( .A(n546), .Y(n543) );
  INVX1 U65 ( .A(wr_dacv[2]), .Y(n335) );
  INVX1 U66 ( .A(n583), .Y(n190) );
  INVX1 U67 ( .A(n518), .Y(n165) );
  INVX1 U68 ( .A(n475), .Y(n187) );
  INVX1 U69 ( .A(n292), .Y(n342) );
  INVX1 U70 ( .A(n344), .Y(n675) );
  INVX1 U71 ( .A(n489), .Y(n688) );
  NAND2XL U72 ( .A(n200), .B(n201), .Y(n348) );
  INVX4 U73 ( .A(n154), .Y(n214) );
  INVX1 U74 ( .A(wr_dacv[16]), .Y(n309) );
  INVX1 U75 ( .A(n550), .Y(n402) );
  AND2X1 U76 ( .A(n543), .B(n551), .Y(N1017) );
  AND2X1 U77 ( .A(n402), .B(n552), .Y(N1004) );
  AND2X1 U78 ( .A(n402), .B(n554), .Y(N1006) );
  AND2X1 U79 ( .A(n551), .B(n556), .Y(N1015) );
  AND2X1 U80 ( .A(n551), .B(n554), .Y(N1018) );
  AND2X1 U81 ( .A(n554), .B(n553), .Y(N1014) );
  AND2X1 U82 ( .A(n552), .B(n551), .Y(N1016) );
  INVXL U83 ( .A(wr_dacv[12]), .Y(n316) );
  INVX1 U84 ( .A(n547), .Y(n553) );
  OR2X1 U85 ( .A(n400), .B(n401), .Y(n549) );
  NAND21X1 U86 ( .B(n401), .A(n400), .Y(n546) );
  INVX1 U87 ( .A(stop), .Y(n61) );
  AND2X1 U88 ( .A(n588), .B(n22), .Y(n583) );
  NAND2X1 U89 ( .A(n685), .B(n700), .Y(sub_395_S2_I7_aco_carry[4]) );
  INVX1 U90 ( .A(n230), .Y(n169) );
  INVX1 U91 ( .A(n473), .Y(n174) );
  NAND21X1 U92 ( .B(n22), .A(n588), .Y(n475) );
  NAND2X1 U93 ( .A(n108), .B(n109), .Y(n292) );
  NAND21X1 U94 ( .B(n108), .A(n109), .Y(n518) );
  OA2222XL U95 ( .A(n681), .B(n473), .C(n517), .D(n265), .E(n687), .F(n424), 
        .G(n690), .H(n475), .Y(n266) );
  INVX1 U96 ( .A(N1430), .Y(n265) );
  NAND21X1 U97 ( .B(n188), .A(n583), .Y(n472) );
  INVX1 U98 ( .A(N1348), .Y(n687) );
  INVX1 U99 ( .A(N1594), .Y(n693) );
  NOR2X1 U100 ( .A(n499), .B(n54), .Y(n622) );
  INVX1 U101 ( .A(n647), .Y(n684) );
  INVX1 U102 ( .A(n516), .Y(n702) );
  INVX1 U103 ( .A(n631), .Y(n697) );
  INVX1 U104 ( .A(n481), .Y(n643) );
  OAI21X1 U105 ( .B(n676), .C(n705), .A(n465), .Y(n344) );
  INVX1 U106 ( .A(n367), .Y(n80) );
  MUX2X1 U107 ( .D0(n483), .D1(n485), .S(n6), .Y(n79) );
  OAI21X1 U108 ( .B(n496), .C(n709), .A(n491), .Y(n489) );
  OA222X1 U109 ( .A(n111), .B(n352), .C(n110), .D(n292), .E(n679), .F(n340), 
        .Y(n112) );
  INVX1 U110 ( .A(N1266), .Y(n690) );
  INVX1 U111 ( .A(n175), .Y(n307) );
  AND4X1 U112 ( .A(n517), .B(n424), .C(n473), .D(n475), .Y(n339) );
  AND4X1 U113 ( .A(n471), .B(n336), .C(n484), .D(n472), .Y(n337) );
  INVX1 U114 ( .A(n507), .Y(n692) );
  INVX1 U115 ( .A(n565), .Y(n699) );
  INVX1 U116 ( .A(n385), .Y(n691) );
  INVX1 U117 ( .A(n349), .Y(n290) );
  NOR2X1 U118 ( .A(n674), .B(n67), .Y(n606) );
  INVX1 U119 ( .A(n351), .Y(n289) );
  NAND2X1 U120 ( .A(n496), .B(n709), .Y(n491) );
  NAND2X1 U121 ( .A(n676), .B(n705), .Y(n465) );
  INVX1 U122 ( .A(n467), .Y(n676) );
  NAND21X1 U123 ( .B(n3), .A(n352), .Y(n340) );
  NAND21X1 U124 ( .B(n682), .A(n199), .Y(n147) );
  INVX1 U125 ( .A(N1307), .Y(n263) );
  INVX1 U126 ( .A(n574), .Y(n338) );
  INVX1 U127 ( .A(n345), .Y(n680) );
  INVX1 U128 ( .A(n298), .Y(n118) );
  INVX1 U129 ( .A(n327), .Y(n678) );
  XNOR2XL U130 ( .A(n19), .B(n575), .Y(n18) );
  OR2X1 U131 ( .A(n571), .B(n573), .Y(n19) );
  INVX1 U132 ( .A(n73), .Y(n111) );
  INVX1 U133 ( .A(n121), .Y(n206) );
  INVX1 U134 ( .A(n682), .Y(n581) );
  INVX1 U135 ( .A(n487), .Y(n679) );
  INVX1 U136 ( .A(n387), .Y(n567) );
  NAND2X1 U137 ( .A(n574), .B(n671), .Y(n528) );
  NAND2X1 U138 ( .A(n671), .B(n338), .Y(n529) );
  INVX1 U139 ( .A(n306), .Y(n698) );
  INVX1 U140 ( .A(n613), .Y(n686) );
  INVX1 U141 ( .A(n572), .Y(n645) );
  XOR2X1 U142 ( .A(n683), .B(n139), .Y(n142) );
  AOI21BBXL U143 ( .B(n572), .C(n87), .A(n573), .Y(n88) );
  INVX1 U144 ( .A(n199), .Y(n139) );
  INVX1 U145 ( .A(n110), .Y(n328) );
  INVX1 U146 ( .A(n288), .Y(n569) );
  INVX1 U147 ( .A(n386), .Y(n568) );
  INVX1 U148 ( .A(n291), .Y(n677) );
  INVX1 U149 ( .A(n86), .Y(n245) );
  OAI211X1 U150 ( .C(n578), .D(n85), .A(n132), .B(n645), .Y(n86) );
  INVX1 U151 ( .A(n571), .Y(n85) );
  XNOR2XL U152 ( .A(n199), .B(n683), .Y(n20) );
  AND2X1 U153 ( .A(n284), .B(n283), .Y(n301) );
  OAI211X1 U154 ( .C(n227), .D(n534), .A(n226), .B(n225), .Y(ps_ptr[1]) );
  AND2X1 U155 ( .A(n113), .B(n112), .Y(n227) );
  OA222X1 U156 ( .A(n20), .B(n348), .C(n671), .D(n353), .E(n30), .F(n347), .Y(
        n225) );
  OA22X1 U157 ( .A(n41), .B(n395), .C(n728), .D(n394), .Y(n368) );
  OA21XL U158 ( .B(n357), .C(n534), .A(n353), .Y(n358) );
  AND4X1 U159 ( .A(n352), .B(n351), .C(n350), .D(n349), .Y(n357) );
  AND3XL U160 ( .A(n348), .B(n347), .C(n346), .Y(n359) );
  OAI31XL U161 ( .A(n343), .B(n526), .C(n342), .D(n341), .Y(n346) );
  INVX1 U162 ( .A(n340), .Y(n343) );
  NAND21X1 U163 ( .B(n32), .A(n541), .Y(n538) );
  NAND21X1 U164 ( .B(n538), .A(n34), .Y(n547) );
  OR2X1 U165 ( .A(n34), .B(n538), .Y(n550) );
  INVX1 U166 ( .A(n542), .Y(n551) );
  NAND32X1 U167 ( .B(n541), .C(n32), .A(n34), .Y(n542) );
  AND2X1 U168 ( .A(n557), .B(n556), .Y(N1019) );
  AND2X1 U169 ( .A(n552), .B(n557), .Y(N1020) );
  OR2X1 U170 ( .A(n35), .B(n398), .Y(n401) );
  INVX1 U171 ( .A(n372), .Y(n374) );
  AND2X1 U172 ( .A(n539), .B(n543), .Y(N1009) );
  AND2X1 U173 ( .A(n539), .B(n554), .Y(N1010) );
  NAND32XL U174 ( .B(mxcyc_done), .C(semi_start), .A(n152), .Y(n378) );
  INVX1 U175 ( .A(n397), .Y(n400) );
  INVX1 U176 ( .A(n396), .Y(n552) );
  NAND32X1 U177 ( .B(n400), .C(n398), .A(n35), .Y(n396) );
  INVX1 U178 ( .A(n399), .Y(n554) );
  NAND32X1 U179 ( .B(n398), .C(n397), .A(n35), .Y(n399) );
  INVX1 U180 ( .A(n559), .Y(n52) );
  NOR21XL U181 ( .B(n562), .A(n586), .Y(n588) );
  NAND32X1 U182 ( .B(n190), .C(n4), .A(n188), .Y(n473) );
  NAND21X1 U183 ( .B(n582), .A(n559), .Y(n230) );
  INVX1 U184 ( .A(n189), .Y(n562) );
  NAND32X1 U185 ( .B(n584), .C(n231), .A(n2), .Y(n189) );
  INVX1 U186 ( .A(n277), .Y(n685) );
  NOR2X1 U187 ( .A(cs_ptr[0]), .B(cs_ptr[1]), .Y(n653) );
  INVX1 U188 ( .A(n563), .Y(n701) );
  NAND2X1 U189 ( .A(n519), .B(n165), .Y(n351) );
  OAI21BBX1 U190 ( .A(n278), .B(n277), .C(sub_395_S2_I7_aco_carry[4]), .Y(n647) );
  OAI21X1 U191 ( .B(n694), .C(n703), .A(sub_395_S2_I11_aco_carry[4]), .Y(n507)
         );
  OA2222XL U192 ( .A(n350), .B(n678), .C(n330), .D(n259), .E(n107), .F(n351), 
        .G(n349), .H(n106), .Y(n113) );
  INVX1 U193 ( .A(n331), .Y(n106) );
  NAND21X1 U194 ( .B(n247), .A(n246), .Y(n248) );
  AO2222XL U195 ( .A(n291), .B(n287), .C(n430), .D(n290), .E(n342), .F(n244), 
        .G(n526), .H(n243), .Y(n247) );
  OA222X1 U196 ( .A(n245), .B(n351), .C(n6), .D(n340), .E(n37), .F(n352), .Y(
        n246) );
  AOI221X1 U197 ( .A(n499), .B(N1339), .C(N1339), .D(n709), .E(n218), .Y(n54)
         );
  NAND32X1 U198 ( .B(n191), .C(n190), .A(n4), .Y(n336) );
  NOR2X1 U199 ( .A(n706), .B(cs_ptr[0]), .Y(n516) );
  NAND21X1 U200 ( .B(n532), .A(n3), .Y(n101) );
  INVX1 U201 ( .A(N1389), .Y(n696) );
  NOR2X1 U202 ( .A(n582), .B(n53), .Y(n508) );
  NOR2X1 U203 ( .A(cs_ptr[1]), .B(n68), .Y(n631) );
  NOR2X1 U204 ( .A(cs_ptr[1]), .B(n66), .Y(n481) );
  INVX1 U205 ( .A(n260), .Y(N1717) );
  INVX1 U206 ( .A(n501), .Y(n709) );
  INVX1 U207 ( .A(n103), .Y(n109) );
  NAND21X1 U208 ( .B(n104), .A(n105), .Y(n103) );
  OAI22AX1 U209 ( .D(n330), .C(n505), .A(n506), .B(n330), .Y(n504) );
  AOI22X1 U210 ( .A(n692), .B(n144), .C(n507), .D(n662), .Y(n506) );
  AOI32X1 U211 ( .A(n666), .B(n693), .C(n692), .D(n507), .E(n661), .Y(n505) );
  NAND2X1 U212 ( .A(n582), .B(n495), .Y(n499) );
  AOI22X1 U213 ( .A(n692), .B(n669), .C(n507), .D(n664), .Y(n513) );
  NAND2X1 U214 ( .A(n622), .B(n501), .Y(sub_395_S2_I5_aco_carry[4]) );
  NAND2X1 U215 ( .A(n694), .B(n703), .Y(sub_395_S2_I11_aco_carry[4]) );
  NAND2X1 U216 ( .A(n179), .B(n180), .Y(sub_395_S2_I14_aco_carry_4_) );
  INVX1 U217 ( .A(n510), .Y(n694) );
  XOR2X1 U218 ( .A(n69), .B(n180), .Y(n565) );
  INVX1 U219 ( .A(n179), .Y(n69) );
  NAND21X1 U220 ( .B(n495), .A(n582), .Y(n682) );
  OR3XL U221 ( .A(n231), .B(n2), .C(n584), .Y(n424) );
  NAND2X1 U222 ( .A(n104), .B(n105), .Y(n349) );
  AOI221X1 U223 ( .A(n674), .B(N1298), .C(n705), .D(N1298), .E(n210), .Y(n67)
         );
  XNOR2XL U224 ( .A(n463), .B(n464), .Y(n456) );
  NAND2X1 U225 ( .A(n465), .B(n466), .Y(n464) );
  XOR2X1 U226 ( .A(n582), .B(n54), .Y(n175) );
  AOI211X1 U227 ( .C(N1257), .D(n703), .A(n598), .B(n205), .Y(n56) );
  OA21X1 U228 ( .B(n566), .C(n582), .A(N1257), .Y(n598) );
  AOI21AX1 U229 ( .B(n658), .C(N1266), .A(n23), .Y(n22) );
  MUX2IX1 U230 ( .D0(n590), .D1(n591), .S(n234), .Y(n23) );
  OR3XL U231 ( .A(n582), .B(n566), .C(n56), .Y(n385) );
  OA2222XL U232 ( .A(n5), .B(n473), .C(n517), .D(n684), .E(n686), .F(n424), 
        .G(n689), .H(n475), .Y(n283) );
  OAI21X1 U233 ( .B(n622), .C(n501), .A(sub_395_S2_I5_aco_carry[4]), .Y(n613)
         );
  OA2222XL U234 ( .A(n456), .B(n350), .C(n693), .D(n259), .E(n18), .F(n351), 
        .G(n432), .H(n349), .Y(n262) );
  NAND2X1 U235 ( .A(n586), .B(n562), .Y(n484) );
  NAND21X1 U236 ( .B(n231), .A(n584), .Y(n471) );
  INVX1 U237 ( .A(n233), .Y(n271) );
  OAI21X1 U238 ( .B(n621), .C(n495), .A(n232), .Y(n233) );
  NOR2X1 U239 ( .A(n54), .B(n683), .Y(n621) );
  INVX1 U240 ( .A(n622), .Y(n232) );
  XNOR2XL U241 ( .A(n180), .B(n178), .Y(n354) );
  OA222X1 U242 ( .A(n260), .B(n352), .C(n406), .D(n292), .E(n367), .F(n340), 
        .Y(n261) );
  XNOR2XL U243 ( .A(n49), .B(n470), .Y(n463) );
  INVX1 U244 ( .A(N1184), .Y(n681) );
  NOR2X1 U245 ( .A(n499), .B(n493), .Y(n496) );
  INVX1 U246 ( .A(n70), .Y(n578) );
  NOR2X1 U247 ( .A(n682), .B(n55), .Y(n635) );
  NAND21X1 U248 ( .B(n294), .A(n293), .Y(n295) );
  OA222X1 U249 ( .A(n352), .B(n699), .C(n680), .D(n292), .E(n688), .F(n340), 
        .Y(n293) );
  AO2222XL U250 ( .A(n290), .B(n596), .C(n289), .D(n288), .E(n526), .F(n507), 
        .G(n344), .H(n287), .Y(n294) );
  INVX1 U251 ( .A(n532), .Y(n352) );
  INVX1 U252 ( .A(n278), .Y(n700) );
  NAND2X1 U253 ( .A(n469), .B(n466), .Y(n467) );
  NAND2X1 U254 ( .A(n635), .B(n707), .Y(sub_395_S2_aco_carry[4]) );
  INVX1 U255 ( .A(n180), .Y(n711) );
  XNOR2XL U256 ( .A(n559), .B(n683), .Y(n24) );
  INVX1 U257 ( .A(n259), .Y(n526) );
  OAI22X1 U258 ( .A(n497), .B(n487), .C(n498), .D(n679), .Y(n483) );
  AOI22X1 U259 ( .A(n688), .B(n140), .C(n489), .D(n141), .Y(n497) );
  AOI22X1 U260 ( .A(n688), .B(n669), .C(n489), .D(n664), .Y(n498) );
  OAI22AX1 U261 ( .D(n28), .C(n592), .A(n593), .B(n28), .Y(n591) );
  AOI22X1 U262 ( .A(n689), .B(n144), .C(n594), .D(n662), .Y(n592) );
  AOI32X1 U263 ( .A(n666), .B(n690), .C(n689), .D(n594), .E(n661), .Y(n593) );
  OAI22X1 U264 ( .A(n486), .B(n487), .C(n488), .D(n679), .Y(n485) );
  AOI22X1 U265 ( .A(n688), .B(n144), .C(n489), .D(n662), .Y(n488) );
  AOI32X1 U266 ( .A(n367), .B(n666), .C(n688), .D(n489), .E(n661), .Y(n486) );
  INVX1 U267 ( .A(n350), .Y(n287) );
  AOI31X1 U268 ( .A(n666), .B(n681), .C(n5), .D(n661), .Y(n634) );
  NAND2X1 U269 ( .A(n605), .B(n606), .Y(sub_395_S2_I4_aco_carry[4]) );
  INVX1 U270 ( .A(n605), .Y(n705) );
  INVX1 U271 ( .A(n221), .Y(n63) );
  AOI21BBXL U272 ( .B(n576), .C(n575), .A(n49), .Y(n571) );
  NOR2X1 U273 ( .A(n673), .B(n708), .Y(n576) );
  OR2X1 U274 ( .A(n138), .B(n25), .Y(n199) );
  AOI21X1 U275 ( .B(n707), .C(n581), .A(n585), .Y(n25) );
  XOR2X1 U276 ( .A(n131), .B(n87), .Y(n574) );
  MUX4X1 U277 ( .D0(n144), .D1(n662), .D2(n119), .D3(n661), .S0(n118), .S1(
        n117), .Y(n122) );
  AND2X1 U278 ( .A(n666), .B(n268), .Y(n119) );
  OAI21BBX1 U279 ( .A(n120), .B(n278), .C(n26), .Y(n268) );
  XNOR2XL U280 ( .A(n555), .B(n208), .Y(n26) );
  NAND21X1 U281 ( .B(n338), .A(n127), .Y(n387) );
  AO21X1 U282 ( .B(n151), .C(n658), .A(n150), .Y(n200) );
  INVX1 U283 ( .A(n272), .Y(n151) );
  MUX2X1 U284 ( .D0(n149), .D1(n148), .S(n252), .Y(n150) );
  MUX4X1 U285 ( .D0(n664), .D1(n669), .D2(n141), .D3(n140), .S0(n27), .S1(n142), .Y(n149) );
  NAND21X1 U286 ( .B(n15), .A(n116), .Y(n121) );
  AO21X1 U287 ( .B(n125), .C(n658), .A(n124), .Y(n212) );
  INVX1 U288 ( .A(n268), .Y(n125) );
  MUX2X1 U289 ( .D0(n123), .D1(n122), .S(n38), .Y(n124) );
  MUX4X1 U290 ( .D0(n669), .D1(n664), .D2(n140), .D3(n141), .S0(n118), .S1(
        n117), .Y(n123) );
  OAI21BX1 U291 ( .C(n707), .B(n1), .A(n412), .Y(n345) );
  AO21X1 U292 ( .B(n66), .C(n728), .A(n481), .Y(n73) );
  OAI21BX1 U293 ( .C(n566), .B(n508), .A(n510), .Y(n243) );
  XOR2X1 U294 ( .A(n115), .B(n700), .Y(n298) );
  XNOR2XL U295 ( .A(n683), .B(n493), .Y(n487) );
  XNOR2XL U296 ( .A(n147), .B(n707), .Y(n27) );
  OAI21X1 U297 ( .B(n406), .C(n97), .A(n96), .Y(n108) );
  MUX2X1 U298 ( .D0(n403), .D1(n404), .S(n95), .Y(n96) );
  INVX1 U299 ( .A(n244), .Y(n95) );
  AOI22AXL U300 ( .A(n328), .B(n407), .D(n328), .C(n408), .Y(n404) );
  OAI21X1 U301 ( .B(n605), .C(n606), .A(sub_395_S2_I4_aco_carry[4]), .Y(n356)
         );
  AOI21X1 U302 ( .B(n728), .C(n68), .A(n631), .Y(n306) );
  XNOR2XL U303 ( .A(n683), .B(n53), .Y(n330) );
  XNOR2XL U304 ( .A(n577), .B(n49), .Y(n575) );
  NOR2X1 U305 ( .A(n645), .B(n708), .Y(n573) );
  NOR2X1 U306 ( .A(n673), .B(n571), .Y(n572) );
  INVX1 U307 ( .A(n231), .Y(n517) );
  NAND2X1 U308 ( .A(n490), .B(n491), .Y(n367) );
  XNOR2XL U309 ( .A(n492), .B(n493), .Y(n490) );
  NAND2X1 U310 ( .A(n411), .B(n412), .Y(n406) );
  XOR2X1 U311 ( .A(n413), .B(n414), .Y(n411) );
  NAND2X1 U312 ( .A(n467), .B(n468), .Y(n291) );
  OAI21BBX1 U313 ( .A(n466), .B(n728), .C(n578), .Y(n468) );
  XNOR2XL U314 ( .A(n15), .B(n56), .Y(n28) );
  INVX1 U315 ( .A(n116), .Y(n208) );
  INVX1 U316 ( .A(n708), .Y(n87) );
  INVX1 U317 ( .A(n115), .Y(n120) );
  INVX1 U318 ( .A(n594), .Y(n689) );
  INVX1 U319 ( .A(n469), .Y(n674) );
  NAND21X1 U320 ( .B(n585), .A(n139), .Y(n272) );
  NAND21X1 U321 ( .B(n574), .A(n127), .Y(n386) );
  AO21X1 U322 ( .B(n708), .C(n645), .A(n573), .Y(n288) );
  XOR2X1 U323 ( .A(n15), .B(n414), .Y(n110) );
  NAND21X1 U324 ( .B(n1), .A(n94), .Y(n244) );
  AO21X1 U325 ( .B(n414), .C(n15), .A(n93), .Y(n94) );
  INVX1 U326 ( .A(n495), .Y(n93) );
  AOI21X1 U327 ( .B(n683), .C(n495), .A(n635), .Y(n29) );
  OA21X1 U328 ( .B(n683), .C(n116), .A(n121), .Y(n117) );
  MUX2X1 U329 ( .D0(n663), .D1(n668), .S(n569), .Y(n84) );
  INVX1 U330 ( .A(n127), .Y(n671) );
  INVX1 U331 ( .A(n582), .Y(n683) );
  NAND2X1 U332 ( .A(n436), .B(n437), .Y(n432) );
  XOR2X1 U333 ( .A(n438), .B(n439), .Y(n436) );
  INVX1 U334 ( .A(n672), .Y(n311) );
  NOR2X1 U335 ( .A(n706), .B(n71), .Y(n640) );
  INVX1 U336 ( .A(n191), .Y(n188) );
  INVX1 U337 ( .A(n173), .Y(n560) );
  NAND21X1 U338 ( .B(n55), .A(n15), .Y(n173) );
  OAI211X1 U339 ( .C(n578), .D(n72), .A(n132), .B(n673), .Y(n228) );
  INVX1 U340 ( .A(n67), .Y(n72) );
  NOR2X1 U341 ( .A(n493), .B(n683), .Y(n494) );
  INVX1 U342 ( .A(n496), .Y(n78) );
  NOR21XL U343 ( .B(n147), .A(n146), .Y(n252) );
  NOR21XL U344 ( .B(n495), .A(n145), .Y(n146) );
  AND2X1 U345 ( .A(n15), .B(n199), .Y(n145) );
  INVX1 U346 ( .A(N1225), .Y(n264) );
  INVX1 U347 ( .A(n269), .Y(n579) );
  OA222X1 U348 ( .A(n203), .B(n517), .C(n209), .D(n484), .E(n202), .F(n475), 
        .Y(n520) );
  XOR2X1 U349 ( .A(sub_395_S2_I4_aco_carry[5]), .B(n210), .Y(n209) );
  XOR2X1 U350 ( .A(sub_395_S2_I3_aco_carry[5]), .B(n205), .Y(n202) );
  XOR2X1 U351 ( .A(sub_395_S2_I7_aco_carry[5]), .B(n204), .Y(n203) );
  NAND21X1 U352 ( .B(cs_ptr[1]), .A(n70), .Y(n132) );
  INVX1 U353 ( .A(n97), .Y(n658) );
  AOI221XL U354 ( .A(n533), .B(n532), .C(n526), .D(n525), .E(n524), .Y(n535)
         );
  XOR2X1 U355 ( .A(n422), .B(n421), .Y(n533) );
  XOR2X1 U356 ( .A(n423), .B(sub_395_S2_I11_aco_carry[5]), .Y(n525) );
  AOI211X1 U357 ( .C(n521), .D(n520), .A(n519), .B(n518), .Y(n524) );
  AOI21X1 U358 ( .B(n208), .C(n15), .A(n206), .Y(n30) );
  INVX1 U359 ( .A(n704), .Y(n564) );
  INVX1 U360 ( .A(n133), .Y(n251) );
  OAI211X1 U361 ( .C(n50), .D(n578), .A(n132), .B(n131), .Y(n133) );
  XOR2X1 U362 ( .A(sub_395_S2_I5_aco_carry[5]), .B(n218), .Y(n211) );
  INVX1 U363 ( .A(n197), .Y(n423) );
  INVX1 U364 ( .A(n219), .Y(n422) );
  NAND21X1 U365 ( .B(n313), .A(n157), .Y(n159) );
  INVX1 U366 ( .A(n304), .Y(n157) );
  NAND21XL U367 ( .B(wr_dacv[14]), .A(n156), .Y(n313) );
  OAI221X1 U368 ( .A(n364), .B(n363), .C(n362), .D(n361), .E(n360), .Y(
        ps_ptr[0]) );
  MUX2X1 U369 ( .D0(n339), .D1(n337), .S(cs_ptr[0]), .Y(n362) );
  MUX2X1 U370 ( .D0(n359), .D1(n358), .S(cs_ptr[0]), .Y(n360) );
  AOI31X1 U371 ( .A(n335), .B(n334), .C(n333), .D(n332), .Y(n364) );
  INVX1 U372 ( .A(n212), .Y(n224) );
  NAND2X1 U373 ( .A(n216), .B(n214), .Y(n353) );
  OAI211X1 U374 ( .C(n255), .D(n361), .A(n254), .B(n253), .Y(ps_ptr[2]) );
  AND2X1 U375 ( .A(n236), .B(n235), .Y(n255) );
  OA222X1 U376 ( .A(n252), .B(n348), .C(n251), .D(n353), .E(n38), .F(n347), 
        .Y(n253) );
  NOR43X1 U377 ( .B(n285), .C(n323), .D(n33), .A(n31), .Y(n275) );
  OAI21X1 U378 ( .B(n50), .C(n286), .A(n297), .Y(n31) );
  OAI31XL U379 ( .A(n164), .B(n320), .C(n319), .D(n242), .Y(n196) );
  AND3X1 U380 ( .A(n162), .B(n323), .C(n161), .Y(n164) );
  INVX1 U381 ( .A(n322), .Y(n162) );
  NAND32X1 U382 ( .B(n302), .C(n324), .A(n160), .Y(n161) );
  OR3XL U383 ( .A(n304), .B(n237), .C(n313), .Y(n256) );
  NAND21XL U384 ( .B(wr_dacv[9]), .A(n656), .Y(n302) );
  OAI22XL U385 ( .A(n12), .B(ps_ptr[2]), .C(n47), .D(ps_ptr[1]), .Y(n366) );
  NAND32XL U386 ( .B(n41), .C(wr_dacv[17]), .A(n303), .Y(n305) );
  NAND21X1 U387 ( .B(n57), .A(n389), .Y(n372) );
  MUX2IX1 U388 ( .D0(n58), .D1(n389), .S(ps_sample), .Y(n32) );
  OAI211X1 U389 ( .C(n384), .D(n383), .A(n382), .B(n398), .Y(N1002) );
  INVX1 U390 ( .A(n381), .Y(n382) );
  INVX1 U391 ( .A(n366), .Y(n376) );
  INVX1 U392 ( .A(n544), .Y(n541) );
  AND3X1 U393 ( .A(n402), .B(n556), .C(n548), .Y(N1003) );
  OAI32X1 U394 ( .A(n550), .B(n549), .C(n548), .D(n547), .E(n546), .Y(N1013)
         );
  INVX1 U395 ( .A(n405), .Y(n539) );
  NAND32X1 U396 ( .B(n34), .C(n32), .A(n544), .Y(n405) );
  NOR3XL U397 ( .A(n238), .B(n302), .C(n324), .Y(n33) );
  AND2X1 U398 ( .A(n556), .B(n540), .Y(N1011) );
  AND2X1 U399 ( .A(n552), .B(n540), .Y(N1012) );
  INVX1 U400 ( .A(n545), .Y(n557) );
  NAND32X1 U401 ( .B(n34), .C(n544), .A(n32), .Y(n545) );
  INVX1 U402 ( .A(n369), .Y(n373) );
  NAND21X1 U403 ( .B(n10), .A(n388), .Y(n369) );
  MUX2IX1 U404 ( .D0(n10), .D1(n388), .S(ps_sample), .Y(n34) );
  AND3X1 U405 ( .A(n539), .B(n556), .C(n548), .Y(N1007) );
  AND3X1 U406 ( .A(n539), .B(n552), .C(n548), .Y(N1008) );
  MUX2X1 U407 ( .D0(n47), .D1(n394), .S(ps_sample), .Y(n397) );
  NAND21X1 U408 ( .B(n381), .A(n380), .Y(n398) );
  MUX2X1 U409 ( .D0(n379), .D1(n378), .S(ps_sample), .Y(n380) );
  AND2X1 U410 ( .A(sampl_begn), .B(n383), .Y(n379) );
  AND2XL U411 ( .A(n558), .B(ps_ptr[2]), .Y(N1033) );
  OR3XL U412 ( .A(n319), .B(n322), .C(n320), .Y(n257) );
  NAND21X1 U413 ( .B(wr_dacv[6]), .A(n155), .Y(n322) );
  INVX1 U414 ( .A(n239), .Y(n323) );
  INVX1 U415 ( .A(n332), .Y(n250) );
  NOR2X1 U416 ( .A(n220), .B(n724), .Y(N957) );
  NOR2X1 U417 ( .A(n14), .B(n712), .Y(N967) );
  NOR2X1 U418 ( .A(n220), .B(n713), .Y(N969) );
  NOR2X1 U419 ( .A(n14), .B(n714), .Y(N966) );
  NOR2X1 U420 ( .A(n220), .B(n723), .Y(N959) );
  NOR2X1 U421 ( .A(n14), .B(n725), .Y(N956) );
  NOR2X1 U422 ( .A(n220), .B(n716), .Y(N968) );
  NOR2X1 U423 ( .A(n14), .B(n720), .Y(N961) );
  NOR2X1 U424 ( .A(n220), .B(n721), .Y(N960) );
  NOR2X1 U425 ( .A(n14), .B(n715), .Y(N971) );
  NOR2X1 U426 ( .A(n220), .B(n719), .Y(N962) );
  NOR2X1 U427 ( .A(n14), .B(n718), .Y(N963) );
  NOR2X1 U428 ( .A(n220), .B(n722), .Y(N958) );
  NOR2X1 U429 ( .A(n14), .B(n717), .Y(N970) );
  NAND21X1 U430 ( .B(n168), .A(n167), .Y(n559) );
  INVX1 U431 ( .A(n204), .Y(n167) );
  AO21X1 U432 ( .B(N1421), .C(n278), .A(n652), .Y(n168) );
  OA21X1 U433 ( .B(n582), .C(n509), .A(N1421), .Y(n652) );
  AO21X1 U434 ( .B(N1430), .C(n658), .A(n171), .Y(n231) );
  MUX4X1 U435 ( .D0(n649), .D1(n648), .D2(n646), .D3(n644), .S0(n24), .S1(n170), .Y(n171) );
  NAND2X1 U436 ( .A(n511), .B(n512), .Y(n649) );
  OA21X1 U437 ( .B(n566), .C(n169), .A(n277), .Y(n170) );
  NAND21X1 U438 ( .B(n509), .A(n169), .Y(n277) );
  NAND21X1 U439 ( .B(n193), .A(n192), .Y(n194) );
  OA2222XL U440 ( .A(n704), .B(n472), .C(n672), .D(n484), .E(n47), .F(n336), 
        .G(n306), .H(n471), .Y(n192) );
  AO2222XL U441 ( .A(n187), .B(n28), .C(n176), .D(n175), .E(n24), .F(n231), 
        .G(n560), .H(n174), .Y(n193) );
  INVX1 U442 ( .A(n424), .Y(n176) );
  OAI221X1 U443 ( .A(n563), .B(n426), .C(n50), .D(n701), .E(n427), .Y(N1421)
         );
  NOR2X1 U444 ( .A(n587), .B(n653), .Y(n563) );
  INVX1 U445 ( .A(n47), .Y(cs_ptr[1]) );
  OAI31XL U446 ( .A(n647), .B(N1430), .C(n410), .D(n409), .Y(n646) );
  NAND2X1 U447 ( .A(n711), .B(n178), .Y(sub_395_S2_I6_aco_carry[4]) );
  XOR3X1 U448 ( .A(n66), .B(sub_395_S2_I14_aco_carry_4_), .C(n65), .Y(n260) );
  INVX1 U449 ( .A(N1708), .Y(n65) );
  XOR2X1 U450 ( .A(n589), .B(n563), .Y(n278) );
  OAI211X1 U451 ( .C(n41), .D(n587), .A(n482), .B(n636), .Y(n495) );
  NAND3X1 U452 ( .A(cs_ptr[1]), .B(n587), .C(cs_ptr[0]), .Y(n636) );
  AO21X1 U453 ( .B(N1717), .C(n77), .A(n76), .Y(n532) );
  INVX1 U454 ( .A(n431), .Y(n77) );
  MUX2BXL U455 ( .D0(n75), .D1(n74), .S(n37), .Y(n76) );
  MUX2X1 U456 ( .D0(n478), .D1(n477), .S(n111), .Y(n75) );
  INVX1 U457 ( .A(n270), .Y(n695) );
  AOI21X1 U458 ( .B(n629), .C(n698), .A(n630), .Y(n625) );
  EORX1 U459 ( .A(n627), .B(n698), .C(n628), .D(n698), .Y(n626) );
  AO21X1 U460 ( .B(N1594), .C(n658), .A(n82), .Y(n100) );
  MUX2X1 U461 ( .D0(n503), .D1(n504), .S(n81), .Y(n82) );
  INVX1 U462 ( .A(n243), .Y(n81) );
  OAI222XL U463 ( .A(n511), .B(n692), .C(n512), .D(n507), .E(n513), .F(n330), 
        .Y(n503) );
  OA2222XL U464 ( .A(n229), .B(n472), .C(n484), .D(n228), .E(n12), .F(n336), 
        .G(n270), .H(n471), .Y(n236) );
  INVX1 U465 ( .A(n276), .Y(n229) );
  OA2222XL U466 ( .A(n29), .B(n473), .C(n7), .D(n517), .E(n271), .F(n424), .G(
        n234), .H(n475), .Y(n235) );
  INVX1 U467 ( .A(n102), .Y(n105) );
  NAND32X1 U468 ( .B(n101), .C(n100), .A(n99), .Y(n102) );
  OA2222XL U469 ( .A(n264), .B(n472), .C(n263), .D(n484), .E(n51), .F(n336), 
        .G(n696), .H(n471), .Y(n267) );
  OAI21X1 U470 ( .B(n58), .C(n701), .A(n222), .Y(n204) );
  XNOR2XL U471 ( .A(n46), .B(cs_ptr[0]), .Y(n36) );
  INVX1 U472 ( .A(n36), .Y(n582) );
  AOI221XL U473 ( .A(n482), .B(N1708), .C(N1708), .D(n711), .E(n219), .Y(n66)
         );
  AOI221XL U474 ( .A(n482), .B(N1380), .C(N1380), .D(n180), .E(n217), .Y(n68)
         );
  OAI221X1 U475 ( .A(n516), .B(n427), .C(n58), .D(n702), .E(n426), .Y(N1585)
         );
  OAI221X1 U476 ( .A(n426), .B(n710), .C(n50), .D(n502), .E(n427), .Y(N1339)
         );
  NAND2X1 U477 ( .A(n508), .B(n509), .Y(n510) );
  INVX1 U478 ( .A(n57), .Y(n49) );
  NOR2X1 U479 ( .A(n643), .B(n12), .Y(n179) );
  AOI211X1 U480 ( .C(N1585), .D(n514), .A(n515), .B(n197), .Y(n53) );
  OA21X1 U481 ( .B(n566), .C(n582), .A(N1585), .Y(n515) );
  NAND2X1 U482 ( .A(n49), .B(n589), .Y(n426) );
  INVX1 U483 ( .A(n44), .Y(cs_ptr[0]) );
  OAI21X1 U484 ( .B(n58), .C(n502), .A(n222), .Y(n218) );
  INVX1 U485 ( .A(n43), .Y(n41) );
  OAI21X1 U486 ( .B(n303), .C(n687), .A(n618), .Y(n609) );
  OAI21X1 U487 ( .B(n620), .C(n233), .A(n44), .Y(n608) );
  NOR2X1 U488 ( .A(n697), .B(n12), .Y(n178) );
  INVX1 U489 ( .A(n43), .Y(n42) );
  INVX1 U490 ( .A(n57), .Y(n50) );
  OAI22X1 U491 ( .A(n418), .B(n684), .C(n419), .D(n647), .Y(n648) );
  OAI22X1 U492 ( .A(n415), .B(n684), .C(n416), .D(n647), .Y(n644) );
  AOI221XL U493 ( .A(n474), .B(n73), .C(n565), .D(n650), .E(n476), .Y(n74) );
  OAI22X1 U494 ( .A(n440), .B(n699), .C(n442), .D(n565), .Y(n474) );
  NOR3XL U495 ( .A(n565), .B(N1717), .C(n435), .Y(n476) );
  INVX1 U496 ( .A(n447), .Y(n706) );
  AOI31X1 U497 ( .A(n354), .B(n696), .C(n651), .D(n650), .Y(n628) );
  INVX1 U498 ( .A(n435), .Y(n651) );
  INVX1 U499 ( .A(n502), .Y(n710) );
  OAI21X1 U500 ( .B(n221), .C(n222), .A(n223), .Y(N1175) );
  OAI21BBX1 U501 ( .A(n728), .B(n587), .C(n482), .Y(n70) );
  OR2X1 U502 ( .A(n101), .B(n99), .Y(n350) );
  NAND32X1 U503 ( .B(n83), .C(n101), .A(n99), .Y(n259) );
  INVX1 U504 ( .A(n100), .Y(n83) );
  OA2222XL U505 ( .A(n472), .B(n280), .C(n484), .D(n279), .E(n10), .F(n336), 
        .G(n354), .H(n471), .Y(n284) );
  INVX1 U506 ( .A(n355), .Y(n280) );
  INVX1 U507 ( .A(n356), .Y(n279) );
  OAI221X1 U508 ( .A(n599), .B(n561), .C(n431), .D(n263), .E(n600), .Y(n586)
         );
  OAI31XL U509 ( .A(n601), .B(n668), .C(n663), .D(n561), .Y(n600) );
  AOI22X1 U510 ( .A(n672), .B(n602), .C(n311), .D(n603), .Y(n599) );
  INVX1 U511 ( .A(n228), .Y(n561) );
  INVX1 U512 ( .A(n172), .Y(n55) );
  NAND32X1 U513 ( .B(n682), .C(n223), .A(n707), .Y(n172) );
  OAI21X1 U514 ( .B(n691), .C(n514), .A(sub_395_S2_I3_aco_carry[4]), .Y(n594)
         );
  XNOR2XL U515 ( .A(n607), .B(n49), .Y(N1298) );
  OAI21X1 U516 ( .B(n469), .C(n463), .A(n58), .Y(n466) );
  AND2X1 U517 ( .A(n500), .B(n222), .Y(n493) );
  OAI21X1 U518 ( .B(n501), .C(n499), .A(n492), .Y(n500) );
  OAI221X1 U519 ( .A(n426), .B(n702), .C(n50), .D(n516), .E(n427), .Y(N1257)
         );
  NOR2X1 U520 ( .A(n46), .B(n578), .Y(n469) );
  NOR2X1 U521 ( .A(n607), .B(n470), .Y(n605) );
  INVX1 U522 ( .A(n580), .Y(n707) );
  NOR2X1 U523 ( .A(n222), .B(n516), .Y(n197) );
  NOR2X1 U524 ( .A(n222), .B(n587), .Y(n219) );
  OAI221X1 U525 ( .A(n502), .B(n427), .C(n58), .D(n710), .E(n426), .Y(n492) );
  OAI21X1 U526 ( .B(n58), .C(n587), .A(n222), .Y(n217) );
  OR2X1 U527 ( .A(n446), .B(n44), .Y(n221) );
  INVX1 U528 ( .A(n509), .Y(n566) );
  INVX1 U529 ( .A(n514), .Y(n703) );
  OAI21X1 U530 ( .B(n440), .C(n354), .A(n442), .Y(n627) );
  OAI22X1 U531 ( .A(n675), .B(n665), .C(n670), .D(n344), .Y(n455) );
  OAI22X1 U532 ( .A(n444), .B(n699), .C(n445), .D(n565), .Y(n478) );
  OAI22X1 U533 ( .A(n479), .B(n699), .C(n480), .D(n565), .Y(n477) );
  OAI21X1 U534 ( .B(n444), .C(n354), .A(n445), .Y(n629) );
  OAI31XL U535 ( .A(n356), .B(N1307), .C(n435), .D(n604), .Y(n602) );
  NOR2X1 U536 ( .A(n589), .B(n447), .Y(n470) );
  NAND2X1 U537 ( .A(n691), .B(n514), .Y(sub_395_S2_I3_aco_carry[4]) );
  NOR2X1 U538 ( .A(n607), .B(n58), .Y(n210) );
  AOI221XL U539 ( .A(N1184), .B(n658), .C(n29), .D(n633), .E(n664), .Y(n632)
         );
  OAI211X1 U540 ( .C(n634), .D(n560), .A(n415), .B(n416), .Y(n633) );
  NAND21X1 U541 ( .B(n126), .A(n577), .Y(n708) );
  AO21X1 U542 ( .B(n555), .C(n114), .A(n138), .Y(n116) );
  NAND32X1 U543 ( .B(n509), .C(n15), .A(n278), .Y(n114) );
  NAND21X1 U544 ( .B(n47), .A(n578), .Y(n673) );
  MUX4X1 U545 ( .D0(n662), .D1(n144), .D2(n661), .D3(n143), .S0(n27), .S1(n142), .Y(n148) );
  INVX1 U546 ( .A(n416), .Y(n144) );
  NAND21X1 U547 ( .B(n509), .A(n206), .Y(n115) );
  OAI221X1 U548 ( .A(n92), .B(n245), .C(n431), .D(n18), .E(n91), .Y(n519) );
  AOI21X1 U549 ( .B(n570), .C(n89), .A(n84), .Y(n92) );
  MUX4X1 U550 ( .D0(n604), .D1(n440), .D2(n90), .D3(n442), .S0(n89), .S1(n88), 
        .Y(n91) );
  INVX1 U551 ( .A(n107), .Y(n89) );
  AOI21X1 U552 ( .B(n12), .C(n697), .A(n178), .Y(n270) );
  OR2X1 U553 ( .A(n51), .B(n673), .Y(n131) );
  NAND21X1 U554 ( .B(n435), .A(n18), .Y(n90) );
  NAND2X1 U555 ( .A(n1), .B(n580), .Y(n412) );
  OAI221X1 U556 ( .A(n701), .B(n427), .C(n58), .D(n563), .E(n426), .Y(n555) );
  OAI21X1 U557 ( .B(n51), .C(n516), .A(n222), .Y(n205) );
  OAI211X1 U558 ( .C(n50), .D(n221), .A(n426), .B(n427), .Y(n413) );
  AOI222XL U559 ( .A(n328), .B(n417), .C(n680), .D(n140), .E(n345), .F(n141), 
        .Y(n403) );
  OAI21X1 U560 ( .B(n418), .C(n680), .A(n419), .Y(n417) );
  AOI21X1 U561 ( .B(n12), .C(n643), .A(n179), .Y(n37) );
  INVX1 U562 ( .A(sub_395_S2_aco_carry[4]), .Y(n281) );
  INVX1 U563 ( .A(n635), .Y(n282) );
  NAND2X1 U564 ( .A(n425), .B(n51), .Y(n414) );
  OAI21X1 U565 ( .B(n682), .C(n707), .A(n413), .Y(n425) );
  OAI22AX1 U566 ( .D(n406), .C(n410), .A(n409), .B(n680), .Y(n408) );
  NAND2X1 U567 ( .A(n589), .B(n446), .Y(n577) );
  OAI21X1 U568 ( .B(n415), .C(n680), .A(n416), .Y(n407) );
  AOI21X1 U569 ( .B(n479), .C(n480), .A(n698), .Y(n630) );
  AOI21X1 U570 ( .B(n511), .C(n512), .A(n28), .Y(n597) );
  NOR21XL U571 ( .B(n607), .A(n49), .Y(n71) );
  XOR2X1 U572 ( .A(n46), .B(n49), .Y(n127) );
  XOR2X1 U573 ( .A(n46), .B(n67), .Y(n672) );
  XOR2X1 U574 ( .A(n46), .B(n571), .Y(n107) );
  NOR21XL U575 ( .B(n385), .A(n166), .Y(n234) );
  AOI21BBXL U576 ( .B(n56), .C(n15), .A(n509), .Y(n166) );
  OAI21X1 U577 ( .B(n432), .C(n431), .A(n98), .Y(n104) );
  MUX2X1 U578 ( .D0(n429), .D1(n428), .S(n430), .Y(n98) );
  AOI221XL U579 ( .A(n331), .B(n433), .C(n596), .D(n650), .E(n434), .Y(n429)
         );
  AOI222XL U580 ( .A(n331), .B(n443), .C(n441), .D(n668), .E(n596), .F(n663), 
        .Y(n428) );
  OAI221X1 U581 ( .A(n637), .B(n276), .C(n431), .D(n264), .E(n638), .Y(n191)
         );
  OAI31XL U582 ( .A(n639), .B(n668), .C(n663), .D(n276), .Y(n638) );
  AOI22X1 U583 ( .A(n704), .B(n641), .C(n564), .D(n603), .Y(n637) );
  AOI21X1 U584 ( .B(n444), .C(n445), .A(n704), .Y(n639) );
  INVX1 U585 ( .A(n441), .Y(n596) );
  INVX1 U586 ( .A(n223), .Y(n585) );
  NAND2X1 U587 ( .A(n222), .B(n448), .Y(n438) );
  OAI21X1 U588 ( .B(n589), .C(n706), .A(n439), .Y(n448) );
  OAI22X1 U589 ( .A(n444), .B(n441), .C(n445), .D(n596), .Y(n443) );
  OAI22X1 U590 ( .A(n440), .B(n441), .C(n442), .D(n596), .Y(n433) );
  OAI21X1 U591 ( .B(n444), .C(n569), .A(n445), .Y(n570) );
  OAI31XL U592 ( .A(n355), .B(N1225), .C(n435), .D(n604), .Y(n641) );
  NAND2X1 U593 ( .A(n447), .B(n438), .Y(n437) );
  NOR21XL U594 ( .B(n272), .A(n410), .Y(n143) );
  AOI21X1 U595 ( .B(n444), .C(n445), .A(n672), .Y(n601) );
  NOR3XL U596 ( .A(n596), .B(n435), .C(n595), .Y(n434) );
  INVX1 U597 ( .A(n432), .Y(n595) );
  NAND2X1 U598 ( .A(n640), .B(n589), .Y(sub_395_S2_I2_aco_carry[4]) );
  NAND2X1 U599 ( .A(n427), .B(n426), .Y(n439) );
  INVX1 U600 ( .A(n222), .Y(n138) );
  NAND21X1 U601 ( .B(n49), .A(n126), .Y(n269) );
  XNOR2XL U602 ( .A(n46), .B(n438), .Y(n331) );
  OAI21X1 U603 ( .B(n640), .C(n589), .A(sub_395_S2_I2_aco_carry[4]), .Y(n355)
         );
  INVX1 U604 ( .A(n410), .Y(n666) );
  OAI211X1 U605 ( .C(n12), .D(n438), .A(n437), .B(n446), .Y(n430) );
  INVX1 U606 ( .A(n409), .Y(n661) );
  INVX1 U607 ( .A(n419), .Y(n669) );
  INVX1 U608 ( .A(n418), .Y(n664) );
  AOI21X1 U609 ( .B(n121), .C(n509), .A(n120), .Y(n38) );
  INVX1 U610 ( .A(n415), .Y(n662) );
  INVX1 U611 ( .A(n604), .Y(n650) );
  MUX2X1 U612 ( .D0(n303), .D1(n308), .S(cs_ptr[0]), .Y(n97) );
  NAND21X1 U613 ( .B(n71), .A(n46), .Y(n704) );
  NAND21X1 U614 ( .B(n640), .A(n446), .Y(n276) );
  OA2222XL U615 ( .A(n215), .B(n473), .C(n207), .D(n472), .E(n213), .F(n471), 
        .G(n211), .H(n424), .Y(n521) );
  XNOR2XL U616 ( .A(sub_395_S2_I2_aco_carry[5]), .B(n51), .Y(n207) );
  XNOR2XL U617 ( .A(sub_395_S2_aco_carry[5]), .B(n585), .Y(n215) );
  XOR2X1 U618 ( .A(sub_395_S2_I6_aco_carry[5]), .B(n217), .Y(n213) );
  INVX1 U619 ( .A(n511), .Y(n141) );
  INVX1 U620 ( .A(n512), .Y(n140) );
  INVX1 U621 ( .A(n479), .Y(n663) );
  INVX1 U622 ( .A(n480), .Y(n668) );
  NAND2X1 U623 ( .A(n440), .B(n442), .Y(n603) );
  INVX1 U624 ( .A(n57), .Y(cs_ptr[4]) );
  INVX1 U625 ( .A(sampl_done), .Y(n383) );
  AND2X1 U626 ( .A(n57), .B(n10), .Y(n391) );
  NAND4X1 U627 ( .A(n725), .B(n714), .C(n712), .D(n716), .Y(n184) );
  NOR4XL U628 ( .A(n181), .B(n182), .C(n183), .D(n184), .Y(sh_hold) );
  NAND4X1 U629 ( .A(n724), .B(n722), .C(n723), .D(n721), .Y(n182) );
  NAND4X1 U630 ( .A(n720), .B(n719), .C(n186), .D(n718), .Y(n181) );
  OR2XL U631 ( .A(wr_dacv[15]), .B(r_dac_en[15]), .Y(n304) );
  INVX1 U632 ( .A(n319), .Y(n321) );
  OAI31XL U633 ( .A(n318), .B(wr_dacv[11]), .C(n8), .D(n317), .Y(n325) );
  AND3X1 U634 ( .A(n654), .B(n316), .C(n315), .Y(n318) );
  OAI211X1 U635 ( .C(n314), .D(n313), .A(n312), .B(n310), .Y(n315) );
  INVX1 U636 ( .A(r_dac_en[13]), .Y(n312) );
  INVXL U637 ( .A(wr_dacv[13]), .Y(n310) );
  NAND43X1 U638 ( .B(r_dac_en[17]), .C(r_dac_en[16]), .D(wr_dacv[17]), .A(n309), .Y(n286) );
  NAND43X1 U639 ( .B(wr_dacv[12]), .C(wr_dacv[13]), .D(r_dac_en[13]), .A(n654), 
        .Y(n237) );
  OR2XL U640 ( .A(wr_dacv[8]), .B(r_dac_en[8]), .Y(n324) );
  NAND21X1 U641 ( .B(n371), .A(n372), .Y(n420) );
  OA22X1 U642 ( .A(n49), .B(n389), .C(n370), .D(n373), .Y(n371) );
  OA222X1 U643 ( .A(n368), .B(n366), .C(n11), .D(n365), .E(cs_ptr[3]), .F(n388), .Y(n370) );
  INVXL U644 ( .A(ps_ptr[2]), .Y(n365) );
  OR2X1 U645 ( .A(n239), .B(n257), .Y(n240) );
  AOI21BX1 U646 ( .C(r_loop), .B(n420), .A(r_semi), .Y(n536) );
  MUX2IX1 U647 ( .D0(cs_mux_5_), .D1(n39), .S(n558), .Y(n537) );
  OAI22XL U648 ( .A(cs_mux_5_), .B(n536), .C(n535), .D(n534), .Y(n39) );
  AO21X1 U649 ( .B(n539), .C(r_comp_swtch), .A(n553), .Y(n540) );
  AO21X1 U650 ( .B(ps_md4ch), .C(n393), .A(n392), .Y(n544) );
  MUX2X1 U651 ( .D0(n391), .D1(n390), .S(ps_sample), .Y(n393) );
  AO21XL U652 ( .B(stop), .C(n377), .A(n177), .Y(n381) );
  INVX1 U653 ( .A(ps_sample), .Y(n377) );
  INVX1 U654 ( .A(n60), .Y(n558) );
  NAND32X1 U655 ( .B(n59), .C(n62), .A(n61), .Y(n60) );
  INVX1 U656 ( .A(n378), .Y(n59) );
  AO21X1 U657 ( .B(n62), .C(n61), .A(n558), .Y(N1030) );
  OR2X1 U658 ( .A(wr_dacv[5]), .B(r_dac_en[5]), .Y(n319) );
  OR2X1 U659 ( .A(wr_dacv[1]), .B(r_dac_en[1]), .Y(n332) );
  OR2X1 U660 ( .A(wr_dacv[4]), .B(r_dac_en[4]), .Y(n320) );
  OR2X1 U661 ( .A(wr_dacv[7]), .B(r_dac_en[7]), .Y(n239) );
  INVX1 U662 ( .A(n163), .Y(n242) );
  NAND43X1 U663 ( .B(r_dac_en[2]), .C(wr_dacv[3]), .D(wr_dacv[2]), .A(n657), 
        .Y(n163) );
  NAND2X1 U664 ( .A(sampl_done), .B(srstz), .Y(n220) );
  INVX1 U665 ( .A(cs_mux_5_), .Y(busy) );
  NOR21XL U666 ( .B(pos_dacis[17]), .A(n220), .Y(N973) );
  NOR21XL U667 ( .B(pos_dacis[16]), .A(n14), .Y(N972) );
  NOR21XL U668 ( .B(pos_dacis[8]), .A(n220), .Y(N964) );
  NOR21XL U669 ( .B(pos_dacis[9]), .A(n14), .Y(N965) );
  OR2X1 U670 ( .A(neg_dacis_9_), .B(pos_dacis[9]), .Y(app_dacis[9]) );
  OR2X1 U671 ( .A(neg_dacis_8_), .B(pos_dacis[8]), .Y(app_dacis[8]) );
  OR2X1 U672 ( .A(neg_dacis_2_), .B(pos_dacis[2]), .Y(app_dacis[2]) );
  OR2X1 U673 ( .A(neg_dacis_3_), .B(pos_dacis[3]), .Y(app_dacis[3]) );
  OR2X1 U674 ( .A(neg_dacis_10_), .B(pos_dacis[10]), .Y(app_dacis[10]) );
  OR2X1 U675 ( .A(neg_dacis_7_), .B(pos_dacis[7]), .Y(app_dacis[7]) );
  OR2X1 U676 ( .A(neg_dacis_5_), .B(pos_dacis[5]), .Y(app_dacis[5]) );
  OR2X1 U677 ( .A(neg_dacis_13_), .B(pos_dacis[13]), .Y(app_dacis[13]) );
  OR2X1 U678 ( .A(neg_dacis_15_), .B(pos_dacis[15]), .Y(app_dacis[15]) );
  OR2X1 U679 ( .A(neg_dacis_6_), .B(pos_dacis[6]), .Y(app_dacis[6]) );
  OR2X1 U680 ( .A(neg_dacis_0_), .B(pos_dacis[0]), .Y(app_dacis[0]) );
  OR2X1 U681 ( .A(neg_dacis_1_), .B(pos_dacis[1]), .Y(app_dacis[1]) );
  OR2X1 U682 ( .A(test_so1), .B(pos_dacis[17]), .Y(app_dacis[17]) );
  OR2X1 U683 ( .A(neg_dacis_11_), .B(pos_dacis[11]), .Y(app_dacis[11]) );
  OR2X1 U684 ( .A(neg_dacis_12_), .B(pos_dacis[12]), .Y(app_dacis[12]) );
  OR2X1 U685 ( .A(neg_dacis_14_), .B(pos_dacis[14]), .Y(app_dacis[14]) );
  OR2X1 U686 ( .A(neg_dacis_4_), .B(pos_dacis[4]), .Y(app_dacis[4]) );
  OR2X1 U687 ( .A(neg_dacis_16_), .B(pos_dacis[16]), .Y(app_dacis[16]) );
  INVX1 U688 ( .A(pos_dacis[14]), .Y(n717) );
  INVX1 U689 ( .A(pos_dacis[2]), .Y(n722) );
  INVX1 U690 ( .A(pos_dacis[7]), .Y(n718) );
  INVX1 U691 ( .A(pos_dacis[6]), .Y(n719) );
  INVX1 U692 ( .A(pos_dacis[15]), .Y(n715) );
  INVX1 U693 ( .A(pos_dacis[4]), .Y(n721) );
  INVX1 U694 ( .A(pos_dacis[12]), .Y(n716) );
  INVX1 U695 ( .A(pos_dacis[5]), .Y(n720) );
  INVX1 U696 ( .A(pos_dacis[0]), .Y(n725) );
  INVX1 U697 ( .A(pos_dacis[3]), .Y(n723) );
  INVX1 U698 ( .A(pos_dacis[10]), .Y(n714) );
  INVX1 U699 ( .A(pos_dacis[13]), .Y(n713) );
  INVX1 U700 ( .A(pos_dacis[11]), .Y(n712) );
  INVX1 U701 ( .A(pos_dacis[1]), .Y(n724) );
  INVX1 U702 ( .A(n728), .Y(n47) );
  OAI22X1 U703 ( .A(n41), .B(n482), .C(n653), .D(cs_ptr[2]), .Y(n509) );
  OAI221X1 U704 ( .A(n587), .B(n427), .C(cs_ptr[2]), .D(n58), .E(n426), .Y(
        N1708) );
  AOI21X1 U705 ( .B(n728), .C(n42), .A(cs_ptr[2]), .Y(n502) );
  INVX1 U706 ( .A(n727), .Y(n589) );
  INVX1 U707 ( .A(cs_ptr[2]), .Y(n587) );
  NAND2X1 U708 ( .A(n727), .B(n49), .Y(n222) );
  NOR2X1 U709 ( .A(cs_ptr[1]), .B(cs_ptr[2]), .Y(n447) );
  OAI221X1 U710 ( .A(cs_ptr[2]), .B(n426), .C(n50), .D(n587), .E(n427), .Y(
        N1380) );
  NAND2X1 U711 ( .A(cs_ptr[2]), .B(n46), .Y(n482) );
  NAND2X1 U712 ( .A(n727), .B(n51), .Y(n427) );
  INVX1 U713 ( .A(n728), .Y(n46) );
  AOI32X1 U714 ( .A(n307), .B(n687), .C(r_dac_en[0]), .D(n175), .E(r_dac_en[2]), .Y(n616) );
  INVX1 U715 ( .A(n726), .Y(n51) );
  OAI2B11X1 U716 ( .D(r_dac_en[16]), .C(n687), .A(n611), .B(n41), .Y(n610) );
  OAI32X1 U717 ( .A(n612), .B(r_dac_en[8]), .C(n686), .D(n613), .E(n614), .Y(
        n611) );
  OAI22X1 U718 ( .A(n271), .B(n617), .C(n655), .D(n307), .Y(n612) );
  OAI22X1 U719 ( .A(n271), .B(n615), .C(n616), .D(n233), .Y(n614) );
  INVX1 U720 ( .A(n726), .Y(n57) );
  AOI22X1 U721 ( .A(n175), .B(n623), .C(n307), .D(n624), .Y(n620) );
  OAI21BBX1 U722 ( .A(n613), .B(n8), .C(n657), .Y(n623) );
  OAI31XL U723 ( .A(n613), .B(N1348), .C(n667), .D(n656), .Y(n624) );
  INVX1 U724 ( .A(n729), .Y(n43) );
  INVX1 U725 ( .A(n729), .Y(n44) );
  XOR2X1 U726 ( .A(n63), .B(n727), .Y(n580) );
  AO21X1 U727 ( .B(n727), .C(n63), .A(n50), .Y(n223) );
  OR2X1 U728 ( .A(n450), .B(n449), .Y(n99) );
  AOI221XL U729 ( .A(n457), .B(n458), .C(n642), .D(r_dac_en[16]), .E(n41), .Y(
        n449) );
  AOI211X1 U730 ( .C(n642), .D(r_dac_en[17]), .A(n451), .B(n44), .Y(n450) );
  INVX1 U731 ( .A(n456), .Y(n642) );
  NAND2X1 U732 ( .A(cs_ptr[1]), .B(cs_ptr[2]), .Y(n446) );
  NOR2X1 U733 ( .A(n706), .B(n727), .Y(n607) );
  OAI222XL U734 ( .A(n452), .B(n678), .C(n453), .D(n327), .E(n677), .F(n454), 
        .Y(n451) );
  AOI22X1 U735 ( .A(n675), .B(r_dac_en[3]), .C(n8), .D(n344), .Y(n452) );
  AOI32X1 U736 ( .A(n456), .B(r_dac_en[1]), .C(n675), .D(r_dac_en[9]), .E(n344), .Y(n453) );
  AOI222XL U737 ( .A(n327), .B(n455), .C(n675), .D(r_dac_en[5]), .E(
        r_dac_en[13]), .F(n344), .Y(n454) );
  AOI21X1 U738 ( .B(n175), .C(r_dac_en[6]), .A(r_dac_en[4]), .Y(n615) );
  AOI21X1 U739 ( .B(n175), .C(r_dac_en[14]), .A(r_dac_en[12]), .Y(n617) );
  INVX1 U740 ( .A(n726), .Y(n58) );
  GEN2XL U742 ( .D(n729), .E(n137), .C(r_dac_en[16]), .B(n579), .A(n136), .Y(
        n216) );
  INVX1 U743 ( .A(n303), .Y(n137) );
  MUX2X1 U744 ( .D0(n135), .D1(n134), .S(n251), .Y(n136) );
  OAI221X1 U745 ( .A(n529), .B(n659), .C(n523), .D(n43), .E(n130), .Y(n134) );
  GEN2XL U746 ( .D(n665), .E(n670), .C(n307), .B(n619), .A(n271), .Y(n618) );
  OAI21X1 U747 ( .B(r_dac_en[5]), .C(r_dac_en[13]), .A(n307), .Y(n619) );
  OAI22BX1 U748 ( .B(r_dac_en[5]), .A(n528), .D(r_dac_en[13]), .C(n529), .Y(
        n530) );
  INVX1 U749 ( .A(n64), .Y(n126) );
  NAND21X1 U750 ( .B(n446), .A(n727), .Y(n64) );
  OAI221X1 U751 ( .A(n386), .B(n156), .C(n387), .D(n155), .E(n128), .Y(n135)
         );
  AOI21BX1 U752 ( .C(n522), .B(n41), .A(n531), .Y(n128) );
  OAI22AX1 U753 ( .D(r_dac_en[4]), .C(n528), .A(n654), .B(n529), .Y(n531) );
  AOI221XL U754 ( .A(n568), .B(r_dac_en[15]), .C(n567), .D(r_dac_en[7]), .E(
        n530), .Y(n522) );
  AOI221XL U755 ( .A(n568), .B(n8), .C(n567), .D(r_dac_en[3]), .E(n527), .Y(
        n523) );
  OAI32X1 U756 ( .A(n528), .B(n579), .C(n667), .D(n656), .E(n529), .Y(n527) );
  OAI211X1 U757 ( .C(n677), .D(n461), .A(n675), .B(n462), .Y(n457) );
  AOI21X1 U758 ( .B(r_dac_en[6]), .C(n327), .A(r_dac_en[4]), .Y(n461) );
  AOI32X1 U759 ( .A(n456), .B(r_dac_en[0]), .C(n678), .D(r_dac_en[2]), .E(n327), .Y(n462) );
  OAI211X1 U760 ( .C(n659), .D(n327), .A(n344), .B(n459), .Y(n458) );
  AOI22X1 U761 ( .A(r_dac_en[10]), .B(n327), .C(n460), .D(n291), .Y(n459) );
  OAI21BBX1 U762 ( .A(n327), .B(r_dac_en[14]), .C(n654), .Y(n460) );
  XNOR2XL U763 ( .A(n437), .B(n727), .Y(n441) );
  NAND2X1 U764 ( .A(r_dac_en[0]), .B(n269), .Y(n129) );
  AOI22X1 U765 ( .A(n42), .B(r_dac_en[12]), .C(n44), .D(n9), .Y(n511) );
  AOI22X1 U766 ( .A(n729), .B(r_dac_en[4]), .C(n44), .D(r_dac_en[5]), .Y(n512)
         );
  AOI22X1 U767 ( .A(n42), .B(r_dac_en[6]), .C(n44), .D(r_dac_en[7]), .Y(n419)
         );
  AOI22X1 U768 ( .A(n42), .B(r_dac_en[10]), .C(n44), .D(n8), .Y(n415) );
  AOI22X1 U769 ( .A(n729), .B(r_dac_en[2]), .C(n44), .D(r_dac_en[3]), .Y(n416)
         );
  AOI22X1 U770 ( .A(n42), .B(r_dac_en[8]), .C(n43), .D(r_dac_en[9]), .Y(n409)
         );
  AOI22X1 U771 ( .A(n729), .B(r_dac_en[14]), .C(n43), .D(r_dac_en[15]), .Y(
        n418) );
  AOI22X1 U772 ( .A(n42), .B(r_dac_en[0]), .C(n43), .D(r_dac_en[1]), .Y(n410)
         );
  AOI22X1 U773 ( .A(cs_ptr[0]), .B(r_dac_en[1]), .C(n44), .D(r_dac_en[0]), .Y(
        n435) );
  AOI22X1 U774 ( .A(cs_ptr[0]), .B(r_dac_en[9]), .C(n43), .D(r_dac_en[8]), .Y(
        n604) );
  AOI21X1 U775 ( .B(n42), .C(r_dac_en[13]), .A(r_dac_en[12]), .Y(n479) );
  AOI21X1 U776 ( .B(n42), .C(r_dac_en[5]), .A(r_dac_en[4]), .Y(n480) );
  AOI21X1 U777 ( .B(n42), .C(r_dac_en[3]), .A(r_dac_en[2]), .Y(n442) );
  AOI21X1 U778 ( .B(n41), .C(n8), .A(r_dac_en[10]), .Y(n440) );
  AOI21X1 U779 ( .B(n41), .C(r_dac_en[15]), .A(r_dac_en[14]), .Y(n444) );
  AOI22X1 U780 ( .A(n729), .B(r_dac_en[7]), .C(n43), .D(r_dac_en[6]), .Y(n445)
         );
  AOI22X1 U781 ( .A(n729), .B(r_dac_en[17]), .C(n43), .D(r_dac_en[16]), .Y(
        n431) );
  INVX1 U782 ( .A(r_dac_en[17]), .Y(n303) );
  INVX1 U783 ( .A(r_dac_en[12]), .Y(n654) );
  INVX1 U784 ( .A(r_dac_en[9]), .Y(n656) );
  INVX1 U785 ( .A(r_dac_en[10]), .Y(n655) );
  INVX1 U786 ( .A(r_dac_en[15]), .Y(n665) );
  INVX1 U787 ( .A(r_dac_en[7]), .Y(n670) );
  INVX1 U788 ( .A(r_dac_en[3]), .Y(n657) );
  INVX1 U789 ( .A(r_dac_en[16]), .Y(n308) );
  INVX1 U790 ( .A(r_dac_en[1]), .Y(n667) );
  INVX1 U791 ( .A(r_dac_en[8]), .Y(n659) );
  INVX1 U792 ( .A(r_dac_en[2]), .Y(n334) );
  INVX1 U793 ( .A(r_dac_en[14]), .Y(n156) );
  INVX1 U794 ( .A(r_dac_en[6]), .Y(n155) );
  NAND4X1 U795 ( .A(n713), .B(n717), .C(n185), .D(n715), .Y(n183) );
  NOR2X1 U796 ( .A(pos_dacis[17]), .B(pos_dacis[16]), .Y(n185) );
  NOR2X1 U797 ( .A(pos_dacis[9]), .B(pos_dacis[8]), .Y(n186) );
  INVX1 U798 ( .A(r_comp_swtch), .Y(n548) );
  AND2XL U799 ( .A(n558), .B(ps_ptr[4]), .Y(N1035) );
  INVXL U800 ( .A(ps_ptr[4]), .Y(n389) );
  AND2XL U801 ( .A(n558), .B(ps_ptr[1]), .Y(N1032) );
  INVXL U802 ( .A(ps_ptr[1]), .Y(n394) );
  AOI32XL U803 ( .A(n250), .B(n249), .C(n17), .D(n341), .E(n248), .Y(n254) );
  AO21XL U804 ( .B(n267), .C(n266), .A(n361), .Y(n274) );
  MUX2XL U805 ( .D0(n11), .D1(ps_ptr[2]), .S(ps_sample), .Y(n392) );
  NAND43X1 U806 ( .B(wr_dacv[10]), .C(wr_dacv[11]), .D(n8), .A(n655), .Y(n238)
         );
  NAND32X2 U807 ( .B(n519), .C(n534), .A(n165), .Y(n361) );
  INVXL U808 ( .A(n258), .Y(n297) );
  NAND21X4 U809 ( .B(n200), .A(n201), .Y(n154) );
  AOI32X1 U810 ( .A(n198), .B(n250), .C(n196), .D(n195), .E(n194), .Y(n226) );
  INVX8 U811 ( .A(srstz), .Y(n62) );
  NAND32X4 U812 ( .B(n212), .C(n216), .A(n214), .Y(n534) );
  MAJ3X1 U813 ( .A(sub_395_S2_I14_aco_carry_4_), .B(n66), .C(N1708), .Y(n421)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dac2sar_a0 ( r_dac_t, r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, 
        auto_sar, busy, stop, sync_i, sampl_begn, sampl_done, sh_rst, 
        dacyc_done, sacyc_done, dac_v, rpt_v, clk, srstz, test_si2, test_si1, 
        test_so1, test_se );
  input [1:0] r_dac_t;
  output [9:0] dac_v;
  output [9:0] rpt_v;
  input r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, auto_sar, busy, stop,
         sync_i, clk, srstz, test_si2, test_si1, test_se;
  output sampl_begn, sampl_done, sh_rst, dacyc_done, sacyc_done, test_so1;
  wire   N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N60, N61, N62, N63, N64, N68, updlo, updup, upd1v, r_lt_up_8_,
         r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, r_lt_up_3_,
         r_lt_up_2_, r_lt_up_1_, r_lt_up_0_, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         net10186, net10192, n133, n24, n25, n26, n27, n11, n19, n20, n21, n22,
         n23, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n57, n58, n59, n60, n61, n62, n63, n64, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n1, n2, n4, n5, n6, n10, n12, n13, n14, n15, n16,
         n17, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3;
  wire   [6:0] dacnt;
  wire   [3:0] sarcyc;
  wire   [9:0] r_lt_lo;
  wire   [9:0] r_avg00;
  wire   [9:0] r_avgup;
  wire   [9:0] r_dacvo;

  INVX1 U33 ( .A(n27), .Y(n25) );
  INVX1 U34 ( .A(n27), .Y(n26) );
  INVX1 U35 ( .A(srstz), .Y(n27) );
  INVX1 U36 ( .A(n27), .Y(n24) );
  glreg_WIDTH10_2 u0_dac1v ( .clk(clk), .arstz(n26), .we(upd1v), .wdat(r_dacvo), .rdat({dac_v[9:1], n133}), .test_si(sarcyc[3]), .test_se(test_se) );
  glreg_WIDTH10_1 u0_lt_lo ( .clk(clk), .arstz(n25), .we(updlo), .wdat({n13, 
        n14, n12, n115, n114, n1, n15, n113, n112, n16}), .rdat(r_lt_lo), 
        .test_si(dac_v[9]), .test_se(test_se) );
  glreg_WIDTH10_0 u0_lt_up ( .clk(clk), .arstz(n24), .we(updup), .wdat(r_avgup), .rdat({test_so1, r_lt_up_8_, r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, 
        r_lt_up_3_, r_lt_up_2_, r_lt_up_1_, r_lt_up_0_}), .test_si(r_lt_lo[9]), 
        .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 clk_gate_dacnt_reg ( .CLK(clk), .EN(N43), 
        .ENCLK(net10186), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 clk_gate_sarcyc_reg ( .CLK(clk), .EN(N60), 
        .ENCLK(net10192), .TE(test_se) );
  dac2sar_a0_DW01_add_0 add_303 ( .A({1'b0, n19, n21, n23, n29, n31, n33, n35, 
        n37, n39, n41}), .B({1'b0, n11, n20, n22, n28, n30, n32, n34, n36, n38, 
        n40}), .CI(1'b0), .SUM({N91, N90, N89, N88, N87, N86, N85, N84, N83, 
        N82, SYNOPSYS_UNCONNECTED_1}), .CO() );
  dac2sar_a0_DW01_add_2 add_296 ( .A({1'b0, r_lt_lo}), .B({1'b0, test_so1, 
        r_lt_up_8_, r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, r_lt_up_3_, 
        r_lt_up_2_, r_lt_up_1_, r_lt_up_0_}), .CI(1'b0), .SUM({r_avg00, 
        SYNOPSYS_UNCONNECTED_2}), .CO() );
  dac2sar_a0_DW01_inc_0 add_276 ( .A(dacnt), .SUM({N42, N41, N40, N39, N38, 
        N37, N36}) );
  dac2sar_a0_DW01_add_1 add_301 ( .A({1'b0, n13, n14, n12, n115, n114, n1, n15, 
        n113, n112, n16}), .B({1'b0, r_avgup}), .CI(1'b0), .SUM({N80, N79, N78, 
        N77, N76, N75, N74, N73, N72, N71, SYNOPSYS_UNCONNECTED_3}), .CO() );
  SDFFQX1 sarcyc_reg_2_ ( .D(N63), .SIN(sarcyc[1]), .SMC(test_se), .C(net10192), .Q(sarcyc[2]) );
  SDFFNQX1 sh_rst_n_reg ( .D(N68), .SIN(test_si1), .SMC(test_se), .XC(clk), 
        .Q(sh_rst) );
  SDFFQX1 sarcyc_reg_1_ ( .D(N62), .SIN(sarcyc[0]), .SMC(test_se), .C(net10192), .Q(sarcyc[1]) );
  SDFFQX1 sarcyc_reg_0_ ( .D(N61), .SIN(dacnt[6]), .SMC(test_se), .C(net10192), 
        .Q(sarcyc[0]) );
  SDFFQX1 dacnt_reg_1_ ( .D(N45), .SIN(dacnt[0]), .SMC(test_se), .C(net10186), 
        .Q(dacnt[1]) );
  SDFFQX1 dacnt_reg_2_ ( .D(N46), .SIN(dacnt[1]), .SMC(test_se), .C(net10186), 
        .Q(dacnt[2]) );
  SDFFQX1 sarcyc_reg_3_ ( .D(N64), .SIN(sarcyc[2]), .SMC(test_se), .C(net10192), .Q(sarcyc[3]) );
  SDFFQX1 dacnt_reg_0_ ( .D(N44), .SIN(test_si2), .SMC(test_se), .C(net10186), 
        .Q(dacnt[0]) );
  SDFFQX1 dacnt_reg_6_ ( .D(N50), .SIN(dacnt[5]), .SMC(test_se), .C(net10186), 
        .Q(dacnt[6]) );
  SDFFQX1 dacnt_reg_3_ ( .D(N47), .SIN(dacnt[2]), .SMC(test_se), .C(net10186), 
        .Q(dacnt[3]) );
  SDFFQX1 dacnt_reg_4_ ( .D(N48), .SIN(dacnt[3]), .SMC(test_se), .C(net10186), 
        .Q(dacnt[4]) );
  SDFFQX1 dacnt_reg_5_ ( .D(N49), .SIN(dacnt[4]), .SMC(test_se), .C(net10186), 
        .Q(dacnt[5]) );
  MUX2X2 U6 ( .D0(N78), .D1(r_avg00[7]), .S(n5), .Y(r_dacvo[7]) );
  MUX2X2 U7 ( .D0(N79), .D1(r_avg00[8]), .S(n5), .Y(r_dacvo[8]) );
  NAND21X1 U8 ( .B(n30), .A(n55), .Y(r_avgup[5]) );
  INVX1 U9 ( .A(n70), .Y(n114) );
  INVX1 U10 ( .A(n68), .Y(n115) );
  INVX1 U11 ( .A(n88), .Y(n112) );
  MUX2X1 U12 ( .D0(N76), .D1(r_avg00[5]), .S(semi_nxt), .Y(r_dacvo[5]) );
  MUX2X1 U13 ( .D0(N77), .D1(r_avg00[6]), .S(semi_nxt), .Y(r_dacvo[6]) );
  MUX2X1 U14 ( .D0(N75), .D1(r_avg00[4]), .S(semi_nxt), .Y(r_dacvo[4]) );
  MUX2X1 U15 ( .D0(N80), .D1(r_avg00[9]), .S(semi_nxt), .Y(r_dacvo[9]) );
  NOR2X1 U16 ( .A(sar_ini), .B(n80), .Y(n1) );
  INVXL U17 ( .A(n133), .Y(n2) );
  INVXL U18 ( .A(n2), .Y(dac_v[0]) );
  INVXL U19 ( .A(n2), .Y(n4) );
  BUFX3 U20 ( .A(semi_nxt), .Y(n5) );
  INVX1 U21 ( .A(n10), .Y(n6) );
  INVX2 U22 ( .A(sar_ini), .Y(n55) );
  BUFXL U23 ( .A(sar_ini), .Y(n10) );
  NAND2X1 U24 ( .A(n120), .B(n55), .Y(r_avgup[4]) );
  NAND2X1 U25 ( .A(n117), .B(n55), .Y(r_avgup[1]) );
  NAND2XL U26 ( .A(n55), .B(n39), .Y(n88) );
  MUX2X1 U27 ( .D0(N73), .D1(r_avg00[2]), .S(semi_nxt), .Y(r_dacvo[2]) );
  NAND2XL U28 ( .A(n116), .B(n55), .Y(r_avgup[0]) );
  NOR2XL U29 ( .A(sar_ini), .B(n81), .Y(n15) );
  NOR2XL U30 ( .A(sar_ini), .B(n84), .Y(n16) );
  NAND2XL U31 ( .A(n118), .B(n55), .Y(r_avgup[2]) );
  NAND2XL U32 ( .A(n119), .B(n55), .Y(r_avgup[3]) );
  NAND2XL U37 ( .A(n123), .B(n6), .Y(r_avgup[7]) );
  OR3XL U38 ( .A(sar_nxt), .B(n10), .C(semi_nxt), .Y(upd1v) );
  INVX1 U39 ( .A(n95), .Y(n99) );
  INVX1 U40 ( .A(n98), .Y(n110) );
  INVX1 U41 ( .A(n90), .Y(n91) );
  OR2X1 U42 ( .A(n99), .B(n52), .Y(N60) );
  MUX2X1 U43 ( .D0(N71), .D1(r_avg00[0]), .S(semi_nxt), .Y(r_dacvo[0]) );
  OR2XL U44 ( .A(sar_ini), .B(n78), .Y(n68) );
  NAND2XL U45 ( .A(n125), .B(n6), .Y(r_avgup[9]) );
  NAND2XL U46 ( .A(n124), .B(n6), .Y(r_avgup[8]) );
  NOR2XL U47 ( .A(sar_ini), .B(n77), .Y(n12) );
  NOR2XL U48 ( .A(n10), .B(n75), .Y(n13) );
  NOR2XL U49 ( .A(sar_ini), .B(n76), .Y(n14) );
  MUX2X1 U50 ( .D0(N74), .D1(r_avg00[3]), .S(semi_nxt), .Y(r_dacvo[3]) );
  NAND21XL U51 ( .B(sar_ini), .A(n31), .Y(n70) );
  NAND2XL U52 ( .A(n122), .B(n55), .Y(r_avgup[6]) );
  MUX2X1 U53 ( .D0(N72), .D1(r_avg00[1]), .S(semi_nxt), .Y(r_dacvo[1]) );
  NOR2X1 U54 ( .A(n64), .B(n130), .Y(sampl_begn) );
  NAND32X1 U55 ( .B(n53), .C(n52), .A(auto_sar), .Y(n95) );
  OR2X1 U56 ( .A(sacyc_done), .B(n54), .Y(n52) );
  NAND21X1 U57 ( .B(n100), .A(n99), .Y(n98) );
  NAND31X1 U58 ( .C(n54), .A(busy), .B(n53), .Y(n90) );
  AND2X1 U59 ( .A(n99), .B(n97), .Y(N61) );
  AND2X1 U60 ( .A(N39), .B(n91), .Y(N47) );
  AND2X1 U61 ( .A(N38), .B(n91), .Y(N46) );
  AND2X1 U62 ( .A(N41), .B(n91), .Y(N49) );
  AND2X1 U63 ( .A(N40), .B(n91), .Y(N48) );
  AND2X1 U64 ( .A(N37), .B(n91), .Y(N45) );
  NAND32X1 U65 ( .B(dacyc_done), .C(n54), .A(n90), .Y(N43) );
  NAND21X1 U66 ( .B(n105), .A(n106), .Y(n60) );
  XNOR2XL U67 ( .A(n132), .B(n106), .Y(n62) );
  INVX1 U68 ( .A(n107), .Y(n127) );
  NOR32XL U69 ( .B(busy), .C(n130), .A(n64), .Y(N68) );
  INVX1 U70 ( .A(n82), .Y(n37) );
  INVX1 U71 ( .A(n118), .Y(n36) );
  INVX1 U72 ( .A(n81), .Y(n35) );
  INVX1 U73 ( .A(n119), .Y(n34) );
  INVX1 U74 ( .A(n80), .Y(n33) );
  INVX1 U75 ( .A(n120), .Y(n32) );
  INVX1 U76 ( .A(n79), .Y(n31) );
  INVX1 U77 ( .A(n121), .Y(n30) );
  INVX1 U78 ( .A(n78), .Y(n29) );
  INVX1 U79 ( .A(n122), .Y(n28) );
  INVX1 U80 ( .A(n123), .Y(n22) );
  INVX1 U81 ( .A(n77), .Y(n23) );
  INVX1 U82 ( .A(n124), .Y(n20) );
  INVX1 U83 ( .A(n76), .Y(n21) );
  INVX1 U84 ( .A(n75), .Y(n19) );
  INVX1 U85 ( .A(n125), .Y(n11) );
  INVX1 U86 ( .A(r_avg00[9]), .Y(n56) );
  INVX1 U87 ( .A(r_avg00[8]), .Y(n65) );
  INVX1 U88 ( .A(r_avg00[0]), .Y(n89) );
  INVX1 U89 ( .A(r_avg00[1]), .Y(n87) );
  INVX1 U90 ( .A(r_avg00[2]), .Y(n73) );
  INVX1 U91 ( .A(r_avg00[3]), .Y(n72) );
  INVX1 U92 ( .A(r_avg00[4]), .Y(n71) );
  INVX1 U93 ( .A(r_avg00[5]), .Y(n69) );
  INVX1 U94 ( .A(r_avg00[6]), .Y(n67) );
  INVX1 U95 ( .A(r_avg00[7]), .Y(n66) );
  INVX1 U96 ( .A(n83), .Y(n39) );
  INVX1 U97 ( .A(n117), .Y(n38) );
  INVX1 U98 ( .A(n116), .Y(n40) );
  INVX1 U99 ( .A(n84), .Y(n41) );
  INVX1 U100 ( .A(n53), .Y(dacyc_done) );
  INVX1 U101 ( .A(n46), .Y(n45) );
  INVX1 U102 ( .A(n46), .Y(n44) );
  AOI22X1 U103 ( .A(n85), .B(n127), .C(n126), .D(n128), .Y(n109) );
  INVX1 U104 ( .A(n85), .Y(n126) );
  NAND21XL U105 ( .B(stop), .A(n26), .Y(n54) );
  MUX2X1 U106 ( .D0(n111), .D1(n110), .S(sarcyc[2]), .Y(N63) );
  AND2X1 U107 ( .A(n100), .B(n99), .Y(n111) );
  ENOX1 U108 ( .A(dac_v[0]), .B(n123), .C(N89), .D(n4), .Y(rpt_v[7]) );
  ENOX1 U109 ( .A(n4), .B(n121), .C(N87), .D(n4), .Y(rpt_v[5]) );
  ENOX1 U110 ( .A(n4), .B(n116), .C(N82), .D(n133), .Y(rpt_v[0]) );
  ENOX1 U111 ( .A(n133), .B(n117), .C(N83), .D(dac_v[0]), .Y(rpt_v[1]) );
  ENOX1 U112 ( .A(n133), .B(n119), .C(N85), .D(dac_v[0]), .Y(rpt_v[3]) );
  ENOX1 U113 ( .A(dac_v[0]), .B(n120), .C(N86), .D(n4), .Y(rpt_v[4]) );
  ENOX1 U114 ( .A(n4), .B(n118), .C(N84), .D(n4), .Y(rpt_v[2]) );
  ENOX1 U115 ( .A(dac_v[0]), .B(n122), .C(N88), .D(dac_v[0]), .Y(rpt_v[6]) );
  ENOX1 U116 ( .A(dac_v[0]), .B(n124), .C(N90), .D(n4), .Y(rpt_v[8]) );
  ENOX1 U117 ( .A(n4), .B(n125), .C(n4), .D(N91), .Y(rpt_v[9]) );
  OA21X1 U118 ( .B(sarcyc[1]), .C(sarcyc[0]), .A(n110), .Y(N62) );
  OAI22X1 U119 ( .A(n96), .B(n95), .C(n98), .D(n94), .Y(N64) );
  MUX2BXL U120 ( .D0(n94), .D1(n93), .S(sarcyc[2]), .Y(n96) );
  AND2X1 U121 ( .A(n100), .B(n94), .Y(n93) );
  AND2X1 U122 ( .A(N36), .B(n91), .Y(N44) );
  AND2X1 U123 ( .A(N42), .B(n91), .Y(N50) );
  AOI21BBXL U124 ( .B(r_dac_t[0]), .C(n105), .A(n107), .Y(n106) );
  NOR41XL U125 ( .D(dacnt[1]), .A(n57), .B(n58), .C(n59), .Y(sampl_done) );
  XNOR2XL U126 ( .A(n127), .B(dacnt[2]), .Y(n58) );
  XNOR2XL U127 ( .A(n60), .B(dacnt[6]), .Y(n59) );
  NAND4X1 U128 ( .A(n61), .B(n62), .C(n63), .D(n130), .Y(n57) );
  XNOR2XL U129 ( .A(n104), .B(dacnt[4]), .Y(n63) );
  OAI21X1 U130 ( .B(r_dac_t[0]), .C(n105), .A(n60), .Y(n104) );
  NOR2X1 U131 ( .A(r_dac_t[1]), .B(n105), .Y(n107) );
  NOR2X1 U132 ( .A(r_dac_t[0]), .B(r_dac_t[1]), .Y(n105) );
  XNOR2XL U133 ( .A(n60), .B(dacnt[5]), .Y(n61) );
  INVX1 U134 ( .A(dacnt[3]), .Y(n132) );
  NOR4XL U135 ( .A(sarcyc[0]), .B(sarcyc[1]), .C(sarcyc[2]), .D(sarcyc[3]), 
        .Y(n85) );
  NAND42X1 U136 ( .C(dacnt[2]), .D(dacnt[1]), .A(n85), .B(n86), .Y(n64) );
  NOR4XL U137 ( .A(dacnt[6]), .B(dacnt[5]), .C(dacnt[4]), .D(dacnt[3]), .Y(n86) );
  INVX1 U138 ( .A(dacnt[0]), .Y(n130) );
  MUX2BXL U139 ( .D0(n87), .D1(r_lt_up_1_), .S(n45), .Y(n117) );
  MUX2BXL U140 ( .D0(n67), .D1(r_lt_up_6_), .S(n45), .Y(n122) );
  MUX2BXL U141 ( .D0(n73), .D1(r_lt_up_2_), .S(n45), .Y(n118) );
  MUX2BXL U142 ( .D0(n72), .D1(r_lt_up_3_), .S(n45), .Y(n119) );
  MUX2BXL U143 ( .D0(n71), .D1(r_lt_up_4_), .S(n45), .Y(n120) );
  MUX2BXL U144 ( .D0(n69), .D1(r_lt_up_5_), .S(n45), .Y(n121) );
  MUX2BXL U145 ( .D0(n66), .D1(r_lt_up_7_), .S(n45), .Y(n123) );
  MUX2BXL U146 ( .D0(n65), .D1(r_lt_up_8_), .S(n45), .Y(n124) );
  MUX2BXL U147 ( .D0(n56), .D1(test_so1), .S(n44), .Y(n125) );
  MUX2BXL U148 ( .D0(n89), .D1(r_lt_up_0_), .S(n45), .Y(n116) );
  MUX2AXL U149 ( .D0(r_lt_lo[0]), .D1(n89), .S(n45), .Y(n84) );
  MUX2AXL U150 ( .D0(r_lt_lo[1]), .D1(n87), .S(n44), .Y(n83) );
  MUX2AXL U151 ( .D0(r_lt_lo[2]), .D1(n73), .S(n44), .Y(n82) );
  MUX2AXL U152 ( .D0(r_lt_lo[3]), .D1(n72), .S(n44), .Y(n81) );
  MUX2AXL U153 ( .D0(r_lt_lo[4]), .D1(n71), .S(n44), .Y(n80) );
  MUX2AXL U154 ( .D0(r_lt_lo[5]), .D1(n69), .S(n44), .Y(n79) );
  MUX2AXL U155 ( .D0(r_lt_lo[6]), .D1(n67), .S(n44), .Y(n78) );
  MUX2AXL U156 ( .D0(r_lt_lo[7]), .D1(n66), .S(n44), .Y(n77) );
  MUX2AXL U157 ( .D0(r_lt_lo[8]), .D1(n65), .S(n44), .Y(n76) );
  MUX2AXL U158 ( .D0(r_lt_lo[9]), .D1(n56), .S(n44), .Y(n75) );
  NAND42X1 U159 ( .C(n50), .D(n102), .A(n49), .B(n48), .Y(n53) );
  AND2X1 U160 ( .A(dacnt[6]), .B(dacnt[5]), .Y(n50) );
  NOR32XL U161 ( .B(dacnt[0]), .C(dacnt[1]), .A(n47), .Y(n49) );
  XNOR2XL U162 ( .A(n109), .B(dacnt[2]), .Y(n48) );
  NOR32XL U163 ( .B(dacyc_done), .C(sarcyc[0]), .A(n17), .Y(n51) );
  XNOR2XL U164 ( .A(n94), .B(r_sar10), .Y(n17) );
  AND3X1 U165 ( .A(n42), .B(n43), .C(n51), .Y(sacyc_done) );
  XOR2X1 U166 ( .A(sarcyc[1]), .B(r_sar10), .Y(n42) );
  XOR2X1 U167 ( .A(sarcyc[2]), .B(r_sar10), .Y(n43) );
  AOI31X1 U168 ( .A(n62), .B(n63), .C(n103), .D(n126), .Y(n102) );
  EORX1 U169 ( .A(n60), .B(n131), .C(n60), .D(dacnt[6]), .Y(n103) );
  INVX1 U170 ( .A(dacnt[5]), .Y(n131) );
  INVX1 U171 ( .A(sync_i), .Y(n46) );
  AND2X1 U172 ( .A(n101), .B(n126), .Y(n47) );
  OAI221X1 U173 ( .A(n129), .B(n132), .C(dacnt[4]), .D(n128), .E(n108), .Y(
        n101) );
  INVX1 U174 ( .A(dacnt[4]), .Y(n129) );
  AOI211X1 U175 ( .C(n132), .D(n128), .A(dacnt[6]), .B(dacnt[5]), .Y(n108) );
  INVX1 U176 ( .A(r_dacyc), .Y(n128) );
  INVX1 U177 ( .A(sarcyc[3]), .Y(n94) );
  INVX1 U178 ( .A(n92), .Y(n100) );
  NAND21X1 U179 ( .B(n97), .A(sarcyc[1]), .Y(n92) );
  INVX1 U180 ( .A(sarcyc[0]), .Y(n97) );
  INVX1 U181 ( .A(n74), .Y(n113) );
  NAND21XL U182 ( .B(sar_ini), .A(n37), .Y(n74) );
  AO21XL U183 ( .B(sar_nxt), .C(sync_i), .A(n10), .Y(updlo) );
  AO21XL U184 ( .B(sar_nxt), .C(n46), .A(n10), .Y(updup) );
endmodule


module dac2sar_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n6, n7, n8, n9, n10, n18, n19, n21, n23, n24, n26, n27, n28, n29,
         n30, n32, n33, n34, n37, n39, n40, n45, n46, n49, n50, n51, n56, n57,
         n58, n59, n60, n63, n64, n65, n68, n70, n71, n72, n73, n74, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130;

  AOI21X1 U25 ( .B(n27), .C(n40), .A(n28), .Y(n26) );
  OAI21X1 U27 ( .B(n29), .C(n37), .A(n30), .Y(n28) );
  NOR2X1 U40 ( .A(A[6]), .B(B[6]), .Y(n34) );
  XOR2X1 U71 ( .A(n117), .B(n8), .Y(SUM[2]) );
  XOR2X1 U77 ( .A(n9), .B(n65), .Y(SUM[1]) );
  AO21X1 U88 ( .B(n129), .C(n39), .A(n40), .Y(n123) );
  AO21X1 U89 ( .B(n129), .C(n71), .A(n49), .Y(n121) );
  AO21X1 U90 ( .B(n129), .C(n32), .A(n33), .Y(n126) );
  OAI21X1 U91 ( .B(n45), .C(n51), .A(n46), .Y(n40) );
  NOR2XL U92 ( .A(n50), .B(n45), .Y(n39) );
  NOR2X1 U93 ( .A(A[1]), .B(B[1]), .Y(n63) );
  NOR2XL U94 ( .A(n34), .B(n29), .Y(n27) );
  NOR2X1 U95 ( .A(A[7]), .B(B[7]), .Y(n29) );
  NAND2X1 U96 ( .A(A[4]), .B(B[4]), .Y(n51) );
  OR2X1 U97 ( .A(n59), .B(n56), .Y(n116) );
  NOR2X1 U98 ( .A(A[2]), .B(B[2]), .Y(n59) );
  AND2X1 U99 ( .A(n119), .B(n120), .Y(n113) );
  AND2X1 U100 ( .A(n39), .B(n27), .Y(n114) );
  OAI21BBX1 U101 ( .A(n129), .B(n114), .C(n26), .Y(n24) );
  NAND2X1 U102 ( .A(A[1]), .B(B[1]), .Y(n64) );
  OAI21BX1 U103 ( .C(n40), .B(n34), .A(n37), .Y(n33) );
  NAND2XL U104 ( .A(A[8]), .B(B[8]), .Y(n23) );
  AOI21BBX1 U105 ( .B(n63), .C(n65), .A(n118), .Y(n117) );
  NOR21XL U106 ( .B(n39), .A(n34), .Y(n32) );
  OR2X1 U107 ( .A(A[8]), .B(B[8]), .Y(n119) );
  OAI21X1 U108 ( .B(n117), .C(n59), .A(n60), .Y(n58) );
  XNOR2XL U109 ( .A(n7), .B(n58), .Y(SUM[3]) );
  INVX1 U110 ( .A(n64), .Y(n118) );
  INVXL U111 ( .A(n50), .Y(n71) );
  NAND2XL U112 ( .A(A[7]), .B(B[7]), .Y(n30) );
  OR2X2 U113 ( .A(A[9]), .B(B[9]), .Y(n120) );
  NAND2XL U114 ( .A(A[9]), .B(B[9]), .Y(n18) );
  NAND2XL U115 ( .A(n119), .B(n23), .Y(n2) );
  AND2XL U116 ( .A(n68), .B(n30), .Y(n127) );
  XOR2XL U117 ( .A(n126), .B(n127), .Y(SUM[7]) );
  XOR2XL U118 ( .A(n121), .B(n122), .Y(SUM[5]) );
  XOR2XL U119 ( .A(n123), .B(n124), .Y(SUM[6]) );
  OAI21BBX1 U120 ( .A(n120), .B(n21), .C(n18), .Y(n115) );
  INVX1 U121 ( .A(n29), .Y(n68) );
  OAI21X1 U122 ( .B(n116), .C(n117), .A(n130), .Y(n129) );
  INVX1 U123 ( .A(n23), .Y(n21) );
  INVXL U124 ( .A(n51), .Y(n49) );
  NOR2XL U125 ( .A(A[4]), .B(B[4]), .Y(n50) );
  NOR2X2 U126 ( .A(A[5]), .B(B[5]), .Y(n45) );
  NAND2X1 U127 ( .A(A[2]), .B(B[2]), .Y(n60) );
  OR2XL U128 ( .A(A[6]), .B(B[6]), .Y(n128) );
  NAND2XL U129 ( .A(A[5]), .B(B[5]), .Y(n46) );
  NAND2XL U130 ( .A(A[6]), .B(B[6]), .Y(n37) );
  NAND2X1 U131 ( .A(A[3]), .B(B[3]), .Y(n57) );
  NAND2X1 U132 ( .A(A[0]), .B(B[0]), .Y(n65) );
  AND2XL U133 ( .A(n70), .B(n46), .Y(n122) );
  AND2XL U134 ( .A(n128), .B(n37), .Y(n124) );
  XNOR2X1 U135 ( .A(n19), .B(n125), .Y(SUM[9]) );
  AND2XL U136 ( .A(n120), .B(n18), .Y(n125) );
  NAND2XL U137 ( .A(n74), .B(n64), .Y(n9) );
  INVXL U138 ( .A(n63), .Y(n74) );
  NAND2XL U139 ( .A(n72), .B(n57), .Y(n7) );
  XNOR2XL U140 ( .A(n6), .B(n129), .Y(SUM[4]) );
  NAND2XL U141 ( .A(n71), .B(n51), .Y(n6) );
  NAND2XL U142 ( .A(n73), .B(n60), .Y(n8) );
  INVXL U143 ( .A(n59), .Y(n73) );
  INVX1 U144 ( .A(n45), .Y(n70) );
  INVX1 U145 ( .A(n56), .Y(n72) );
  NOR2X1 U146 ( .A(A[3]), .B(B[3]), .Y(n56) );
  XNOR2XL U147 ( .A(n2), .B(n24), .Y(SUM[8]) );
  AOI21XL U148 ( .B(n24), .C(n113), .A(n115), .Y(n10) );
  AOI21X1 U149 ( .B(n24), .C(n119), .A(n21), .Y(n19) );
  OA21X1 U150 ( .B(n56), .C(n60), .A(n57), .Y(n130) );
  INVXL U151 ( .A(n10), .Y(SUM[10]) );
endmodule


module dac2sar_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module dac2sar_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module dac2sar_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10209;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10209), .TE(test_se) );
  SDFFRQXL mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10209), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10227;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10227), .TE(test_se) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10227), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10245;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10245), .TE(test_se) );
  SDFFRQXL mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[9]) );
  SDFFRQXL mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[8]) );
  SDFFRQXL mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[7]) );
  SDFFRQXL mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[4]) );
  SDFFRQXL mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[6]) );
  SDFFRQXL mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[5]) );
  SDFFRQXL mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[2]) );
  SDFFRQXL mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[3]) );
  SDFFRQXL mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[0]) );
  SDFFRQXL mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10245), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_00000012 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [17:0] wdat;
  output [17:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10263, n1, n2, n3;

  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(arstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_glreg_00000012 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10263), .TE(test_se) );
  SDFFRQX1 mem_reg_14_ ( .D(wdat[14]), .SIN(rdat[13]), .SMC(test_se), .C(
        net10263), .XR(n1), .Q(rdat[14]) );
  SDFFRQX1 mem_reg_11_ ( .D(wdat[11]), .SIN(rdat[10]), .SMC(test_se), .C(
        net10263), .XR(n1), .Q(rdat[11]) );
  SDFFRQX1 mem_reg_10_ ( .D(wdat[10]), .SIN(rdat[9]), .SMC(test_se), .C(
        net10263), .XR(n1), .Q(rdat[10]) );
  SDFFRQX1 mem_reg_16_ ( .D(wdat[16]), .SIN(rdat[15]), .SMC(test_se), .C(
        net10263), .XR(n1), .Q(rdat[16]) );
  SDFFRQX1 mem_reg_17_ ( .D(wdat[17]), .SIN(rdat[16]), .SMC(test_se), .C(
        net10263), .XR(n1), .Q(rdat[17]) );
  SDFFRQX1 mem_reg_13_ ( .D(wdat[13]), .SIN(rdat[12]), .SMC(test_se), .C(
        net10263), .XR(n1), .Q(rdat[13]) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10263), .XR(n1), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_12_ ( .D(wdat[12]), .SIN(rdat[11]), .SMC(test_se), .C(
        net10263), .XR(n1), .Q(rdat[12]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10263), .XR(n1), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10263), .XR(n2), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10263), .XR(n2), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10263), .XR(n2), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10263), .XR(n2), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10263), .XR(n2), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10263), .XR(n2), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10263), .XR(n2), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10263), .XR(n2), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_15_ ( .D(wdat[15]), .SIN(rdat[14]), .SMC(test_se), .C(
        net10263), .XR(n1), .Q(rdat[15]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_00000012 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( i_cc, i_cc_49, i_sqlch, r_sqlch, 
        r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, 
        r_fiforst, r_unlock, r_first, r_last, r_set_cpmsgid, r_rdy, r_wdat, 
        r_rdat, r_txnumk, r_txendk, r_txshrt, r_auto_discard, r_txauto, 
        r_rxords_ena, r_spec, r_dat_spec, r_auto_gdcrc, r_rxdb_opt, r_pshords, 
        r_dat_portrole, r_dat_datarole, r_discard, pid_goidle, pid_gobusy, 
        pff_ack, pff_rdat, pff_rxpart, prx_rcvinf, pff_obsd, pff_ptr, 
        pff_empty, pff_full, ptx_ack, ptx_cc, ptx_oe, prx_setsta, prx_rst, 
        prl_c0set, prl_cany0, prl_cany0r, prl_cany0w, prl_discard, 
        prl_GCTxDone, prl_cany0adr, prl_cpmsgid, prx_fifowdat, ptx_fsm, 
        prl_fsm, prx_fsm, prx_adpn, dbgpo, clk, srstz, test_si, test_so, 
        test_se );
  input [1:0] r_sqlch;
  input [7:0] r_wdat;
  input [7:0] r_rdat;
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [6:0] r_rxords_ena;
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [1:0] r_auto_gdcrc;
  input [1:0] r_rxdb_opt;
  output [1:0] pff_ack;
  output [7:0] pff_rdat;
  output [15:0] pff_rxpart;
  output [4:0] prx_rcvinf;
  output [5:0] pff_ptr;
  output [6:0] prx_setsta;
  output [1:0] prx_rst;
  output [7:0] prl_cany0adr;
  output [2:0] prl_cpmsgid;
  output [7:0] prx_fifowdat;
  output [2:0] ptx_fsm;
  output [3:0] prl_fsm;
  output [3:0] prx_fsm;
  output [5:0] prx_adpn;
  output [31:0] dbgpo;
  input i_cc, i_cc_49, i_sqlch, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4,
         r_fifopsh, r_fifopop, r_fiforst, r_unlock, r_first, r_last,
         r_set_cpmsgid, r_rdy, r_txendk, r_txshrt, r_auto_discard, r_pshords,
         r_dat_portrole, r_dat_datarole, r_discard, clk, srstz, test_si,
         test_se;
  output pid_goidle, pid_gobusy, pff_obsd, pff_empty, pff_full, ptx_ack,
         ptx_cc, ptx_oe, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_discard, prl_GCTxDone, test_so;
  wire   n107, rx_pshords, auto_rx_gdcrc, prx_trans, prx_fiforst, pcc_rxgood,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd, x_trans, ptx_goidle,
         c0_txendk, mux_one, ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4,
         crcstart, crcshfi4, crcshfo4, prl_idle, lockena, fifosrstz,
         fifopop_pff, fifopsh_pff, pff_txreq, pff_one, obsd, prl_last,
         prl_txreq, fifopop_prl, fifopsh_prl, prx_gdmsgrcvd, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, d_sqlch, net10281, n106, n58, n59, n60,
         n61, n55, n56, n57, n62, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n4, n6, n7, n10, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n63, n64, n65, n66, n67, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;
  wire   [1:0] prx_cccnt;
  wire   [3:0] prx_crcsidat;
  wire   [4:0] c0_txnumk;
  wire   [6:0] c0_txauto;
  wire   [7:0] mux_rdat;
  wire   [3:0] ptx_crcsidat;
  wire   [3:0] crc32_3_0;
  wire   [3:0] crcsidat;
  wire   [55:0] pff_dat_7_1;
  wire   [47:16] pff_c0dat;
  wire   [7:0] prl_rdat;
  wire   [4:0] prl_txauto;
  wire   [1:0] d_cc;
  wire   [8:0] cclow_cnt;

  phyrx_a0 u0_phyrx ( .i_cc(i_cc), .ptx_txact(n6), .r_adprx_en(r_adprx_en), 
        .r_adp2nd(r_adp2nd), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), 
        .r_rxdb_opt(r_rxdb_opt), .r_ords_ena(r_rxords_ena), .r_pshords(
        rx_pshords), .r_rgdcrc(auto_rx_gdcrc), .prx_cccnt(prx_cccnt), 
        .prx_rst(prx_rst), .prx_setsta({prx_setsta[6:1], 
        SYNOPSYS_UNCONNECTED_1}), .prx_idle(), .prx_d_cc(prx_rcvinf[3]), 
        .prx_bmc(dbgpo[18]), .prx_trans(prx_trans), .prx_fiforst(prx_fiforst), 
        .prx_fifopsh(dbgpo[29]), .prx_fifowdat(prx_fifowdat), .pff_txreq(n10), 
        .pid_gobusy(pid_gobusy), .pid_goidle(pid_goidle), .pid_ccidle(
        prx_rcvinf[4]), .pcc_rxgood(pcc_rxgood), .prx_crcstart(prx_crcstart), 
        .prx_crcshfi4(prx_crcshfi4), .prx_crcsidat(prx_crcsidat), .prx_rxcode(
        dbgpo[28:24]), .prx_adpn(prx_adpn), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_eoprcvd(prx_eoprcvd), .prx_fsm(prx_fsm), .clk(clk), .srstz(srstz), 
        .test_si(n60), .test_so(n59), .test_se(test_se) );
  phyidd_a0 u0_phyidd ( .i_trans(x_trans), .i_goidle(ptx_goidle), .o_ccidle(
        prx_rcvinf[4]), .o_goidle(pid_goidle), .o_gobusy(pid_gobusy), .clk(clk), .srstz(n35), .test_si(pff_ptr[5]), .test_so(n60), .test_se(test_se) );
  phytx_a0 u0_phytx ( .r_txnumk(c0_txnumk), .r_txendk(c0_txendk), .r_txshrt(
        r_txshrt), .r_txauto(c0_txauto), .prx_cccnt(prx_cccnt), .ptx_txact(
        n106), .ptx_cc(ptx_cc), .ptx_goidle(ptx_goidle), .ptx_fifopop(
        dbgpo[30]), .ptx_pspyld(), .i_rdat(mux_rdat), .i_txreq(n10), .i_one(
        mux_one), .ptx_crcstart(ptx_crcstart), .ptx_crcshfi4(ptx_crcshfi4), 
        .ptx_crcshfo4(ptx_crcshfo4), .ptx_crcsidat(ptx_crcsidat), .ptx_fsm(
        ptx_fsm), .pcc_crc30(crc32_3_0), .clk(clk), .srstz(n35), .test_si(n59), 
        .test_se(test_se) );
  phycrc_a0 u0_phycrc ( .crc32_3_0(crc32_3_0), .rx_good(pcc_rxgood), 
        .i_shfidat(crcsidat), .i_start(crcstart), .i_shfi4(crcshfi4), 
        .i_shfo4(crcshfo4), .clk(clk), .test_si(d_cc[1]), .test_so(n61), 
        .test_se(test_se) );
  phyff_DEPTH_NUM34_DEPTH_NBT6 u0_phyff ( .r_psh(r_fifopsh), .r_pop(r_fifopop), 
        .prx_psh(fifopsh_pff), .ptx_pop(fifopop_pff), .r_last(r_last), 
        .r_unlock(r_unlock), .i_lockena(lockena), .r_fiforst(r_fiforst), 
        .i_ccidle(prx_rcvinf[4]), .r_wdat(r_wdat), .prx_wdat(prx_fifowdat), 
        .txreq(pff_txreq), .ffack(pff_ack), .rdat0(pff_rdat), .full(pff_full), 
        .empty(pff_empty), .one(pff_one), .half(), .obsd(obsd), .dat_7_1(
        pff_dat_7_1), .ptr(pff_ptr), .fifowdat(dbgpo[7:0]), .fifopsh(dbgpo[16]), .clk(clk), .srstz(fifosrstz), .test_si(n61), .test_se(test_se) );
  updprl_a0 u0_updprl ( .r_spec(r_spec), .r_dat_spec(r_dat_spec), 
        .r_auto_txgdcrc(r_auto_gdcrc[0]), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_auto_discard(r_auto_discard), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_dat_cpmsgid(r_wdat[2:0]), .r_rdat(
        r_rdat), .r_rdy(r_rdy), .pid_ccidle(prx_rcvinf[4]), .r_discard(
        r_discard), .ptx_ack(ptx_goidle), .ptx_txact(n6), .ptx_fifopop(
        fifopop_prl), .prx_fifopsh(fifopsh_prl), .prx_gdmsgrcvd(prx_gdmsgrcvd), 
        .prx_eoprcvd(prx_eoprcvd), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_fifowdat(prx_fifowdat), .pff_c0dat({pff_c0dat, pff_rxpart}), 
        .prl_rdat(prl_rdat), .prl_txauto({SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, prl_txauto[4], SYNOPSYS_UNCONNECTED_4, 
        prl_txauto[2:0]}), .prl_last(prl_last), .prl_txreq(prl_txreq), 
        .prl_c0set(prl_c0set), .prl_cany0(n107), .prl_cany0r(prl_cany0r), 
        .prl_cany0w(prl_cany0w), .prl_idle(prl_idle), .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_fsm(prl_fsm), .prl_cpmsgid(prl_cpmsgid), 
        .prl_cany0adr(prl_cany0adr), .clk(clk), .srstz(n35), .test_si(n58), 
        .test_so(test_so), .test_se(test_se) );
  dbnc_WIDTH3 u0_sqlch_db ( .o_dbc(d_sqlch), .o_chg(), .i_org(i_sqlch), .clk(
        clk), .rstz(n35), .test_si(ptx_cc), .test_so(n58), .test_se(test_se)
         );
  SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 clk_gate_cclow_cnt_reg ( 
        .CLK(clk), .EN(N34), .ENCLK(net10281), .TE(test_se) );
  SDFFSQX1 d_cc_reg_0_ ( .D(i_cc_49), .SIN(cclow_cnt[8]), .SMC(test_se), .C(
        clk), .XS(srstz), .Q(d_cc[0]) );
  SDFFSQX1 d_cc_reg_1_ ( .D(d_cc[0]), .SIN(d_cc[0]), .SMC(test_se), .C(clk), 
        .XS(srstz), .Q(d_cc[1]) );
  SDFFQX1 cclow_cnt_reg_1_ ( .D(N36), .SIN(cclow_cnt[0]), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[1]) );
  SDFFQX1 cclow_cnt_reg_3_ ( .D(N38), .SIN(cclow_cnt[2]), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[3]) );
  SDFFQX1 cclow_cnt_reg_8_ ( .D(n101), .SIN(cclow_cnt[7]), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[8]) );
  SDFFQX1 cclow_cnt_reg_4_ ( .D(N39), .SIN(cclow_cnt[3]), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[4]) );
  SDFFQX1 cclow_cnt_reg_5_ ( .D(N40), .SIN(cclow_cnt[4]), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[5]) );
  SDFFQX1 cclow_cnt_reg_6_ ( .D(N41), .SIN(cclow_cnt[5]), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[6]) );
  SDFFQX1 cclow_cnt_reg_2_ ( .D(N37), .SIN(cclow_cnt[1]), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[2]) );
  SDFFQX1 cclow_cnt_reg_7_ ( .D(N42), .SIN(cclow_cnt[6]), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[7]) );
  SDFFQX1 cclow_cnt_reg_0_ ( .D(N35), .SIN(test_si), .SMC(test_se), .C(
        net10281), .Q(cclow_cnt[0]) );
  INVX1 U3 ( .A(1'b1), .Y(dbgpo[31]) );
  AND2XL U5 ( .A(r_txnumk[2]), .B(prl_idle), .Y(c0_txnumk[2]) );
  AND2X1 U6 ( .A(n33), .B(n40), .Y(rx_pshords) );
  MUX2IX1 U7 ( .D0(n44), .D1(n93), .S(n38), .Y(pff_rxpart[7]) );
  INVX1 U8 ( .A(n106), .Y(n4) );
  INVX1 U9 ( .A(n4), .Y(ptx_oe) );
  INVX1 U10 ( .A(n4), .Y(n6) );
  INVX1 U11 ( .A(n107), .Y(n7) );
  INVX1 U12 ( .A(n7), .Y(prl_cany0) );
  BUFX3 U13 ( .A(prx_fsm[3]), .Y(dbgpo[23]) );
  BUFX3 U14 ( .A(prx_rcvinf[4]), .Y(dbgpo[19]) );
  BUFX3 U15 ( .A(prx_fsm[0]), .Y(dbgpo[20]) );
  BUFX3 U16 ( .A(prx_fsm[1]), .Y(dbgpo[21]) );
  BUFX3 U17 ( .A(prx_fsm[2]), .Y(dbgpo[22]) );
  BUFX3 U18 ( .A(pff_rdat[4]), .Y(dbgpo[12]) );
  BUFX3 U19 ( .A(pff_rdat[2]), .Y(dbgpo[10]) );
  BUFX3 U20 ( .A(pff_rdat[7]), .Y(dbgpo[15]) );
  BUFX3 U21 ( .A(pff_rdat[0]), .Y(dbgpo[8]) );
  BUFX3 U22 ( .A(pff_rdat[3]), .Y(dbgpo[11]) );
  BUFX3 U23 ( .A(pff_rdat[1]), .Y(dbgpo[9]) );
  BUFX3 U24 ( .A(pff_rdat[6]), .Y(dbgpo[14]) );
  BUFX3 U25 ( .A(pff_rdat[5]), .Y(dbgpo[13]) );
  INVX1 U26 ( .A(prl_idle), .Y(n34) );
  MUX2X2 U27 ( .D0(prl_last), .D1(pff_one), .S(n33), .Y(mux_one) );
  AND2X1 U28 ( .A(r_txnumk[1]), .B(prl_idle), .Y(c0_txnumk[1]) );
  MUX2XL U29 ( .D0(prl_txreq), .D1(pff_txreq), .S(n32), .Y(n10) );
  AND2XL U30 ( .A(dbgpo[29]), .B(n33), .Y(fifopsh_pff) );
  AND2XL U31 ( .A(r_txendk), .B(n33), .Y(c0_txendk) );
  MUX2XL U32 ( .D0(prl_rdat[1]), .D1(pff_rdat[1]), .S(n33), .Y(mux_rdat[1]) );
  MUX2XL U33 ( .D0(prl_rdat[5]), .D1(pff_rdat[5]), .S(n33), .Y(mux_rdat[5]) );
  AND2XL U34 ( .A(r_txauto[6]), .B(n33), .Y(c0_txauto[6]) );
  AO22XL U35 ( .A(ptx_crcsidat[3]), .B(n6), .C(prx_crcsidat[3]), .D(n4), .Y(
        crcsidat[3]) );
  MUX2XL U36 ( .D0(prl_txauto[0]), .D1(r_txauto[0]), .S(n32), .Y(c0_txauto[0])
         );
  MUX2XL U37 ( .D0(prl_txauto[2]), .D1(r_txauto[2]), .S(n32), .Y(c0_txauto[2])
         );
  MUX2XL U38 ( .D0(prl_txauto[1]), .D1(r_txauto[1]), .S(n32), .Y(c0_txauto[1])
         );
  MUX2XL U39 ( .D0(prl_txauto[4]), .D1(r_txauto[4]), .S(n32), .Y(c0_txauto[4])
         );
  NAND21XL U40 ( .B(r_txauto[3]), .A(n32), .Y(c0_txauto[3]) );
  NAND21XL U41 ( .B(r_txauto[5]), .A(n32), .Y(c0_txauto[5]) );
  INVX1 U42 ( .A(n34), .Y(n32) );
  INVX1 U43 ( .A(n34), .Y(n33) );
  AND2X1 U44 ( .A(dbgpo[30]), .B(n34), .Y(fifopop_prl) );
  NOR21XL U45 ( .B(ptx_crcshfo4), .A(n4), .Y(crcshfo4) );
  AND2X1 U46 ( .A(prx_setsta[3]), .B(n62), .Y(prx_gdmsgrcvd) );
  NOR2X1 U47 ( .A(prx_fiforst), .B(n36), .Y(fifosrstz) );
  AND2XL U48 ( .A(dbgpo[30]), .B(prl_idle), .Y(fifopop_pff) );
  MUX2X1 U49 ( .D0(pff_dat_7_1[18]), .D1(pff_dat_7_1[34]), .S(n39), .Y(
        pff_c0dat[26]) );
  MUX2X1 U50 ( .D0(pff_dat_7_1[17]), .D1(pff_dat_7_1[33]), .S(n39), .Y(
        pff_c0dat[25]) );
  MUX2X1 U51 ( .D0(pff_dat_7_1[15]), .D1(pff_dat_7_1[31]), .S(n39), .Y(
        pff_c0dat[23]) );
  INVX1 U52 ( .A(n36), .Y(n35) );
  AND2X2 U53 ( .A(dbgpo[29]), .B(n34), .Y(fifopsh_prl) );
  INVX1 U54 ( .A(n43), .Y(n40) );
  AO22X1 U55 ( .A(ptx_crcstart), .B(n6), .C(prx_crcstart), .D(n4), .Y(crcstart) );
  AO22X1 U56 ( .A(ptx_crcshfi4), .B(ptx_oe), .C(prx_crcshfi4), .D(n4), .Y(
        crcshfi4) );
  MUX2X1 U57 ( .D0(pff_dat_7_1[11]), .D1(pff_dat_7_1[27]), .S(n38), .Y(
        pff_c0dat[19]) );
  NAND42X1 U58 ( .C(pff_rxpart[14]), .D(pff_rxpart[13]), .A(n53), .B(n52), .Y(
        n62) );
  AND3X1 U59 ( .A(n51), .B(pff_rxpart[0]), .C(n50), .Y(n52) );
  NOR32XL U60 ( .B(n49), .C(n48), .A(n47), .Y(n53) );
  NAND21X1 U61 ( .B(pff_rxpart[4]), .A(n46), .Y(n47) );
  INVX1 U62 ( .A(n43), .Y(n38) );
  INVX1 U63 ( .A(pff_rxpart[12]), .Y(n46) );
  INVX1 U64 ( .A(pff_rxpart[2]), .Y(n48) );
  INVX1 U65 ( .A(pff_rxpart[3]), .Y(n49) );
  MUX2IX1 U66 ( .D0(n92), .D1(n87), .S(n39), .Y(pff_c0dat[24]) );
  MUX2IX1 U67 ( .D0(n95), .D1(n67), .S(n39), .Y(pff_c0dat[21]) );
  MUX2BXL U68 ( .D0(pff_dat_7_1[21]), .D1(n66), .S(n39), .Y(pff_c0dat[29]) );
  INVX1 U69 ( .A(n43), .Y(n39) );
  MUX2X1 U70 ( .D0(pff_dat_7_1[20]), .D1(pff_dat_7_1[36]), .S(n39), .Y(
        pff_c0dat[28]) );
  MUX2X1 U71 ( .D0(pff_dat_7_1[19]), .D1(pff_dat_7_1[35]), .S(n39), .Y(
        pff_c0dat[27]) );
  INVX1 U72 ( .A(n43), .Y(n41) );
  INVX1 U73 ( .A(n51), .Y(pff_rxpart[15]) );
  INVX1 U74 ( .A(n43), .Y(n42) );
  MUX2IX1 U75 ( .D0(n94), .D1(n65), .S(n39), .Y(pff_c0dat[22]) );
  MUX2BXL U76 ( .D0(pff_dat_7_1[12]), .D1(n83), .S(n39), .Y(pff_c0dat[20]) );
  INVX1 U77 ( .A(n50), .Y(pff_rxpart[1]) );
  INVX1 U78 ( .A(srstz), .Y(n36) );
  INVX1 U79 ( .A(n72), .Y(n103) );
  INVX1 U80 ( .A(n76), .Y(n105) );
  INVX1 U81 ( .A(n74), .Y(n104) );
  MUX2X1 U82 ( .D0(prl_rdat[7]), .D1(pff_rdat[7]), .S(n32), .Y(mux_rdat[7]) );
  MUX2X1 U83 ( .D0(prl_rdat[4]), .D1(pff_rdat[4]), .S(n33), .Y(mux_rdat[4]) );
  MUX2X1 U84 ( .D0(prl_rdat[6]), .D1(pff_rdat[6]), .S(n32), .Y(mux_rdat[6]) );
  AND2X1 U85 ( .A(r_txnumk[0]), .B(prl_idle), .Y(c0_txnumk[0]) );
  AND2XL U86 ( .A(r_txnumk[3]), .B(prl_idle), .Y(c0_txnumk[3]) );
  MUX2X1 U87 ( .D0(prl_rdat[0]), .D1(pff_rdat[0]), .S(n33), .Y(mux_rdat[0]) );
  MUX2X1 U88 ( .D0(prl_rdat[3]), .D1(pff_rdat[3]), .S(n33), .Y(mux_rdat[3]) );
  MUX2X1 U89 ( .D0(prl_rdat[2]), .D1(pff_rdat[2]), .S(n32), .Y(mux_rdat[2]) );
  AND2XL U90 ( .A(r_txnumk[4]), .B(prl_idle), .Y(c0_txnumk[4]) );
  INVX1 U91 ( .A(r_pshords), .Y(n43) );
  BUFX3 U92 ( .A(prx_rcvinf[3]), .Y(dbgpo[17]) );
  AOI21AXL U93 ( .B(n6), .C(prl_idle), .A(r_first), .Y(lockena) );
  INVX1 U94 ( .A(n45), .Y(pff_rxpart[8]) );
  MUX2AXL U95 ( .D0(pff_dat_7_1[0]), .D1(n92), .S(n37), .Y(n45) );
  MUX2BXL U96 ( .D0(pff_rdat[6]), .D1(n94), .S(n37), .Y(pff_rxpart[6]) );
  MUX2BXL U97 ( .D0(pff_rdat[5]), .D1(n95), .S(n38), .Y(pff_rxpart[5]) );
  NOR21XL U98 ( .B(obsd), .A(prx_setsta[6]), .Y(pff_obsd) );
  MUX2X1 U99 ( .D0(pff_rdat[2]), .D1(pff_dat_7_1[10]), .S(n37), .Y(
        pff_rxpart[2]) );
  MUX2X1 U100 ( .D0(pff_rdat[3]), .D1(pff_dat_7_1[11]), .S(n38), .Y(
        pff_rxpart[3]) );
  MUX2X1 U101 ( .D0(pff_dat_7_1[4]), .D1(pff_dat_7_1[20]), .S(n38), .Y(
        pff_rxpart[12]) );
  MUX2IX1 U102 ( .D0(pff_rdat[1]), .D1(pff_dat_7_1[9]), .S(n37), .Y(n50) );
  MUX2IX1 U103 ( .D0(pff_dat_7_1[7]), .D1(pff_dat_7_1[23]), .S(n37), .Y(n51)
         );
  MUX2X1 U104 ( .D0(pff_dat_7_1[5]), .D1(pff_dat_7_1[21]), .S(n38), .Y(
        pff_rxpart[13]) );
  MUX2X1 U105 ( .D0(pff_dat_7_1[6]), .D1(pff_dat_7_1[22]), .S(n38), .Y(
        pff_rxpart[14]) );
  MUX2X1 U106 ( .D0(pff_rdat[4]), .D1(pff_dat_7_1[12]), .S(n37), .Y(
        pff_rxpart[4]) );
  INVX1 U107 ( .A(n43), .Y(n37) );
  MUX2X1 U108 ( .D0(pff_rdat[0]), .D1(pff_dat_7_1[8]), .S(n37), .Y(
        pff_rxpart[0]) );
  NOR21XL U109 ( .B(r_auto_gdcrc[1]), .A(n62), .Y(auto_rx_gdcrc) );
  ENOX1 U110 ( .A(n41), .B(n63), .C(pff_dat_7_1[55]), .D(n42), .Y(
        pff_c0dat[47]) );
  ENOX1 U111 ( .A(n41), .B(n66), .C(pff_dat_7_1[53]), .D(n42), .Y(
        pff_c0dat[45]) );
  MUX2BXL U112 ( .D0(pff_dat_7_1[9]), .D1(n100), .S(n38), .Y(pff_c0dat[17]) );
  MUX2BXL U113 ( .D0(pff_dat_7_1[23]), .D1(n63), .S(n40), .Y(pff_c0dat[31]) );
  ENOX1 U114 ( .A(n41), .B(n86), .C(pff_dat_7_1[49]), .D(n42), .Y(
        pff_c0dat[41]) );
  ENOX1 U115 ( .A(n41), .B(n64), .C(pff_dat_7_1[47]), .D(n42), .Y(
        pff_c0dat[39]) );
  ENOX1 U116 ( .A(n40), .B(n65), .C(pff_dat_7_1[46]), .D(n42), .Y(
        pff_c0dat[38]) );
  ENOX1 U117 ( .A(n40), .B(n100), .C(pff_dat_7_1[41]), .D(r_pshords), .Y(
        pff_c0dat[33]) );
  MUX2X1 U118 ( .D0(pff_dat_7_1[22]), .D1(pff_dat_7_1[38]), .S(n40), .Y(
        pff_c0dat[30]) );
  MUX2X1 U119 ( .D0(pff_dat_7_1[8]), .D1(pff_dat_7_1[24]), .S(n38), .Y(
        pff_c0dat[16]) );
  MUX2X1 U120 ( .D0(pff_dat_7_1[10]), .D1(pff_dat_7_1[26]), .S(n38), .Y(
        pff_c0dat[18]) );
  ENOX1 U121 ( .A(n41), .B(n98), .C(pff_dat_7_1[51]), .D(n42), .Y(
        pff_c0dat[43]) );
  ENOX1 U122 ( .A(n41), .B(n99), .C(pff_dat_7_1[50]), .D(n42), .Y(
        pff_c0dat[42]) );
  ENOX1 U123 ( .A(n41), .B(n97), .C(pff_dat_7_1[52]), .D(n42), .Y(
        pff_c0dat[44]) );
  ENOX1 U124 ( .A(n40), .B(n88), .C(pff_dat_7_1[40]), .D(n41), .Y(
        pff_c0dat[32]) );
  ENOX1 U125 ( .A(n40), .B(n67), .C(pff_dat_7_1[45]), .D(r_pshords), .Y(
        pff_c0dat[37]) );
  ENOX1 U126 ( .A(n40), .B(n84), .C(pff_dat_7_1[43]), .D(r_pshords), .Y(
        pff_c0dat[35]) );
  ENOX1 U127 ( .A(n40), .B(n83), .C(pff_dat_7_1[44]), .D(r_pshords), .Y(
        pff_c0dat[36]) );
  INVX1 U128 ( .A(pff_dat_7_1[26]), .Y(n85) );
  INVX1 U129 ( .A(pff_dat_7_1[24]), .Y(n88) );
  INVX1 U130 ( .A(pff_dat_7_1[29]), .Y(n67) );
  INVX1 U131 ( .A(pff_dat_7_1[32]), .Y(n87) );
  INVX1 U132 ( .A(pff_dat_7_1[38]), .Y(n96) );
  INVX1 U133 ( .A(pff_dat_7_1[35]), .Y(n98) );
  INVX1 U134 ( .A(pff_dat_7_1[36]), .Y(n97) );
  INVX1 U135 ( .A(pff_dat_7_1[34]), .Y(n99) );
  INVX1 U136 ( .A(pff_dat_7_1[25]), .Y(n100) );
  INVX1 U137 ( .A(pff_dat_7_1[27]), .Y(n84) );
  INVX1 U138 ( .A(pff_dat_7_1[37]), .Y(n66) );
  INVX1 U139 ( .A(pff_dat_7_1[39]), .Y(n63) );
  INVX1 U140 ( .A(pff_dat_7_1[31]), .Y(n64) );
  INVX1 U141 ( .A(pff_dat_7_1[33]), .Y(n86) );
  INVX1 U142 ( .A(pff_dat_7_1[30]), .Y(n65) );
  INVX1 U143 ( .A(pff_dat_7_1[28]), .Y(n83) );
  INVX1 U144 ( .A(pff_dat_7_1[16]), .Y(n92) );
  INVX1 U145 ( .A(pff_dat_7_1[19]), .Y(n89) );
  INVX1 U146 ( .A(pff_dat_7_1[17]), .Y(n91) );
  INVX1 U147 ( .A(pff_dat_7_1[18]), .Y(n90) );
  ENOX1 U148 ( .A(n40), .B(n85), .C(pff_dat_7_1[42]), .D(n42), .Y(
        pff_c0dat[34]) );
  INVX1 U149 ( .A(pff_dat_7_1[14]), .Y(n94) );
  INVX1 U150 ( .A(pff_dat_7_1[15]), .Y(n93) );
  INVX1 U151 ( .A(pff_dat_7_1[13]), .Y(n95) );
  ENOX1 U152 ( .A(n41), .B(n96), .C(pff_dat_7_1[54]), .D(n42), .Y(
        pff_c0dat[46]) );
  ENOX1 U153 ( .A(n41), .B(n87), .C(pff_dat_7_1[48]), .D(r_pshords), .Y(
        pff_c0dat[40]) );
  NOR21XL U154 ( .B(ptx_goidle), .A(prl_cany0), .Y(ptx_ack) );
  AOI31X1 U155 ( .A(d_sqlch), .B(n55), .C(r_sqlch[0]), .D(n54), .Y(x_trans) );
  OAI21X1 U156 ( .B(n6), .C(prx_fsm[3]), .A(r_sqlch[1]), .Y(n55) );
  INVX1 U157 ( .A(prx_trans), .Y(n54) );
  NOR4XL U158 ( .A(n56), .B(n57), .C(cclow_cnt[5]), .D(cclow_cnt[4]), .Y(
        prx_setsta[0]) );
  OR3XL U159 ( .A(cclow_cnt[7]), .B(cclow_cnt[6]), .C(cclow_cnt[8]), .Y(n57)
         );
  NAND43X1 U160 ( .B(cclow_cnt[3]), .C(cclow_cnt[1]), .D(cclow_cnt[2]), .A(
        cclow_cnt[0]), .Y(n56) );
  OAI211X1 U161 ( .C(cclow_cnt[8]), .D(n69), .A(n35), .B(n82), .Y(n72) );
  XNOR2XL U162 ( .A(d_cc[1]), .B(d_cc[0]), .Y(n82) );
  GEN2XL U163 ( .D(cclow_cnt[1]), .E(cclow_cnt[0]), .C(n80), .B(n103), .A(n70), 
        .Y(N36) );
  GEN2XL U164 ( .D(cclow_cnt[4]), .E(n75), .C(n76), .B(n103), .A(n70), .Y(N39)
         );
  GEN2XL U165 ( .D(cclow_cnt[6]), .E(n104), .C(n73), .B(n103), .A(n70), .Y(N41) );
  GEN2XL U166 ( .D(cclow_cnt[5]), .E(n105), .C(n74), .B(n103), .A(n70), .Y(N40) );
  NAND21X1 U167 ( .B(cclow_cnt[2]), .A(n80), .Y(n78) );
  NAND21X1 U168 ( .B(cclow_cnt[7]), .A(n73), .Y(n69) );
  NOR2X1 U169 ( .A(n75), .B(cclow_cnt[4]), .Y(n76) );
  NOR2X1 U170 ( .A(n105), .B(cclow_cnt[5]), .Y(n74) );
  NOR2X1 U171 ( .A(n104), .B(cclow_cnt[6]), .Y(n73) );
  NOR2X1 U172 ( .A(cclow_cnt[1]), .B(cclow_cnt[0]), .Y(n80) );
  AOI21X1 U173 ( .B(n69), .C(n71), .A(n72), .Y(N42) );
  NAND21X1 U174 ( .B(n73), .A(cclow_cnt[7]), .Y(n71) );
  AOI21X1 U175 ( .B(n78), .C(n79), .A(n72), .Y(N37) );
  NAND21X1 U176 ( .B(n80), .A(cclow_cnt[2]), .Y(n79) );
  AOI21X1 U178 ( .B(n75), .C(n77), .A(n72), .Y(N38) );
  NAND2X1 U179 ( .A(cclow_cnt[3]), .B(n78), .Y(n77) );
  OR2X1 U180 ( .A(n78), .B(cclow_cnt[3]), .Y(n75) );
  NOR2X1 U181 ( .A(cclow_cnt[0]), .B(n72), .Y(N35) );
  INVX1 U182 ( .A(n68), .Y(n101) );
  AOI31X1 U183 ( .A(n103), .B(n69), .C(cclow_cnt[8]), .D(n70), .Y(n68) );
  MUX2BXL U184 ( .D0(pff_dat_7_1[2]), .D1(n90), .S(n37), .Y(pff_rxpart[10]) );
  MUX2BXL U185 ( .D0(pff_dat_7_1[1]), .D1(n91), .S(n37), .Y(pff_rxpart[9]) );
  NAND31X1 U186 ( .C(n70), .A(n72), .B(n81), .Y(N34) );
  AOI21X1 U187 ( .B(d_cc[0]), .C(n102), .A(n36), .Y(n81) );
  NOR3XL U188 ( .A(n36), .B(d_cc[0]), .C(n102), .Y(n70) );
  MUX2BXL U189 ( .D0(pff_dat_7_1[3]), .D1(n89), .S(n37), .Y(pff_rxpart[11]) );
  INVX1 U190 ( .A(d_cc[1]), .Y(n102) );
  INVX1 U191 ( .A(pff_rdat[7]), .Y(n44) );
  AO22XL U192 ( .A(ptx_crcsidat[0]), .B(n6), .C(prx_crcsidat[0]), .D(n4), .Y(
        crcsidat[0]) );
  AO22XL U193 ( .A(ptx_crcsidat[2]), .B(n6), .C(prx_crcsidat[2]), .D(n4), .Y(
        crcsidat[2]) );
  AO22XL U194 ( .A(ptx_crcsidat[1]), .B(n6), .C(prx_crcsidat[1]), .D(n4), .Y(
        crcsidat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_1_, db_cnt_0_, N14, N15, N16, N17, net10299, n8, n1,
         n2, n3, n4, n5;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N14), 
        .ENCLK(net10299), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N17), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net10299), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N16), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net10299), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N15), .SIN(o_dbc), .SMC(test_se), .C(net10299), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n8), .SIN(d_org_0_), .SMC(test_se), .C(net10299), 
        .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n2), .A(n1), .Y(n4) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U5 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n8) );
  NOR2X1 U6 ( .A(n1), .B(n2), .Y(o_chg) );
  NAND3X1 U7 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(test_so), .Y(n1) );
  NOR2X1 U8 ( .A(n5), .B(n4), .Y(N16) );
  XNOR2XL U9 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n5) );
  NOR2X1 U10 ( .A(db_cnt_0_), .B(n4), .Y(N15) );
  NOR2X1 U11 ( .A(n3), .B(n4), .Y(N17) );
  AOI21X1 U12 ( .B(db_cnt_1_), .C(db_cnt_0_), .A(test_so), .Y(n3) );
  NAND43X1 U13 ( .B(test_so), .C(db_cnt_0_), .D(db_cnt_1_), .A(n2), .Y(N14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updprl_a0 ( r_spec, r_dat_spec, r_auto_txgdcrc, r_dat_portrole, 
        r_dat_datarole, r_auto_discard, r_set_cpmsgid, r_dat_cpmsgid, r_rdat, 
        r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact, ptx_fifopop, 
        prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, prx_rcvdords, prx_fifowdat, 
        pff_c0dat, prl_rdat, prl_txauto, prl_last, prl_txreq, prl_c0set, 
        prl_cany0, prl_cany0r, prl_cany0w, prl_idle, prl_discard, prl_GCTxDone, 
        prl_fsm, prl_cpmsgid, prl_cany0adr, clk, srstz, test_si, test_so, 
        test_se );
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [2:0] r_dat_cpmsgid;
  input [7:0] r_rdat;
  input [2:0] prx_rcvdords;
  input [7:0] prx_fifowdat;
  input [47:0] pff_c0dat;
  output [7:0] prl_rdat;
  output [6:0] prl_txauto;
  output [3:0] prl_fsm;
  output [2:0] prl_cpmsgid;
  output [7:0] prl_cany0adr;
  input r_auto_txgdcrc, r_dat_portrole, r_dat_datarole, r_auto_discard,
         r_set_cpmsgid, r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact,
         ptx_fifopop, prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, clk, srstz,
         test_si, test_se;
  output prl_last, prl_txreq, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_idle, prl_discard, prl_GCTxDone, test_so;
  wire   sendgdcrc, stoptimer, N41, c0_iop, N113, N114, N115, N116, N117, N118,
         N119, N120, N151, N152, N153, N154, N155, N156, N157, N158, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N189, N190, N191,
         N192, N193, N194, N196, N203, N204, N205, N206, net10322, net10328,
         net10333, net10338, net10343, n99, n100, n37, n39, n51, n56, n57, n58,
         n59, n67, n68, n72, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n98, n101, n7, n8, n9, n10, n11, n13,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n38, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n52, n53, n54, n55, n60, n61, n62, n63, n64, n65,
         n66, n69, n70, n71, n73, n74, n75, n76, n77, n78, n79, n80, n97, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156;
  wire   [1:0] PrlTo;
  wire   [8:0] c0_cnt;
  wire   [7:0] txbuf;

  PrlTimer_1112a0 u0_PrlTimer ( .to(PrlTo), .restart(sendgdcrc), .stop(
        stoptimer), .clk(clk), .srstz(n17), .test_si(txbuf[7]), .test_so(
        test_so), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_0 clk_gate_txbuf_reg ( .CLK(clk), .EN(N41), 
        .ENCLK(net10322), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_4 clk_gate_c0_adr_reg ( .CLK(clk), .EN(N194), 
        .ENCLK(net10328), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_3 clk_gate_cs_prcl_reg ( .CLK(clk), .EN(N189), 
        .ENCLK(net10333), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_2 clk_gate_c0_cnt_reg ( .CLK(clk), .EN(N196), 
        .ENCLK(net10338), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_1 clk_gate_CpMsgId_reg ( .CLK(clk), .EN(N203), 
        .ENCLK(net10343), .TE(test_se) );
  updprl_a0_DW01_inc_0 r328 ( .A(prl_cany0adr), .SUM({N120, N119, N118, N117, 
        N116, N115, N114, N113}) );
  SDFFQX1 c0_iop_reg ( .D(n99), .SIN(c0_cnt[8]), .SMC(test_se), .C(net10333), 
        .Q(c0_iop) );
  SDFFQX1 canyon_m0_reg ( .D(n100), .SIN(c0_iop), .SMC(test_se), .C(clk), .Q(
        prl_cany0) );
  SDFFQX1 c0_adr_reg_2_ ( .D(N153), .SIN(prl_cany0adr[1]), .SMC(test_se), .C(
        net10328), .Q(prl_cany0adr[2]) );
  SDFFQX1 c0_adr_reg_1_ ( .D(N152), .SIN(prl_cany0adr[0]), .SMC(test_se), .C(
        net10328), .Q(prl_cany0adr[1]) );
  SDFFQX1 c0_adr_reg_3_ ( .D(N154), .SIN(prl_cany0adr[2]), .SMC(test_se), .C(
        net10328), .Q(prl_cany0adr[3]) );
  SDFFQX1 c0_adr_reg_4_ ( .D(N155), .SIN(prl_cany0adr[3]), .SMC(test_se), .C(
        net10328), .Q(prl_cany0adr[4]) );
  SDFFQX1 c0_adr_reg_5_ ( .D(N156), .SIN(prl_cany0adr[4]), .SMC(test_se), .C(
        net10328), .Q(prl_cany0adr[5]) );
  SDFFQX1 c0_adr_reg_6_ ( .D(N157), .SIN(prl_cany0adr[5]), .SMC(test_se), .C(
        net10328), .Q(prl_cany0adr[6]) );
  SDFFQX1 c0_adr_reg_0_ ( .D(N151), .SIN(prl_cpmsgid[2]), .SMC(test_se), .C(
        net10328), .Q(prl_cany0adr[0]) );
  SDFFQX1 c0_adr_reg_7_ ( .D(N158), .SIN(prl_cany0adr[6]), .SMC(test_se), .C(
        net10328), .Q(prl_cany0adr[7]) );
  SDFFQX1 txbuf_reg_4_ ( .D(r_rdat[4]), .SIN(txbuf[3]), .SMC(test_se), .C(
        net10322), .Q(txbuf[4]) );
  SDFFQX1 txbuf_reg_1_ ( .D(r_rdat[1]), .SIN(txbuf[0]), .SMC(test_se), .C(
        net10322), .Q(txbuf[1]) );
  SDFFQX1 txbuf_reg_7_ ( .D(r_rdat[7]), .SIN(txbuf[6]), .SMC(test_se), .C(
        net10322), .Q(txbuf[7]) );
  SDFFQX1 CpMsgId_reg_0_ ( .D(N204), .SIN(test_si), .SMC(test_se), .C(net10343), .Q(prl_cpmsgid[0]) );
  SDFFQX1 CpMsgId_reg_2_ ( .D(N206), .SIN(prl_cpmsgid[1]), .SMC(test_se), .C(
        net10343), .Q(prl_cpmsgid[2]) );
  SDFFQX1 c0_cnt_reg_5_ ( .D(N170), .SIN(c0_cnt[4]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[5]) );
  SDFFQX1 c0_cnt_reg_7_ ( .D(N172), .SIN(c0_cnt[6]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[7]) );
  SDFFQX1 c0_cnt_reg_6_ ( .D(N171), .SIN(c0_cnt[5]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[6]) );
  SDFFQX1 c0_cnt_reg_4_ ( .D(N169), .SIN(c0_cnt[3]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[4]) );
  SDFFQX1 c0_cnt_reg_3_ ( .D(N168), .SIN(c0_cnt[2]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[3]) );
  SDFFQX1 c0_cnt_reg_2_ ( .D(N167), .SIN(c0_cnt[1]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[2]) );
  SDFFQX1 c0_cnt_reg_1_ ( .D(N166), .SIN(c0_cnt[0]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[1]) );
  SDFFQX1 cs_prcl_reg_2_ ( .D(N192), .SIN(prl_fsm[1]), .SMC(test_se), .C(
        net10333), .Q(prl_fsm[2]) );
  SDFFQXL txbuf_reg_5_ ( .D(r_rdat[5]), .SIN(txbuf[4]), .SMC(test_se), .C(
        net10322), .Q(txbuf[5]) );
  SDFFQXL txbuf_reg_2_ ( .D(r_rdat[2]), .SIN(txbuf[1]), .SMC(test_se), .C(
        net10322), .Q(txbuf[2]) );
  SDFFQXL txbuf_reg_6_ ( .D(r_rdat[6]), .SIN(txbuf[5]), .SMC(test_se), .C(
        net10322), .Q(txbuf[6]) );
  SDFFQXL txbuf_reg_3_ ( .D(r_rdat[3]), .SIN(txbuf[2]), .SMC(test_se), .C(
        net10322), .Q(txbuf[3]) );
  SDFFQXL c0_cnt_reg_8_ ( .D(N173), .SIN(c0_cnt[7]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[8]) );
  SDFFQXL CpMsgId_reg_1_ ( .D(N205), .SIN(prl_cpmsgid[0]), .SMC(test_se), .C(
        net10343), .Q(prl_cpmsgid[1]) );
  SDFFQX1 txbuf_reg_0_ ( .D(r_rdat[0]), .SIN(prl_fsm[3]), .SMC(test_se), .C(
        net10322), .Q(txbuf[0]) );
  SDFFQX1 cs_prcl_reg_1_ ( .D(N191), .SIN(prl_fsm[0]), .SMC(test_se), .C(
        net10333), .Q(prl_fsm[1]) );
  SDFFQX1 cs_prcl_reg_0_ ( .D(N190), .SIN(prl_cany0), .SMC(test_se), .C(
        net10333), .Q(prl_fsm[0]) );
  SDFFQX1 cs_prcl_reg_3_ ( .D(N193), .SIN(prl_fsm[2]), .SMC(test_se), .C(
        net10333), .Q(prl_fsm[3]) );
  SDFFQX1 c0_cnt_reg_0_ ( .D(N165), .SIN(prl_cany0adr[7]), .SMC(test_se), .C(
        net10338), .Q(c0_cnt[0]) );
  INVX1 U3 ( .A(1'b0), .Y(prl_txauto[3]) );
  INVX1 U5 ( .A(1'b0), .Y(prl_txauto[5]) );
  INVX1 U7 ( .A(1'b1), .Y(prl_txauto[6]) );
  INVX3 U9 ( .A(prx_fifopsh), .Y(n30) );
  INVX1 U10 ( .A(prl_fsm[1]), .Y(n23) );
  NAND21X1 U11 ( .B(n77), .A(n75), .Y(n65) );
  AND2X1 U12 ( .A(n10), .B(n114), .Y(n9) );
  INVX1 U13 ( .A(n119), .Y(n124) );
  INVX1 U14 ( .A(n122), .Y(n118) );
  INVX1 U15 ( .A(n131), .Y(n121) );
  INVX1 U16 ( .A(n127), .Y(n130) );
  INVX1 U17 ( .A(n115), .Y(n111) );
  INVX1 U18 ( .A(n112), .Y(n126) );
  NAND3X1 U19 ( .A(prx_fifopsh), .B(n8), .C(n141), .Y(n7) );
  AND3X4 U20 ( .A(prx_fifopsh), .B(n8), .C(n141), .Y(prl_cany0w) );
  INVX1 U21 ( .A(n109), .Y(n8) );
  INVX1 U22 ( .A(prl_fsm[2]), .Y(n25) );
  INVX1 U23 ( .A(prl_fsm[3]), .Y(n19) );
  INVX1 U24 ( .A(c0_cnt[8]), .Y(n10) );
  NAND32X1 U25 ( .B(prl_fsm[2]), .C(n24), .A(n23), .Y(n103) );
  OAI211XL U26 ( .C(n18), .D(n75), .A(n105), .B(n79), .Y(N192) );
  INVXL U27 ( .A(n75), .Y(n40) );
  NAND21X1 U28 ( .B(prl_txauto[4]), .A(ptx_fifopop), .Y(n31) );
  INVXL U29 ( .A(prl_txauto[4]), .Y(n41) );
  INVXL U30 ( .A(n109), .Y(n133) );
  OR2XL U31 ( .A(n140), .B(n22), .Y(n132) );
  AOI31XL U32 ( .A(n67), .B(n146), .C(n78), .D(n77), .Y(n97) );
  AO21XL U33 ( .B(n103), .C(n102), .A(n18), .Y(n104) );
  AOI22XL U34 ( .A(n98), .B(n133), .C(n41), .D(ptx_ack), .Y(n20) );
  NAND32XL U35 ( .B(n25), .C(n24), .A(n23), .Y(n73) );
  OR2XL U36 ( .A(n140), .B(n24), .Y(n71) );
  NAND32XL U37 ( .B(n25), .C(n22), .A(n23), .Y(n33) );
  OAI22AXL U38 ( .D(txbuf[6]), .C(n65), .A(n61), .B(n102), .Y(prl_rdat[6]) );
  INVXL U39 ( .A(n65), .Y(n49) );
  OAI22XL U40 ( .A(n65), .B(n46), .C(n75), .D(n45), .Y(prl_rdat[2]) );
  INVXL U41 ( .A(txbuf[2]), .Y(n46) );
  OAI22XL U42 ( .A(n65), .B(n48), .C(n75), .D(n47), .Y(prl_rdat[3]) );
  INVXL U43 ( .A(txbuf[3]), .Y(n48) );
  OAI221XL U44 ( .A(n65), .B(n42), .C(r_dat_portrole), .D(n75), .E(n102), .Y(
        prl_rdat[0]) );
  INVXL U45 ( .A(txbuf[0]), .Y(n42) );
  OAI22XL U46 ( .A(n65), .B(n44), .C(n75), .D(n43), .Y(prl_rdat[1]) );
  INVXL U47 ( .A(txbuf[1]), .Y(n44) );
  NAND42XL U48 ( .C(n102), .D(r_dat_datarole), .A(n52), .B(n50), .Y(n53) );
  INVXL U49 ( .A(r_spec[0]), .Y(n60) );
  INVXL U50 ( .A(prl_cpmsgid[2]), .Y(n47) );
  INVXL U51 ( .A(prl_cpmsgid[1]), .Y(n45) );
  NAND21XL U52 ( .B(n23), .A(prl_fsm[2]), .Y(n140) );
  BUFXL U53 ( .A(prx_rcvdords[0]), .Y(prl_txauto[0]) );
  BUFXL U54 ( .A(prx_rcvdords[2]), .Y(prl_txauto[2]) );
  BUFXL U55 ( .A(prx_rcvdords[1]), .Y(prl_txauto[1]) );
  NAND32XL U56 ( .B(prl_fsm[2]), .C(n22), .A(n23), .Y(n76) );
  AOI21XL U57 ( .B(c0_cnt[8]), .C(n116), .A(n9), .Y(n13) );
  OAI22XL U58 ( .A(n155), .B(n132), .C(c0_cnt[0]), .D(n109), .Y(N165) );
  INVX1 U59 ( .A(r_discard), .Y(n69) );
  INVX1 U60 ( .A(n18), .Y(n17) );
  NOR21XL U61 ( .B(prx_gdmsgrcvd), .A(r_set_cpmsgid), .Y(n57) );
  NAND32X1 U62 ( .B(r_set_cpmsgid), .C(prx_gdmsgrcvd), .A(n17), .Y(N203) );
  INVX1 U63 ( .A(srstz), .Y(n18) );
  INVX1 U64 ( .A(n102), .Y(n77) );
  INVX1 U65 ( .A(n51), .Y(prl_c0set) );
  NAND21X1 U66 ( .B(n106), .A(n138), .Y(n79) );
  INVX1 U67 ( .A(n106), .Y(n142) );
  INVX1 U68 ( .A(n72), .Y(n147) );
  INVX1 U69 ( .A(n149), .Y(n136) );
  OR3XL U70 ( .A(pff_c0dat[26]), .B(pff_c0dat[25]), .C(pff_c0dat[23]), .Y(n89)
         );
  NOR2X1 U71 ( .A(n152), .B(n73), .Y(n11) );
  INVX1 U72 ( .A(prx_fifowdat[3]), .Y(n156) );
  INVX1 U73 ( .A(n71), .Y(n107) );
  NAND21X1 U74 ( .B(n133), .A(n132), .Y(n139) );
  INVX1 U75 ( .A(n132), .Y(n128) );
  INVX1 U76 ( .A(n33), .Y(n138) );
  NAND32X1 U77 ( .B(n23), .C(n22), .A(n25), .Y(n75) );
  NAND32X1 U78 ( .B(n23), .C(n24), .A(n25), .Y(n102) );
  AO21X1 U79 ( .B(n9), .C(n41), .A(n40), .Y(prl_last) );
  INVX1 U80 ( .A(n103), .Y(prl_idle) );
  INVX1 U81 ( .A(n116), .Y(n114) );
  OAI22X1 U82 ( .A(n39), .B(n76), .C(ptx_txact), .D(prl_txauto[4]), .Y(
        prl_txreq) );
  OAI211X1 U83 ( .C(n18), .D(n97), .A(n80), .B(n79), .Y(N191) );
  INVX1 U84 ( .A(n76), .Y(n78) );
  NOR2X1 U85 ( .A(r_discard), .B(n68), .Y(n67) );
  NAND5XL U86 ( .A(n142), .B(n70), .C(n29), .D(n28), .E(n27), .Y(N189) );
  AOI211XL U87 ( .C(ptx_fifopop), .D(n65), .A(n26), .B(n11), .Y(n27) );
  AO21X1 U88 ( .B(n39), .C(n69), .A(n76), .Y(n29) );
  NAND2X1 U89 ( .A(n58), .B(n17), .Y(N205) );
  AOI22X1 U90 ( .A(pff_c0dat[10]), .B(n57), .C(r_dat_cpmsgid[1]), .D(
        r_set_cpmsgid), .Y(n58) );
  NAND2X1 U91 ( .A(n56), .B(n17), .Y(N206) );
  AOI22X1 U92 ( .A(pff_c0dat[11]), .B(n57), .C(r_set_cpmsgid), .D(
        r_dat_cpmsgid[2]), .Y(n56) );
  NAND2X1 U93 ( .A(n59), .B(n17), .Y(N204) );
  AOI22X1 U94 ( .A(pff_c0dat[9]), .B(n57), .C(r_dat_cpmsgid[0]), .D(
        r_set_cpmsgid), .Y(n59) );
  NAND4X1 U95 ( .A(n81), .B(n82), .C(n83), .D(n84), .Y(n51) );
  NOR4XL U96 ( .A(n88), .B(n89), .C(pff_c0dat[22]), .D(pff_c0dat[20]), .Y(n83)
         );
  NOR4XL U97 ( .A(n85), .B(n86), .C(pff_c0dat[36]), .D(pff_c0dat[34]), .Y(n84)
         );
  NOR42XL U98 ( .C(pff_c0dat[46]), .D(pff_c0dat[40]), .A(n94), .B(n95), .Y(n81) );
  NOR42XL U99 ( .C(pff_c0dat[1]), .D(pff_c0dat[19]), .A(n91), .B(n92), .Y(n82)
         );
  NAND3X1 U100 ( .A(pff_c0dat[12]), .B(pff_c0dat[0]), .C(pff_c0dat[17]), .Y(
        n92) );
  NAND42X1 U101 ( .C(pff_c0dat[14]), .D(pff_c0dat[13]), .A(prx_gdmsgrcvd), .B(
        n93), .Y(n91) );
  OAI21BBXL U102 ( .A(sendgdcrc), .B(prl_idle), .C(n32), .Y(n26) );
  NAND32X1 U103 ( .B(n21), .C(n18), .A(n20), .Y(n106) );
  INVX1 U104 ( .A(n74), .Y(n105) );
  OAI31XL U105 ( .A(n18), .B(n151), .C(n73), .D(n80), .Y(n74) );
  NAND42X1 U106 ( .C(n71), .D(n106), .A(n147), .B(n155), .Y(n80) );
  AOI21AX1 U107 ( .B(n151), .C(n51), .A(n142), .Y(n100) );
  OAI211X1 U108 ( .C(n106), .D(n132), .A(n105), .B(n104), .Y(N190) );
  NAND4X1 U109 ( .A(n156), .B(n149), .C(n154), .D(n101), .Y(n72) );
  NAND32X1 U110 ( .B(pff_c0dat[28]), .C(pff_c0dat[27]), .A(n90), .Y(n88) );
  NOR3XL U111 ( .A(pff_c0dat[29]), .B(pff_c0dat[32]), .C(pff_c0dat[31]), .Y(
        n90) );
  INVX1 U112 ( .A(n148), .Y(n135) );
  INVX1 U113 ( .A(n150), .Y(n134) );
  AO22X1 U114 ( .A(N119), .B(n139), .C(n138), .D(n134), .Y(N157) );
  AO22X1 U115 ( .A(N118), .B(n139), .C(n138), .D(n135), .Y(N156) );
  AO22X1 U116 ( .A(N117), .B(n139), .C(n138), .D(n136), .Y(N155) );
  INVX1 U117 ( .A(ptx_ack), .Y(n152) );
  NAND21X1 U118 ( .B(n76), .A(n68), .Y(n70) );
  INVX1 U119 ( .A(n39), .Y(n146) );
  AO22X1 U120 ( .A(N114), .B(n139), .C(n138), .D(n145), .Y(N152) );
  AO22X1 U121 ( .A(N115), .B(n139), .C(n138), .D(n137), .Y(N153) );
  AO22X1 U122 ( .A(N116), .B(n139), .C(n138), .D(prx_fifowdat[3]), .Y(N154) );
  INVX1 U123 ( .A(n154), .Y(n137) );
  OAI22X1 U124 ( .A(n66), .B(n102), .C(n65), .D(n64), .Y(prl_rdat[7]) );
  INVX1 U125 ( .A(txbuf[7]), .Y(n64) );
  MUX2BXL U126 ( .D0(n63), .D1(r_dat_spec[1]), .S(n62), .Y(n66) );
  AND2X1 U127 ( .A(txbuf[4]), .B(n49), .Y(prl_rdat[4]) );
  MUX2BXL U128 ( .D0(n60), .D1(r_dat_spec[0]), .S(n62), .Y(n61) );
  NAND21X1 U129 ( .B(prl_fsm[0]), .A(n19), .Y(n24) );
  NAND21XL U130 ( .B(prl_fsm[3]), .A(prl_fsm[0]), .Y(n22) );
  NAND21X1 U131 ( .B(c0_cnt[7]), .A(n111), .Y(n116) );
  NAND21X1 U132 ( .B(c0_cnt[2]), .A(n124), .Y(n122) );
  NAND21X1 U133 ( .B(c0_cnt[3]), .A(n118), .Y(n131) );
  NAND21X1 U134 ( .B(c0_cnt[4]), .A(n121), .Y(n127) );
  NAND21X1 U135 ( .B(c0_cnt[5]), .A(n130), .Y(n112) );
  NAND21X1 U136 ( .B(c0_cnt[6]), .A(n126), .Y(n115) );
  OR2X1 U137 ( .A(c0_cnt[0]), .B(c0_cnt[1]), .Y(n119) );
  NAND21X1 U138 ( .B(n54), .A(n53), .Y(prl_rdat[5]) );
  NOR21XL U139 ( .B(txbuf[5]), .A(n65), .Y(n54) );
  INVX1 U140 ( .A(n55), .Y(n62) );
  NAND21X1 U141 ( .B(n63), .A(r_spec[0]), .Y(n55) );
  INVX1 U142 ( .A(r_spec[1]), .Y(n63) );
  NAND21XL U143 ( .B(n109), .A(prl_fsm[0]), .Y(prl_txauto[4]) );
  NOR21XL U144 ( .B(prx_rcvdords[0]), .A(prx_rcvdords[1]), .Y(n52) );
  INVX1 U145 ( .A(prx_rcvdords[2]), .Y(n50) );
  INVX1 U146 ( .A(prl_cpmsgid[0]), .Y(n43) );
  INVXL U147 ( .A(prl_fsm[0]), .Y(n141) );
  OAI21BX1 U148 ( .C(PrlTo[0]), .B(r_auto_discard), .A(n37), .Y(stoptimer) );
  AND3X1 U149 ( .A(n70), .B(n39), .C(n69), .Y(n37) );
  NAND21X1 U150 ( .B(r_rdy), .A(n38), .Y(N41) );
  OAI21BBX1 U151 ( .A(r_auto_txgdcrc), .B(prx_gdmsgrcvd), .C(n51), .Y(
        sendgdcrc) );
  INVX1 U152 ( .A(c0_iop), .Y(n35) );
  AOI31XL U153 ( .A(n32), .B(n7), .C(n31), .D(n106), .Y(n36) );
  INVX1 U154 ( .A(n79), .Y(n34) );
  AOI21BBXL U155 ( .B(pid_ccidle), .C(prx_eoprcvd), .A(prl_fsm[0]), .Y(n98) );
  MUX2X1 U156 ( .D0(c0_iop), .D1(n145), .S(n144), .Y(n99) );
  AND4X1 U157 ( .A(n147), .B(n143), .C(n142), .D(n141), .Y(n144) );
  INVX1 U158 ( .A(n140), .Y(n143) );
  OA21X1 U159 ( .B(n128), .C(n108), .A(n142), .Y(N193) );
  AND3X1 U160 ( .A(prx_fifowdat[0]), .B(n147), .C(n107), .Y(n108) );
  NAND42X1 U161 ( .C(pff_c0dat[47]), .D(pff_c0dat[45]), .A(n151), .B(n87), .Y(
        n85) );
  NOR3XL U162 ( .A(pff_c0dat[42]), .B(pff_c0dat[44]), .C(pff_c0dat[43]), .Y(
        n87) );
  OR3XL U163 ( .A(pff_c0dat[41]), .B(pff_c0dat[39]), .C(pff_c0dat[38]), .Y(n86) );
  NAND4X1 U164 ( .A(pff_c0dat[33]), .B(pff_c0dat[30]), .C(n96), .D(
        pff_c0dat[2]), .Y(n94) );
  AND2X1 U168 ( .A(pff_c0dat[24]), .B(pff_c0dat[21]), .Y(n96) );
  NOR3XL U169 ( .A(pff_c0dat[15]), .B(pff_c0dat[18]), .C(pff_c0dat[16]), .Y(
        n93) );
  NAND3X1 U170 ( .A(pff_c0dat[37]), .B(pff_c0dat[35]), .C(pff_c0dat[3]), .Y(
        n95) );
  INVX1 U171 ( .A(prl_cany0), .Y(n151) );
  GEN2XL U172 ( .D(c0_cnt[4]), .E(n131), .C(n130), .B(n133), .A(n129), .Y(N169) );
  AND2X1 U173 ( .A(n128), .B(n136), .Y(n129) );
  AO22X1 U174 ( .A(N120), .B(n139), .C(n138), .D(prx_fifowdat[7]), .Y(N158) );
  GEN2XL U175 ( .D(c0_cnt[5]), .E(n127), .C(n126), .B(n133), .A(n125), .Y(N170) );
  AND2X1 U176 ( .A(n128), .B(n135), .Y(n125) );
  GEN2XL U177 ( .D(c0_cnt[6]), .E(n112), .C(n111), .B(n133), .A(n110), .Y(N171) );
  AND2X1 U178 ( .A(n128), .B(n134), .Y(n110) );
  GEN2XL U179 ( .D(c0_cnt[7]), .E(n115), .C(n114), .B(n133), .A(n113), .Y(N172) );
  AND2X1 U180 ( .A(n128), .B(prx_fifowdat[7]), .Y(n113) );
  NAND2X1 U181 ( .A(pid_ccidle), .B(PrlTo[0]), .Y(n39) );
  AND2X1 U182 ( .A(n11), .B(n151), .Y(prl_GCTxDone) );
  AND2X1 U183 ( .A(r_auto_discard), .B(PrlTo[1]), .Y(n68) );
  INVX1 U184 ( .A(n70), .Y(prl_discard) );
  INVX1 U185 ( .A(prx_fifowdat[2]), .Y(n154) );
  NAND21X1 U186 ( .B(n132), .A(pid_ccidle), .Y(n32) );
  NOR21XL U187 ( .B(n133), .A(n13), .Y(N173) );
  GEN2XL U188 ( .D(c0_cnt[0]), .E(c0_cnt[1]), .C(n124), .B(n133), .A(n123), 
        .Y(N166) );
  AND2X1 U189 ( .A(n128), .B(n145), .Y(n123) );
  GEN2XL U190 ( .D(c0_cnt[2]), .E(n119), .C(n118), .B(n133), .A(n117), .Y(N167) );
  AND2X1 U191 ( .A(n128), .B(n137), .Y(n117) );
  GEN2XL U192 ( .D(c0_cnt[3]), .E(n122), .C(n121), .B(n133), .A(n120), .Y(N168) );
  AND2X1 U193 ( .A(n128), .B(prx_fifowdat[3]), .Y(n120) );
  INVX1 U194 ( .A(prx_fifowdat[0]), .Y(n155) );
  AO22X1 U195 ( .A(N113), .B(n139), .C(n138), .D(prx_fifowdat[0]), .Y(N151) );
  INVX1 U196 ( .A(n153), .Y(n145) );
  INVX1 U197 ( .A(prx_fifowdat[1]), .Y(n153) );
  INVXL U198 ( .A(prx_fifowdat[4]), .Y(n149) );
  INVXL U199 ( .A(prx_fifowdat[6]), .Y(n150) );
  INVXL U200 ( .A(prx_fifowdat[5]), .Y(n148) );
  NOR3XL U201 ( .A(prx_fifowdat[5]), .B(prx_fifowdat[7]), .C(prx_fifowdat[6]), 
        .Y(n101) );
  AND2XL U202 ( .A(n142), .B(prl_cany0r), .Y(N196) );
  INVXL U203 ( .A(prl_cany0r), .Y(n38) );
  OAI22X1 U204 ( .A(n30), .B(n132), .C(n9), .D(n31), .Y(prl_cany0r) );
  NAND32XL U205 ( .B(prl_fsm[2]), .C(n19), .A(n23), .Y(n109) );
  AO21XL U206 ( .B(n33), .C(n71), .A(n30), .Y(n28) );
  AO22XL U207 ( .A(n36), .B(n35), .C(n34), .D(prx_fifopsh), .Y(N194) );
  AND3X1 U208 ( .A(prx_fifopsh), .B(n72), .C(n107), .Y(n21) );
endmodule


module updprl_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module PrlTimer_1112a0 ( to, restart, stop, clk, srstz, test_si, test_so, 
        test_se );
  output [1:0] to;
  input restart, stop, clk, srstz, test_si, test_se;
  output test_so;
  wire   timer_10_, timer_9_, timer_8_, timer_7_, timer_6_, timer_5_, timer_4_,
         timer_3_, timer_2_, timer_1_, timer_0_, ena, N4, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, net10360, n7, n8, n9, n10, n11, n12, n13, n1,
         n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 clk_gate_timer_reg ( .CLK(clk), .EN(N18), .ENCLK(net10360), .TE(test_se) );
  PrlTimer_1112a0_DW01_inc_0 add_25 ( .A({test_so, timer_10_, timer_9_, 
        timer_8_, timer_7_, timer_6_, timer_5_, timer_4_, timer_3_, timer_2_, 
        timer_1_, timer_0_}), .SUM({N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, N4}) );
  SDFFQX1 ena_reg ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .Q(ena) );
  SDFFQX1 timer_reg_1_ ( .D(N20), .SIN(timer_0_), .SMC(test_se), .C(net10360), 
        .Q(timer_1_) );
  SDFFQX1 timer_reg_2_ ( .D(N21), .SIN(timer_1_), .SMC(test_se), .C(net10360), 
        .Q(timer_2_) );
  SDFFQX1 timer_reg_0_ ( .D(N19), .SIN(ena), .SMC(test_se), .C(net10360), .Q(
        timer_0_) );
  SDFFQX1 timer_reg_11_ ( .D(N30), .SIN(timer_10_), .SMC(test_se), .C(net10360), .Q(test_so) );
  SDFFQX1 timer_reg_9_ ( .D(N28), .SIN(timer_8_), .SMC(test_se), .C(net10360), 
        .Q(timer_9_) );
  SDFFQX1 timer_reg_10_ ( .D(N29), .SIN(timer_9_), .SMC(test_se), .C(net10360), 
        .Q(timer_10_) );
  SDFFQX1 timer_reg_7_ ( .D(N26), .SIN(timer_6_), .SMC(test_se), .C(net10360), 
        .Q(timer_7_) );
  SDFFQX1 timer_reg_6_ ( .D(N25), .SIN(timer_5_), .SMC(test_se), .C(net10360), 
        .Q(timer_6_) );
  SDFFQX1 timer_reg_8_ ( .D(N27), .SIN(timer_7_), .SMC(test_se), .C(net10360), 
        .Q(timer_8_) );
  SDFFQX1 timer_reg_3_ ( .D(N22), .SIN(timer_2_), .SMC(test_se), .C(net10360), 
        .Q(timer_3_) );
  SDFFQX1 timer_reg_4_ ( .D(N23), .SIN(timer_3_), .SMC(test_se), .C(net10360), 
        .Q(timer_4_) );
  SDFFQX1 timer_reg_5_ ( .D(N24), .SIN(timer_4_), .SMC(test_se), .C(net10360), 
        .Q(timer_5_) );
  BUFX3 U3 ( .A(n11), .Y(n1) );
  NOR21XL U4 ( .B(N9), .A(n11), .Y(N24) );
  NOR21XL U5 ( .B(N7), .A(n11), .Y(N22) );
  NOR21XL U6 ( .B(N8), .A(n11), .Y(N23) );
  NOR21XL U7 ( .B(N13), .A(n11), .Y(N28) );
  NOR21XL U8 ( .B(N12), .A(n11), .Y(N27) );
  NOR21XL U9 ( .B(N11), .A(n11), .Y(N26) );
  NOR21XL U10 ( .B(N10), .A(n11), .Y(N25) );
  NOR21XL U11 ( .B(N14), .A(n11), .Y(N29) );
  NOR21XL U12 ( .B(N6), .A(n11), .Y(N21) );
  NOR21XL U13 ( .B(N5), .A(n1), .Y(N20) );
  NAND31X1 U14 ( .C(restart), .A(n1), .B(srstz), .Y(N18) );
  NAND3X1 U15 ( .A(srstz), .B(ena), .C(n12), .Y(n11) );
  NOR3XL U16 ( .A(to[1]), .B(stop), .C(restart), .Y(n12) );
  NOR21XL U17 ( .B(N15), .A(n1), .Y(N30) );
  NOR21XL U18 ( .B(N4), .A(n1), .Y(N19) );
  INVX1 U19 ( .A(n10), .Y(n2) );
  AOI31X1 U20 ( .A(srstz), .B(n3), .C(ena), .D(restart), .Y(n10) );
  INVX1 U21 ( .A(stop), .Y(n3) );
  INVX1 U22 ( .A(n7), .Y(to[0]) );
  AOI211X1 U23 ( .C(n4), .D(timer_9_), .A(timer_10_), .B(test_so), .Y(n7) );
  INVX1 U24 ( .A(n8), .Y(n4) );
  AOI211X1 U25 ( .C(timer_6_), .D(n9), .A(timer_8_), .B(timer_7_), .Y(n8) );
  AO21X1 U26 ( .B(timer_4_), .C(timer_3_), .A(timer_5_), .Y(n9) );
  OAI31XL U27 ( .A(timer_10_), .B(timer_9_), .C(timer_8_), .D(test_so), .Y(n13) );
  INVX1 U28 ( .A(n13), .Y(to[1]) );
endmodule


module PrlTimer_1112a0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyff_DEPTH_NUM34_DEPTH_NBT6 ( r_psh, r_pop, prx_psh, ptx_pop, r_last, 
        r_unlock, i_lockena, r_fiforst, i_ccidle, r_wdat, prx_wdat, txreq, 
        ffack, rdat0, full, empty, one, half, obsd, dat_7_1, ptr, fifowdat, 
        fifopsh, clk, srstz, test_si, test_se );
  input [7:0] r_wdat;
  input [7:0] prx_wdat;
  output [1:0] ffack;
  output [7:0] rdat0;
  output [55:0] dat_7_1;
  output [5:0] ptr;
  output [7:0] fifowdat;
  input r_psh, r_pop, prx_psh, ptx_pop, r_last, r_unlock, i_lockena, r_fiforst,
         i_ccidle, clk, srstz, test_si, test_se;
  output txreq, full, empty, one, half, obsd, fifopsh;
  wire   ps_locked, locked, mem_8__7_, mem_8__6_, mem_8__5_, mem_8__4_,
         mem_8__3_, mem_8__2_, mem_8__1_, mem_8__0_, mem_9__7_, mem_9__6_,
         mem_9__5_, mem_9__4_, mem_9__3_, mem_9__2_, mem_9__1_, mem_9__0_,
         mem_10__7_, mem_10__6_, mem_10__5_, mem_10__4_, mem_10__3_,
         mem_10__2_, mem_10__1_, mem_10__0_, mem_11__7_, mem_11__6_,
         mem_11__5_, mem_11__4_, mem_11__3_, mem_11__2_, mem_11__1_,
         mem_11__0_, mem_12__7_, mem_12__6_, mem_12__5_, mem_12__4_,
         mem_12__3_, mem_12__2_, mem_12__1_, mem_12__0_, mem_13__7_,
         mem_13__6_, mem_13__5_, mem_13__4_, mem_13__3_, mem_13__2_,
         mem_13__1_, mem_13__0_, mem_14__7_, mem_14__6_, mem_14__5_,
         mem_14__4_, mem_14__3_, mem_14__2_, mem_14__1_, mem_14__0_,
         mem_15__7_, mem_15__6_, mem_15__5_, mem_15__4_, mem_15__3_,
         mem_15__2_, mem_15__1_, mem_15__0_, mem_16__7_, mem_16__6_,
         mem_16__5_, mem_16__4_, mem_16__3_, mem_16__2_, mem_16__1_,
         mem_16__0_, mem_17__7_, mem_17__6_, mem_17__5_, mem_17__4_,
         mem_17__3_, mem_17__2_, mem_17__1_, mem_17__0_, mem_18__7_,
         mem_18__6_, mem_18__5_, mem_18__4_, mem_18__3_, mem_18__2_,
         mem_18__1_, mem_18__0_, mem_19__7_, mem_19__6_, mem_19__5_,
         mem_19__4_, mem_19__3_, mem_19__2_, mem_19__1_, mem_19__0_,
         mem_20__7_, mem_20__6_, mem_20__5_, mem_20__4_, mem_20__3_,
         mem_20__2_, mem_20__1_, mem_20__0_, mem_21__7_, mem_21__6_,
         mem_21__5_, mem_21__4_, mem_21__3_, mem_21__2_, mem_21__1_,
         mem_21__0_, mem_22__7_, mem_22__6_, mem_22__5_, mem_22__4_,
         mem_22__3_, mem_22__2_, mem_22__1_, mem_22__0_, mem_23__7_,
         mem_23__6_, mem_23__5_, mem_23__4_, mem_23__3_, mem_23__2_,
         mem_23__1_, mem_23__0_, mem_24__7_, mem_24__6_, mem_24__5_,
         mem_24__4_, mem_24__3_, mem_24__2_, mem_24__1_, mem_24__0_,
         mem_25__7_, mem_25__6_, mem_25__5_, mem_25__4_, mem_25__3_,
         mem_25__2_, mem_25__1_, mem_25__0_, mem_26__7_, mem_26__6_,
         mem_26__5_, mem_26__4_, mem_26__3_, mem_26__2_, mem_26__1_,
         mem_26__0_, mem_27__7_, mem_27__6_, mem_27__5_, mem_27__4_,
         mem_27__3_, mem_27__2_, mem_27__1_, mem_27__0_, mem_28__7_,
         mem_28__6_, mem_28__5_, mem_28__4_, mem_28__3_, mem_28__2_,
         mem_28__1_, mem_28__0_, mem_29__7_, mem_29__6_, mem_29__5_,
         mem_29__4_, mem_29__3_, mem_29__2_, mem_29__1_, mem_29__0_,
         mem_30__7_, mem_30__6_, mem_30__5_, mem_30__4_, mem_30__3_,
         mem_30__2_, mem_30__1_, mem_30__0_, mem_31__7_, mem_31__6_,
         mem_31__5_, mem_31__4_, mem_31__3_, mem_31__2_, mem_31__1_,
         mem_31__0_, mem_32__7_, mem_32__6_, mem_32__5_, mem_32__4_,
         mem_32__3_, mem_32__2_, mem_32__1_, mem_32__0_, mem_33__7_,
         mem_33__6_, mem_33__5_, mem_33__4_, mem_33__3_, mem_33__2_,
         mem_33__1_, mem_33__0_, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1053, N1054, N1055,
         N1056, N1057, N1058, N1059, net10378, net10384, net10389, net10394,
         net10399, net10404, net10409, net10414, net10419, net10424, net10429,
         net10434, net10439, net10444, net10449, net10454, net10459, net10464,
         net10469, net10474, net10479, net10484, net10489, net10494, net10499,
         net10504, net10509, net10514, net10519, net10524, net10529, net10534,
         net10539, net10544, net10549, n44, n45, n47, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38,
         n39, n41, n42, n43, n46, n48, n113, n220, n439, n480, n482, n483,
         n484, n485, n486, n488, n489, n490, n491, n492, n493, n494, n496,
         n497, n498, n499, n500, n501, n502, n504, n505, n506, n507, n508,
         n509, n510, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551;

  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 clk_gate_mem_reg_0_ ( 
        .CLK(clk), .EN(N1022), .ENCLK(net10378), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 clk_gate_mem_reg_1_ ( 
        .CLK(clk), .EN(N1013), .ENCLK(net10384), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 clk_gate_mem_reg_2_ ( 
        .CLK(clk), .EN(N1004), .ENCLK(net10389), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 clk_gate_mem_reg_3_ ( 
        .CLK(clk), .EN(N995), .ENCLK(net10394), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 clk_gate_mem_reg_4_ ( 
        .CLK(clk), .EN(N986), .ENCLK(net10399), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 clk_gate_mem_reg_5_ ( 
        .CLK(clk), .EN(N977), .ENCLK(net10404), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 clk_gate_mem_reg_6_ ( 
        .CLK(clk), .EN(N968), .ENCLK(net10409), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 clk_gate_mem_reg_7_ ( 
        .CLK(clk), .EN(N959), .ENCLK(net10414), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 clk_gate_mem_reg_8_ ( 
        .CLK(clk), .EN(N950), .ENCLK(net10419), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 clk_gate_mem_reg_9_ ( 
        .CLK(clk), .EN(N941), .ENCLK(net10424), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 clk_gate_mem_reg_10_ ( 
        .CLK(clk), .EN(N932), .ENCLK(net10429), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 clk_gate_mem_reg_11_ ( 
        .CLK(clk), .EN(N923), .ENCLK(net10434), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 clk_gate_mem_reg_12_ ( 
        .CLK(clk), .EN(N914), .ENCLK(net10439), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 clk_gate_mem_reg_13_ ( 
        .CLK(clk), .EN(N905), .ENCLK(net10444), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 clk_gate_mem_reg_14_ ( 
        .CLK(clk), .EN(N896), .ENCLK(net10449), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 clk_gate_mem_reg_15_ ( 
        .CLK(clk), .EN(N887), .ENCLK(net10454), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 clk_gate_mem_reg_16_ ( 
        .CLK(clk), .EN(N878), .ENCLK(net10459), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 clk_gate_mem_reg_17_ ( 
        .CLK(clk), .EN(N869), .ENCLK(net10464), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 clk_gate_mem_reg_18_ ( 
        .CLK(clk), .EN(N860), .ENCLK(net10469), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 clk_gate_mem_reg_19_ ( 
        .CLK(clk), .EN(N851), .ENCLK(net10474), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 clk_gate_mem_reg_20_ ( 
        .CLK(clk), .EN(N842), .ENCLK(net10479), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 clk_gate_mem_reg_21_ ( 
        .CLK(clk), .EN(N833), .ENCLK(net10484), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 clk_gate_mem_reg_22_ ( 
        .CLK(clk), .EN(N824), .ENCLK(net10489), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 clk_gate_mem_reg_23_ ( 
        .CLK(clk), .EN(N815), .ENCLK(net10494), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 clk_gate_mem_reg_24_ ( 
        .CLK(clk), .EN(N806), .ENCLK(net10499), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 clk_gate_mem_reg_25_ ( 
        .CLK(clk), .EN(N797), .ENCLK(net10504), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 clk_gate_mem_reg_26_ ( 
        .CLK(clk), .EN(N788), .ENCLK(net10509), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 clk_gate_mem_reg_27_ ( 
        .CLK(clk), .EN(N779), .ENCLK(net10514), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 clk_gate_mem_reg_28_ ( 
        .CLK(clk), .EN(N770), .ENCLK(net10519), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 clk_gate_mem_reg_29_ ( 
        .CLK(clk), .EN(N761), .ENCLK(net10524), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 clk_gate_mem_reg_30_ ( 
        .CLK(clk), .EN(N752), .ENCLK(net10529), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 clk_gate_mem_reg_31_ ( 
        .CLK(clk), .EN(N743), .ENCLK(net10534), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 clk_gate_mem_reg_32_ ( 
        .CLK(clk), .EN(N734), .ENCLK(net10539), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 clk_gate_mem_reg_33_ ( 
        .CLK(clk), .EN(N733), .ENCLK(net10544), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 clk_gate_pshptr_reg ( 
        .CLK(clk), .EN(N1053), .ENCLK(net10549), .TE(test_se) );
  SDFFQX1 mem_reg_33__7_ ( .D(fifowdat[7]), .SIN(mem_33__6_), .SMC(test_se), 
        .C(net10544), .Q(mem_33__7_) );
  SDFFQX1 mem_reg_32__7_ ( .D(N742), .SIN(mem_32__6_), .SMC(test_se), .C(
        net10539), .Q(mem_32__7_) );
  SDFFQX1 mem_reg_31__7_ ( .D(N751), .SIN(mem_31__6_), .SMC(test_se), .C(
        net10534), .Q(mem_31__7_) );
  SDFFQX1 mem_reg_30__7_ ( .D(N760), .SIN(mem_30__6_), .SMC(test_se), .C(
        net10529), .Q(mem_30__7_) );
  SDFFQX1 mem_reg_29__7_ ( .D(N769), .SIN(mem_29__6_), .SMC(test_se), .C(
        net10524), .Q(mem_29__7_) );
  SDFFQX1 mem_reg_28__7_ ( .D(N778), .SIN(mem_28__6_), .SMC(test_se), .C(
        net10519), .Q(mem_28__7_) );
  SDFFQX1 mem_reg_33__6_ ( .D(fifowdat[6]), .SIN(mem_33__5_), .SMC(test_se), 
        .C(net10544), .Q(mem_33__6_) );
  SDFFQX1 mem_reg_32__6_ ( .D(N741), .SIN(mem_32__5_), .SMC(test_se), .C(
        net10539), .Q(mem_32__6_) );
  SDFFQX1 mem_reg_31__6_ ( .D(N750), .SIN(mem_31__5_), .SMC(test_se), .C(
        net10534), .Q(mem_31__6_) );
  SDFFQX1 mem_reg_30__6_ ( .D(N759), .SIN(mem_30__5_), .SMC(test_se), .C(
        net10529), .Q(mem_30__6_) );
  SDFFQX1 mem_reg_29__6_ ( .D(N768), .SIN(mem_29__5_), .SMC(test_se), .C(
        net10524), .Q(mem_29__6_) );
  SDFFQX1 mem_reg_28__6_ ( .D(N777), .SIN(mem_28__5_), .SMC(test_se), .C(
        net10519), .Q(mem_28__6_) );
  SDFFQX1 mem_reg_33__5_ ( .D(fifowdat[5]), .SIN(mem_33__4_), .SMC(test_se), 
        .C(net10544), .Q(mem_33__5_) );
  SDFFQX1 mem_reg_32__5_ ( .D(N740), .SIN(mem_32__4_), .SMC(test_se), .C(
        net10539), .Q(mem_32__5_) );
  SDFFQX1 mem_reg_31__5_ ( .D(N749), .SIN(mem_31__4_), .SMC(test_se), .C(
        net10534), .Q(mem_31__5_) );
  SDFFQX1 mem_reg_30__5_ ( .D(N758), .SIN(mem_30__4_), .SMC(test_se), .C(
        net10529), .Q(mem_30__5_) );
  SDFFQX1 mem_reg_29__5_ ( .D(N767), .SIN(mem_29__4_), .SMC(test_se), .C(
        net10524), .Q(mem_29__5_) );
  SDFFQX1 mem_reg_28__5_ ( .D(N776), .SIN(mem_28__4_), .SMC(test_se), .C(
        net10519), .Q(mem_28__5_) );
  SDFFQX1 mem_reg_33__4_ ( .D(fifowdat[4]), .SIN(mem_33__3_), .SMC(test_se), 
        .C(net10544), .Q(mem_33__4_) );
  SDFFQX1 mem_reg_32__4_ ( .D(N739), .SIN(mem_32__3_), .SMC(test_se), .C(
        net10539), .Q(mem_32__4_) );
  SDFFQX1 mem_reg_31__4_ ( .D(N748), .SIN(mem_31__3_), .SMC(test_se), .C(
        net10534), .Q(mem_31__4_) );
  SDFFQX1 mem_reg_30__4_ ( .D(N757), .SIN(mem_30__3_), .SMC(test_se), .C(
        net10529), .Q(mem_30__4_) );
  SDFFQX1 mem_reg_29__4_ ( .D(N766), .SIN(mem_29__3_), .SMC(test_se), .C(
        net10524), .Q(mem_29__4_) );
  SDFFQX1 mem_reg_28__4_ ( .D(N775), .SIN(mem_28__3_), .SMC(test_se), .C(
        net10519), .Q(mem_28__4_) );
  SDFFQX1 mem_reg_33__3_ ( .D(fifowdat[3]), .SIN(mem_33__2_), .SMC(test_se), 
        .C(net10544), .Q(mem_33__3_) );
  SDFFQX1 mem_reg_32__3_ ( .D(N738), .SIN(mem_32__2_), .SMC(test_se), .C(
        net10539), .Q(mem_32__3_) );
  SDFFQX1 mem_reg_31__3_ ( .D(N747), .SIN(mem_31__2_), .SMC(test_se), .C(
        net10534), .Q(mem_31__3_) );
  SDFFQX1 mem_reg_30__3_ ( .D(N756), .SIN(mem_30__2_), .SMC(test_se), .C(
        net10529), .Q(mem_30__3_) );
  SDFFQX1 mem_reg_29__3_ ( .D(N765), .SIN(mem_29__2_), .SMC(test_se), .C(
        net10524), .Q(mem_29__3_) );
  SDFFQX1 mem_reg_28__3_ ( .D(N774), .SIN(mem_28__2_), .SMC(test_se), .C(
        net10519), .Q(mem_28__3_) );
  SDFFQX1 mem_reg_33__2_ ( .D(fifowdat[2]), .SIN(mem_33__1_), .SMC(test_se), 
        .C(net10544), .Q(mem_33__2_) );
  SDFFQX1 mem_reg_32__2_ ( .D(N737), .SIN(mem_32__1_), .SMC(test_se), .C(
        net10539), .Q(mem_32__2_) );
  SDFFQX1 mem_reg_31__2_ ( .D(N746), .SIN(mem_31__1_), .SMC(test_se), .C(
        net10534), .Q(mem_31__2_) );
  SDFFQX1 mem_reg_30__2_ ( .D(N755), .SIN(mem_30__1_), .SMC(test_se), .C(
        net10529), .Q(mem_30__2_) );
  SDFFQX1 mem_reg_29__2_ ( .D(N764), .SIN(mem_29__1_), .SMC(test_se), .C(
        net10524), .Q(mem_29__2_) );
  SDFFQX1 mem_reg_28__2_ ( .D(N773), .SIN(mem_28__1_), .SMC(test_se), .C(
        net10519), .Q(mem_28__2_) );
  SDFFQX1 mem_reg_33__1_ ( .D(fifowdat[1]), .SIN(mem_33__0_), .SMC(test_se), 
        .C(net10544), .Q(mem_33__1_) );
  SDFFQX1 mem_reg_32__1_ ( .D(N736), .SIN(mem_32__0_), .SMC(test_se), .C(
        net10539), .Q(mem_32__1_) );
  SDFFQX1 mem_reg_31__1_ ( .D(N745), .SIN(mem_31__0_), .SMC(test_se), .C(
        net10534), .Q(mem_31__1_) );
  SDFFQX1 mem_reg_30__1_ ( .D(N754), .SIN(mem_30__0_), .SMC(test_se), .C(
        net10529), .Q(mem_30__1_) );
  SDFFQX1 mem_reg_29__1_ ( .D(N763), .SIN(mem_29__0_), .SMC(test_se), .C(
        net10524), .Q(mem_29__1_) );
  SDFFQX1 mem_reg_28__1_ ( .D(N772), .SIN(mem_28__0_), .SMC(test_se), .C(
        net10519), .Q(mem_28__1_) );
  SDFFQX1 mem_reg_33__0_ ( .D(fifowdat[0]), .SIN(mem_32__7_), .SMC(test_se), 
        .C(net10544), .Q(mem_33__0_) );
  SDFFQX1 mem_reg_32__0_ ( .D(N735), .SIN(mem_31__7_), .SMC(test_se), .C(
        net10539), .Q(mem_32__0_) );
  SDFFQX1 mem_reg_31__0_ ( .D(N744), .SIN(mem_30__7_), .SMC(test_se), .C(
        net10534), .Q(mem_31__0_) );
  SDFFQX1 mem_reg_30__0_ ( .D(N753), .SIN(mem_29__7_), .SMC(test_se), .C(
        net10529), .Q(mem_30__0_) );
  SDFFQX1 mem_reg_29__0_ ( .D(N762), .SIN(mem_28__7_), .SMC(test_se), .C(
        net10524), .Q(mem_29__0_) );
  SDFFQX1 mem_reg_28__0_ ( .D(N771), .SIN(mem_27__7_), .SMC(test_se), .C(
        net10519), .Q(mem_28__0_) );
  SDFFQX1 mem_reg_27__7_ ( .D(N787), .SIN(mem_27__6_), .SMC(test_se), .C(
        net10514), .Q(mem_27__7_) );
  SDFFQX1 mem_reg_26__7_ ( .D(N796), .SIN(mem_26__6_), .SMC(test_se), .C(
        net10509), .Q(mem_26__7_) );
  SDFFQX1 mem_reg_25__7_ ( .D(N805), .SIN(mem_25__6_), .SMC(test_se), .C(
        net10504), .Q(mem_25__7_) );
  SDFFQX1 mem_reg_24__7_ ( .D(N814), .SIN(mem_24__6_), .SMC(test_se), .C(
        net10499), .Q(mem_24__7_) );
  SDFFQX1 mem_reg_23__7_ ( .D(N823), .SIN(mem_23__6_), .SMC(test_se), .C(
        net10494), .Q(mem_23__7_) );
  SDFFQX1 mem_reg_22__7_ ( .D(N832), .SIN(mem_22__6_), .SMC(test_se), .C(
        net10489), .Q(mem_22__7_) );
  SDFFQX1 mem_reg_21__7_ ( .D(N841), .SIN(mem_21__6_), .SMC(test_se), .C(
        net10484), .Q(mem_21__7_) );
  SDFFQX1 mem_reg_20__7_ ( .D(N850), .SIN(mem_20__6_), .SMC(test_se), .C(
        net10479), .Q(mem_20__7_) );
  SDFFQX1 mem_reg_19__7_ ( .D(N859), .SIN(mem_19__6_), .SMC(test_se), .C(
        net10474), .Q(mem_19__7_) );
  SDFFQX1 mem_reg_18__7_ ( .D(N868), .SIN(mem_18__6_), .SMC(test_se), .C(
        net10469), .Q(mem_18__7_) );
  SDFFQX1 mem_reg_17__7_ ( .D(N877), .SIN(mem_17__6_), .SMC(test_se), .C(
        net10464), .Q(mem_17__7_) );
  SDFFQX1 mem_reg_16__7_ ( .D(N886), .SIN(mem_16__6_), .SMC(test_se), .C(
        net10459), .Q(mem_16__7_) );
  SDFFQX1 mem_reg_15__7_ ( .D(N895), .SIN(mem_15__6_), .SMC(test_se), .C(
        net10454), .Q(mem_15__7_) );
  SDFFQX1 mem_reg_14__7_ ( .D(N904), .SIN(mem_14__6_), .SMC(test_se), .C(
        net10449), .Q(mem_14__7_) );
  SDFFQX1 mem_reg_13__7_ ( .D(N913), .SIN(mem_13__6_), .SMC(test_se), .C(
        net10444), .Q(mem_13__7_) );
  SDFFQX1 mem_reg_12__7_ ( .D(N922), .SIN(mem_12__6_), .SMC(test_se), .C(
        net10439), .Q(mem_12__7_) );
  SDFFQX1 mem_reg_11__7_ ( .D(N931), .SIN(mem_11__6_), .SMC(test_se), .C(
        net10434), .Q(mem_11__7_) );
  SDFFQX1 mem_reg_10__7_ ( .D(N940), .SIN(mem_10__6_), .SMC(test_se), .C(
        net10429), .Q(mem_10__7_) );
  SDFFQX1 mem_reg_9__7_ ( .D(N949), .SIN(mem_9__6_), .SMC(test_se), .C(
        net10424), .Q(mem_9__7_) );
  SDFFQX1 mem_reg_8__7_ ( .D(N958), .SIN(mem_8__6_), .SMC(test_se), .C(
        net10419), .Q(mem_8__7_) );
  SDFFQX1 mem_reg_27__6_ ( .D(N786), .SIN(mem_27__5_), .SMC(test_se), .C(
        net10514), .Q(mem_27__6_) );
  SDFFQX1 mem_reg_26__6_ ( .D(N795), .SIN(mem_26__5_), .SMC(test_se), .C(
        net10509), .Q(mem_26__6_) );
  SDFFQX1 mem_reg_25__6_ ( .D(N804), .SIN(mem_25__5_), .SMC(test_se), .C(
        net10504), .Q(mem_25__6_) );
  SDFFQX1 mem_reg_24__6_ ( .D(N813), .SIN(mem_24__5_), .SMC(test_se), .C(
        net10499), .Q(mem_24__6_) );
  SDFFQX1 mem_reg_23__6_ ( .D(N822), .SIN(mem_23__5_), .SMC(test_se), .C(
        net10494), .Q(mem_23__6_) );
  SDFFQX1 mem_reg_22__6_ ( .D(N831), .SIN(mem_22__5_), .SMC(test_se), .C(
        net10489), .Q(mem_22__6_) );
  SDFFQX1 mem_reg_21__6_ ( .D(N840), .SIN(mem_21__5_), .SMC(test_se), .C(
        net10484), .Q(mem_21__6_) );
  SDFFQX1 mem_reg_20__6_ ( .D(N849), .SIN(mem_20__5_), .SMC(test_se), .C(
        net10479), .Q(mem_20__6_) );
  SDFFQX1 mem_reg_19__6_ ( .D(N858), .SIN(mem_19__5_), .SMC(test_se), .C(
        net10474), .Q(mem_19__6_) );
  SDFFQX1 mem_reg_18__6_ ( .D(N867), .SIN(mem_18__5_), .SMC(test_se), .C(
        net10469), .Q(mem_18__6_) );
  SDFFQX1 mem_reg_17__6_ ( .D(N876), .SIN(mem_17__5_), .SMC(test_se), .C(
        net10464), .Q(mem_17__6_) );
  SDFFQX1 mem_reg_16__6_ ( .D(N885), .SIN(mem_16__5_), .SMC(test_se), .C(
        net10459), .Q(mem_16__6_) );
  SDFFQX1 mem_reg_15__6_ ( .D(N894), .SIN(mem_15__5_), .SMC(test_se), .C(
        net10454), .Q(mem_15__6_) );
  SDFFQX1 mem_reg_14__6_ ( .D(N903), .SIN(mem_14__5_), .SMC(test_se), .C(
        net10449), .Q(mem_14__6_) );
  SDFFQX1 mem_reg_13__6_ ( .D(N912), .SIN(mem_13__5_), .SMC(test_se), .C(
        net10444), .Q(mem_13__6_) );
  SDFFQX1 mem_reg_12__6_ ( .D(N921), .SIN(mem_12__5_), .SMC(test_se), .C(
        net10439), .Q(mem_12__6_) );
  SDFFQX1 mem_reg_11__6_ ( .D(N930), .SIN(mem_11__5_), .SMC(test_se), .C(
        net10434), .Q(mem_11__6_) );
  SDFFQX1 mem_reg_10__6_ ( .D(N939), .SIN(mem_10__5_), .SMC(test_se), .C(
        net10429), .Q(mem_10__6_) );
  SDFFQX1 mem_reg_9__6_ ( .D(N948), .SIN(mem_9__5_), .SMC(test_se), .C(
        net10424), .Q(mem_9__6_) );
  SDFFQX1 mem_reg_8__6_ ( .D(N957), .SIN(mem_8__5_), .SMC(test_se), .C(
        net10419), .Q(mem_8__6_) );
  SDFFQX1 mem_reg_27__5_ ( .D(N785), .SIN(mem_27__4_), .SMC(test_se), .C(
        net10514), .Q(mem_27__5_) );
  SDFFQX1 mem_reg_26__5_ ( .D(N794), .SIN(mem_26__4_), .SMC(test_se), .C(
        net10509), .Q(mem_26__5_) );
  SDFFQX1 mem_reg_25__5_ ( .D(N803), .SIN(mem_25__4_), .SMC(test_se), .C(
        net10504), .Q(mem_25__5_) );
  SDFFQX1 mem_reg_24__5_ ( .D(N812), .SIN(mem_24__4_), .SMC(test_se), .C(
        net10499), .Q(mem_24__5_) );
  SDFFQX1 mem_reg_23__5_ ( .D(N821), .SIN(mem_23__4_), .SMC(test_se), .C(
        net10494), .Q(mem_23__5_) );
  SDFFQX1 mem_reg_22__5_ ( .D(N830), .SIN(mem_22__4_), .SMC(test_se), .C(
        net10489), .Q(mem_22__5_) );
  SDFFQX1 mem_reg_21__5_ ( .D(N839), .SIN(mem_21__4_), .SMC(test_se), .C(
        net10484), .Q(mem_21__5_) );
  SDFFQX1 mem_reg_20__5_ ( .D(N848), .SIN(mem_20__4_), .SMC(test_se), .C(
        net10479), .Q(mem_20__5_) );
  SDFFQX1 mem_reg_19__5_ ( .D(N857), .SIN(mem_19__4_), .SMC(test_se), .C(
        net10474), .Q(mem_19__5_) );
  SDFFQX1 mem_reg_18__5_ ( .D(N866), .SIN(mem_18__4_), .SMC(test_se), .C(
        net10469), .Q(mem_18__5_) );
  SDFFQX1 mem_reg_17__5_ ( .D(N875), .SIN(mem_17__4_), .SMC(test_se), .C(
        net10464), .Q(mem_17__5_) );
  SDFFQX1 mem_reg_16__5_ ( .D(N884), .SIN(mem_16__4_), .SMC(test_se), .C(
        net10459), .Q(mem_16__5_) );
  SDFFQX1 mem_reg_15__5_ ( .D(N893), .SIN(mem_15__4_), .SMC(test_se), .C(
        net10454), .Q(mem_15__5_) );
  SDFFQX1 mem_reg_14__5_ ( .D(N902), .SIN(mem_14__4_), .SMC(test_se), .C(
        net10449), .Q(mem_14__5_) );
  SDFFQX1 mem_reg_13__5_ ( .D(N911), .SIN(mem_13__4_), .SMC(test_se), .C(
        net10444), .Q(mem_13__5_) );
  SDFFQX1 mem_reg_12__5_ ( .D(N920), .SIN(mem_12__4_), .SMC(test_se), .C(
        net10439), .Q(mem_12__5_) );
  SDFFQX1 mem_reg_11__5_ ( .D(N929), .SIN(mem_11__4_), .SMC(test_se), .C(
        net10434), .Q(mem_11__5_) );
  SDFFQX1 mem_reg_10__5_ ( .D(N938), .SIN(mem_10__4_), .SMC(test_se), .C(
        net10429), .Q(mem_10__5_) );
  SDFFQX1 mem_reg_9__5_ ( .D(N947), .SIN(mem_9__4_), .SMC(test_se), .C(
        net10424), .Q(mem_9__5_) );
  SDFFQX1 mem_reg_8__5_ ( .D(N956), .SIN(mem_8__4_), .SMC(test_se), .C(
        net10419), .Q(mem_8__5_) );
  SDFFQX1 mem_reg_27__4_ ( .D(N784), .SIN(mem_27__3_), .SMC(test_se), .C(
        net10514), .Q(mem_27__4_) );
  SDFFQX1 mem_reg_26__4_ ( .D(N793), .SIN(mem_26__3_), .SMC(test_se), .C(
        net10509), .Q(mem_26__4_) );
  SDFFQX1 mem_reg_25__4_ ( .D(N802), .SIN(mem_25__3_), .SMC(test_se), .C(
        net10504), .Q(mem_25__4_) );
  SDFFQX1 mem_reg_24__4_ ( .D(N811), .SIN(mem_24__3_), .SMC(test_se), .C(
        net10499), .Q(mem_24__4_) );
  SDFFQX1 mem_reg_23__4_ ( .D(N820), .SIN(mem_23__3_), .SMC(test_se), .C(
        net10494), .Q(mem_23__4_) );
  SDFFQX1 mem_reg_22__4_ ( .D(N829), .SIN(mem_22__3_), .SMC(test_se), .C(
        net10489), .Q(mem_22__4_) );
  SDFFQX1 mem_reg_21__4_ ( .D(N838), .SIN(mem_21__3_), .SMC(test_se), .C(
        net10484), .Q(mem_21__4_) );
  SDFFQX1 mem_reg_20__4_ ( .D(N847), .SIN(mem_20__3_), .SMC(test_se), .C(
        net10479), .Q(mem_20__4_) );
  SDFFQX1 mem_reg_19__4_ ( .D(N856), .SIN(mem_19__3_), .SMC(test_se), .C(
        net10474), .Q(mem_19__4_) );
  SDFFQX1 mem_reg_18__4_ ( .D(N865), .SIN(mem_18__3_), .SMC(test_se), .C(
        net10469), .Q(mem_18__4_) );
  SDFFQX1 mem_reg_17__4_ ( .D(N874), .SIN(mem_17__3_), .SMC(test_se), .C(
        net10464), .Q(mem_17__4_) );
  SDFFQX1 mem_reg_16__4_ ( .D(N883), .SIN(mem_16__3_), .SMC(test_se), .C(
        net10459), .Q(mem_16__4_) );
  SDFFQX1 mem_reg_15__4_ ( .D(N892), .SIN(mem_15__3_), .SMC(test_se), .C(
        net10454), .Q(mem_15__4_) );
  SDFFQX1 mem_reg_14__4_ ( .D(N901), .SIN(mem_14__3_), .SMC(test_se), .C(
        net10449), .Q(mem_14__4_) );
  SDFFQX1 mem_reg_13__4_ ( .D(N910), .SIN(mem_13__3_), .SMC(test_se), .C(
        net10444), .Q(mem_13__4_) );
  SDFFQX1 mem_reg_12__4_ ( .D(N919), .SIN(mem_12__3_), .SMC(test_se), .C(
        net10439), .Q(mem_12__4_) );
  SDFFQX1 mem_reg_11__4_ ( .D(N928), .SIN(mem_11__3_), .SMC(test_se), .C(
        net10434), .Q(mem_11__4_) );
  SDFFQX1 mem_reg_10__4_ ( .D(N937), .SIN(mem_10__3_), .SMC(test_se), .C(
        net10429), .Q(mem_10__4_) );
  SDFFQX1 mem_reg_9__4_ ( .D(N946), .SIN(mem_9__3_), .SMC(test_se), .C(
        net10424), .Q(mem_9__4_) );
  SDFFQX1 mem_reg_8__4_ ( .D(N955), .SIN(mem_8__3_), .SMC(test_se), .C(
        net10419), .Q(mem_8__4_) );
  SDFFQX1 mem_reg_27__3_ ( .D(N783), .SIN(mem_27__2_), .SMC(test_se), .C(
        net10514), .Q(mem_27__3_) );
  SDFFQX1 mem_reg_26__3_ ( .D(N792), .SIN(mem_26__2_), .SMC(test_se), .C(
        net10509), .Q(mem_26__3_) );
  SDFFQX1 mem_reg_25__3_ ( .D(N801), .SIN(mem_25__2_), .SMC(test_se), .C(
        net10504), .Q(mem_25__3_) );
  SDFFQX1 mem_reg_24__3_ ( .D(N810), .SIN(mem_24__2_), .SMC(test_se), .C(
        net10499), .Q(mem_24__3_) );
  SDFFQX1 mem_reg_23__3_ ( .D(N819), .SIN(mem_23__2_), .SMC(test_se), .C(
        net10494), .Q(mem_23__3_) );
  SDFFQX1 mem_reg_22__3_ ( .D(N828), .SIN(mem_22__2_), .SMC(test_se), .C(
        net10489), .Q(mem_22__3_) );
  SDFFQX1 mem_reg_21__3_ ( .D(N837), .SIN(mem_21__2_), .SMC(test_se), .C(
        net10484), .Q(mem_21__3_) );
  SDFFQX1 mem_reg_20__3_ ( .D(N846), .SIN(mem_20__2_), .SMC(test_se), .C(
        net10479), .Q(mem_20__3_) );
  SDFFQX1 mem_reg_19__3_ ( .D(N855), .SIN(mem_19__2_), .SMC(test_se), .C(
        net10474), .Q(mem_19__3_) );
  SDFFQX1 mem_reg_18__3_ ( .D(N864), .SIN(mem_18__2_), .SMC(test_se), .C(
        net10469), .Q(mem_18__3_) );
  SDFFQX1 mem_reg_17__3_ ( .D(N873), .SIN(mem_17__2_), .SMC(test_se), .C(
        net10464), .Q(mem_17__3_) );
  SDFFQX1 mem_reg_16__3_ ( .D(N882), .SIN(mem_16__2_), .SMC(test_se), .C(
        net10459), .Q(mem_16__3_) );
  SDFFQX1 mem_reg_15__3_ ( .D(N891), .SIN(mem_15__2_), .SMC(test_se), .C(
        net10454), .Q(mem_15__3_) );
  SDFFQX1 mem_reg_14__3_ ( .D(N900), .SIN(mem_14__2_), .SMC(test_se), .C(
        net10449), .Q(mem_14__3_) );
  SDFFQX1 mem_reg_13__3_ ( .D(N909), .SIN(mem_13__2_), .SMC(test_se), .C(
        net10444), .Q(mem_13__3_) );
  SDFFQX1 mem_reg_12__3_ ( .D(N918), .SIN(mem_12__2_), .SMC(test_se), .C(
        net10439), .Q(mem_12__3_) );
  SDFFQX1 mem_reg_11__3_ ( .D(N927), .SIN(mem_11__2_), .SMC(test_se), .C(
        net10434), .Q(mem_11__3_) );
  SDFFQX1 mem_reg_10__3_ ( .D(N936), .SIN(mem_10__2_), .SMC(test_se), .C(
        net10429), .Q(mem_10__3_) );
  SDFFQX1 mem_reg_9__3_ ( .D(N945), .SIN(mem_9__2_), .SMC(test_se), .C(
        net10424), .Q(mem_9__3_) );
  SDFFQX1 mem_reg_8__3_ ( .D(N954), .SIN(mem_8__2_), .SMC(test_se), .C(
        net10419), .Q(mem_8__3_) );
  SDFFQX1 mem_reg_27__2_ ( .D(N782), .SIN(mem_27__1_), .SMC(test_se), .C(
        net10514), .Q(mem_27__2_) );
  SDFFQX1 mem_reg_26__2_ ( .D(N791), .SIN(mem_26__1_), .SMC(test_se), .C(
        net10509), .Q(mem_26__2_) );
  SDFFQX1 mem_reg_25__2_ ( .D(N800), .SIN(mem_25__1_), .SMC(test_se), .C(
        net10504), .Q(mem_25__2_) );
  SDFFQX1 mem_reg_24__2_ ( .D(N809), .SIN(mem_24__1_), .SMC(test_se), .C(
        net10499), .Q(mem_24__2_) );
  SDFFQX1 mem_reg_23__2_ ( .D(N818), .SIN(mem_23__1_), .SMC(test_se), .C(
        net10494), .Q(mem_23__2_) );
  SDFFQX1 mem_reg_22__2_ ( .D(N827), .SIN(mem_22__1_), .SMC(test_se), .C(
        net10489), .Q(mem_22__2_) );
  SDFFQX1 mem_reg_21__2_ ( .D(N836), .SIN(mem_21__1_), .SMC(test_se), .C(
        net10484), .Q(mem_21__2_) );
  SDFFQX1 mem_reg_20__2_ ( .D(N845), .SIN(mem_20__1_), .SMC(test_se), .C(
        net10479), .Q(mem_20__2_) );
  SDFFQX1 mem_reg_19__2_ ( .D(N854), .SIN(mem_19__1_), .SMC(test_se), .C(
        net10474), .Q(mem_19__2_) );
  SDFFQX1 mem_reg_18__2_ ( .D(N863), .SIN(mem_18__1_), .SMC(test_se), .C(
        net10469), .Q(mem_18__2_) );
  SDFFQX1 mem_reg_17__2_ ( .D(N872), .SIN(mem_17__1_), .SMC(test_se), .C(
        net10464), .Q(mem_17__2_) );
  SDFFQX1 mem_reg_16__2_ ( .D(N881), .SIN(mem_16__1_), .SMC(test_se), .C(
        net10459), .Q(mem_16__2_) );
  SDFFQX1 mem_reg_15__2_ ( .D(N890), .SIN(mem_15__1_), .SMC(test_se), .C(
        net10454), .Q(mem_15__2_) );
  SDFFQX1 mem_reg_14__2_ ( .D(N899), .SIN(mem_14__1_), .SMC(test_se), .C(
        net10449), .Q(mem_14__2_) );
  SDFFQX1 mem_reg_13__2_ ( .D(N908), .SIN(mem_13__1_), .SMC(test_se), .C(
        net10444), .Q(mem_13__2_) );
  SDFFQX1 mem_reg_12__2_ ( .D(N917), .SIN(mem_12__1_), .SMC(test_se), .C(
        net10439), .Q(mem_12__2_) );
  SDFFQX1 mem_reg_11__2_ ( .D(N926), .SIN(mem_11__1_), .SMC(test_se), .C(
        net10434), .Q(mem_11__2_) );
  SDFFQX1 mem_reg_10__2_ ( .D(N935), .SIN(mem_10__1_), .SMC(test_se), .C(
        net10429), .Q(mem_10__2_) );
  SDFFQX1 mem_reg_9__2_ ( .D(N944), .SIN(mem_9__1_), .SMC(test_se), .C(
        net10424), .Q(mem_9__2_) );
  SDFFQX1 mem_reg_8__2_ ( .D(N953), .SIN(mem_8__1_), .SMC(test_se), .C(
        net10419), .Q(mem_8__2_) );
  SDFFQX1 mem_reg_27__1_ ( .D(N781), .SIN(mem_27__0_), .SMC(test_se), .C(
        net10514), .Q(mem_27__1_) );
  SDFFQX1 mem_reg_26__1_ ( .D(N790), .SIN(mem_26__0_), .SMC(test_se), .C(
        net10509), .Q(mem_26__1_) );
  SDFFQX1 mem_reg_25__1_ ( .D(N799), .SIN(mem_25__0_), .SMC(test_se), .C(
        net10504), .Q(mem_25__1_) );
  SDFFQX1 mem_reg_24__1_ ( .D(N808), .SIN(mem_24__0_), .SMC(test_se), .C(
        net10499), .Q(mem_24__1_) );
  SDFFQX1 mem_reg_23__1_ ( .D(N817), .SIN(mem_23__0_), .SMC(test_se), .C(
        net10494), .Q(mem_23__1_) );
  SDFFQX1 mem_reg_22__1_ ( .D(N826), .SIN(mem_22__0_), .SMC(test_se), .C(
        net10489), .Q(mem_22__1_) );
  SDFFQX1 mem_reg_21__1_ ( .D(N835), .SIN(mem_21__0_), .SMC(test_se), .C(
        net10484), .Q(mem_21__1_) );
  SDFFQX1 mem_reg_20__1_ ( .D(N844), .SIN(mem_20__0_), .SMC(test_se), .C(
        net10479), .Q(mem_20__1_) );
  SDFFQX1 mem_reg_19__1_ ( .D(N853), .SIN(mem_19__0_), .SMC(test_se), .C(
        net10474), .Q(mem_19__1_) );
  SDFFQX1 mem_reg_18__1_ ( .D(N862), .SIN(mem_18__0_), .SMC(test_se), .C(
        net10469), .Q(mem_18__1_) );
  SDFFQX1 mem_reg_17__1_ ( .D(N871), .SIN(mem_17__0_), .SMC(test_se), .C(
        net10464), .Q(mem_17__1_) );
  SDFFQX1 mem_reg_16__1_ ( .D(N880), .SIN(mem_16__0_), .SMC(test_se), .C(
        net10459), .Q(mem_16__1_) );
  SDFFQX1 mem_reg_15__1_ ( .D(N889), .SIN(mem_15__0_), .SMC(test_se), .C(
        net10454), .Q(mem_15__1_) );
  SDFFQX1 mem_reg_14__1_ ( .D(N898), .SIN(mem_14__0_), .SMC(test_se), .C(
        net10449), .Q(mem_14__1_) );
  SDFFQX1 mem_reg_13__1_ ( .D(N907), .SIN(mem_13__0_), .SMC(test_se), .C(
        net10444), .Q(mem_13__1_) );
  SDFFQX1 mem_reg_12__1_ ( .D(N916), .SIN(mem_12__0_), .SMC(test_se), .C(
        net10439), .Q(mem_12__1_) );
  SDFFQX1 mem_reg_11__1_ ( .D(N925), .SIN(mem_11__0_), .SMC(test_se), .C(
        net10434), .Q(mem_11__1_) );
  SDFFQX1 mem_reg_10__1_ ( .D(N934), .SIN(mem_10__0_), .SMC(test_se), .C(
        net10429), .Q(mem_10__1_) );
  SDFFQX1 mem_reg_9__1_ ( .D(N943), .SIN(mem_9__0_), .SMC(test_se), .C(
        net10424), .Q(mem_9__1_) );
  SDFFQX1 mem_reg_8__1_ ( .D(N952), .SIN(mem_8__0_), .SMC(test_se), .C(
        net10419), .Q(mem_8__1_) );
  SDFFQX1 mem_reg_27__0_ ( .D(N780), .SIN(mem_26__7_), .SMC(test_se), .C(
        net10514), .Q(mem_27__0_) );
  SDFFQX1 mem_reg_26__0_ ( .D(N789), .SIN(mem_25__7_), .SMC(test_se), .C(
        net10509), .Q(mem_26__0_) );
  SDFFQX1 mem_reg_25__0_ ( .D(N798), .SIN(mem_24__7_), .SMC(test_se), .C(
        net10504), .Q(mem_25__0_) );
  SDFFQX1 mem_reg_24__0_ ( .D(N807), .SIN(mem_23__7_), .SMC(test_se), .C(
        net10499), .Q(mem_24__0_) );
  SDFFQX1 mem_reg_23__0_ ( .D(N816), .SIN(mem_22__7_), .SMC(test_se), .C(
        net10494), .Q(mem_23__0_) );
  SDFFQX1 mem_reg_22__0_ ( .D(N825), .SIN(mem_21__7_), .SMC(test_se), .C(
        net10489), .Q(mem_22__0_) );
  SDFFQX1 mem_reg_21__0_ ( .D(N834), .SIN(mem_20__7_), .SMC(test_se), .C(
        net10484), .Q(mem_21__0_) );
  SDFFQX1 mem_reg_20__0_ ( .D(N843), .SIN(mem_19__7_), .SMC(test_se), .C(
        net10479), .Q(mem_20__0_) );
  SDFFQX1 mem_reg_19__0_ ( .D(N852), .SIN(mem_18__7_), .SMC(test_se), .C(
        net10474), .Q(mem_19__0_) );
  SDFFQX1 mem_reg_18__0_ ( .D(N861), .SIN(mem_17__7_), .SMC(test_se), .C(
        net10469), .Q(mem_18__0_) );
  SDFFQX1 mem_reg_17__0_ ( .D(N870), .SIN(mem_16__7_), .SMC(test_se), .C(
        net10464), .Q(mem_17__0_) );
  SDFFQX1 mem_reg_16__0_ ( .D(N879), .SIN(mem_15__7_), .SMC(test_se), .C(
        net10459), .Q(mem_16__0_) );
  SDFFQX1 mem_reg_15__0_ ( .D(N888), .SIN(mem_14__7_), .SMC(test_se), .C(
        net10454), .Q(mem_15__0_) );
  SDFFQX1 mem_reg_14__0_ ( .D(N897), .SIN(mem_13__7_), .SMC(test_se), .C(
        net10449), .Q(mem_14__0_) );
  SDFFQX1 mem_reg_13__0_ ( .D(N906), .SIN(mem_12__7_), .SMC(test_se), .C(
        net10444), .Q(mem_13__0_) );
  SDFFQX1 mem_reg_12__0_ ( .D(N915), .SIN(mem_11__7_), .SMC(test_se), .C(
        net10439), .Q(mem_12__0_) );
  SDFFQX1 mem_reg_11__0_ ( .D(N924), .SIN(mem_10__7_), .SMC(test_se), .C(
        net10434), .Q(mem_11__0_) );
  SDFFQX1 mem_reg_10__0_ ( .D(N933), .SIN(mem_9__7_), .SMC(test_se), .C(
        net10429), .Q(mem_10__0_) );
  SDFFQX1 mem_reg_9__0_ ( .D(N942), .SIN(mem_8__7_), .SMC(test_se), .C(
        net10424), .Q(mem_9__0_) );
  SDFFQX1 mem_reg_8__0_ ( .D(N951), .SIN(dat_7_1[55]), .SMC(test_se), .C(
        net10419), .Q(mem_8__0_) );
  SDFFQX1 mem_reg_1__3_ ( .D(N1017), .SIN(dat_7_1[2]), .SMC(test_se), .C(
        net10384), .Q(dat_7_1[3]) );
  SDFFQX1 mem_reg_1__2_ ( .D(N1016), .SIN(dat_7_1[1]), .SMC(test_se), .C(
        net10384), .Q(dat_7_1[2]) );
  SDFFQX1 mem_reg_1__1_ ( .D(N1015), .SIN(dat_7_1[0]), .SMC(test_se), .C(
        net10384), .Q(dat_7_1[1]) );
  SDFFQX1 mem_reg_1__0_ ( .D(N1014), .SIN(rdat0[7]), .SMC(test_se), .C(
        net10384), .Q(dat_7_1[0]) );
  SDFFQX1 locked_reg ( .D(ps_locked), .SIN(test_si), .SMC(test_se), .C(clk), 
        .Q(locked) );
  SDFFQX1 mem_reg_7__6_ ( .D(N966), .SIN(dat_7_1[53]), .SMC(test_se), .C(
        net10414), .Q(dat_7_1[54]) );
  SDFFQX1 mem_reg_7__0_ ( .D(N960), .SIN(dat_7_1[47]), .SMC(test_se), .C(
        net10414), .Q(dat_7_1[48]) );
  SDFFQX1 mem_reg_7__7_ ( .D(N967), .SIN(dat_7_1[54]), .SMC(test_se), .C(
        net10414), .Q(dat_7_1[55]) );
  SDFFQX1 mem_reg_6__7_ ( .D(N976), .SIN(dat_7_1[46]), .SMC(test_se), .C(
        net10409), .Q(dat_7_1[47]) );
  SDFFQX1 mem_reg_6__6_ ( .D(N975), .SIN(dat_7_1[45]), .SMC(test_se), .C(
        net10409), .Q(dat_7_1[46]) );
  SDFFQX1 mem_reg_7__5_ ( .D(N965), .SIN(dat_7_1[52]), .SMC(test_se), .C(
        net10414), .Q(dat_7_1[53]) );
  SDFFQX1 mem_reg_6__5_ ( .D(N974), .SIN(dat_7_1[44]), .SMC(test_se), .C(
        net10409), .Q(dat_7_1[45]) );
  SDFFQX1 mem_reg_6__4_ ( .D(N973), .SIN(dat_7_1[43]), .SMC(test_se), .C(
        net10409), .Q(dat_7_1[44]) );
  SDFFQX1 mem_reg_7__3_ ( .D(N963), .SIN(dat_7_1[50]), .SMC(test_se), .C(
        net10414), .Q(dat_7_1[51]) );
  SDFFQX1 mem_reg_6__3_ ( .D(N972), .SIN(dat_7_1[42]), .SMC(test_se), .C(
        net10409), .Q(dat_7_1[43]) );
  SDFFQX1 mem_reg_6__2_ ( .D(N971), .SIN(dat_7_1[41]), .SMC(test_se), .C(
        net10409), .Q(dat_7_1[42]) );
  SDFFQX1 mem_reg_7__1_ ( .D(N961), .SIN(dat_7_1[48]), .SMC(test_se), .C(
        net10414), .Q(dat_7_1[49]) );
  SDFFQX1 mem_reg_6__0_ ( .D(N969), .SIN(dat_7_1[39]), .SMC(test_se), .C(
        net10409), .Q(dat_7_1[40]) );
  SDFFQX1 mem_reg_7__4_ ( .D(N964), .SIN(dat_7_1[51]), .SMC(test_se), .C(
        net10414), .Q(dat_7_1[52]) );
  SDFFQX1 mem_reg_7__2_ ( .D(N962), .SIN(dat_7_1[49]), .SMC(test_se), .C(
        net10414), .Q(dat_7_1[50]) );
  SDFFQX1 mem_reg_6__1_ ( .D(N970), .SIN(dat_7_1[40]), .SMC(test_se), .C(
        net10409), .Q(dat_7_1[41]) );
  SDFFQX1 mem_reg_5__7_ ( .D(N985), .SIN(dat_7_1[38]), .SMC(test_se), .C(
        net10404), .Q(dat_7_1[39]) );
  SDFFQX1 mem_reg_4__7_ ( .D(N994), .SIN(dat_7_1[30]), .SMC(test_se), .C(
        net10399), .Q(dat_7_1[31]) );
  SDFFQX1 mem_reg_4__6_ ( .D(N993), .SIN(dat_7_1[29]), .SMC(test_se), .C(
        net10399), .Q(dat_7_1[30]) );
  SDFFQX1 mem_reg_5__5_ ( .D(N983), .SIN(dat_7_1[36]), .SMC(test_se), .C(
        net10404), .Q(dat_7_1[37]) );
  SDFFQX1 mem_reg_4__5_ ( .D(N992), .SIN(dat_7_1[28]), .SMC(test_se), .C(
        net10399), .Q(dat_7_1[29]) );
  SDFFQX1 mem_reg_4__4_ ( .D(N991), .SIN(dat_7_1[27]), .SMC(test_se), .C(
        net10399), .Q(dat_7_1[28]) );
  SDFFQX1 mem_reg_4__3_ ( .D(N990), .SIN(dat_7_1[26]), .SMC(test_se), .C(
        net10399), .Q(dat_7_1[27]) );
  SDFFQX1 mem_reg_4__2_ ( .D(N989), .SIN(dat_7_1[25]), .SMC(test_se), .C(
        net10399), .Q(dat_7_1[26]) );
  SDFFQX1 mem_reg_5__1_ ( .D(N979), .SIN(dat_7_1[32]), .SMC(test_se), .C(
        net10404), .Q(dat_7_1[33]) );
  SDFFQX1 mem_reg_5__0_ ( .D(N978), .SIN(dat_7_1[31]), .SMC(test_se), .C(
        net10404), .Q(dat_7_1[32]) );
  SDFFQX1 mem_reg_4__0_ ( .D(N987), .SIN(dat_7_1[23]), .SMC(test_se), .C(
        net10399), .Q(dat_7_1[24]) );
  SDFFQX1 mem_reg_3__3_ ( .D(N999), .SIN(dat_7_1[18]), .SMC(test_se), .C(
        net10394), .Q(dat_7_1[19]) );
  SDFFQX1 mem_reg_3__2_ ( .D(N998), .SIN(dat_7_1[17]), .SMC(test_se), .C(
        net10394), .Q(dat_7_1[18]) );
  SDFFQX1 mem_reg_3__1_ ( .D(N997), .SIN(dat_7_1[16]), .SMC(test_se), .C(
        net10394), .Q(dat_7_1[17]) );
  SDFFQX1 mem_reg_3__0_ ( .D(N996), .SIN(dat_7_1[15]), .SMC(test_se), .C(
        net10394), .Q(dat_7_1[16]) );
  SDFFQX1 mem_reg_2__7_ ( .D(N1012), .SIN(dat_7_1[14]), .SMC(test_se), .C(
        net10389), .Q(dat_7_1[15]) );
  SDFFQX1 mem_reg_2__6_ ( .D(N1011), .SIN(dat_7_1[13]), .SMC(test_se), .C(
        net10389), .Q(dat_7_1[14]) );
  SDFFQX1 mem_reg_2__5_ ( .D(N1010), .SIN(dat_7_1[12]), .SMC(test_se), .C(
        net10389), .Q(dat_7_1[13]) );
  SDFFQX1 mem_reg_5__6_ ( .D(N984), .SIN(dat_7_1[37]), .SMC(test_se), .C(
        net10404), .Q(dat_7_1[38]) );
  SDFFQX1 mem_reg_5__4_ ( .D(N982), .SIN(dat_7_1[35]), .SMC(test_se), .C(
        net10404), .Q(dat_7_1[36]) );
  SDFFQX1 mem_reg_5__3_ ( .D(N981), .SIN(dat_7_1[34]), .SMC(test_se), .C(
        net10404), .Q(dat_7_1[35]) );
  SDFFQX1 mem_reg_5__2_ ( .D(N980), .SIN(dat_7_1[33]), .SMC(test_se), .C(
        net10404), .Q(dat_7_1[34]) );
  SDFFQX1 mem_reg_4__1_ ( .D(N988), .SIN(dat_7_1[24]), .SMC(test_se), .C(
        net10399), .Q(dat_7_1[25]) );
  SDFFQX1 mem_reg_1__7_ ( .D(N1021), .SIN(dat_7_1[6]), .SMC(test_se), .C(
        net10384), .Q(dat_7_1[7]) );
  SDFFQX1 mem_reg_1__6_ ( .D(N1020), .SIN(dat_7_1[5]), .SMC(test_se), .C(
        net10384), .Q(dat_7_1[6]) );
  SDFFQX1 mem_reg_1__5_ ( .D(N1019), .SIN(dat_7_1[4]), .SMC(test_se), .C(
        net10384), .Q(dat_7_1[5]) );
  SDFFQX1 mem_reg_1__4_ ( .D(N1018), .SIN(dat_7_1[3]), .SMC(test_se), .C(
        net10384), .Q(dat_7_1[4]) );
  SDFFQX1 mem_reg_3__6_ ( .D(N1002), .SIN(dat_7_1[21]), .SMC(test_se), .C(
        net10394), .Q(dat_7_1[22]) );
  SDFFQX1 mem_reg_3__5_ ( .D(N1001), .SIN(dat_7_1[20]), .SMC(test_se), .C(
        net10394), .Q(dat_7_1[21]) );
  SDFFQX1 mem_reg_3__4_ ( .D(N1000), .SIN(dat_7_1[19]), .SMC(test_se), .C(
        net10394), .Q(dat_7_1[20]) );
  SDFFQX1 mem_reg_2__4_ ( .D(N1009), .SIN(dat_7_1[11]), .SMC(test_se), .C(
        net10389), .Q(dat_7_1[12]) );
  SDFFQX1 mem_reg_2__3_ ( .D(N1008), .SIN(dat_7_1[10]), .SMC(test_se), .C(
        net10389), .Q(dat_7_1[11]) );
  SDFFQX1 mem_reg_3__7_ ( .D(N1003), .SIN(dat_7_1[22]), .SMC(test_se), .C(
        net10394), .Q(dat_7_1[23]) );
  SDFFQX1 mem_reg_2__1_ ( .D(N1006), .SIN(dat_7_1[8]), .SMC(test_se), .C(
        net10389), .Q(dat_7_1[9]) );
  SDFFQX1 mem_reg_2__0_ ( .D(N1005), .SIN(dat_7_1[7]), .SMC(test_se), .C(
        net10389), .Q(dat_7_1[8]) );
  SDFFQX1 mem_reg_2__2_ ( .D(N1007), .SIN(dat_7_1[9]), .SMC(test_se), .C(
        net10389), .Q(dat_7_1[10]) );
  SDFFQX1 mem_reg_0__2_ ( .D(N1025), .SIN(rdat0[1]), .SMC(test_se), .C(
        net10378), .Q(rdat0[2]) );
  SDFFQX1 mem_reg_0__4_ ( .D(N1027), .SIN(rdat0[3]), .SMC(test_se), .C(
        net10378), .Q(rdat0[4]) );
  SDFFQX1 mem_reg_0__3_ ( .D(N1026), .SIN(rdat0[2]), .SMC(test_se), .C(
        net10378), .Q(rdat0[3]) );
  SDFFQX1 mem_reg_0__5_ ( .D(N1028), .SIN(rdat0[4]), .SMC(test_se), .C(
        net10378), .Q(rdat0[5]) );
  SDFFQX1 mem_reg_0__1_ ( .D(N1024), .SIN(rdat0[0]), .SMC(test_se), .C(
        net10378), .Q(rdat0[1]) );
  SDFFQX1 mem_reg_0__7_ ( .D(N1030), .SIN(rdat0[6]), .SMC(test_se), .C(
        net10378), .Q(rdat0[7]) );
  SDFFQX1 mem_reg_0__6_ ( .D(N1029), .SIN(rdat0[5]), .SMC(test_se), .C(
        net10378), .Q(rdat0[6]) );
  SDFFQX1 mem_reg_0__0_ ( .D(N1023), .SIN(locked), .SMC(test_se), .C(net10378), 
        .Q(rdat0[0]) );
  SDFFQX1 pshptr_reg_0_ ( .D(N1054), .SIN(mem_33__7_), .SMC(test_se), .C(
        net10549), .Q(ptr[0]) );
  SDFFQX1 pshptr_reg_4_ ( .D(N1058), .SIN(ptr[3]), .SMC(test_se), .C(net10549), 
        .Q(ptr[4]) );
  SDFFQX1 pshptr_reg_3_ ( .D(N1057), .SIN(ptr[2]), .SMC(test_se), .C(net10549), 
        .Q(ptr[3]) );
  SDFFQX1 pshptr_reg_2_ ( .D(N1056), .SIN(ptr[1]), .SMC(test_se), .C(net10549), 
        .Q(ptr[2]) );
  SDFFQX1 pshptr_reg_1_ ( .D(N1055), .SIN(ptr[0]), .SMC(test_se), .C(net10549), 
        .Q(ptr[1]) );
  SDFFQX1 pshptr_reg_5_ ( .D(N1059), .SIN(ptr[4]), .SMC(test_se), .C(net10549), 
        .Q(ptr[5]) );
  NAND2X1 U3 ( .A(n526), .B(n542), .Y(n1) );
  NAND2X1 U4 ( .A(n539), .B(n526), .Y(n2) );
  BUFX3 U5 ( .A(n125), .Y(n3) );
  INVX1 U6 ( .A(n528), .Y(n4) );
  BUFX3 U7 ( .A(n219), .Y(n5) );
  NOR3XL U8 ( .A(ptr[3]), .B(ptr[2]), .C(ptr[1]), .Y(n6) );
  INVXL U9 ( .A(n517), .Y(n514) );
  OAI21BBXL U10 ( .A(n6), .B(n515), .C(ptr[5]), .Y(n522) );
  NAND32XL U11 ( .B(ptr[4]), .C(n517), .A(n516), .Y(n519) );
  NAND2XL U12 ( .A(ptr[2]), .B(n442), .Y(n173) );
  NAND2XL U13 ( .A(ptr[5]), .B(n442), .Y(n346) );
  NAND2XL U14 ( .A(ptr[1]), .B(n442), .Y(n380) );
  NAND2XL U15 ( .A(ptr[3]), .B(n442), .Y(n208) );
  NAND2XL U16 ( .A(ptr[0]), .B(n442), .Y(n381) );
  AOI21XL U17 ( .B(one), .C(r_pop), .A(n547), .Y(n7) );
  INVX1 U18 ( .A(n507), .Y(n505) );
  INVX1 U19 ( .A(n507), .Y(n506) );
  INVX1 U20 ( .A(n507), .Y(n504) );
  INVX1 U21 ( .A(n51), .Y(n507) );
  INVX1 U22 ( .A(n20), .Y(n19) );
  INVX1 U23 ( .A(n20), .Y(n18) );
  INVX1 U24 ( .A(n28), .Y(n27) );
  INVX1 U25 ( .A(n28), .Y(n26) );
  INVX1 U26 ( .A(n36), .Y(n35) );
  INVX1 U27 ( .A(n36), .Y(n34) );
  INVX1 U28 ( .A(n46), .Y(n43) );
  INVX1 U29 ( .A(n46), .Y(n42) );
  NOR21XL U30 ( .B(n49), .A(n11), .Y(n53) );
  NOR21XL U31 ( .B(n163), .A(n8), .Y(n165) );
  NOR21XL U32 ( .B(n347), .A(n10), .Y(n349) );
  INVX1 U33 ( .A(n28), .Y(n25) );
  INVX1 U34 ( .A(n76), .Y(n28) );
  INVX1 U35 ( .A(n36), .Y(n33) );
  INVX1 U36 ( .A(n73), .Y(n36) );
  INVX1 U37 ( .A(n46), .Y(n41) );
  INVX1 U38 ( .A(n69), .Y(n46) );
  INVX1 U39 ( .A(n483), .Y(n480) );
  INVX1 U40 ( .A(n491), .Y(n489) );
  INVX1 U41 ( .A(n499), .Y(n497) );
  INVX1 U42 ( .A(n483), .Y(n482) );
  INVX1 U43 ( .A(n491), .Y(n490) );
  INVX1 U44 ( .A(n499), .Y(n498) );
  INVX1 U45 ( .A(n20), .Y(n17) );
  INVX1 U46 ( .A(n79), .Y(n20) );
  NAND2X1 U47 ( .A(fifowdat[3]), .B(n11), .Y(n51) );
  INVX1 U48 ( .A(n423), .Y(n534) );
  INVX1 U49 ( .A(r_psh), .Y(n546) );
  NOR21XL U50 ( .B(n102), .A(n8), .Y(n104) );
  AND2X1 U51 ( .A(n112), .B(n64), .Y(n102) );
  INVX1 U52 ( .A(fifowdat[3]), .Y(n510) );
  INVX1 U53 ( .A(fifowdat[3]), .Y(n509) );
  INVX1 U54 ( .A(fifowdat[3]), .Y(n508) );
  NOR21XL U55 ( .B(srstz), .A(r_fiforst), .Y(n442) );
  NOR21XL U56 ( .B(n443), .A(n10), .Y(n445) );
  NOR21XL U57 ( .B(n465), .A(n10), .Y(n467) );
  NOR21XL U58 ( .B(n66), .A(n8), .Y(n70) );
  NOR21XL U59 ( .B(n89), .A(n8), .Y(n91) );
  NOR21XL U60 ( .B(n115), .A(n8), .Y(n117) );
  NOR21XL U61 ( .B(n455), .A(n11), .Y(n457) );
  NOR21XL U62 ( .B(n127), .A(n8), .Y(n129) );
  NOR21XL U63 ( .B(n140), .A(n8), .Y(n142) );
  NOR21XL U64 ( .B(n152), .A(n8), .Y(n154) );
  NOR21XL U65 ( .B(n174), .A(n8), .Y(n176) );
  NOR21XL U66 ( .B(n186), .A(n8), .Y(n188) );
  NOR21XL U67 ( .B(n209), .A(n9), .Y(n211) );
  NOR21XL U68 ( .B(n221), .A(n9), .Y(n223) );
  NOR21XL U69 ( .B(n232), .A(n9), .Y(n234) );
  NOR21XL U70 ( .B(n244), .A(n9), .Y(n246) );
  NOR21XL U71 ( .B(n255), .A(n9), .Y(n257) );
  NOR21XL U72 ( .B(n266), .A(n9), .Y(n268) );
  NOR21XL U73 ( .B(n278), .A(n9), .Y(n280) );
  NOR21XL U74 ( .B(n300), .A(n9), .Y(n302) );
  NOR21XL U75 ( .B(n311), .A(n9), .Y(n313) );
  NOR21XL U76 ( .B(n322), .A(n10), .Y(n324) );
  NOR21XL U77 ( .B(n334), .A(n10), .Y(n336) );
  NOR21XL U78 ( .B(n358), .A(n10), .Y(n360) );
  NOR21XL U79 ( .B(n370), .A(n10), .Y(n372) );
  AOI21BBXL U80 ( .B(n86), .C(n64), .A(n63), .Y(n49) );
  AOI21BBXL U81 ( .B(n86), .C(n310), .A(n357), .Y(n347) );
  AOI21BBXL U82 ( .B(n86), .C(n125), .A(n530), .Y(n163) );
  INVX1 U83 ( .A(n16), .Y(n11) );
  NOR2X1 U84 ( .A(n441), .B(n538), .Y(n423) );
  NAND2X1 U85 ( .A(n539), .B(n526), .Y(n310) );
  NAND2X1 U86 ( .A(n526), .B(n542), .Y(n64) );
  INVX1 U87 ( .A(n422), .Y(n535) );
  INVX1 U88 ( .A(n16), .Y(n12) );
  INVX1 U89 ( .A(n491), .Y(n488) );
  INVX1 U90 ( .A(n58), .Y(n491) );
  INVX1 U91 ( .A(n499), .Y(n496) );
  INVX1 U92 ( .A(n55), .Y(n499) );
  INVX1 U93 ( .A(n483), .Y(n439) );
  INVX1 U94 ( .A(n61), .Y(n483) );
  NAND2X1 U95 ( .A(fifowdat[4]), .B(n12), .Y(n79) );
  NAND2X1 U96 ( .A(fifowdat[5]), .B(n11), .Y(n76) );
  NAND2X1 U97 ( .A(fifowdat[6]), .B(n11), .Y(n73) );
  NAND2X1 U98 ( .A(fifowdat[7]), .B(n11), .Y(n69) );
  NAND2X1 U99 ( .A(n546), .B(n548), .Y(n47) );
  NOR21XL U100 ( .B(n197), .A(n9), .Y(n199) );
  NOR21XL U101 ( .B(n289), .A(n10), .Y(n291) );
  NOR21XL U102 ( .B(n382), .A(n10), .Y(n384) );
  NOR21XL U103 ( .B(n404), .A(n11), .Y(n406) );
  INVX1 U104 ( .A(n15), .Y(n8) );
  INVX1 U105 ( .A(n15), .Y(n9) );
  INVX1 U106 ( .A(n15), .Y(n10) );
  AND2X1 U107 ( .A(n63), .B(n434), .Y(n475) );
  INVX1 U108 ( .A(n15), .Y(n13) );
  INVX1 U109 ( .A(n16), .Y(n14) );
  OAI22X1 U110 ( .A(n543), .B(n14), .C(n3), .D(n114), .Y(N887) );
  OAI22X1 U111 ( .A(n542), .B(n14), .C(n64), .D(n114), .Y(N959) );
  OAI22X1 U112 ( .A(n86), .B(n310), .C(n368), .D(n13), .Y(N770) );
  OAI22X1 U113 ( .A(n86), .B(n125), .C(n184), .D(n13), .Y(N914) );
  OAI22X1 U114 ( .A(n86), .B(n1), .C(n85), .D(n14), .Y(N986) );
  NAND2X1 U115 ( .A(n542), .B(n114), .Y(n112) );
  INVX1 U116 ( .A(n434), .Y(n531) );
  INVX1 U117 ( .A(n345), .Y(n539) );
  NAND2X1 U118 ( .A(n441), .B(n442), .Y(N1053) );
  INVX1 U119 ( .A(fifowdat[4]), .Y(n23) );
  INVX1 U120 ( .A(fifowdat[4]), .Y(n22) );
  INVX1 U121 ( .A(fifowdat[5]), .Y(n31) );
  INVX1 U122 ( .A(fifowdat[5]), .Y(n30) );
  INVX1 U123 ( .A(fifowdat[6]), .Y(n39) );
  INVX1 U124 ( .A(fifowdat[6]), .Y(n38) );
  INVX1 U125 ( .A(fifowdat[7]), .Y(n220) );
  INVX1 U126 ( .A(fifowdat[7]), .Y(n113) );
  INVX1 U127 ( .A(fifowdat[4]), .Y(n21) );
  INVX1 U128 ( .A(fifowdat[5]), .Y(n29) );
  INVX1 U129 ( .A(fifowdat[6]), .Y(n37) );
  INVX1 U130 ( .A(fifowdat[7]), .Y(n48) );
  INVX1 U131 ( .A(n50), .Y(fifowdat[3]) );
  AOI21BBXL U132 ( .B(n1), .C(n65), .A(n475), .Y(n465) );
  AOI21BBXL U133 ( .B(n64), .C(n84), .A(n85), .Y(n66) );
  AOI21BBXL U134 ( .B(n1), .C(n99), .A(n87), .Y(n89) );
  AOI21BBXL U135 ( .B(n125), .C(n126), .A(n542), .Y(n115) );
  AOI21BBXL U136 ( .B(n64), .C(n150), .A(n527), .Y(n455) );
  AOI21BBXL U137 ( .B(n125), .C(n150), .A(n139), .Y(n140) );
  AOI21BBXL U138 ( .B(n126), .C(n2), .A(n540), .Y(n300) );
  AOI21BBXL U139 ( .B(n137), .C(n310), .A(n321), .Y(n311) );
  AOI21BBXL U140 ( .B(n150), .C(n2), .A(n332), .Y(n322) );
  AOI21BBXL U141 ( .B(n65), .C(n310), .A(n344), .Y(n334) );
  AOI21BBXL U142 ( .B(n84), .C(n2), .A(n368), .Y(n358) );
  AOI21BBXL U143 ( .B(n99), .C(n310), .A(n369), .Y(n370) );
  AOI21BBXL U144 ( .B(n1), .C(n137), .A(n453), .Y(n443) );
  AOI21BBXL U145 ( .B(n125), .C(n137), .A(n138), .Y(n127) );
  AOI21BBXL U146 ( .B(n65), .C(n125), .A(n162), .Y(n152) );
  AOI21BBXL U147 ( .B(n84), .C(n125), .A(n184), .Y(n174) );
  AOI21BBXL U148 ( .B(n99), .C(n125), .A(n185), .Y(n186) );
  AOI21BBXL U149 ( .B(n126), .C(n219), .A(n543), .Y(n209) );
  AOI21BBXL U150 ( .B(n137), .C(n219), .A(n231), .Y(n221) );
  AOI21BBXL U151 ( .B(n150), .C(n219), .A(n242), .Y(n232) );
  AOI21BBXL U152 ( .B(n65), .C(n219), .A(n254), .Y(n244) );
  AOI21BBXL U153 ( .B(n86), .C(n219), .A(n529), .Y(n255) );
  AOI21BBXL U154 ( .B(n84), .C(n219), .A(n276), .Y(n266) );
  AOI21BBXL U155 ( .B(n99), .C(n219), .A(n277), .Y(n278) );
  XNOR2XL U156 ( .A(n536), .B(n538), .Y(n441) );
  NOR2X1 U157 ( .A(n440), .B(n441), .Y(n422) );
  NAND3X1 U158 ( .A(n526), .B(n543), .C(n545), .Y(n125) );
  INVX1 U159 ( .A(n520), .Y(n526) );
  INVX1 U160 ( .A(n440), .Y(n538) );
  INVX1 U161 ( .A(n537), .Y(n16) );
  NAND2X1 U162 ( .A(fifowdat[0]), .B(n11), .Y(n61) );
  NAND2X1 U163 ( .A(fifowdat[1]), .B(n11), .Y(n58) );
  NAND2X1 U164 ( .A(fifowdat[2]), .B(n11), .Y(n55) );
  INVX1 U165 ( .A(r_pop), .Y(n548) );
  NOR21XL U166 ( .B(n393), .A(n10), .Y(n395) );
  NOR21XL U167 ( .B(n87), .A(n88), .Y(n85) );
  AND2X1 U168 ( .A(n414), .B(n415), .Y(n404) );
  AND2X1 U169 ( .A(n207), .B(n125), .Y(n197) );
  AND2X1 U170 ( .A(n299), .B(n219), .Y(n289) );
  AND2X1 U171 ( .A(n392), .B(n2), .Y(n382) );
  OAI21X1 U172 ( .B(n101), .C(n196), .A(n100), .Y(n185) );
  OAI21X1 U173 ( .B(n101), .C(n544), .A(n288), .Y(n369) );
  MUX2X1 U174 ( .D0(n525), .D1(n524), .S(n532), .Y(N1054) );
  AND2X1 U175 ( .A(full), .B(n422), .Y(n524) );
  OAI22X1 U176 ( .A(n534), .B(empty), .C(n535), .D(full), .Y(n525) );
  NAND32X1 U177 ( .B(n520), .C(n346), .A(n512), .Y(n415) );
  INVX1 U178 ( .A(n137), .Y(n512) );
  AOI21X1 U179 ( .B(n533), .C(n545), .A(n151), .Y(n139) );
  AOI21X1 U180 ( .B(n101), .C(n541), .A(n288), .Y(n277) );
  AOI21X1 U181 ( .B(n531), .C(n545), .A(n151), .Y(n162) );
  AOI21X1 U182 ( .B(n533), .C(n541), .A(n243), .Y(n242) );
  AOI21X1 U183 ( .B(n531), .C(n541), .A(n243), .Y(n254) );
  AOI21AX1 U184 ( .B(n532), .C(n545), .A(n139), .Y(n138) );
  AOI21AX1 U185 ( .B(n88), .C(n541), .A(n277), .Y(n276) );
  AOI21AX1 U186 ( .B(n88), .C(n545), .A(n185), .Y(n184) );
  AOI21AX1 U187 ( .B(n88), .C(n539), .A(n369), .Y(n368) );
  NAND2X1 U188 ( .A(n541), .B(n545), .Y(n345) );
  NOR2X1 U189 ( .A(n100), .B(n528), .Y(n63) );
  NOR2X1 U190 ( .A(n532), .B(n533), .Y(n438) );
  NAND2X1 U191 ( .A(n532), .B(n533), .Y(n434) );
  NOR2X1 U192 ( .A(n100), .B(n101), .Y(n87) );
  INVX1 U193 ( .A(n196), .Y(n543) );
  INVX1 U194 ( .A(n100), .Y(n542) );
  NOR3XL U195 ( .A(n545), .B(n541), .C(n126), .Y(n416) );
  NOR2X1 U196 ( .A(n454), .B(n532), .Y(n453) );
  OAI22X1 U197 ( .A(n424), .B(n534), .C(n425), .D(n535), .Y(N1058) );
  XNOR2XL U198 ( .A(n420), .B(n541), .Y(n424) );
  XNOR2XL U199 ( .A(n421), .B(n541), .Y(n425) );
  INVX1 U200 ( .A(n151), .Y(n530) );
  INVX1 U201 ( .A(n243), .Y(n529) );
  INVX1 U202 ( .A(n288), .Y(n540) );
  INVX1 U203 ( .A(n537), .Y(n15) );
  NAND3X1 U204 ( .A(n416), .B(n526), .C(n544), .Y(n403) );
  INVX1 U205 ( .A(n454), .Y(n527) );
  OAI21X1 U206 ( .B(n544), .C(n126), .A(n288), .Y(n321) );
  OAI21X1 U207 ( .B(n544), .C(n528), .A(n288), .Y(n357) );
  OAI31XL U208 ( .A(n126), .B(n544), .C(n545), .D(n196), .Y(n231) );
  AOI21X1 U209 ( .B(n533), .C(n539), .A(n333), .Y(n332) );
  AOI21X1 U210 ( .B(n531), .C(n539), .A(n333), .Y(n344) );
  NAND2X1 U211 ( .A(n101), .B(n532), .Y(n114) );
  NAND2X1 U212 ( .A(n528), .B(n438), .Y(n86) );
  NOR2X1 U213 ( .A(n429), .B(n545), .Y(n420) );
  OAI22X1 U214 ( .A(n63), .B(n14), .C(n1), .D(n65), .Y(N995) );
  OAI22X1 U215 ( .A(n65), .B(n3), .C(n12), .D(n530), .Y(N923) );
  OAI22X1 U216 ( .A(n453), .B(n14), .C(n64), .D(n126), .Y(N1022) );
  OAI22X1 U217 ( .A(n137), .B(n2), .C(n332), .D(n13), .Y(N797) );
  OAI22X1 U218 ( .A(n84), .B(n5), .C(n277), .D(n13), .Y(N833) );
  OAI22X1 U219 ( .A(n86), .B(n5), .C(n276), .D(n13), .Y(N842) );
  OAI22X1 U220 ( .A(n65), .B(n5), .C(n529), .D(n13), .Y(N851) );
  OAI22X1 U221 ( .A(n150), .B(n5), .C(n254), .D(n13), .Y(N860) );
  OAI22X1 U222 ( .A(n137), .B(n5), .C(n242), .D(n13), .Y(N869) );
  OAI22X1 U223 ( .A(n3), .B(n150), .C(n162), .D(n13), .Y(N932) );
  OAI22X1 U224 ( .A(n3), .B(n137), .C(n139), .D(n13), .Y(N941) );
  OAI22X1 U225 ( .A(n3), .B(n126), .C(n138), .D(n14), .Y(N950) );
  OAI22X1 U226 ( .A(n1), .B(n84), .C(n87), .D(n14), .Y(N977) );
  OAI22X1 U227 ( .A(n150), .B(n310), .C(n344), .D(n12), .Y(N788) );
  OAI22X1 U228 ( .A(n12), .B(n369), .C(n84), .D(n2), .Y(N761) );
  OAI22X1 U229 ( .A(n65), .B(n2), .C(n12), .D(n357), .Y(N779) );
  OAI22X1 U230 ( .A(n126), .B(n310), .C(n12), .D(n321), .Y(N806) );
  OAI22X1 U231 ( .A(n475), .B(n14), .C(n1), .D(n150), .Y(N1004) );
  OAI22X1 U232 ( .A(n126), .B(n5), .C(n12), .D(n231), .Y(N878) );
  OAI22X1 U233 ( .A(n84), .B(n3), .C(n12), .D(n185), .Y(N905) );
  OAI22X1 U234 ( .A(n540), .B(n14), .C(n114), .D(n219), .Y(N815) );
  OAI22X1 U235 ( .A(n527), .B(n14), .C(n64), .D(n137), .Y(N1013) );
  INVX1 U236 ( .A(n521), .Y(n433) );
  NAND21X1 U237 ( .B(empty), .A(n438), .Y(n521) );
  ENOX1 U238 ( .A(n64), .B(n99), .C(n112), .D(n15), .Y(N968) );
  ENOX1 U239 ( .A(n99), .B(n2), .C(n392), .D(n15), .Y(N752) );
  ENOX1 U240 ( .A(n99), .B(n5), .C(n299), .D(n15), .Y(N824) );
  ENOX1 U241 ( .A(n99), .B(n3), .C(n207), .D(n15), .Y(N896) );
  OAI21BBX1 U242 ( .A(n15), .B(n414), .C(n403), .Y(N734) );
  INVX1 U243 ( .A(n77), .Y(fifowdat[4]) );
  INVX1 U244 ( .A(n74), .Y(fifowdat[5]) );
  OAI22X1 U245 ( .A(prx_wdat[3]), .B(n549), .C(r_wdat[3]), .D(prx_psh), .Y(n50) );
  INVX1 U246 ( .A(fifowdat[0]), .Y(n486) );
  INVX1 U247 ( .A(fifowdat[0]), .Y(n485) );
  INVX1 U248 ( .A(fifowdat[1]), .Y(n494) );
  INVX1 U249 ( .A(fifowdat[1]), .Y(n493) );
  INVX1 U250 ( .A(fifowdat[2]), .Y(n502) );
  INVX1 U251 ( .A(fifowdat[2]), .Y(n501) );
  INVX1 U252 ( .A(fifowdat[0]), .Y(n484) );
  INVX1 U253 ( .A(fifowdat[1]), .Y(n492) );
  INVX1 U254 ( .A(fifowdat[2]), .Y(n500) );
  INVX1 U255 ( .A(n67), .Y(fifowdat[7]) );
  INVX1 U256 ( .A(n71), .Y(fifowdat[6]) );
  INVX1 U257 ( .A(prx_psh), .Y(n549) );
  INVX1 U258 ( .A(ptx_pop), .Y(n550) );
  AND3X1 U259 ( .A(ptr[4]), .B(ptr[0]), .C(n514), .Y(half) );
  INVX1 U260 ( .A(n518), .Y(one) );
  NAND32X1 U261 ( .B(n517), .C(n516), .A(n515), .Y(n518) );
  INVX1 U262 ( .A(n522), .Y(full) );
  INVX1 U263 ( .A(n519), .Y(empty) );
  NOR3XL U264 ( .A(n551), .B(n44), .C(n45), .Y(txreq) );
  NAND21X1 U265 ( .B(n536), .A(n522), .Y(n520) );
  OAI21X1 U266 ( .B(n44), .C(n548), .A(n550), .Y(n440) );
  NAND21X1 U267 ( .B(n538), .A(n519), .Y(n537) );
  NAND3X1 U268 ( .A(n526), .B(n208), .C(n541), .Y(n219) );
  OAI21X1 U269 ( .B(n429), .C(n534), .A(n431), .Y(N1056) );
  AOI32X1 U270 ( .A(n430), .B(n4), .C(n422), .D(n528), .E(n432), .Y(n431) );
  OAI22X1 U271 ( .A(n433), .B(n534), .C(n430), .D(n535), .Y(n432) );
  OAI21BBX1 U272 ( .A(n420), .B(n423), .C(n427), .Y(N1057) );
  AOI32X1 U273 ( .A(n426), .B(n208), .C(n422), .D(n545), .E(n428), .Y(n427) );
  ENOX1 U274 ( .A(n426), .B(n535), .C(n429), .D(n423), .Y(n428) );
  INVX1 U275 ( .A(fifopsh), .Y(n536) );
  OAI21X1 U276 ( .B(n44), .C(n546), .A(n549), .Y(fifopsh) );
  NOR21XL U277 ( .B(n403), .A(n346), .Y(n393) );
  NOR21XL U278 ( .B(n430), .A(n4), .Y(n426) );
  OAI21X1 U279 ( .B(n173), .C(n265), .A(n540), .Y(n243) );
  AOI21X1 U280 ( .B(n173), .C(n543), .A(n542), .Y(n151) );
  INVX1 U281 ( .A(n381), .Y(n532) );
  NOR2X1 U282 ( .A(n380), .B(n173), .Y(n101) );
  NAND2X1 U283 ( .A(n543), .B(n208), .Y(n100) );
  NAND2X1 U284 ( .A(n346), .B(n345), .Y(n288) );
  NAND2X1 U285 ( .A(n265), .B(n346), .Y(n196) );
  NAND2X1 U286 ( .A(n63), .B(n380), .Y(n454) );
  NAND2X1 U287 ( .A(n438), .B(n173), .Y(n126) );
  INVX1 U288 ( .A(n208), .Y(n545) );
  INVX1 U289 ( .A(n265), .Y(n541) );
  INVX1 U290 ( .A(n380), .Y(n533) );
  INVX1 U291 ( .A(n523), .Y(n430) );
  NAND21X1 U292 ( .B(n434), .A(n522), .Y(n523) );
  NOR2X1 U293 ( .A(n346), .B(n416), .Y(n414) );
  NAND2X1 U294 ( .A(n418), .B(n419), .Y(N1059) );
  GEN2XL U295 ( .D(n420), .E(n265), .C(n534), .B(n535), .A(n346), .Y(n419) );
  AOI33X1 U296 ( .A(n421), .B(n541), .C(n422), .D(n420), .E(n543), .F(n423), 
        .Y(n418) );
  NAND3X1 U297 ( .A(n435), .B(n436), .C(n437), .Y(N1055) );
  OAI21X1 U298 ( .B(n433), .C(n531), .A(n423), .Y(n435) );
  OAI211X1 U299 ( .C(n381), .D(full), .A(n533), .B(n422), .Y(n437) );
  NAND43X1 U300 ( .B(full), .C(n381), .D(n535), .A(n380), .Y(n436) );
  NOR21XL U301 ( .B(n426), .A(n208), .Y(n421) );
  NAND3X1 U302 ( .A(n380), .B(n173), .C(n532), .Y(n137) );
  NOR2X1 U303 ( .A(n381), .B(n173), .Y(n88) );
  INVX1 U304 ( .A(n346), .Y(n544) );
  NAND3X1 U305 ( .A(n381), .B(n173), .C(n533), .Y(n150) );
  OAI21X1 U306 ( .B(n208), .C(n114), .A(n543), .Y(n207) );
  OAI21X1 U307 ( .B(n114), .C(n265), .A(n540), .Y(n299) );
  OAI21X1 U308 ( .B(n114), .C(n345), .A(n346), .Y(n392) );
  OAI21X1 U309 ( .B(n173), .C(n345), .A(n346), .Y(n333) );
  NAND2X1 U310 ( .A(n531), .B(n173), .Y(n65) );
  NAND2X1 U311 ( .A(n88), .B(n380), .Y(n84) );
  NAND2X1 U312 ( .A(n101), .B(n381), .Y(n99) );
  OAI22X1 U313 ( .A(n12), .B(n346), .C(n114), .D(n310), .Y(N743) );
  OAI31XL U314 ( .A(n536), .B(n12), .C(n522), .D(n415), .Y(N733) );
  INVX1 U315 ( .A(n173), .Y(n528) );
  NAND2X1 U316 ( .A(n433), .B(n4), .Y(n429) );
  INVX1 U317 ( .A(n45), .Y(n547) );
  OAI22X1 U318 ( .A(prx_wdat[7]), .B(n549), .C(r_wdat[7]), .D(prx_psh), .Y(n67) );
  INVX1 U319 ( .A(n60), .Y(fifowdat[0]) );
  INVX1 U320 ( .A(n57), .Y(fifowdat[1]) );
  INVX1 U321 ( .A(n54), .Y(fifowdat[2]) );
  NAND21X1 U322 ( .B(ptr[5]), .A(n6), .Y(n517) );
  INVX1 U323 ( .A(ptr[4]), .Y(n515) );
  INVX1 U324 ( .A(ptr[0]), .Y(n516) );
  NOR43XL U325 ( .B(n550), .C(n442), .D(n549), .A(n481), .Y(ps_locked) );
  AOI21X1 U326 ( .B(i_lockena), .C(n47), .A(locked), .Y(n481) );
  NOR2X1 U327 ( .A(r_unlock), .B(ps_locked), .Y(n44) );
  AO2222XL U328 ( .A(r_pop), .B(empty), .C(r_psh), .D(full), .E(n47), .F(n44), 
        .G(n551), .H(n547), .Y(ffack[1]) );
  OAI211X1 U329 ( .C(n443), .D(n484), .A(n452), .B(n61), .Y(N1023) );
  NAND2X1 U330 ( .A(dat_7_1[0]), .B(n445), .Y(n452) );
  OAI211X1 U331 ( .C(n443), .D(n500), .A(n450), .B(n55), .Y(N1025) );
  NAND2X1 U332 ( .A(dat_7_1[2]), .B(n445), .Y(n450) );
  OAI211X1 U333 ( .C(n443), .D(n508), .A(n449), .B(n51), .Y(N1026) );
  NAND2X1 U334 ( .A(dat_7_1[3]), .B(n445), .Y(n449) );
  OAI211X1 U335 ( .C(n443), .D(n21), .A(n448), .B(n17), .Y(N1027) );
  NAND2X1 U336 ( .A(dat_7_1[4]), .B(n445), .Y(n448) );
  OAI211X1 U337 ( .C(n443), .D(n37), .A(n446), .B(n33), .Y(N1029) );
  NAND2X1 U338 ( .A(dat_7_1[6]), .B(n445), .Y(n446) );
  OAI211X1 U339 ( .C(n443), .D(n48), .A(n444), .B(n41), .Y(N1030) );
  NAND2X1 U340 ( .A(dat_7_1[7]), .B(n445), .Y(n444) );
  OAI211X1 U341 ( .C(n443), .D(n492), .A(n451), .B(n58), .Y(N1024) );
  NAND2X1 U342 ( .A(dat_7_1[1]), .B(n445), .Y(n451) );
  OAI211X1 U343 ( .C(n443), .D(n29), .A(n447), .B(n25), .Y(N1028) );
  NAND2X1 U344 ( .A(dat_7_1[5]), .B(n445), .Y(n447) );
  OAI211X1 U345 ( .C(n465), .D(n484), .A(n474), .B(n61), .Y(N1005) );
  NAND2X1 U346 ( .A(dat_7_1[16]), .B(n467), .Y(n474) );
  OAI211X1 U347 ( .C(n465), .D(n492), .A(n488), .B(n473), .Y(N1006) );
  NAND2X1 U348 ( .A(dat_7_1[17]), .B(n467), .Y(n473) );
  OAI211X1 U349 ( .C(n465), .D(n500), .A(n496), .B(n472), .Y(N1007) );
  NAND2X1 U350 ( .A(dat_7_1[18]), .B(n467), .Y(n472) );
  OAI211X1 U351 ( .C(n465), .D(n508), .A(n504), .B(n471), .Y(N1008) );
  NAND2X1 U352 ( .A(dat_7_1[19]), .B(n467), .Y(n471) );
  OAI211X1 U353 ( .C(n465), .D(n21), .A(n470), .B(n17), .Y(N1009) );
  NAND2X1 U354 ( .A(dat_7_1[20]), .B(n467), .Y(n470) );
  OAI211X1 U355 ( .C(n49), .D(n21), .A(n479), .B(n17), .Y(N1000) );
  NAND2X1 U356 ( .A(dat_7_1[28]), .B(n53), .Y(n479) );
  OAI211X1 U357 ( .C(n49), .D(n29), .A(n25), .B(n478), .Y(N1001) );
  NAND2X1 U358 ( .A(dat_7_1[29]), .B(n53), .Y(n478) );
  OAI211X1 U359 ( .C(n49), .D(n37), .A(n33), .B(n477), .Y(N1002) );
  NAND2X1 U360 ( .A(dat_7_1[30]), .B(n53), .Y(n477) );
  OAI211X1 U361 ( .C(n49), .D(n48), .A(n41), .B(n476), .Y(N1003) );
  NAND2X1 U362 ( .A(dat_7_1[31]), .B(n53), .Y(n476) );
  OAI211X1 U363 ( .C(n455), .D(n21), .A(n460), .B(n17), .Y(N1018) );
  NAND2X1 U364 ( .A(dat_7_1[12]), .B(n457), .Y(n460) );
  OAI211X1 U365 ( .C(n455), .D(n29), .A(n459), .B(n25), .Y(N1019) );
  NAND2X1 U366 ( .A(dat_7_1[13]), .B(n457), .Y(n459) );
  OAI211X1 U367 ( .C(n455), .D(n37), .A(n458), .B(n33), .Y(N1020) );
  NAND2X1 U368 ( .A(dat_7_1[14]), .B(n457), .Y(n458) );
  OAI211X1 U369 ( .C(n455), .D(n48), .A(n456), .B(n41), .Y(N1021) );
  NAND2X1 U370 ( .A(dat_7_1[15]), .B(n457), .Y(n456) );
  OAI211X1 U371 ( .C(n102), .D(n494), .A(n110), .B(n488), .Y(N970) );
  NAND2X1 U372 ( .A(dat_7_1[49]), .B(n104), .Y(n110) );
  OAI211X1 U373 ( .C(n115), .D(n502), .A(n122), .B(n496), .Y(N962) );
  NAND2X1 U374 ( .A(mem_8__2_), .B(n117), .Y(n122) );
  OAI211X1 U375 ( .C(n115), .D(n23), .A(n120), .B(n19), .Y(N964) );
  NAND2X1 U376 ( .A(mem_8__4_), .B(n117), .Y(n120) );
  OAI211X1 U377 ( .C(n465), .D(n29), .A(n469), .B(n25), .Y(N1010) );
  NAND2X1 U378 ( .A(dat_7_1[21]), .B(n467), .Y(n469) );
  OAI211X1 U379 ( .C(n465), .D(n37), .A(n468), .B(n33), .Y(N1011) );
  NAND2X1 U380 ( .A(dat_7_1[22]), .B(n467), .Y(n468) );
  OAI211X1 U381 ( .C(n465), .D(n48), .A(n466), .B(n41), .Y(N1012) );
  NAND2X1 U382 ( .A(dat_7_1[23]), .B(n467), .Y(n466) );
  OAI211X1 U383 ( .C(n102), .D(n486), .A(n111), .B(n439), .Y(N969) );
  NAND2X1 U384 ( .A(dat_7_1[48]), .B(n104), .Y(n111) );
  OAI211X1 U385 ( .C(n115), .D(n486), .A(n124), .B(n439), .Y(N960) );
  NAND2X1 U386 ( .A(mem_8__0_), .B(n117), .Y(n124) );
  OAI211X1 U387 ( .C(n115), .D(n494), .A(n123), .B(n488), .Y(N961) );
  NAND2X1 U388 ( .A(mem_8__1_), .B(n117), .Y(n123) );
  OAI211X1 U389 ( .C(n102), .D(n502), .A(n109), .B(n496), .Y(N971) );
  NAND2X1 U390 ( .A(dat_7_1[50]), .B(n104), .Y(n109) );
  OAI211X1 U391 ( .C(n102), .D(n510), .A(n108), .B(n504), .Y(N972) );
  NAND2X1 U392 ( .A(dat_7_1[51]), .B(n104), .Y(n108) );
  OAI211X1 U393 ( .C(n115), .D(n510), .A(n121), .B(n504), .Y(N963) );
  NAND2X1 U394 ( .A(mem_8__3_), .B(n117), .Y(n121) );
  OAI211X1 U395 ( .C(n115), .D(n31), .A(n119), .B(n27), .Y(N965) );
  NAND2X1 U396 ( .A(mem_8__5_), .B(n117), .Y(n119) );
  OAI211X1 U397 ( .C(n115), .D(n39), .A(n118), .B(n35), .Y(N966) );
  NAND2X1 U398 ( .A(mem_8__6_), .B(n117), .Y(n118) );
  OAI211X1 U399 ( .C(n115), .D(n220), .A(n116), .B(n43), .Y(N967) );
  NAND2X1 U400 ( .A(mem_8__7_), .B(n117), .Y(n116) );
  OAI211X1 U401 ( .C(n455), .D(n484), .A(n464), .B(n61), .Y(N1014) );
  NAND2X1 U402 ( .A(dat_7_1[8]), .B(n457), .Y(n464) );
  OAI211X1 U403 ( .C(n455), .D(n492), .A(n463), .B(n488), .Y(N1015) );
  NAND2X1 U404 ( .A(dat_7_1[9]), .B(n457), .Y(n463) );
  OAI211X1 U405 ( .C(n455), .D(n500), .A(n462), .B(n496), .Y(N1016) );
  NAND2X1 U406 ( .A(dat_7_1[10]), .B(n457), .Y(n462) );
  OAI211X1 U407 ( .C(n455), .D(n508), .A(n461), .B(n504), .Y(N1017) );
  NAND2X1 U408 ( .A(dat_7_1[11]), .B(n457), .Y(n461) );
  OAI211X1 U409 ( .C(n127), .D(n486), .A(n136), .B(n439), .Y(N951) );
  NAND2X1 U410 ( .A(mem_9__0_), .B(n129), .Y(n136) );
  OAI211X1 U411 ( .C(n140), .D(n486), .A(n149), .B(n439), .Y(N942) );
  NAND2X1 U412 ( .A(mem_10__0_), .B(n142), .Y(n149) );
  OAI211X1 U413 ( .C(n152), .D(n486), .A(n161), .B(n439), .Y(N933) );
  NAND2X1 U414 ( .A(mem_11__0_), .B(n154), .Y(n161) );
  OAI211X1 U415 ( .C(n163), .D(n486), .A(n172), .B(n439), .Y(N924) );
  NAND2X1 U416 ( .A(mem_12__0_), .B(n165), .Y(n172) );
  OAI211X1 U417 ( .C(n174), .D(n486), .A(n183), .B(n439), .Y(N915) );
  NAND2X1 U418 ( .A(mem_13__0_), .B(n176), .Y(n183) );
  OAI211X1 U419 ( .C(n186), .D(n486), .A(n195), .B(n480), .Y(N906) );
  NAND2X1 U420 ( .A(mem_14__0_), .B(n188), .Y(n195) );
  OAI211X1 U421 ( .C(n197), .D(n486), .A(n206), .B(n480), .Y(N897) );
  NAND2X1 U422 ( .A(mem_15__0_), .B(n199), .Y(n206) );
  OAI211X1 U423 ( .C(n209), .D(n486), .A(n218), .B(n480), .Y(N888) );
  NAND2X1 U424 ( .A(mem_16__0_), .B(n211), .Y(n218) );
  OAI211X1 U425 ( .C(n221), .D(n485), .A(n230), .B(n480), .Y(N879) );
  NAND2X1 U426 ( .A(mem_17__0_), .B(n223), .Y(n230) );
  OAI211X1 U427 ( .C(n232), .D(n485), .A(n241), .B(n480), .Y(N870) );
  NAND2X1 U428 ( .A(mem_18__0_), .B(n234), .Y(n241) );
  OAI211X1 U429 ( .C(n244), .D(n485), .A(n253), .B(n480), .Y(N861) );
  NAND2X1 U430 ( .A(mem_19__0_), .B(n246), .Y(n253) );
  OAI211X1 U431 ( .C(n255), .D(n485), .A(n264), .B(n480), .Y(N852) );
  NAND2X1 U432 ( .A(mem_20__0_), .B(n257), .Y(n264) );
  OAI211X1 U433 ( .C(n266), .D(n485), .A(n275), .B(n480), .Y(N843) );
  NAND2X1 U434 ( .A(mem_21__0_), .B(n268), .Y(n275) );
  OAI211X1 U435 ( .C(n278), .D(n485), .A(n287), .B(n480), .Y(N834) );
  NAND2X1 U436 ( .A(mem_22__0_), .B(n280), .Y(n287) );
  OAI211X1 U437 ( .C(n289), .D(n485), .A(n298), .B(n480), .Y(N825) );
  NAND2X1 U438 ( .A(mem_23__0_), .B(n291), .Y(n298) );
  OAI211X1 U439 ( .C(n300), .D(n485), .A(n309), .B(n482), .Y(N816) );
  NAND2X1 U440 ( .A(mem_24__0_), .B(n302), .Y(n309) );
  OAI211X1 U441 ( .C(n311), .D(n485), .A(n320), .B(n482), .Y(N807) );
  NAND2X1 U442 ( .A(mem_25__0_), .B(n313), .Y(n320) );
  OAI211X1 U443 ( .C(n322), .D(n485), .A(n331), .B(n482), .Y(N798) );
  NAND2X1 U444 ( .A(mem_26__0_), .B(n324), .Y(n331) );
  OAI211X1 U445 ( .C(n334), .D(n484), .A(n343), .B(n482), .Y(N789) );
  NAND2X1 U446 ( .A(mem_27__0_), .B(n336), .Y(n343) );
  OAI211X1 U447 ( .C(n347), .D(n484), .A(n356), .B(n482), .Y(N780) );
  NAND2X1 U448 ( .A(mem_28__0_), .B(n349), .Y(n356) );
  OAI211X1 U449 ( .C(n127), .D(n494), .A(n135), .B(n488), .Y(N952) );
  NAND2X1 U450 ( .A(mem_9__1_), .B(n129), .Y(n135) );
  OAI211X1 U451 ( .C(n140), .D(n494), .A(n148), .B(n488), .Y(N943) );
  NAND2X1 U452 ( .A(mem_10__1_), .B(n142), .Y(n148) );
  OAI211X1 U453 ( .C(n152), .D(n494), .A(n160), .B(n488), .Y(N934) );
  NAND2X1 U454 ( .A(mem_11__1_), .B(n154), .Y(n160) );
  OAI211X1 U455 ( .C(n163), .D(n494), .A(n171), .B(n489), .Y(N925) );
  NAND2X1 U456 ( .A(mem_12__1_), .B(n165), .Y(n171) );
  OAI211X1 U457 ( .C(n174), .D(n494), .A(n182), .B(n489), .Y(N916) );
  NAND2X1 U458 ( .A(mem_13__1_), .B(n176), .Y(n182) );
  OAI211X1 U459 ( .C(n186), .D(n494), .A(n194), .B(n489), .Y(N907) );
  NAND2X1 U460 ( .A(mem_14__1_), .B(n188), .Y(n194) );
  OAI211X1 U461 ( .C(n197), .D(n494), .A(n205), .B(n489), .Y(N898) );
  NAND2X1 U462 ( .A(mem_15__1_), .B(n199), .Y(n205) );
  OAI211X1 U463 ( .C(n209), .D(n494), .A(n217), .B(n489), .Y(N889) );
  NAND2X1 U464 ( .A(mem_16__1_), .B(n211), .Y(n217) );
  OAI211X1 U465 ( .C(n221), .D(n493), .A(n229), .B(n489), .Y(N880) );
  NAND2X1 U466 ( .A(mem_17__1_), .B(n223), .Y(n229) );
  OAI211X1 U467 ( .C(n232), .D(n493), .A(n240), .B(n489), .Y(N871) );
  NAND2X1 U468 ( .A(mem_18__1_), .B(n234), .Y(n240) );
  OAI211X1 U469 ( .C(n244), .D(n493), .A(n252), .B(n489), .Y(N862) );
  NAND2X1 U470 ( .A(mem_19__1_), .B(n246), .Y(n252) );
  OAI211X1 U471 ( .C(n255), .D(n493), .A(n263), .B(n489), .Y(N853) );
  NAND2X1 U472 ( .A(mem_20__1_), .B(n257), .Y(n263) );
  OAI211X1 U473 ( .C(n266), .D(n493), .A(n274), .B(n489), .Y(N844) );
  NAND2X1 U474 ( .A(mem_21__1_), .B(n268), .Y(n274) );
  OAI211X1 U475 ( .C(n278), .D(n493), .A(n286), .B(n490), .Y(N835) );
  NAND2X1 U476 ( .A(mem_22__1_), .B(n280), .Y(n286) );
  OAI211X1 U477 ( .C(n289), .D(n493), .A(n297), .B(n490), .Y(N826) );
  NAND2X1 U478 ( .A(mem_23__1_), .B(n291), .Y(n297) );
  OAI211X1 U479 ( .C(n300), .D(n493), .A(n308), .B(n490), .Y(N817) );
  NAND2X1 U480 ( .A(mem_24__1_), .B(n302), .Y(n308) );
  OAI211X1 U481 ( .C(n311), .D(n493), .A(n319), .B(n490), .Y(N808) );
  NAND2X1 U482 ( .A(mem_25__1_), .B(n313), .Y(n319) );
  OAI211X1 U483 ( .C(n322), .D(n493), .A(n330), .B(n490), .Y(N799) );
  NAND2X1 U484 ( .A(mem_26__1_), .B(n324), .Y(n330) );
  OAI211X1 U485 ( .C(n334), .D(n492), .A(n342), .B(n490), .Y(N790) );
  NAND2X1 U486 ( .A(mem_27__1_), .B(n336), .Y(n342) );
  OAI211X1 U487 ( .C(n347), .D(n492), .A(n355), .B(n490), .Y(N781) );
  NAND2X1 U488 ( .A(mem_28__1_), .B(n349), .Y(n355) );
  OAI211X1 U489 ( .C(n127), .D(n502), .A(n134), .B(n496), .Y(N953) );
  NAND2X1 U490 ( .A(mem_9__2_), .B(n129), .Y(n134) );
  OAI211X1 U491 ( .C(n140), .D(n502), .A(n147), .B(n496), .Y(N944) );
  NAND2X1 U492 ( .A(mem_10__2_), .B(n142), .Y(n147) );
  OAI211X1 U493 ( .C(n152), .D(n502), .A(n159), .B(n496), .Y(N935) );
  NAND2X1 U494 ( .A(mem_11__2_), .B(n154), .Y(n159) );
  OAI211X1 U495 ( .C(n163), .D(n502), .A(n170), .B(n497), .Y(N926) );
  NAND2X1 U496 ( .A(mem_12__2_), .B(n165), .Y(n170) );
  OAI211X1 U497 ( .C(n174), .D(n502), .A(n181), .B(n497), .Y(N917) );
  NAND2X1 U498 ( .A(mem_13__2_), .B(n176), .Y(n181) );
  OAI211X1 U499 ( .C(n186), .D(n502), .A(n193), .B(n497), .Y(N908) );
  NAND2X1 U500 ( .A(mem_14__2_), .B(n188), .Y(n193) );
  OAI211X1 U501 ( .C(n197), .D(n502), .A(n204), .B(n497), .Y(N899) );
  NAND2X1 U502 ( .A(mem_15__2_), .B(n199), .Y(n204) );
  OAI211X1 U503 ( .C(n209), .D(n502), .A(n216), .B(n497), .Y(N890) );
  NAND2X1 U504 ( .A(mem_16__2_), .B(n211), .Y(n216) );
  OAI211X1 U505 ( .C(n221), .D(n501), .A(n228), .B(n497), .Y(N881) );
  NAND2X1 U506 ( .A(mem_17__2_), .B(n223), .Y(n228) );
  OAI211X1 U507 ( .C(n232), .D(n501), .A(n239), .B(n497), .Y(N872) );
  NAND2X1 U508 ( .A(mem_18__2_), .B(n234), .Y(n239) );
  OAI211X1 U509 ( .C(n244), .D(n501), .A(n251), .B(n497), .Y(N863) );
  NAND2X1 U510 ( .A(mem_19__2_), .B(n246), .Y(n251) );
  OAI211X1 U511 ( .C(n255), .D(n501), .A(n262), .B(n497), .Y(N854) );
  NAND2X1 U512 ( .A(mem_20__2_), .B(n257), .Y(n262) );
  OAI211X1 U513 ( .C(n266), .D(n501), .A(n273), .B(n497), .Y(N845) );
  NAND2X1 U514 ( .A(mem_21__2_), .B(n268), .Y(n273) );
  OAI211X1 U515 ( .C(n278), .D(n501), .A(n285), .B(n498), .Y(N836) );
  NAND2X1 U516 ( .A(mem_22__2_), .B(n280), .Y(n285) );
  OAI211X1 U517 ( .C(n289), .D(n501), .A(n296), .B(n498), .Y(N827) );
  NAND2X1 U518 ( .A(mem_23__2_), .B(n291), .Y(n296) );
  OAI211X1 U519 ( .C(n300), .D(n501), .A(n307), .B(n498), .Y(N818) );
  NAND2X1 U520 ( .A(mem_24__2_), .B(n302), .Y(n307) );
  OAI211X1 U521 ( .C(n311), .D(n501), .A(n318), .B(n498), .Y(N809) );
  NAND2X1 U522 ( .A(mem_25__2_), .B(n313), .Y(n318) );
  OAI211X1 U523 ( .C(n322), .D(n501), .A(n329), .B(n498), .Y(N800) );
  NAND2X1 U524 ( .A(mem_26__2_), .B(n324), .Y(n329) );
  OAI211X1 U525 ( .C(n334), .D(n500), .A(n341), .B(n498), .Y(N791) );
  NAND2X1 U526 ( .A(mem_27__2_), .B(n336), .Y(n341) );
  OAI211X1 U527 ( .C(n347), .D(n500), .A(n354), .B(n498), .Y(N782) );
  NAND2X1 U528 ( .A(mem_28__2_), .B(n349), .Y(n354) );
  OAI211X1 U529 ( .C(n127), .D(n510), .A(n133), .B(n504), .Y(N954) );
  NAND2X1 U530 ( .A(mem_9__3_), .B(n129), .Y(n133) );
  OAI211X1 U531 ( .C(n140), .D(n510), .A(n146), .B(n504), .Y(N945) );
  NAND2X1 U532 ( .A(mem_10__3_), .B(n142), .Y(n146) );
  OAI211X1 U533 ( .C(n152), .D(n510), .A(n158), .B(n504), .Y(N936) );
  NAND2X1 U534 ( .A(mem_11__3_), .B(n154), .Y(n158) );
  OAI211X1 U535 ( .C(n163), .D(n510), .A(n169), .B(n505), .Y(N927) );
  NAND2X1 U536 ( .A(mem_12__3_), .B(n165), .Y(n169) );
  OAI211X1 U537 ( .C(n174), .D(n510), .A(n180), .B(n505), .Y(N918) );
  NAND2X1 U538 ( .A(mem_13__3_), .B(n176), .Y(n180) );
  OAI211X1 U539 ( .C(n186), .D(n510), .A(n192), .B(n505), .Y(N909) );
  NAND2X1 U540 ( .A(mem_14__3_), .B(n188), .Y(n192) );
  OAI211X1 U541 ( .C(n197), .D(n510), .A(n203), .B(n505), .Y(N900) );
  NAND2X1 U542 ( .A(mem_15__3_), .B(n199), .Y(n203) );
  OAI211X1 U543 ( .C(n209), .D(n510), .A(n215), .B(n505), .Y(N891) );
  NAND2X1 U544 ( .A(mem_16__3_), .B(n211), .Y(n215) );
  OAI211X1 U545 ( .C(n221), .D(n509), .A(n227), .B(n505), .Y(N882) );
  NAND2X1 U546 ( .A(mem_17__3_), .B(n223), .Y(n227) );
  OAI211X1 U547 ( .C(n232), .D(n509), .A(n238), .B(n505), .Y(N873) );
  NAND2X1 U548 ( .A(mem_18__3_), .B(n234), .Y(n238) );
  OAI211X1 U549 ( .C(n244), .D(n509), .A(n250), .B(n505), .Y(N864) );
  NAND2X1 U550 ( .A(mem_19__3_), .B(n246), .Y(n250) );
  OAI211X1 U551 ( .C(n255), .D(n509), .A(n261), .B(n505), .Y(N855) );
  NAND2X1 U552 ( .A(mem_20__3_), .B(n257), .Y(n261) );
  OAI211X1 U553 ( .C(n266), .D(n509), .A(n272), .B(n505), .Y(N846) );
  NAND2X1 U554 ( .A(mem_21__3_), .B(n268), .Y(n272) );
  OAI211X1 U555 ( .C(n278), .D(n509), .A(n284), .B(n506), .Y(N837) );
  NAND2X1 U556 ( .A(mem_22__3_), .B(n280), .Y(n284) );
  OAI211X1 U557 ( .C(n289), .D(n509), .A(n295), .B(n506), .Y(N828) );
  NAND2X1 U558 ( .A(mem_23__3_), .B(n291), .Y(n295) );
  OAI211X1 U559 ( .C(n300), .D(n509), .A(n306), .B(n506), .Y(N819) );
  NAND2X1 U560 ( .A(mem_24__3_), .B(n302), .Y(n306) );
  OAI211X1 U561 ( .C(n311), .D(n509), .A(n317), .B(n506), .Y(N810) );
  NAND2X1 U562 ( .A(mem_25__3_), .B(n313), .Y(n317) );
  OAI211X1 U563 ( .C(n322), .D(n509), .A(n328), .B(n506), .Y(N801) );
  NAND2X1 U564 ( .A(mem_26__3_), .B(n324), .Y(n328) );
  OAI211X1 U565 ( .C(n334), .D(n508), .A(n340), .B(n506), .Y(N792) );
  NAND2X1 U566 ( .A(mem_27__3_), .B(n336), .Y(n340) );
  OAI211X1 U567 ( .C(n347), .D(n508), .A(n353), .B(n506), .Y(N783) );
  NAND2X1 U568 ( .A(mem_28__3_), .B(n349), .Y(n353) );
  OAI211X1 U569 ( .C(n127), .D(n23), .A(n132), .B(n19), .Y(N955) );
  NAND2X1 U570 ( .A(mem_9__4_), .B(n129), .Y(n132) );
  OAI211X1 U571 ( .C(n140), .D(n23), .A(n145), .B(n19), .Y(N946) );
  NAND2X1 U572 ( .A(mem_10__4_), .B(n142), .Y(n145) );
  OAI211X1 U573 ( .C(n152), .D(n23), .A(n157), .B(n19), .Y(N937) );
  NAND2X1 U574 ( .A(mem_11__4_), .B(n154), .Y(n157) );
  OAI211X1 U575 ( .C(n163), .D(n23), .A(n168), .B(n19), .Y(N928) );
  NAND2X1 U576 ( .A(mem_12__4_), .B(n165), .Y(n168) );
  OAI211X1 U577 ( .C(n174), .D(n23), .A(n179), .B(n19), .Y(N919) );
  NAND2X1 U578 ( .A(mem_13__4_), .B(n176), .Y(n179) );
  OAI211X1 U579 ( .C(n186), .D(n23), .A(n191), .B(n19), .Y(N910) );
  NAND2X1 U580 ( .A(mem_14__4_), .B(n188), .Y(n191) );
  OAI211X1 U581 ( .C(n197), .D(n23), .A(n202), .B(n19), .Y(N901) );
  NAND2X1 U582 ( .A(mem_15__4_), .B(n199), .Y(n202) );
  OAI211X1 U583 ( .C(n209), .D(n23), .A(n214), .B(n19), .Y(N892) );
  NAND2X1 U584 ( .A(mem_16__4_), .B(n211), .Y(n214) );
  OAI211X1 U585 ( .C(n221), .D(n23), .A(n226), .B(n19), .Y(N883) );
  NAND2X1 U586 ( .A(mem_17__4_), .B(n223), .Y(n226) );
  OAI211X1 U587 ( .C(n232), .D(n22), .A(n237), .B(n18), .Y(N874) );
  NAND2X1 U588 ( .A(mem_18__4_), .B(n234), .Y(n237) );
  OAI211X1 U589 ( .C(n244), .D(n22), .A(n249), .B(n18), .Y(N865) );
  NAND2X1 U590 ( .A(mem_19__4_), .B(n246), .Y(n249) );
  OAI211X1 U591 ( .C(n255), .D(n22), .A(n260), .B(n18), .Y(N856) );
  NAND2X1 U592 ( .A(mem_20__4_), .B(n257), .Y(n260) );
  OAI211X1 U593 ( .C(n266), .D(n22), .A(n271), .B(n18), .Y(N847) );
  NAND2X1 U594 ( .A(mem_21__4_), .B(n268), .Y(n271) );
  OAI211X1 U595 ( .C(n278), .D(n22), .A(n283), .B(n18), .Y(N838) );
  NAND2X1 U596 ( .A(mem_22__4_), .B(n280), .Y(n283) );
  OAI211X1 U597 ( .C(n289), .D(n22), .A(n294), .B(n18), .Y(N829) );
  NAND2X1 U598 ( .A(mem_23__4_), .B(n291), .Y(n294) );
  OAI211X1 U599 ( .C(n300), .D(n22), .A(n305), .B(n18), .Y(N820) );
  NAND2X1 U600 ( .A(mem_24__4_), .B(n302), .Y(n305) );
  OAI211X1 U601 ( .C(n311), .D(n22), .A(n316), .B(n18), .Y(N811) );
  NAND2X1 U602 ( .A(mem_25__4_), .B(n313), .Y(n316) );
  OAI211X1 U603 ( .C(n322), .D(n22), .A(n327), .B(n18), .Y(N802) );
  NAND2X1 U604 ( .A(mem_26__4_), .B(n324), .Y(n327) );
  OAI211X1 U605 ( .C(n334), .D(n22), .A(n339), .B(n18), .Y(N793) );
  NAND2X1 U606 ( .A(mem_27__4_), .B(n336), .Y(n339) );
  OAI211X1 U607 ( .C(n347), .D(n21), .A(n352), .B(n17), .Y(N784) );
  NAND2X1 U608 ( .A(mem_28__4_), .B(n349), .Y(n352) );
  OAI211X1 U609 ( .C(n127), .D(n31), .A(n131), .B(n27), .Y(N956) );
  NAND2X1 U610 ( .A(mem_9__5_), .B(n129), .Y(n131) );
  OAI211X1 U611 ( .C(n140), .D(n31), .A(n144), .B(n27), .Y(N947) );
  NAND2X1 U612 ( .A(mem_10__5_), .B(n142), .Y(n144) );
  OAI211X1 U613 ( .C(n152), .D(n31), .A(n156), .B(n27), .Y(N938) );
  NAND2X1 U614 ( .A(mem_11__5_), .B(n154), .Y(n156) );
  OAI211X1 U615 ( .C(n163), .D(n31), .A(n167), .B(n27), .Y(N929) );
  NAND2X1 U616 ( .A(mem_12__5_), .B(n165), .Y(n167) );
  OAI211X1 U617 ( .C(n174), .D(n31), .A(n178), .B(n27), .Y(N920) );
  NAND2X1 U618 ( .A(mem_13__5_), .B(n176), .Y(n178) );
  OAI211X1 U619 ( .C(n186), .D(n31), .A(n190), .B(n27), .Y(N911) );
  NAND2X1 U620 ( .A(mem_14__5_), .B(n188), .Y(n190) );
  OAI211X1 U621 ( .C(n197), .D(n31), .A(n201), .B(n27), .Y(N902) );
  NAND2X1 U622 ( .A(mem_15__5_), .B(n199), .Y(n201) );
  OAI211X1 U623 ( .C(n209), .D(n31), .A(n213), .B(n27), .Y(N893) );
  NAND2X1 U624 ( .A(mem_16__5_), .B(n211), .Y(n213) );
  OAI211X1 U625 ( .C(n221), .D(n31), .A(n225), .B(n27), .Y(N884) );
  NAND2X1 U626 ( .A(mem_17__5_), .B(n223), .Y(n225) );
  OAI211X1 U627 ( .C(n232), .D(n30), .A(n236), .B(n26), .Y(N875) );
  NAND2X1 U628 ( .A(mem_18__5_), .B(n234), .Y(n236) );
  OAI211X1 U629 ( .C(n244), .D(n30), .A(n248), .B(n26), .Y(N866) );
  NAND2X1 U630 ( .A(mem_19__5_), .B(n246), .Y(n248) );
  OAI211X1 U631 ( .C(n255), .D(n30), .A(n259), .B(n26), .Y(N857) );
  NAND2X1 U632 ( .A(mem_20__5_), .B(n257), .Y(n259) );
  OAI211X1 U633 ( .C(n266), .D(n30), .A(n270), .B(n26), .Y(N848) );
  NAND2X1 U634 ( .A(mem_21__5_), .B(n268), .Y(n270) );
  OAI211X1 U635 ( .C(n278), .D(n30), .A(n282), .B(n26), .Y(N839) );
  NAND2X1 U636 ( .A(mem_22__5_), .B(n280), .Y(n282) );
  OAI211X1 U637 ( .C(n289), .D(n30), .A(n293), .B(n26), .Y(N830) );
  NAND2X1 U638 ( .A(mem_23__5_), .B(n291), .Y(n293) );
  OAI211X1 U639 ( .C(n300), .D(n30), .A(n304), .B(n26), .Y(N821) );
  NAND2X1 U640 ( .A(mem_24__5_), .B(n302), .Y(n304) );
  OAI211X1 U641 ( .C(n311), .D(n30), .A(n315), .B(n26), .Y(N812) );
  NAND2X1 U642 ( .A(mem_25__5_), .B(n313), .Y(n315) );
  OAI211X1 U643 ( .C(n322), .D(n30), .A(n326), .B(n26), .Y(N803) );
  NAND2X1 U644 ( .A(mem_26__5_), .B(n324), .Y(n326) );
  OAI211X1 U645 ( .C(n334), .D(n30), .A(n338), .B(n26), .Y(N794) );
  NAND2X1 U646 ( .A(mem_27__5_), .B(n336), .Y(n338) );
  OAI211X1 U647 ( .C(n347), .D(n29), .A(n351), .B(n25), .Y(N785) );
  NAND2X1 U648 ( .A(mem_28__5_), .B(n349), .Y(n351) );
  OAI211X1 U649 ( .C(n127), .D(n39), .A(n130), .B(n35), .Y(N957) );
  NAND2X1 U650 ( .A(mem_9__6_), .B(n129), .Y(n130) );
  OAI211X1 U651 ( .C(n140), .D(n39), .A(n143), .B(n35), .Y(N948) );
  NAND2X1 U652 ( .A(mem_10__6_), .B(n142), .Y(n143) );
  OAI211X1 U653 ( .C(n152), .D(n39), .A(n155), .B(n35), .Y(N939) );
  NAND2X1 U654 ( .A(mem_11__6_), .B(n154), .Y(n155) );
  OAI211X1 U655 ( .C(n163), .D(n39), .A(n166), .B(n35), .Y(N930) );
  NAND2X1 U656 ( .A(mem_12__6_), .B(n165), .Y(n166) );
  OAI211X1 U657 ( .C(n174), .D(n39), .A(n177), .B(n35), .Y(N921) );
  NAND2X1 U658 ( .A(mem_13__6_), .B(n176), .Y(n177) );
  OAI211X1 U659 ( .C(n186), .D(n39), .A(n189), .B(n35), .Y(N912) );
  NAND2X1 U660 ( .A(mem_14__6_), .B(n188), .Y(n189) );
  OAI211X1 U661 ( .C(n197), .D(n39), .A(n200), .B(n35), .Y(N903) );
  NAND2X1 U662 ( .A(mem_15__6_), .B(n199), .Y(n200) );
  OAI211X1 U663 ( .C(n209), .D(n39), .A(n212), .B(n35), .Y(N894) );
  NAND2X1 U664 ( .A(mem_16__6_), .B(n211), .Y(n212) );
  OAI211X1 U665 ( .C(n221), .D(n39), .A(n224), .B(n35), .Y(N885) );
  NAND2X1 U666 ( .A(mem_17__6_), .B(n223), .Y(n224) );
  OAI211X1 U667 ( .C(n232), .D(n38), .A(n235), .B(n34), .Y(N876) );
  NAND2X1 U668 ( .A(mem_18__6_), .B(n234), .Y(n235) );
  OAI211X1 U669 ( .C(n244), .D(n38), .A(n247), .B(n34), .Y(N867) );
  NAND2X1 U670 ( .A(mem_19__6_), .B(n246), .Y(n247) );
  OAI211X1 U671 ( .C(n255), .D(n38), .A(n258), .B(n34), .Y(N858) );
  NAND2X1 U672 ( .A(mem_20__6_), .B(n257), .Y(n258) );
  OAI211X1 U673 ( .C(n266), .D(n38), .A(n269), .B(n34), .Y(N849) );
  NAND2X1 U674 ( .A(mem_21__6_), .B(n268), .Y(n269) );
  OAI211X1 U675 ( .C(n278), .D(n38), .A(n281), .B(n34), .Y(N840) );
  NAND2X1 U676 ( .A(mem_22__6_), .B(n280), .Y(n281) );
  OAI211X1 U677 ( .C(n289), .D(n38), .A(n292), .B(n34), .Y(N831) );
  NAND2X1 U678 ( .A(mem_23__6_), .B(n291), .Y(n292) );
  OAI211X1 U679 ( .C(n300), .D(n38), .A(n303), .B(n34), .Y(N822) );
  NAND2X1 U680 ( .A(mem_24__6_), .B(n302), .Y(n303) );
  OAI211X1 U681 ( .C(n311), .D(n38), .A(n314), .B(n34), .Y(N813) );
  NAND2X1 U682 ( .A(mem_25__6_), .B(n313), .Y(n314) );
  OAI211X1 U683 ( .C(n322), .D(n38), .A(n325), .B(n34), .Y(N804) );
  NAND2X1 U684 ( .A(mem_26__6_), .B(n324), .Y(n325) );
  OAI211X1 U685 ( .C(n334), .D(n38), .A(n337), .B(n34), .Y(N795) );
  NAND2X1 U686 ( .A(mem_27__6_), .B(n336), .Y(n337) );
  OAI211X1 U687 ( .C(n347), .D(n37), .A(n350), .B(n33), .Y(N786) );
  NAND2X1 U688 ( .A(mem_28__6_), .B(n349), .Y(n350) );
  OAI211X1 U689 ( .C(n127), .D(n220), .A(n128), .B(n43), .Y(N958) );
  NAND2X1 U690 ( .A(mem_9__7_), .B(n129), .Y(n128) );
  OAI211X1 U691 ( .C(n140), .D(n220), .A(n141), .B(n43), .Y(N949) );
  NAND2X1 U692 ( .A(mem_10__7_), .B(n142), .Y(n141) );
  OAI211X1 U693 ( .C(n152), .D(n220), .A(n153), .B(n43), .Y(N940) );
  NAND2X1 U694 ( .A(mem_11__7_), .B(n154), .Y(n153) );
  OAI211X1 U695 ( .C(n163), .D(n220), .A(n164), .B(n43), .Y(N931) );
  NAND2X1 U696 ( .A(mem_12__7_), .B(n165), .Y(n164) );
  OAI211X1 U697 ( .C(n174), .D(n220), .A(n175), .B(n43), .Y(N922) );
  NAND2X1 U698 ( .A(mem_13__7_), .B(n176), .Y(n175) );
  OAI211X1 U699 ( .C(n186), .D(n220), .A(n187), .B(n43), .Y(N913) );
  NAND2X1 U700 ( .A(mem_14__7_), .B(n188), .Y(n187) );
  OAI211X1 U701 ( .C(n197), .D(n220), .A(n198), .B(n43), .Y(N904) );
  NAND2X1 U702 ( .A(mem_15__7_), .B(n199), .Y(n198) );
  OAI211X1 U703 ( .C(n209), .D(n220), .A(n210), .B(n43), .Y(N895) );
  NAND2X1 U704 ( .A(mem_16__7_), .B(n211), .Y(n210) );
  OAI211X1 U705 ( .C(n221), .D(n220), .A(n222), .B(n43), .Y(N886) );
  NAND2X1 U706 ( .A(mem_17__7_), .B(n223), .Y(n222) );
  OAI211X1 U707 ( .C(n232), .D(n113), .A(n233), .B(n42), .Y(N877) );
  NAND2X1 U708 ( .A(mem_18__7_), .B(n234), .Y(n233) );
  OAI211X1 U709 ( .C(n244), .D(n113), .A(n245), .B(n42), .Y(N868) );
  NAND2X1 U710 ( .A(mem_19__7_), .B(n246), .Y(n245) );
  OAI211X1 U711 ( .C(n255), .D(n113), .A(n256), .B(n42), .Y(N859) );
  NAND2X1 U712 ( .A(mem_20__7_), .B(n257), .Y(n256) );
  OAI211X1 U713 ( .C(n266), .D(n113), .A(n267), .B(n42), .Y(N850) );
  NAND2X1 U714 ( .A(mem_21__7_), .B(n268), .Y(n267) );
  OAI211X1 U715 ( .C(n278), .D(n113), .A(n279), .B(n42), .Y(N841) );
  NAND2X1 U716 ( .A(mem_22__7_), .B(n280), .Y(n279) );
  OAI211X1 U717 ( .C(n289), .D(n113), .A(n290), .B(n42), .Y(N832) );
  NAND2X1 U718 ( .A(mem_23__7_), .B(n291), .Y(n290) );
  OAI211X1 U719 ( .C(n300), .D(n113), .A(n301), .B(n42), .Y(N823) );
  NAND2X1 U720 ( .A(mem_24__7_), .B(n302), .Y(n301) );
  OAI211X1 U721 ( .C(n311), .D(n113), .A(n312), .B(n42), .Y(N814) );
  NAND2X1 U722 ( .A(mem_25__7_), .B(n313), .Y(n312) );
  OAI211X1 U723 ( .C(n322), .D(n113), .A(n323), .B(n42), .Y(N805) );
  NAND2X1 U724 ( .A(mem_26__7_), .B(n324), .Y(n323) );
  OAI211X1 U725 ( .C(n334), .D(n113), .A(n335), .B(n42), .Y(N796) );
  NAND2X1 U726 ( .A(mem_27__7_), .B(n336), .Y(n335) );
  OAI211X1 U727 ( .C(n347), .D(n48), .A(n348), .B(n41), .Y(N787) );
  NAND2X1 U728 ( .A(mem_28__7_), .B(n349), .Y(n348) );
  OAI211X1 U729 ( .C(n358), .D(n484), .A(n367), .B(n482), .Y(N771) );
  NAND2X1 U730 ( .A(mem_29__0_), .B(n360), .Y(n367) );
  OAI211X1 U731 ( .C(n370), .D(n484), .A(n379), .B(n482), .Y(N762) );
  NAND2X1 U732 ( .A(mem_30__0_), .B(n372), .Y(n379) );
  OAI211X1 U733 ( .C(n382), .D(n484), .A(n391), .B(n482), .Y(N753) );
  NAND2X1 U734 ( .A(mem_31__0_), .B(n384), .Y(n391) );
  OAI211X1 U735 ( .C(n393), .D(n484), .A(n402), .B(n482), .Y(N744) );
  NAND2X1 U736 ( .A(mem_32__0_), .B(n395), .Y(n402) );
  OAI211X1 U737 ( .C(n404), .D(n484), .A(n413), .B(n482), .Y(N735) );
  NAND2X1 U738 ( .A(mem_33__0_), .B(n406), .Y(n413) );
  OAI211X1 U739 ( .C(n358), .D(n492), .A(n366), .B(n490), .Y(N772) );
  NAND2X1 U740 ( .A(mem_29__1_), .B(n360), .Y(n366) );
  OAI211X1 U741 ( .C(n370), .D(n492), .A(n378), .B(n490), .Y(N763) );
  NAND2X1 U742 ( .A(mem_30__1_), .B(n372), .Y(n378) );
  OAI211X1 U743 ( .C(n382), .D(n492), .A(n390), .B(n490), .Y(N754) );
  NAND2X1 U744 ( .A(mem_31__1_), .B(n384), .Y(n390) );
  OAI211X1 U745 ( .C(n393), .D(n492), .A(n401), .B(n58), .Y(N745) );
  NAND2X1 U746 ( .A(mem_32__1_), .B(n395), .Y(n401) );
  OAI211X1 U747 ( .C(n404), .D(n492), .A(n412), .B(n58), .Y(N736) );
  NAND2X1 U748 ( .A(mem_33__1_), .B(n406), .Y(n412) );
  OAI211X1 U749 ( .C(n358), .D(n500), .A(n365), .B(n498), .Y(N773) );
  NAND2X1 U750 ( .A(mem_29__2_), .B(n360), .Y(n365) );
  OAI211X1 U751 ( .C(n370), .D(n500), .A(n377), .B(n498), .Y(N764) );
  NAND2X1 U752 ( .A(mem_30__2_), .B(n372), .Y(n377) );
  OAI211X1 U753 ( .C(n382), .D(n500), .A(n389), .B(n498), .Y(N755) );
  NAND2X1 U754 ( .A(mem_31__2_), .B(n384), .Y(n389) );
  OAI211X1 U755 ( .C(n393), .D(n500), .A(n400), .B(n55), .Y(N746) );
  NAND2X1 U756 ( .A(mem_32__2_), .B(n395), .Y(n400) );
  OAI211X1 U757 ( .C(n404), .D(n500), .A(n411), .B(n55), .Y(N737) );
  NAND2X1 U758 ( .A(mem_33__2_), .B(n406), .Y(n411) );
  OAI211X1 U759 ( .C(n358), .D(n508), .A(n364), .B(n506), .Y(N774) );
  NAND2X1 U760 ( .A(mem_29__3_), .B(n360), .Y(n364) );
  OAI211X1 U761 ( .C(n370), .D(n508), .A(n376), .B(n506), .Y(N765) );
  NAND2X1 U762 ( .A(mem_30__3_), .B(n372), .Y(n376) );
  OAI211X1 U763 ( .C(n382), .D(n508), .A(n388), .B(n506), .Y(N756) );
  NAND2X1 U764 ( .A(mem_31__3_), .B(n384), .Y(n388) );
  OAI211X1 U765 ( .C(n393), .D(n508), .A(n399), .B(n51), .Y(N747) );
  NAND2X1 U766 ( .A(mem_32__3_), .B(n395), .Y(n399) );
  OAI211X1 U767 ( .C(n404), .D(n508), .A(n410), .B(n51), .Y(N738) );
  NAND2X1 U768 ( .A(mem_33__3_), .B(n406), .Y(n410) );
  OAI211X1 U769 ( .C(n358), .D(n21), .A(n363), .B(n17), .Y(N775) );
  NAND2X1 U770 ( .A(mem_29__4_), .B(n360), .Y(n363) );
  OAI211X1 U771 ( .C(n370), .D(n21), .A(n375), .B(n17), .Y(N766) );
  NAND2X1 U772 ( .A(mem_30__4_), .B(n372), .Y(n375) );
  OAI211X1 U773 ( .C(n382), .D(n21), .A(n387), .B(n17), .Y(N757) );
  NAND2X1 U774 ( .A(mem_31__4_), .B(n384), .Y(n387) );
  OAI211X1 U775 ( .C(n393), .D(n21), .A(n398), .B(n17), .Y(N748) );
  NAND2X1 U776 ( .A(mem_32__4_), .B(n395), .Y(n398) );
  OAI211X1 U777 ( .C(n404), .D(n21), .A(n409), .B(n17), .Y(N739) );
  NAND2X1 U778 ( .A(mem_33__4_), .B(n406), .Y(n409) );
  OAI211X1 U779 ( .C(n358), .D(n29), .A(n362), .B(n25), .Y(N776) );
  NAND2X1 U780 ( .A(mem_29__5_), .B(n360), .Y(n362) );
  OAI211X1 U781 ( .C(n370), .D(n29), .A(n374), .B(n25), .Y(N767) );
  NAND2X1 U782 ( .A(mem_30__5_), .B(n372), .Y(n374) );
  OAI211X1 U783 ( .C(n382), .D(n29), .A(n386), .B(n25), .Y(N758) );
  NAND2X1 U784 ( .A(mem_31__5_), .B(n384), .Y(n386) );
  OAI211X1 U785 ( .C(n393), .D(n29), .A(n397), .B(n25), .Y(N749) );
  NAND2X1 U786 ( .A(mem_32__5_), .B(n395), .Y(n397) );
  OAI211X1 U787 ( .C(n404), .D(n29), .A(n408), .B(n25), .Y(N740) );
  NAND2X1 U788 ( .A(mem_33__5_), .B(n406), .Y(n408) );
  OAI211X1 U789 ( .C(n358), .D(n37), .A(n361), .B(n33), .Y(N777) );
  NAND2X1 U790 ( .A(mem_29__6_), .B(n360), .Y(n361) );
  OAI211X1 U791 ( .C(n370), .D(n37), .A(n373), .B(n33), .Y(N768) );
  NAND2X1 U792 ( .A(mem_30__6_), .B(n372), .Y(n373) );
  OAI211X1 U793 ( .C(n382), .D(n37), .A(n385), .B(n33), .Y(N759) );
  NAND2X1 U794 ( .A(mem_31__6_), .B(n384), .Y(n385) );
  OAI211X1 U795 ( .C(n393), .D(n37), .A(n396), .B(n33), .Y(N750) );
  NAND2X1 U796 ( .A(mem_32__6_), .B(n395), .Y(n396) );
  OAI211X1 U797 ( .C(n404), .D(n37), .A(n407), .B(n33), .Y(N741) );
  NAND2X1 U798 ( .A(mem_33__6_), .B(n406), .Y(n407) );
  OAI211X1 U799 ( .C(n358), .D(n48), .A(n359), .B(n41), .Y(N778) );
  NAND2X1 U800 ( .A(mem_29__7_), .B(n360), .Y(n359) );
  OAI211X1 U801 ( .C(n370), .D(n48), .A(n371), .B(n41), .Y(N769) );
  NAND2X1 U802 ( .A(mem_30__7_), .B(n372), .Y(n371) );
  OAI211X1 U803 ( .C(n382), .D(n48), .A(n383), .B(n41), .Y(N760) );
  NAND2X1 U804 ( .A(mem_31__7_), .B(n384), .Y(n383) );
  OAI211X1 U805 ( .C(n393), .D(n48), .A(n394), .B(n41), .Y(N751) );
  NAND2X1 U806 ( .A(mem_32__7_), .B(n395), .Y(n394) );
  OAI211X1 U807 ( .C(n404), .D(n48), .A(n405), .B(n41), .Y(N742) );
  NAND2X1 U808 ( .A(mem_33__7_), .B(n406), .Y(n405) );
  OAI211X1 U809 ( .C(n66), .D(n57), .A(n82), .B(n488), .Y(N988) );
  NAND2X1 U810 ( .A(dat_7_1[33]), .B(n70), .Y(n82) );
  OAI211X1 U811 ( .C(n89), .D(n54), .A(n96), .B(n496), .Y(N980) );
  NAND2X1 U812 ( .A(dat_7_1[42]), .B(n91), .Y(n96) );
  OAI211X1 U813 ( .C(n89), .D(n50), .A(n95), .B(n504), .Y(N981) );
  NAND2X1 U814 ( .A(dat_7_1[43]), .B(n91), .Y(n95) );
  OAI211X1 U815 ( .C(n89), .D(n77), .A(n94), .B(n79), .Y(N982) );
  NAND2X1 U816 ( .A(dat_7_1[44]), .B(n91), .Y(n94) );
  OAI211X1 U817 ( .C(n89), .D(n71), .A(n92), .B(n73), .Y(N984) );
  NAND2X1 U818 ( .A(dat_7_1[46]), .B(n91), .Y(n92) );
  OAI211X1 U819 ( .C(n49), .D(n60), .A(n439), .B(n62), .Y(N996) );
  NAND2X1 U820 ( .A(dat_7_1[24]), .B(n53), .Y(n62) );
  OAI211X1 U821 ( .C(n49), .D(n57), .A(n488), .B(n59), .Y(N997) );
  NAND2X1 U822 ( .A(dat_7_1[25]), .B(n53), .Y(n59) );
  OAI211X1 U823 ( .C(n49), .D(n54), .A(n496), .B(n56), .Y(N998) );
  NAND2X1 U824 ( .A(dat_7_1[26]), .B(n53), .Y(n56) );
  OAI211X1 U825 ( .C(n49), .D(n50), .A(n504), .B(n52), .Y(N999) );
  NAND2X1 U826 ( .A(dat_7_1[27]), .B(n53), .Y(n52) );
  OAI211X1 U827 ( .C(n66), .D(n60), .A(n83), .B(n439), .Y(N987) );
  NAND2X1 U828 ( .A(dat_7_1[32]), .B(n70), .Y(n83) );
  OAI211X1 U829 ( .C(n89), .D(n60), .A(n98), .B(n439), .Y(N978) );
  NAND2X1 U830 ( .A(dat_7_1[40]), .B(n91), .Y(n98) );
  OAI211X1 U831 ( .C(n89), .D(n57), .A(n97), .B(n488), .Y(N979) );
  NAND2X1 U832 ( .A(dat_7_1[41]), .B(n91), .Y(n97) );
  OAI211X1 U833 ( .C(n66), .D(n54), .A(n81), .B(n496), .Y(N989) );
  NAND2X1 U834 ( .A(dat_7_1[34]), .B(n70), .Y(n81) );
  OAI211X1 U835 ( .C(n66), .D(n50), .A(n80), .B(n504), .Y(N990) );
  NAND2X1 U836 ( .A(dat_7_1[35]), .B(n70), .Y(n80) );
  OAI211X1 U837 ( .C(n66), .D(n77), .A(n78), .B(n79), .Y(N991) );
  NAND2X1 U838 ( .A(dat_7_1[36]), .B(n70), .Y(n78) );
  OAI211X1 U839 ( .C(n66), .D(n74), .A(n75), .B(n76), .Y(N992) );
  NAND2X1 U840 ( .A(dat_7_1[37]), .B(n70), .Y(n75) );
  OAI211X1 U841 ( .C(n89), .D(n74), .A(n93), .B(n76), .Y(N983) );
  NAND2X1 U842 ( .A(dat_7_1[45]), .B(n91), .Y(n93) );
  OAI211X1 U843 ( .C(n66), .D(n71), .A(n72), .B(n73), .Y(N993) );
  NAND2X1 U844 ( .A(dat_7_1[38]), .B(n70), .Y(n72) );
  OAI211X1 U845 ( .C(n66), .D(n67), .A(n68), .B(n69), .Y(N994) );
  NAND2X1 U846 ( .A(dat_7_1[39]), .B(n70), .Y(n68) );
  OAI211X1 U847 ( .C(n89), .D(n67), .A(n90), .B(n69), .Y(N985) );
  NAND2X1 U848 ( .A(dat_7_1[47]), .B(n91), .Y(n90) );
  OAI211X1 U849 ( .C(n102), .D(n77), .A(n107), .B(n79), .Y(N973) );
  NAND2X1 U850 ( .A(dat_7_1[52]), .B(n104), .Y(n107) );
  OAI211X1 U851 ( .C(n102), .D(n74), .A(n106), .B(n76), .Y(N974) );
  NAND2X1 U852 ( .A(dat_7_1[53]), .B(n104), .Y(n106) );
  OAI211X1 U853 ( .C(n102), .D(n71), .A(n105), .B(n73), .Y(N975) );
  NAND2X1 U854 ( .A(dat_7_1[54]), .B(n104), .Y(n105) );
  OAI211X1 U855 ( .C(n102), .D(n67), .A(n103), .B(n69), .Y(N976) );
  NAND2X1 U856 ( .A(dat_7_1[55]), .B(n104), .Y(n103) );
  NOR2X1 U857 ( .A(n7), .B(n44), .Y(ffack[0]) );
  NAND2X1 U858 ( .A(ptr[4]), .B(n442), .Y(n265) );
  NAND2X1 U859 ( .A(r_psh), .B(r_last), .Y(n45) );
  OAI22X1 U860 ( .A(prx_wdat[0]), .B(n549), .C(r_wdat[0]), .D(prx_psh), .Y(n60) );
  OAI22X1 U861 ( .A(prx_wdat[1]), .B(n549), .C(r_wdat[1]), .D(prx_psh), .Y(n57) );
  OAI22X1 U862 ( .A(prx_wdat[2]), .B(n549), .C(r_wdat[2]), .D(prx_psh), .Y(n54) );
  AND2X1 U863 ( .A(n519), .B(n513), .Y(obsd) );
  INVX1 U864 ( .A(srstz), .Y(n513) );
  INVX1 U865 ( .A(i_ccidle), .Y(n551) );
  OAI22XL U866 ( .A(prx_wdat[4]), .B(n549), .C(r_wdat[4]), .D(prx_psh), .Y(n77) );
  OAI22XL U867 ( .A(prx_wdat[6]), .B(n549), .C(r_wdat[6]), .D(prx_psh), .Y(n71) );
  OAI22XL U868 ( .A(prx_wdat[5]), .B(n549), .C(r_wdat[5]), .D(prx_psh), .Y(n74) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phycrc_a0 ( crc32_3_0, rx_good, i_shfidat, i_start, i_shfi4, i_shfo4, 
        clk, test_si, test_so, test_se );
  output [3:0] crc32_3_0;
  input [3:0] i_shfidat;
  input i_start, i_shfi4, i_shfo4, clk, test_si, test_se;
  output rx_good, test_so;
  wire   crc32_r_30_, crc32_r_29_, crc32_r_28_, crc32_r_27_, crc32_r_26_,
         crc32_r_25_, crc32_r_24_, crc32_r_23_, crc32_r_22_, crc32_r_21_,
         crc32_r_20_, crc32_r_19_, crc32_r_18_, crc32_r_17_, crc32_r_16_,
         crc32_r_15_, crc32_r_14_, crc32_r_13_, crc32_r_12_, crc32_r_11_,
         crc32_r_10_, crc32_r_9_, crc32_r_8_, crc32_r_7_, crc32_r_6_,
         crc32_r_5_, crc32_r_4_, crc32_r_3_, crc32_r_2_, crc32_r_1_,
         crc32_r_0_, N188, N189, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, net10566, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n58, n121, n122, n123, n124, n125, n126, n127;

  SNPS_CLOCK_GATE_HIGH_phycrc_a0 clk_gate_crc32_r_reg ( .CLK(clk), .EN(N188), 
        .ENCLK(net10566), .TE(test_se) );
  SDFFQX1 crc32_r_reg_26_ ( .D(N215), .SIN(crc32_r_25_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_26_) );
  SDFFQX1 crc32_r_reg_16_ ( .D(N205), .SIN(crc32_r_15_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_16_) );
  SDFFQX1 crc32_r_reg_27_ ( .D(N216), .SIN(crc32_r_26_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_27_) );
  SDFFQX1 crc32_r_reg_17_ ( .D(N206), .SIN(crc32_r_16_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_17_) );
  SDFFQX1 crc32_r_reg_8_ ( .D(N197), .SIN(crc32_r_7_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_8_) );
  SDFFQX1 crc32_r_reg_5_ ( .D(N194), .SIN(crc32_r_4_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_5_) );
  SDFFQX1 crc32_r_reg_4_ ( .D(N193), .SIN(crc32_r_3_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_4_) );
  SDFFQX1 crc32_r_reg_0_ ( .D(N189), .SIN(test_si), .SMC(test_se), .C(net10566), .Q(crc32_r_0_) );
  SDFFQX1 crc32_r_reg_1_ ( .D(N190), .SIN(crc32_r_0_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_1_) );
  SDFFQX1 crc32_r_reg_10_ ( .D(N199), .SIN(crc32_r_9_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_10_) );
  SDFFQX1 crc32_r_reg_6_ ( .D(N195), .SIN(crc32_r_5_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_6_) );
  SDFFQX1 crc32_r_reg_11_ ( .D(N200), .SIN(crc32_r_10_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_11_) );
  SDFFQX1 crc32_r_reg_15_ ( .D(N204), .SIN(crc32_r_14_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_15_) );
  SDFFQX1 crc32_r_reg_12_ ( .D(N201), .SIN(crc32_r_11_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_12_) );
  SDFFQX1 crc32_r_reg_14_ ( .D(N203), .SIN(crc32_r_13_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_14_) );
  SDFFQX1 crc32_r_reg_18_ ( .D(N207), .SIN(crc32_r_17_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_18_) );
  SDFFQX1 crc32_r_reg_25_ ( .D(N214), .SIN(crc32_r_24_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_25_) );
  SDFFQX1 crc32_r_reg_3_ ( .D(N192), .SIN(crc32_r_2_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_3_) );
  SDFFQX1 crc32_r_reg_24_ ( .D(N213), .SIN(crc32_r_23_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_24_) );
  SDFFQX1 crc32_r_reg_20_ ( .D(N209), .SIN(crc32_r_19_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_20_) );
  SDFFQX1 crc32_r_reg_9_ ( .D(N198), .SIN(crc32_r_8_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_9_) );
  SDFFQX1 crc32_r_reg_21_ ( .D(N210), .SIN(crc32_r_20_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_21_) );
  SDFFQX1 crc32_r_reg_7_ ( .D(N196), .SIN(crc32_r_6_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_7_) );
  SDFFQX1 crc32_r_reg_22_ ( .D(N211), .SIN(crc32_r_21_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_22_) );
  SDFFQX1 crc32_r_reg_2_ ( .D(N191), .SIN(crc32_r_1_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_2_) );
  SDFFQX1 crc32_r_reg_13_ ( .D(N202), .SIN(crc32_r_12_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_13_) );
  SDFFQX1 crc32_r_reg_23_ ( .D(N212), .SIN(crc32_r_22_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_23_) );
  SDFFQX1 crc32_r_reg_28_ ( .D(N217), .SIN(crc32_r_27_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_28_) );
  SDFFQX1 crc32_r_reg_29_ ( .D(N218), .SIN(crc32_r_28_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_29_) );
  SDFFQX1 crc32_r_reg_19_ ( .D(N208), .SIN(crc32_r_18_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_19_) );
  SDFFQX1 crc32_r_reg_31_ ( .D(N220), .SIN(crc32_r_30_), .SMC(test_se), .C(
        net10566), .Q(test_so) );
  SDFFQX1 crc32_r_reg_30_ ( .D(N219), .SIN(crc32_r_29_), .SMC(test_se), .C(
        net10566), .Q(crc32_r_30_) );
  INVX1 U3 ( .A(n18), .Y(n1) );
  XNOR2XL U4 ( .A(i_shfidat[2]), .B(n119), .Y(n56) );
  INVX1 U5 ( .A(n17), .Y(n2) );
  XNOR2XL U6 ( .A(i_shfidat[3]), .B(n120), .Y(n71) );
  INVX1 U7 ( .A(n19), .Y(n3) );
  XNOR2XL U8 ( .A(i_shfidat[1]), .B(n117), .Y(n51) );
  INVX1 U9 ( .A(n15), .Y(n4) );
  XNOR2XL U10 ( .A(i_shfidat[0]), .B(n114), .Y(n62) );
  INVX1 U11 ( .A(n62), .Y(n5) );
  INVX1 U12 ( .A(n62), .Y(n6) );
  AND2X1 U13 ( .A(i_shfo4), .B(n12), .Y(n60) );
  INVX1 U14 ( .A(n60), .Y(n7) );
  INVX1 U15 ( .A(n60), .Y(n8) );
  INVX1 U16 ( .A(n78), .Y(n9) );
  INVX1 U17 ( .A(n78), .Y(n10) );
  INVX1 U18 ( .A(n78), .Y(n16) );
  INVX1 U19 ( .A(n11), .Y(n12) );
  NAND2X1 U20 ( .A(n12), .B(n7), .Y(N188) );
  INVX1 U21 ( .A(n11), .Y(n14) );
  INVX1 U22 ( .A(n11), .Y(n13) );
  NAND2X1 U23 ( .A(i_start), .B(n19), .Y(n49) );
  NAND21X1 U24 ( .B(n81), .A(n80), .Y(n63) );
  OAI21X1 U25 ( .B(n14), .C(n115), .A(n9), .Y(N191) );
  XNOR2XL U26 ( .A(n17), .B(n116), .Y(n115) );
  XNOR2XL U27 ( .A(n18), .B(n19), .Y(n116) );
  INVX1 U28 ( .A(i_start), .Y(n15) );
  NOR2X1 U29 ( .A(i_shfi4), .B(n12), .Y(n78) );
  AND2X1 U30 ( .A(n80), .B(n16), .Y(n48) );
  NOR2X1 U31 ( .A(n12), .B(n4), .Y(n52) );
  OR2X1 U32 ( .A(i_start), .B(i_shfi4), .Y(n11) );
  NAND21X1 U33 ( .B(n12), .A(n81), .Y(n46) );
  OAI21X1 U34 ( .B(n14), .C(n118), .A(n10), .Y(N190) );
  XNOR2XL U35 ( .A(n17), .B(n18), .Y(n118) );
  AOI21X1 U36 ( .B(n18), .C(n4), .A(n78), .Y(n55) );
  AOI21X1 U37 ( .B(n17), .C(n4), .A(n78), .Y(n74) );
  OAI21X1 U38 ( .B(n14), .C(n17), .A(n16), .Y(N189) );
  INVX1 U39 ( .A(n51), .Y(n19) );
  AOI21AX1 U40 ( .B(n15), .C(n51), .A(n49), .Y(n68) );
  NOR2X1 U41 ( .A(n5), .B(i_start), .Y(n81) );
  NAND2X1 U42 ( .A(i_start), .B(n5), .Y(n80) );
  OAI21X1 U43 ( .B(n14), .C(n112), .A(n9), .Y(N192) );
  XNOR2XL U44 ( .A(n18), .B(n113), .Y(n112) );
  XNOR2XL U45 ( .A(n19), .B(n6), .Y(n113) );
  INVX1 U46 ( .A(n56), .Y(n18) );
  INVX1 U47 ( .A(n71), .Y(n17) );
  OAI21BX1 U48 ( .C(n7), .B(n6), .A(N188), .Y(n47) );
  OAI21X1 U49 ( .B(n14), .C(n3), .A(n7), .Y(n53) );
  OAI21X1 U50 ( .B(n14), .C(n56), .A(n7), .Y(n57) );
  OAI21X1 U51 ( .B(n14), .C(n71), .A(n7), .Y(n75) );
  NOR4XL U52 ( .A(n26), .B(n30), .C(n24), .D(n32), .Y(n41) );
  NOR4XL U53 ( .A(n33), .B(n25), .C(n34), .D(n29), .Y(n40) );
  NOR4XL U54 ( .A(n20), .B(n28), .C(n31), .D(n27), .Y(n38) );
  NOR2X1 U55 ( .A(crc32_r_30_), .B(i_start), .Y(n117) );
  OAI221X1 U56 ( .A(n13), .B(n87), .C(n27), .D(n7), .E(n9), .Y(N201) );
  XNOR2XL U57 ( .A(n88), .B(n71), .Y(n87) );
  XNOR2XL U58 ( .A(n89), .B(n18), .Y(n88) );
  AOI22X1 U59 ( .A(n68), .B(n27), .C(n51), .D(crc32_r_8_), .Y(n89) );
  NOR2X1 U60 ( .A(test_so), .B(i_start), .Y(n114) );
  OAI221X1 U61 ( .A(n13), .B(n106), .C(n29), .D(n7), .E(n10), .Y(N194) );
  XNOR2XL U62 ( .A(n107), .B(n71), .Y(n106) );
  XNOR2XL U63 ( .A(n56), .B(n108), .Y(n107) );
  OAI22X1 U64 ( .A(n29), .B(n6), .C(crc32_r_1_), .D(n63), .Y(n108) );
  OAI221X1 U65 ( .A(n13), .B(n98), .C(n20), .D(n7), .E(n16), .Y(N197) );
  XNOR2XL U66 ( .A(n99), .B(n71), .Y(n98) );
  XNOR2XL U67 ( .A(n56), .B(n100), .Y(n99) );
  OAI22X1 U68 ( .A(n20), .B(n6), .C(crc32_r_4_), .D(n63), .Y(n100) );
  OAI221X1 U69 ( .A(n13), .B(n90), .C(n8), .D(n122), .E(n9), .Y(N200) );
  XNOR2XL U70 ( .A(n91), .B(n71), .Y(n90) );
  XNOR2XL U71 ( .A(n56), .B(n92), .Y(n91) );
  OAI22X1 U72 ( .A(n6), .B(n122), .C(crc32_r_7_), .D(n63), .Y(n92) );
  OAI221X1 U73 ( .A(n12), .B(n84), .C(n8), .D(n35), .E(n10), .Y(N202) );
  XNOR2XL U74 ( .A(n85), .B(n56), .Y(n84) );
  XNOR2XL U75 ( .A(n51), .B(n86), .Y(n85) );
  OAI22X1 U76 ( .A(n6), .B(n35), .C(crc32_r_9_), .D(n63), .Y(n86) );
  OAI221X1 U77 ( .A(n13), .B(n101), .C(n21), .D(n7), .E(n16), .Y(N196) );
  XNOR2XL U78 ( .A(n102), .B(n71), .Y(n101) );
  XNOR2XL U79 ( .A(n51), .B(n103), .Y(n102) );
  OAI22X1 U80 ( .A(n21), .B(n5), .C(crc32_r_3_), .D(n63), .Y(n103) );
  OAI221X1 U81 ( .A(n13), .B(n93), .C(n31), .D(n7), .E(n9), .Y(N199) );
  XNOR2XL U82 ( .A(n94), .B(n71), .Y(n93) );
  XNOR2XL U83 ( .A(n51), .B(n95), .Y(n94) );
  OAI22X1 U84 ( .A(n31), .B(n5), .C(crc32_r_6_), .D(n63), .Y(n95) );
  OAI221X1 U85 ( .A(n13), .B(n109), .C(n26), .D(n8), .E(n10), .Y(N193) );
  XNOR2XL U86 ( .A(n110), .B(n71), .Y(n109) );
  XNOR2XL U87 ( .A(n51), .B(n111), .Y(n110) );
  OAI22X1 U88 ( .A(n26), .B(n6), .C(crc32_r_0_), .D(n63), .Y(n111) );
  OAI221X1 U89 ( .A(n12), .B(n64), .C(n8), .D(n58), .E(n16), .Y(N214) );
  XNOR2XL U90 ( .A(n19), .B(n65), .Y(n64) );
  OAI22X1 U91 ( .A(n6), .B(n58), .C(crc32_r_21_), .D(n63), .Y(n65) );
  INVX1 U92 ( .A(crc32_r_21_), .Y(n58) );
  OAI221X1 U93 ( .A(n13), .B(n59), .C(n123), .D(n8), .E(n9), .Y(N215) );
  XNOR2XL U94 ( .A(n17), .B(n61), .Y(n59) );
  OAI22X1 U95 ( .A(n6), .B(n123), .C(crc32_r_22_), .D(n63), .Y(n61) );
  INVX1 U96 ( .A(crc32_r_22_), .Y(n123) );
  OAI221X1 U97 ( .A(n12), .B(n82), .C(n30), .D(n8), .E(n10), .Y(N203) );
  XNOR2XL U98 ( .A(n19), .B(n83), .Y(n82) );
  OAI22X1 U99 ( .A(n30), .B(n6), .C(crc32_r_10_), .D(n63), .Y(n83) );
  OAI221X1 U100 ( .A(n13), .B(n96), .C(n28), .D(n8), .E(n16), .Y(N198) );
  XNOR2XL U101 ( .A(n97), .B(n56), .Y(n96) );
  AOI22X1 U102 ( .A(n68), .B(n28), .C(n51), .D(crc32_r_5_), .Y(n97) );
  OAI221X1 U103 ( .A(n13), .B(n104), .C(n8), .D(n125), .E(n9), .Y(N195) );
  XNOR2XL U104 ( .A(n105), .B(n56), .Y(n104) );
  AOI22X1 U105 ( .A(n68), .B(n125), .C(crc32_r_2_), .D(n51), .Y(n105) );
  INVX1 U106 ( .A(crc32_r_2_), .Y(n125) );
  OAI221X1 U107 ( .A(n12), .B(n66), .C(n8), .D(n121), .E(n10), .Y(N213) );
  XNOR2XL U108 ( .A(n67), .B(n56), .Y(n66) );
  AOI22X1 U109 ( .A(n68), .B(n121), .C(crc32_r_20_), .D(n51), .Y(n67) );
  INVX1 U110 ( .A(crc32_r_20_), .Y(n121) );
  NOR2X1 U111 ( .A(crc32_r_29_), .B(i_start), .Y(n119) );
  NAND2X1 U112 ( .A(n73), .B(n74), .Y(N211) );
  AOI32X1 U113 ( .A(n52), .B(n34), .C(n2), .D(crc32_r_18_), .E(n75), .Y(n73)
         );
  NAND2X1 U114 ( .A(n77), .B(n55), .Y(N206) );
  AOI32X1 U115 ( .A(n52), .B(n124), .C(n1), .D(crc32_r_13_), .E(n57), .Y(n77)
         );
  INVX1 U116 ( .A(crc32_r_13_), .Y(n124) );
  NAND2X1 U117 ( .A(n54), .B(n55), .Y(N216) );
  AOI32X1 U118 ( .A(n52), .B(n126), .C(n1), .D(crc32_r_23_), .E(n57), .Y(n54)
         );
  INVX1 U119 ( .A(crc32_r_23_), .Y(n126) );
  NAND2X1 U120 ( .A(n79), .B(n74), .Y(N205) );
  AOI32X1 U121 ( .A(n52), .B(n32), .C(n2), .D(crc32_r_12_), .E(n75), .Y(n79)
         );
  OAI221X1 U122 ( .A(crc32_r_15_), .B(n46), .C(n25), .D(n47), .E(n48), .Y(N208) );
  OAI221X1 U123 ( .A(crc32_r_25_), .B(n46), .C(n22), .D(n47), .E(n48), .Y(N218) );
  INVX1 U124 ( .A(crc32_r_25_), .Y(n22) );
  OAI221X1 U125 ( .A(crc32_r_11_), .B(n46), .C(n24), .D(n47), .E(n48), .Y(N204) );
  OAI221X1 U126 ( .A(n12), .B(n69), .C(n8), .D(n127), .E(n16), .Y(N212) );
  INVX1 U127 ( .A(crc32_r_19_), .Y(n127) );
  XNOR2XL U128 ( .A(n70), .B(n71), .Y(n69) );
  XNOR2XL U129 ( .A(n72), .B(n56), .Y(n70) );
  NOR2X1 U130 ( .A(crc32_r_28_), .B(i_start), .Y(n120) );
  NAND3X1 U131 ( .A(n49), .B(n10), .C(n50), .Y(N217) );
  AOI32X1 U132 ( .A(n3), .B(n23), .C(n52), .D(crc32_r_24_), .E(n53), .Y(n50)
         );
  INVX1 U133 ( .A(crc32_r_24_), .Y(n23) );
  NAND3X1 U134 ( .A(n49), .B(n16), .C(n76), .Y(N207) );
  AOI32X1 U135 ( .A(n3), .B(n33), .C(n52), .D(crc32_r_14_), .E(n53), .Y(n76)
         );
  OAI21BBX1 U136 ( .A(N188), .B(crc32_r_26_), .C(n15), .Y(N219) );
  OAI21BBX1 U137 ( .A(N188), .B(crc32_r_27_), .C(n15), .Y(N220) );
  OAI21BBX1 U138 ( .A(N188), .B(crc32_r_16_), .C(n15), .Y(N209) );
  OAI21BBX1 U139 ( .A(N188), .B(crc32_r_17_), .C(n15), .Y(N210) );
  NOR2X1 U140 ( .A(crc32_r_19_), .B(i_start), .Y(n72) );
  INVX1 U141 ( .A(crc32_r_28_), .Y(crc32_3_0[3]) );
  INVX1 U142 ( .A(crc32_r_29_), .Y(crc32_3_0[2]) );
  AND4X1 U143 ( .A(crc32_r_24_), .B(crc32_r_25_), .C(crc32_r_26_), .D(
        crc32_r_3_), .Y(n39) );
  NOR2X1 U144 ( .A(n36), .B(n37), .Y(rx_good) );
  NAND4X1 U145 ( .A(n42), .B(n43), .C(n44), .D(n45), .Y(n36) );
  NAND4X1 U146 ( .A(n38), .B(n39), .C(n40), .D(n41), .Y(n37) );
  NOR4XL U147 ( .A(crc32_r_21_), .B(crc32_r_20_), .C(crc32_r_19_), .D(
        crc32_r_17_), .Y(n43) );
  NOR4XL U148 ( .A(crc32_r_9_), .B(crc32_r_7_), .C(crc32_r_2_), .D(crc32_r_29_), .Y(n45) );
  NOR4XL U149 ( .A(crc32_r_28_), .B(crc32_r_27_), .C(crc32_r_23_), .D(
        crc32_r_22_), .Y(n44) );
  NOR4XL U150 ( .A(crc32_r_16_), .B(crc32_r_13_), .C(crc32_3_0[1]), .D(
        crc32_3_0[0]), .Y(n42) );
  INVX1 U151 ( .A(crc32_r_30_), .Y(crc32_3_0[1]) );
  INVX1 U152 ( .A(test_so), .Y(crc32_3_0[0]) );
  INVX1 U153 ( .A(crc32_r_6_), .Y(n31) );
  INVX1 U154 ( .A(crc32_r_1_), .Y(n29) );
  INVX1 U155 ( .A(crc32_r_10_), .Y(n30) );
  INVX1 U156 ( .A(crc32_r_4_), .Y(n20) );
  INVX1 U157 ( .A(crc32_r_0_), .Y(n26) );
  INVX1 U158 ( .A(crc32_r_8_), .Y(n27) );
  INVX1 U159 ( .A(crc32_r_5_), .Y(n28) );
  INVX1 U160 ( .A(crc32_r_18_), .Y(n34) );
  INVX1 U161 ( .A(crc32_r_12_), .Y(n32) );
  INVX1 U162 ( .A(crc32_r_14_), .Y(n33) );
  INVX1 U163 ( .A(crc32_r_11_), .Y(n24) );
  INVX1 U164 ( .A(crc32_r_15_), .Y(n25) );
  INVX1 U165 ( .A(crc32_r_7_), .Y(n122) );
  INVX1 U166 ( .A(crc32_r_9_), .Y(n35) );
  INVX1 U167 ( .A(crc32_r_3_), .Y(n21) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phycrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phytx_a0 ( r_txnumk, r_txendk, r_txshrt, r_txauto, prx_cccnt, ptx_txact, 
        ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, i_rdat, i_txreq, i_one, 
        ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4, ptx_crcsidat, ptx_fsm, 
        pcc_crc30, clk, srstz, test_si, test_se );
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [1:0] prx_cccnt;
  input [7:0] i_rdat;
  output [3:0] ptx_crcsidat;
  output [2:0] ptx_fsm;
  input [3:0] pcc_crc30;
  input r_txendk, r_txshrt, i_txreq, i_one, clk, srstz, test_si, test_se;
  output ptx_txact, ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, ptx_crcstart,
         ptx_crcshfi4, ptx_crcshfo4;
  wire   hinib, N251, N254, N255, N264, N265, N266, N268, N269, N270, N271,
         N272, N273, N297, N298, N299, net10588, net10594, n237, n238, n69,
         n70, n95, n96, n102, n113, n114, n116, n119, n120, n136, n137, n138,
         n139, n140, n152, n153, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n97, n98, n99, n100,
         n101, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n115, n117, n118, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267;
  wire   [4:0] bytcnt;
  wire   [3:0] bitcnt;
  wire   [4:2] add_104_carry;

  HAD1X1 add_104_U1_1_2 ( .A(bytcnt[2]), .B(add_104_carry[2]), .CO(
        add_104_carry[3]), .SO(N265) );
  HAD1X1 add_104_U1_1_3 ( .A(bytcnt[3]), .B(add_104_carry[3]), .CO(
        add_104_carry[4]), .SO(N266) );
  SNPS_CLOCK_GATE_HIGH_phytx_a0_0 clk_gate_bitcnt_reg ( .CLK(clk), .EN(N251), 
        .ENCLK(net10588), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phytx_a0_1 clk_gate_bytcnt_reg ( .CLK(clk), .EN(N268), 
        .ENCLK(net10594), .TE(test_se) );
  SDFFQX1 ptx_cc_reg ( .D(n238), .SIN(n2), .SMC(test_se), .C(clk), .Q(ptx_cc)
         );
  SDFFQX1 bitcnt_reg_3_ ( .D(N255), .SIN(bitcnt[2]), .SMC(test_se), .C(
        net10588), .Q(bitcnt[3]) );
  SDFFQX1 bitcnt_reg_0_ ( .D(n254), .SIN(test_si), .SMC(test_se), .C(net10588), 
        .Q(bitcnt[0]) );
  SDFFQX1 bitcnt_reg_2_ ( .D(N254), .SIN(bitcnt[1]), .SMC(test_se), .C(
        net10588), .Q(bitcnt[2]) );
  SDFFQX1 bitcnt_reg_1_ ( .D(n256), .SIN(bitcnt[0]), .SMC(test_se), .C(
        net10588), .Q(bitcnt[1]) );
  SDFFQX1 bytcnt_reg_4_ ( .D(N273), .SIN(bytcnt[3]), .SMC(test_se), .C(
        net10594), .Q(bytcnt[4]) );
  SDFFQX1 cs_txph_reg_1_ ( .D(N298), .SIN(ptx_fsm[0]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[1]) );
  SDFFQX1 cs_txph_reg_0_ ( .D(N297), .SIN(bytcnt[4]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[0]) );
  SDFFQX1 cs_txph_reg_2_ ( .D(N299), .SIN(ptx_fsm[1]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[2]) );
  SDFFQX1 bytcnt_reg_2_ ( .D(N271), .SIN(bytcnt[1]), .SMC(test_se), .C(
        net10594), .Q(bytcnt[2]) );
  SDFFQX1 bytcnt_reg_1_ ( .D(N270), .SIN(n3), .SMC(test_se), .C(net10594), .Q(
        bytcnt[1]) );
  SDFFQX1 bytcnt_reg_3_ ( .D(N272), .SIN(bytcnt[2]), .SMC(test_se), .C(
        net10594), .Q(bytcnt[3]) );
  SDFFQX1 hinib_reg ( .D(n237), .SIN(ptx_fsm[2]), .SMC(test_se), .C(net10588), 
        .Q(hinib) );
  SDFFQX1 bytcnt_reg_0_ ( .D(N269), .SIN(bitcnt[3]), .SMC(test_se), .C(
        net10594), .Q(bytcnt[0]) );
  HAD1XL add_104_U1_1_1 ( .A(bytcnt[1]), .B(bytcnt[0]), .CO(add_104_carry[2]), 
        .SO(N264) );
  NAND21X1 U3 ( .B(n27), .A(n26), .Y(n31) );
  NOR21XL U4 ( .B(r_txnumk[3]), .A(bytcnt[3]), .Y(n24) );
  GEN2XL U5 ( .D(n205), .E(n216), .C(n170), .B(n159), .A(n158), .Y(n162) );
  INVX1 U6 ( .A(n115), .Y(n63) );
  INVX1 U7 ( .A(n235), .Y(n200) );
  NAND21X1 U8 ( .B(n161), .A(n39), .Y(n191) );
  XOR2X1 U9 ( .A(n191), .B(bitcnt[1]), .Y(n235) );
  AOI21X1 U10 ( .B(n161), .C(n72), .A(n89), .Y(n1) );
  INVX1 U11 ( .A(n211), .Y(n2) );
  MUX2X1 U12 ( .D0(n133), .D1(n44), .S(hinib), .Y(n134) );
  MUX2BXL U13 ( .D0(n157), .D1(i_rdat[7]), .S(hinib), .Y(n160) );
  INVX1 U14 ( .A(n54), .Y(n3) );
  OAI22X1 U15 ( .A(bytcnt[1]), .B(n28), .C(bytcnt[0]), .D(n29), .Y(n22) );
  NAND5XL U16 ( .A(bytcnt[0]), .B(n63), .C(n62), .D(n61), .E(n60), .Y(n74) );
  INVX1 U17 ( .A(r_txnumk[0]), .Y(n29) );
  NAND3X1 U18 ( .A(n56), .B(n55), .C(n22), .Y(n23) );
  INVX1 U19 ( .A(i_one), .Y(n80) );
  MUX2IXL U20 ( .D0(i_rdat[7]), .D1(i_rdat[5]), .S(n221), .Y(n11) );
  INVXL U21 ( .A(n78), .Y(n232) );
  NAND32XL U22 ( .B(n77), .C(n78), .A(n112), .Y(n50) );
  NAND21XL U23 ( .B(n80), .A(n123), .Y(n97) );
  NAND21XL U24 ( .B(n233), .A(n115), .Y(n53) );
  NAND21X1 U25 ( .B(n170), .A(n38), .Y(n39) );
  AOI31XL U26 ( .A(n47), .B(n46), .C(n76), .D(n125), .Y(n49) );
  NAND42XL U27 ( .C(n29), .D(n28), .A(r_txnumk[2]), .B(r_txnumk[3]), .Y(n30)
         );
  AND2XL U28 ( .A(r_txnumk[2]), .B(n62), .Y(n25) );
  OA22XL U29 ( .A(r_txnumk[0]), .B(n54), .C(r_txnumk[4]), .D(n60), .Y(n58) );
  INVXL U30 ( .A(n52), .Y(n233) );
  NAND2XL U31 ( .A(i_rdat[6]), .B(n201), .Y(n10) );
  NAND21XL U32 ( .B(n77), .A(n106), .Y(n84) );
  GEN2XL U33 ( .D(n138), .E(n259), .C(n209), .B(n213), .A(n154), .Y(n163) );
  INVXL U34 ( .A(n106), .Y(n98) );
  MUX2AXL U35 ( .D0(n4), .D1(n222), .S(n18), .Y(n223) );
  AOI21X1 U36 ( .B(n221), .C(n220), .A(n219), .Y(n4) );
  OA21XL U37 ( .B(n198), .C(n173), .A(n172), .Y(n174) );
  NAND32XL U38 ( .B(n126), .C(n125), .A(n130), .Y(n218) );
  NAND21XL U39 ( .B(n52), .A(n164), .Y(n43) );
  INVXL U40 ( .A(n126), .Y(ptx_crcsidat[0]) );
  OAI211XL U41 ( .C(n198), .D(n184), .A(n183), .B(n182), .Y(n189) );
  NAND21XL U42 ( .B(r_txnumk[2]), .A(bytcnt[2]), .Y(n55) );
  NAND32X1 U43 ( .B(n25), .C(n24), .A(n23), .Y(n26) );
  OAI211XL U44 ( .C(n123), .D(n122), .A(n255), .B(n121), .Y(n153) );
  NOR2XL U45 ( .A(n3), .B(n153), .Y(N269) );
  AND3XL U46 ( .A(n112), .B(n233), .C(n232), .Y(n242) );
  AOI211XL U47 ( .C(n14), .D(n240), .A(n239), .B(i_txreq), .Y(n241) );
  AOI31XL U48 ( .A(n119), .B(n261), .C(n95), .D(bytcnt[0]), .Y(n114) );
  NAND21XL U49 ( .B(n95), .A(bytcnt[0]), .Y(n132) );
  OAI211XL U50 ( .C(hinib), .D(bytcnt[0]), .A(n138), .B(n148), .Y(n166) );
  AOI22XL U51 ( .A(n120), .B(bytcnt[0]), .C(n113), .D(n138), .Y(n137) );
  INVXL U52 ( .A(bytcnt[0]), .Y(n54) );
  NAND2XL U53 ( .A(bytcnt[0]), .B(hinib), .Y(n138) );
  INVX1 U54 ( .A(n21), .Y(n20) );
  INVX1 U55 ( .A(n249), .Y(n253) );
  NAND21X1 U56 ( .B(n253), .A(n51), .Y(N251) );
  INVX1 U57 ( .A(n141), .Y(n169) );
  INVX1 U58 ( .A(n181), .Y(n151) );
  INVX1 U59 ( .A(n178), .Y(n180) );
  INVX1 U60 ( .A(srstz), .Y(n21) );
  INVX1 U61 ( .A(n79), .Y(n123) );
  NAND21X1 U62 ( .B(n232), .A(n90), .Y(n79) );
  INVX1 U63 ( .A(i_txreq), .Y(n112) );
  INVX1 U64 ( .A(n243), .Y(n107) );
  NAND21X1 U65 ( .B(n230), .A(n51), .Y(n249) );
  INVX1 U66 ( .A(n50), .Y(n51) );
  AND2X1 U67 ( .A(n243), .B(n20), .Y(N297) );
  AND2X1 U68 ( .A(n244), .B(n20), .Y(N298) );
  AND2X1 U69 ( .A(n135), .B(n53), .Y(ptx_crcshfo4) );
  NAND21X1 U70 ( .B(n141), .A(n187), .Y(n181) );
  NAND21X1 U71 ( .B(n206), .A(n215), .Y(n141) );
  NAND21X1 U72 ( .B(n202), .A(n203), .Y(n178) );
  NAND21X1 U73 ( .B(n207), .A(n215), .Y(n204) );
  MUX2X1 U74 ( .D0(n171), .D1(n178), .S(n208), .Y(n172) );
  AND2X1 U75 ( .A(n181), .B(n204), .Y(n171) );
  AO21X1 U76 ( .B(n203), .C(n207), .A(n181), .Y(n182) );
  INVX1 U77 ( .A(n128), .Y(n215) );
  NAND32XL U78 ( .B(n127), .C(n191), .A(n176), .Y(n128) );
  OAI22X1 U79 ( .A(n205), .B(n204), .C(n203), .D(n202), .Y(n217) );
  AND2X1 U80 ( .A(n151), .B(n155), .Y(n154) );
  INVX1 U81 ( .A(n124), .Y(n130) );
  NAND21XL U82 ( .B(n161), .A(n191), .Y(n124) );
  AND2X1 U83 ( .A(n245), .B(n20), .Y(N299) );
  NOR21XL U84 ( .B(n138), .A(n116), .Y(n146) );
  INVX1 U85 ( .A(n198), .Y(n225) );
  AO21X1 U86 ( .B(n208), .C(n207), .A(n206), .Y(n214) );
  INVX1 U87 ( .A(n155), .Y(n205) );
  INVX1 U88 ( .A(n139), .Y(n260) );
  INVX1 U89 ( .A(n120), .Y(n261) );
  NAND21X1 U90 ( .B(n203), .A(n208), .Y(n185) );
  INVX1 U91 ( .A(n116), .Y(n263) );
  INVX1 U92 ( .A(n96), .Y(n259) );
  NOR43XL U93 ( .B(n95), .C(n119), .D(n139), .A(n6), .Y(n5) );
  OR3XL U94 ( .A(n259), .B(n113), .C(n263), .Y(n6) );
  INVX1 U95 ( .A(n117), .Y(n135) );
  AOI21BX1 U96 ( .C(n138), .B(n259), .A(n113), .Y(n165) );
  INVX1 U97 ( .A(n176), .Y(n213) );
  INVX1 U98 ( .A(n245), .Y(n105) );
  NAND21X1 U99 ( .B(n125), .A(n37), .Y(n38) );
  NAND21X1 U100 ( .B(ptx_crcsidat[1]), .A(n35), .Y(n37) );
  MUX2IX1 U101 ( .D0(n34), .D1(ptx_crcsidat[2]), .S(ptx_crcsidat[3]), .Y(n35)
         );
  INVX1 U102 ( .A(n134), .Y(ptx_crcsidat[2]) );
  NAND21X1 U103 ( .B(n134), .A(n126), .Y(n34) );
  NAND32X1 U104 ( .B(n230), .C(n234), .A(n14), .Y(n115) );
  NAND32X1 U105 ( .B(n248), .C(n48), .A(n200), .Y(n234) );
  OAI31XL U106 ( .A(n49), .B(n170), .C(n52), .D(n115), .Y(n78) );
  NAND21X1 U107 ( .B(n123), .A(n106), .Y(ptx_fifopop) );
  INVX1 U108 ( .A(n160), .Y(ptx_crcsidat[3]) );
  INVX1 U109 ( .A(i_rdat[6]), .Y(n44) );
  INVX1 U110 ( .A(n129), .Y(ptx_crcsidat[1]) );
  INVX1 U111 ( .A(i_rdat[4]), .Y(n46) );
  INVX1 U112 ( .A(i_rdat[5]), .Y(n47) );
  INVX1 U113 ( .A(r_txnumk[1]), .Y(n28) );
  INVX1 U114 ( .A(r_txauto[6]), .Y(n125) );
  INVX1 U115 ( .A(n118), .Y(n161) );
  INVX1 U116 ( .A(n45), .Y(n76) );
  NAND21X1 U117 ( .B(i_rdat[7]), .A(n44), .Y(n45) );
  NAND21X1 U118 ( .B(n93), .A(prx_cccnt[0]), .Y(n230) );
  INVX1 U119 ( .A(ptx_txact), .Y(n93) );
  NAND32X1 U120 ( .B(n101), .C(n88), .A(n82), .Y(n176) );
  INVX1 U121 ( .A(n104), .Y(n90) );
  OAI221X1 U122 ( .A(n1), .B(n88), .C(n118), .D(n5), .E(n87), .Y(n243) );
  AOI211X1 U123 ( .C(n257), .D(n86), .A(n85), .B(n84), .Y(n87) );
  INVX1 U124 ( .A(r_txauto[5]), .Y(n257) );
  OAI22X1 U125 ( .A(n117), .B(n91), .C(r_txauto[4]), .D(n97), .Y(n86) );
  NOR21XL U126 ( .B(N264), .A(n153), .Y(N270) );
  NOR21XL U127 ( .B(N266), .A(n153), .Y(N272) );
  NOR21XL U128 ( .B(N265), .A(n153), .Y(N271) );
  AOI211X1 U129 ( .C(n5), .D(n258), .A(ptx_txact), .B(n112), .Y(n85) );
  NAND2X1 U130 ( .A(n255), .B(n153), .Y(N268) );
  AO21X1 U131 ( .B(n266), .C(n253), .A(n254), .Y(n251) );
  OAI211X1 U132 ( .C(n103), .D(n101), .A(n100), .B(n99), .Y(n244) );
  AOI221XL U133 ( .A(n135), .B(n91), .C(n90), .D(n97), .E(n89), .Y(n103) );
  OA22X1 U134 ( .A(n98), .B(n176), .C(n97), .D(n94), .Y(n99) );
  AOI32X1 U135 ( .A(n258), .B(i_txreq), .C(n93), .D(n161), .E(n92), .Y(n100)
         );
  INVX1 U136 ( .A(n247), .Y(n254) );
  OAI32X1 U137 ( .A(n249), .B(n248), .C(bitcnt[1]), .D(n266), .E(n247), .Y(
        n256) );
  INVX1 U138 ( .A(n246), .Y(n250) );
  NAND32X1 U139 ( .B(n266), .C(n248), .A(n253), .Y(n246) );
  AND4XL U140 ( .A(n170), .B(n59), .C(n58), .D(n57), .Y(ptx_crcstart) );
  AND3XL U141 ( .A(n90), .B(n170), .C(n53), .Y(ptx_crcshfi4) );
  AND4X1 U142 ( .A(n233), .B(n90), .C(n56), .D(n55), .Y(n57) );
  NAND21X1 U143 ( .B(n66), .A(n67), .Y(n91) );
  OAI211X1 U144 ( .C(n83), .D(n82), .A(n81), .B(n97), .Y(n245) );
  INVX1 U145 ( .A(n84), .Y(n81) );
  AND2X1 U146 ( .A(n1), .B(n117), .Y(n83) );
  INVX1 U147 ( .A(n218), .Y(n219) );
  AO2222XL U148 ( .A(n217), .B(n216), .C(n215), .D(n214), .E(i_rdat[4]), .F(
        n225), .G(n213), .H(n212), .Y(n220) );
  OR4X1 U149 ( .A(n164), .B(n163), .C(n162), .D(n222), .Y(n196) );
  NAND43X1 U150 ( .B(n190), .C(n222), .D(n189), .A(n188), .Y(n194) );
  GEN2XL U151 ( .D(n187), .E(n203), .C(n186), .B(n185), .A(n204), .Y(n188) );
  AND3X1 U152 ( .A(n180), .B(n216), .C(n179), .Y(n190) );
  MUX2IX1 U153 ( .D0(n7), .D1(n8), .S(n9), .Y(n228) );
  AOI21X1 U154 ( .B(n225), .C(n224), .A(n223), .Y(n7) );
  MUX4IX1 U155 ( .D0(n197), .D1(n196), .D2(n195), .D3(n194), .S0(n18), .S1(
        n193), .Y(n8) );
  XNOR2XL U156 ( .A(n252), .B(n227), .Y(n9) );
  MUX2IX1 U157 ( .D0(n10), .D1(n11), .S(n18), .Y(n224) );
  NAND21XL U158 ( .B(n170), .A(n169), .Y(n202) );
  INVX1 U159 ( .A(n201), .Y(n221) );
  INVX1 U160 ( .A(n71), .Y(n89) );
  NAND43X1 U161 ( .B(n90), .C(n161), .D(ptx_goidle), .A(n68), .Y(n71) );
  AOI31X1 U162 ( .A(n213), .B(n67), .C(n66), .D(n135), .Y(n68) );
  INVX1 U163 ( .A(n74), .Y(n67) );
  INVX1 U164 ( .A(n92), .Y(n72) );
  OAI22X1 U165 ( .A(n198), .B(n157), .C(n204), .D(n216), .Y(n158) );
  AND2X1 U166 ( .A(n169), .B(n156), .Y(n159) );
  OAI211X1 U167 ( .C(n177), .D(n176), .A(n175), .B(n174), .Y(n195) );
  AND3X1 U168 ( .A(n167), .B(n166), .C(n165), .Y(n177) );
  INVX1 U169 ( .A(n168), .Y(n175) );
  NAND21X1 U170 ( .B(r_txauto[6]), .A(n130), .Y(n198) );
  NAND31X1 U171 ( .C(n161), .A(n12), .B(n218), .Y(n222) );
  NAND3XL U172 ( .A(r_txauto[6]), .B(n160), .C(n191), .Y(n12) );
  INVX1 U173 ( .A(n43), .Y(n77) );
  NAND3X1 U174 ( .A(r_txauto[2]), .B(r_txauto[1]), .C(r_txauto[0]), .Y(n116)
         );
  NAND32X1 U175 ( .B(n168), .C(n145), .A(n144), .Y(n197) );
  OAI221X1 U176 ( .A(n204), .B(n156), .C(n198), .D(n133), .E(n183), .Y(n145)
         );
  AOI32X1 U177 ( .A(n151), .B(n207), .C(n179), .D(n169), .E(n143), .Y(n144) );
  MUX2X1 U178 ( .D0(n203), .D1(n142), .S(n208), .Y(n143) );
  INVXL U179 ( .A(n170), .Y(n207) );
  INVX1 U180 ( .A(n186), .Y(n206) );
  AND2XL U181 ( .A(n216), .B(n170), .Y(n142) );
  NAND32X1 U182 ( .B(r_txauto[0]), .C(r_txauto[1]), .A(r_txauto[2]), .Y(n119)
         );
  NAND21X1 U183 ( .B(n208), .A(n156), .Y(n155) );
  NAND21X1 U184 ( .B(n164), .A(n218), .Y(n168) );
  AO21X1 U185 ( .B(n266), .C(n248), .A(n226), .Y(n227) );
  NOR3XL U186 ( .A(n264), .B(r_txauto[0]), .C(n262), .Y(n113) );
  INVX1 U187 ( .A(n179), .Y(n208) );
  INVX1 U188 ( .A(n156), .Y(n203) );
  INVX1 U189 ( .A(r_txauto[2]), .Y(n262) );
  NAND2X1 U190 ( .A(r_txauto[1]), .B(n262), .Y(n139) );
  NOR2X1 U191 ( .A(n139), .B(r_txauto[0]), .Y(n120) );
  INVX1 U192 ( .A(r_txauto[1]), .Y(n264) );
  INVX1 U193 ( .A(n216), .Y(n187) );
  NAND3X1 U194 ( .A(r_txauto[2]), .B(n264), .C(r_txauto[0]), .Y(n95) );
  AND2X1 U195 ( .A(n260), .B(r_txauto[0]), .Y(n147) );
  NAND3X1 U196 ( .A(n264), .B(n262), .C(r_txauto[0]), .Y(n96) );
  NAND32X1 U197 ( .B(n101), .C(n82), .A(n88), .Y(n117) );
  INVX1 U198 ( .A(n138), .Y(n267) );
  INVX1 U199 ( .A(n64), .Y(n127) );
  INVX1 U200 ( .A(r_txauto[4]), .Y(n94) );
  INVX1 U201 ( .A(r_txauto[3]), .Y(n258) );
  AND4X1 U202 ( .A(n105), .B(n107), .C(n244), .D(n104), .Y(ptx_pspyld) );
  MUX2X1 U203 ( .D0(n184), .D1(n47), .S(hinib), .Y(n129) );
  EORX1 U204 ( .A(n13), .B(r_txnumk[4]), .C(bytcnt[4]), .D(n31), .Y(n32) );
  NAND3X1 U205 ( .A(bytcnt[4]), .B(n31), .C(n30), .Y(n13) );
  MUX2X1 U206 ( .D0(n173), .D1(n46), .S(hinib), .Y(n126) );
  XOR2XL U207 ( .A(n191), .B(bitcnt[0]), .Y(n236) );
  NAND21X1 U208 ( .B(r_txnumk[1]), .A(bytcnt[1]), .Y(n56) );
  NAND21X1 U209 ( .B(r_txnumk[3]), .A(bytcnt[3]), .Y(n59) );
  NAND6XL U210 ( .A(n184), .B(n133), .C(n157), .D(n76), .E(n173), .F(n75), .Y(
        n106) );
  NOR6XL U211 ( .A(i_rdat[5]), .B(i_rdat[4]), .C(bytcnt[1]), .D(n176), .E(n74), 
        .F(n73), .Y(n75) );
  NAND5XL U212 ( .A(bitcnt[2]), .B(n41), .C(n200), .D(n40), .E(n48), .Y(n52)
         );
  INVX1 U213 ( .A(n230), .Y(n41) );
  INVX1 U214 ( .A(n236), .Y(n40) );
  INVX1 U215 ( .A(bytcnt[3]), .Y(n61) );
  INVX1 U216 ( .A(n59), .Y(n27) );
  NAND21X1 U217 ( .B(n80), .A(r_txendk), .Y(n73) );
  XNOR2XL U218 ( .A(n191), .B(bitcnt[2]), .Y(n14) );
  INVX1 U219 ( .A(i_rdat[1]), .Y(n184) );
  INVX1 U220 ( .A(i_rdat[0]), .Y(n173) );
  INVX1 U221 ( .A(i_rdat[3]), .Y(n157) );
  INVX1 U222 ( .A(i_rdat[2]), .Y(n133) );
  INVX1 U223 ( .A(bytcnt[2]), .Y(n62) );
  NAND32X1 U224 ( .B(ptx_fsm[2]), .C(n88), .A(n101), .Y(n118) );
  NAND32X1 U225 ( .B(ptx_fsm[2]), .C(n101), .A(n88), .Y(n104) );
  INVX1 U226 ( .A(ptx_fsm[0]), .Y(n88) );
  INVX1 U227 ( .A(ptx_fsm[1]), .Y(n101) );
  NAND32X1 U228 ( .B(ptx_fsm[1]), .C(ptx_fsm[2]), .A(n88), .Y(ptx_txact) );
  INVX1 U229 ( .A(bitcnt[0]), .Y(n248) );
  INVX1 U230 ( .A(bitcnt[3]), .Y(n48) );
  INVX1 U231 ( .A(bytcnt[4]), .Y(n60) );
  INVX1 U232 ( .A(ptx_fsm[2]), .Y(n82) );
  NAND5XL U233 ( .A(bytcnt[4]), .B(bytcnt[2]), .C(bytcnt[3]), .D(bytcnt[0]), 
        .E(bytcnt[1]), .Y(n121) );
  AOI31XL U234 ( .A(n176), .B(n118), .C(n117), .D(n115), .Y(n122) );
  NOR21XL U235 ( .B(n112), .A(n111), .Y(n255) );
  NAND31X1 U236 ( .C(n110), .A(n109), .B(n108), .Y(n111) );
  NOR21XL U237 ( .B(n245), .A(ptx_fsm[2]), .Y(n110) );
  XNOR2XL U238 ( .A(ptx_fsm[1]), .B(n244), .Y(n109) );
  XOR2X1 U239 ( .A(ptx_fsm[0]), .B(n107), .Y(n108) );
  NOR2X1 U240 ( .A(n152), .B(n153), .Y(N273) );
  XNOR2XL U241 ( .A(bytcnt[4]), .B(add_104_carry[4]), .Y(n152) );
  NAND21X1 U242 ( .B(bitcnt[0]), .A(n253), .Y(n247) );
  MUX2IX1 U243 ( .D0(n15), .D1(n16), .S(bitcnt[3]), .Y(N255) );
  NAND2X1 U244 ( .A(n250), .B(bitcnt[2]), .Y(n15) );
  AOI21X1 U245 ( .B(n253), .C(n252), .A(n251), .Y(n16) );
  MUX2X1 U246 ( .D0(n250), .D1(n251), .S(bitcnt[2]), .Y(N254) );
  OAI21X1 U247 ( .B(n265), .C(n69), .A(n70), .Y(n238) );
  OAI21X1 U248 ( .B(n21), .C(n265), .A(n69), .Y(n70) );
  NAND32X1 U249 ( .B(n21), .C(i_txreq), .A(n231), .Y(n69) );
  INVX1 U250 ( .A(ptx_cc), .Y(n265) );
  MUX2X1 U251 ( .D0(n242), .D1(n2), .S(n241), .Y(n237) );
  INVXL U252 ( .A(n234), .Y(n240) );
  MUX2BXL U253 ( .D0(bitcnt[1]), .D1(n17), .S(n2), .Y(n201) );
  XNOR2XL U254 ( .A(n200), .B(n199), .Y(n17) );
  OAI21BBXL U255 ( .A(r_txshrt), .B(n63), .C(n91), .Y(n92) );
  AND2X1 U256 ( .A(n192), .B(bitcnt[0]), .Y(n199) );
  INVXL U257 ( .A(n191), .Y(n192) );
  MUX2BXL U258 ( .D0(n230), .D1(n229), .S(prx_cccnt[1]), .Y(n231) );
  AND2X1 U259 ( .A(n228), .B(ptx_txact), .Y(n229) );
  NAND43X1 U260 ( .B(n114), .C(n150), .D(n149), .A(n166), .Y(n209) );
  AND2X1 U261 ( .A(n113), .B(n267), .Y(n149) );
  MUX2X1 U262 ( .D0(n147), .D1(n146), .S(hinib), .Y(n150) );
  MUX2BXL U263 ( .D0(n160), .D1(pcc_crc30[3]), .S(n135), .Y(n186) );
  XNOR2XL U264 ( .A(n226), .B(bitcnt[0]), .Y(n18) );
  MUX2BXL U265 ( .D0(n266), .D1(n19), .S(n2), .Y(n193) );
  XNOR2XL U266 ( .A(n235), .B(n199), .Y(n19) );
  NAND21XL U267 ( .B(n191), .A(hinib), .Y(n226) );
  OAI211X1 U268 ( .C(n95), .D(n211), .A(n96), .B(n210), .Y(n212) );
  INVX1 U269 ( .A(hinib), .Y(n211) );
  INVX1 U270 ( .A(n209), .Y(n210) );
  MUX2X1 U271 ( .D0(ptx_crcsidat[0]), .D1(pcc_crc30[0]), .S(n135), .Y(n179) );
  MUX2BXL U272 ( .D0(n129), .D1(pcc_crc30[1]), .S(n135), .Y(n156) );
  MUX2BXL U273 ( .D0(n134), .D1(pcc_crc30[2]), .S(n135), .Y(n216) );
  GEN2XL U274 ( .D(n132), .E(n116), .C(n2), .B(n131), .A(n176), .Y(n183) );
  AND2X1 U275 ( .A(n136), .B(n137), .Y(n131) );
  AOI31X1 U276 ( .A(r_txauto[0]), .B(hinib), .C(n260), .D(n140), .Y(n136) );
  AOI21X1 U277 ( .B(n116), .C(n119), .A(n138), .Y(n140) );
  INVX1 U278 ( .A(n119), .Y(n148) );
  MUX2X1 U279 ( .D0(n116), .D1(n95), .S(n2), .Y(n167) );
  NOR5XL U280 ( .A(n102), .B(bitcnt[3]), .C(n236), .D(n252), .E(n235), .Y(n239) );
  NOR2X1 U281 ( .A(ptx_fsm[1]), .B(ptx_fsm[0]), .Y(n102) );
  INVX1 U282 ( .A(n65), .Y(ptx_goidle) );
  NAND43X1 U283 ( .B(ptx_cc), .C(n64), .D(n230), .A(ptx_fsm[0]), .Y(n65) );
  NAND21X1 U284 ( .B(ptx_fsm[1]), .A(ptx_fsm[2]), .Y(n64) );
  INVX1 U285 ( .A(n42), .Y(n164) );
  NAND21X1 U286 ( .B(ptx_fsm[0]), .A(n127), .Y(n42) );
  INVX1 U287 ( .A(bitcnt[1]), .Y(n266) );
  INVX1 U288 ( .A(bytcnt[1]), .Y(n66) );
  INVX1 U289 ( .A(bitcnt[2]), .Y(n252) );
  AO21X4 U290 ( .B(n32), .C(n73), .A(n104), .Y(n170) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyidd_a0 ( i_trans, i_goidle, o_ccidle, o_goidle, o_gobusy, clk, srstz, 
        test_si, test_so, test_se );
  input i_trans, i_goidle, clk, srstz, test_si, test_se;
  output o_ccidle, o_goidle, o_gobusy, test_so;
  wire   n30, ttranwin_6_, ttranwin_5_, ttranwin_4_, ttranwin_3_, ttranwin_2_,
         ttranwin_1_, ttranwin_0_, N11, N12, N13, N14, N15, N16, N17, N18, N46,
         N47, N48, N49, N50, N51, N52, N53, N55, N56, N57, N58, N59, N60, N61,
         N62, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, net10611, net10617, net10622, n55, n56,
         n57, n18, n19, n20, n21, n22, n23, n24, n25, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n58, n2, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n26, n27, n28, n29;
  wire   [1:0] ntrancnt;
  wire   [7:0] trans0;
  wire   [7:0] ttranwin_minus;
  wire   [7:0] trans1;

  SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 clk_gate_trans1_reg ( .CLK(clk), .EN(N90), 
        .ENCLK(net10611), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 clk_gate_trans0_reg ( .CLK(clk), .EN(N91), 
        .ENCLK(net10617), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 clk_gate_ttranwin_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net10622), .TE(test_se) );
  phyidd_a0_DW01_sub_0 sub_47 ( .A(trans1), .B(trans0), .CI(1'b0), .DIFF({N53, 
        N52, N51, N50, N49, N48, N47, N46}), .CO() );
  phyidd_a0_DW01_sub_1 sub_24 ( .A({n25, n24, n23, n22, n21, n20, n19, n18}), 
        .B(trans0), .CI(1'b0), .DIFF(ttranwin_minus), .CO() );
  phyidd_a0_DW01_inc_0 add_23 ( .A({test_so, ttranwin_6_, ttranwin_5_, 
        ttranwin_4_, ttranwin_3_, ttranwin_2_, ttranwin_1_, ttranwin_0_}), 
        .SUM({N18, N17, N16, N15, N14, N13, N12, N11}) );
  SDFFQX1 trans1_reg_7_ ( .D(N80), .SIN(trans1[6]), .SMC(test_se), .C(net10611), .Q(trans1[7]) );
  SDFFQX1 trans0_reg_7_ ( .D(N62), .SIN(trans0[6]), .SMC(test_se), .C(net10617), .Q(trans0[7]) );
  SDFFQX1 trans1_reg_6_ ( .D(N79), .SIN(trans1[5]), .SMC(test_se), .C(net10611), .Q(trans1[6]) );
  SDFFQX1 trans1_reg_5_ ( .D(N78), .SIN(trans1[4]), .SMC(test_se), .C(net10611), .Q(trans1[5]) );
  SDFFQX1 trans0_reg_6_ ( .D(N61), .SIN(trans0[5]), .SMC(test_se), .C(net10617), .Q(trans0[6]) );
  SDFFQX1 trans1_reg_4_ ( .D(N77), .SIN(trans1[3]), .SMC(test_se), .C(net10611), .Q(trans1[4]) );
  SDFFQX1 ntrancnt_reg_1_ ( .D(n56), .SIN(ntrancnt[0]), .SMC(test_se), .C(clk), 
        .Q(ntrancnt[1]) );
  SDFFQX1 ntrancnt_reg_0_ ( .D(n57), .SIN(n30), .SMC(test_se), .C(clk), .Q(
        ntrancnt[0]) );
  SDFFQX1 trans0_reg_5_ ( .D(N60), .SIN(trans0[4]), .SMC(test_se), .C(net10617), .Q(trans0[5]) );
  SDFFQX1 trans0_reg_4_ ( .D(N59), .SIN(trans0[3]), .SMC(test_se), .C(net10617), .Q(trans0[4]) );
  SDFFQX1 trans1_reg_3_ ( .D(N76), .SIN(trans1[2]), .SMC(test_se), .C(net10611), .Q(trans1[3]) );
  SDFFQX1 trans1_reg_2_ ( .D(N75), .SIN(trans1[1]), .SMC(test_se), .C(net10611), .Q(trans1[2]) );
  SDFFQX1 trans0_reg_3_ ( .D(N58), .SIN(trans0[2]), .SMC(test_se), .C(net10617), .Q(trans0[3]) );
  SDFFQX1 trans1_reg_1_ ( .D(N74), .SIN(trans1[0]), .SMC(test_se), .C(net10611), .Q(trans1[1]) );
  SDFFQX1 trans1_reg_0_ ( .D(N73), .SIN(trans0[7]), .SMC(test_se), .C(net10611), .Q(trans1[0]) );
  SDFFQX1 trans0_reg_2_ ( .D(N57), .SIN(trans0[1]), .SMC(test_se), .C(net10617), .Q(trans0[2]) );
  SDFFQX1 trans0_reg_1_ ( .D(N56), .SIN(trans0[0]), .SMC(test_se), .C(net10617), .Q(trans0[1]) );
  SDFFQX1 ttranwin_reg_7_ ( .D(N89), .SIN(ttranwin_6_), .SMC(test_se), .C(
        net10622), .Q(test_so) );
  SDFFQX1 ttranwin_reg_6_ ( .D(N88), .SIN(ttranwin_5_), .SMC(test_se), .C(
        net10622), .Q(ttranwin_6_) );
  SDFFQX1 trans0_reg_0_ ( .D(N55), .SIN(ntrancnt[1]), .SMC(test_se), .C(
        net10617), .Q(trans0[0]) );
  SDFFQX1 ttranwin_reg_5_ ( .D(N87), .SIN(ttranwin_4_), .SMC(test_se), .C(
        net10622), .Q(ttranwin_5_) );
  SDFFQX1 ttranwin_reg_4_ ( .D(N86), .SIN(ttranwin_3_), .SMC(test_se), .C(
        net10622), .Q(ttranwin_4_) );
  SDFFQX1 ttranwin_reg_1_ ( .D(N83), .SIN(ttranwin_0_), .SMC(test_se), .C(
        net10622), .Q(ttranwin_1_) );
  SDFFQX1 ttranwin_reg_2_ ( .D(N84), .SIN(ttranwin_1_), .SMC(test_se), .C(
        net10622), .Q(ttranwin_2_) );
  SDFFQX1 ttranwin_reg_3_ ( .D(N85), .SIN(ttranwin_2_), .SMC(test_se), .C(
        net10622), .Q(ttranwin_3_) );
  SDFFQX1 ttranwin_reg_0_ ( .D(N82), .SIN(trans1[7]), .SMC(test_se), .C(
        net10622), .Q(ttranwin_0_) );
  SDFFQX1 ccidle_reg ( .D(n55), .SIN(test_si), .SMC(test_se), .C(clk), .Q(n30)
         );
  INVX1 U5 ( .A(n29), .Y(o_ccidle) );
  NAND2X1 U6 ( .A(ntrancnt[0]), .B(n13), .Y(n2) );
  NAND2X1 U7 ( .A(ntrancnt[1]), .B(n14), .Y(n5) );
  INVX1 U8 ( .A(n52), .Y(n8) );
  INVX1 U9 ( .A(srstz), .Y(n6) );
  INVX1 U10 ( .A(n47), .Y(o_goidle) );
  OAI22X1 U11 ( .A(n8), .B(n11), .C(n49), .D(n33), .Y(N87) );
  OAI22X1 U12 ( .A(n8), .B(n10), .C(n32), .D(n49), .Y(N88) );
  NOR3XL U13 ( .A(n6), .B(o_goidle), .C(o_gobusy), .Y(n46) );
  OAI22X1 U14 ( .A(n8), .B(n15), .C(n49), .D(n34), .Y(N86) );
  NOR2X1 U15 ( .A(n12), .B(n48), .Y(n52) );
  OAI22X1 U16 ( .A(n8), .B(n16), .C(n49), .D(n35), .Y(N85) );
  OAI22X1 U17 ( .A(n8), .B(n17), .C(n49), .D(n36), .Y(N84) );
  OAI22X1 U18 ( .A(n8), .B(n26), .C(n49), .D(n37), .Y(N83) );
  INVX1 U19 ( .A(n45), .Y(n12) );
  NAND2X1 U20 ( .A(N12), .B(n44), .Y(n37) );
  OAI22X1 U21 ( .A(n12), .B(n9), .C(n31), .D(n5), .Y(N80) );
  OAI22X1 U22 ( .A(n8), .B(n9), .C(n31), .D(n49), .Y(N89) );
  INVX1 U23 ( .A(n38), .Y(n18) );
  AOI21X1 U24 ( .B(n28), .C(n29), .A(i_goidle), .Y(n47) );
  INVX1 U25 ( .A(ttranwin_minus[5]), .Y(n11) );
  INVX1 U26 ( .A(ttranwin_minus[6]), .Y(n10) );
  NAND2X1 U27 ( .A(N13), .B(n44), .Y(n36) );
  NAND2X1 U28 ( .A(N14), .B(n44), .Y(n35) );
  OAI22X1 U29 ( .A(n12), .B(n11), .C(n5), .D(n33), .Y(N78) );
  OAI22X1 U30 ( .A(n12), .B(n10), .C(n32), .D(n42), .Y(N79) );
  NOR3XL U31 ( .A(n7), .B(n42), .C(n29), .Y(o_gobusy) );
  INVX1 U32 ( .A(ttranwin_minus[4]), .Y(n15) );
  NOR2X1 U33 ( .A(N17), .B(n28), .Y(n32) );
  NAND2X1 U34 ( .A(N16), .B(n44), .Y(n33) );
  NAND2X1 U35 ( .A(N15), .B(n44), .Y(n34) );
  OAI221X1 U36 ( .A(i_trans), .B(n44), .C(n45), .D(n39), .E(n46), .Y(n40) );
  OAI22X1 U37 ( .A(n12), .B(n15), .C(n42), .D(n34), .Y(N77) );
  OAI22X1 U38 ( .A(n13), .B(n40), .C(n41), .D(n39), .Y(n56) );
  AND2X1 U39 ( .A(n42), .B(n2), .Y(n41) );
  INVX1 U40 ( .A(i_trans), .Y(n7) );
  ENOX1 U41 ( .A(n32), .B(n43), .C(N52), .D(n45), .Y(N61) );
  INVX1 U42 ( .A(n44), .Y(n28) );
  NAND2X1 U43 ( .A(n46), .B(i_trans), .Y(n39) );
  AOI31X1 U44 ( .A(n50), .B(n7), .C(n44), .D(n51), .Y(n49) );
  INVX1 U45 ( .A(ttranwin_minus[2]), .Y(n17) );
  INVX1 U46 ( .A(ttranwin_minus[3]), .Y(n16) );
  AOI21X1 U47 ( .B(n5), .C(n43), .A(n48), .Y(n51) );
  OAI22X1 U48 ( .A(n8), .B(n27), .C(n49), .D(n38), .Y(N82) );
  OAI22X1 U49 ( .A(n12), .B(n17), .C(n5), .D(n36), .Y(N75) );
  OAI22X1 U50 ( .A(n12), .B(n16), .C(n42), .D(n35), .Y(N76) );
  NAND2X1 U51 ( .A(n50), .B(i_trans), .Y(n48) );
  ENOX1 U52 ( .A(n43), .B(n33), .C(N51), .D(n45), .Y(N60) );
  OAI211X1 U53 ( .C(i_trans), .D(n28), .A(n50), .B(n53), .Y(N81) );
  NOR2X1 U54 ( .A(n52), .B(n51), .Y(n53) );
  INVX1 U55 ( .A(ttranwin_minus[1]), .Y(n26) );
  OAI22X1 U56 ( .A(n12), .B(n27), .C(n5), .D(n38), .Y(N73) );
  OAI22X1 U57 ( .A(n12), .B(n26), .C(n42), .D(n37), .Y(N74) );
  OAI21X1 U58 ( .B(n43), .C(n48), .A(n8), .Y(N91) );
  OAI21X1 U59 ( .B(n5), .C(n48), .A(n8), .Y(N90) );
  ENOX1 U60 ( .A(n2), .B(n35), .C(N49), .D(n45), .Y(N58) );
  ENOX1 U61 ( .A(n43), .B(n34), .C(N50), .D(n45), .Y(N59) );
  OAI211X1 U62 ( .C(o_gobusy), .D(n29), .A(n47), .B(srstz), .Y(n55) );
  ENOX1 U63 ( .A(n2), .B(n37), .C(N47), .D(n45), .Y(N56) );
  ENOX1 U64 ( .A(n43), .B(n36), .C(N48), .D(n45), .Y(N57) );
  NOR2X1 U65 ( .A(n14), .B(n13), .Y(n45) );
  INVX1 U66 ( .A(n36), .Y(n20) );
  INVX1 U67 ( .A(n35), .Y(n21) );
  INVX1 U68 ( .A(n34), .Y(n22) );
  INVX1 U69 ( .A(n33), .Y(n23) );
  INVX1 U70 ( .A(n37), .Y(n19) );
  INVX1 U71 ( .A(n32), .Y(n24) );
  NAND4X1 U72 ( .A(test_so), .B(ttranwin_6_), .C(n54), .D(n58), .Y(n44) );
  NOR2X1 U73 ( .A(ttranwin_1_), .B(ttranwin_0_), .Y(n54) );
  NOR4XL U74 ( .A(ttranwin_5_), .B(ttranwin_4_), .C(ttranwin_3_), .D(
        ttranwin_2_), .Y(n58) );
  NAND2X1 U75 ( .A(N11), .B(n44), .Y(n38) );
  INVX1 U76 ( .A(ttranwin_minus[7]), .Y(n9) );
  INVX1 U77 ( .A(n31), .Y(n25) );
  ENOX1 U78 ( .A(n31), .B(n2), .C(N53), .D(n45), .Y(N62) );
  OAI22X1 U79 ( .A(ntrancnt[0]), .B(n39), .C(n14), .D(n40), .Y(n57) );
  NOR2X1 U80 ( .A(N18), .B(n28), .Y(n31) );
  INVX1 U81 ( .A(n30), .Y(n29) );
  AOI31X1 U82 ( .A(n30), .B(n14), .C(i_trans), .D(n6), .Y(n50) );
  NAND2X1 U83 ( .A(ntrancnt[1]), .B(n14), .Y(n42) );
  INVX1 U84 ( .A(ttranwin_minus[0]), .Y(n27) );
  INVX1 U85 ( .A(ntrancnt[0]), .Y(n14) );
  NAND2X1 U86 ( .A(ntrancnt[0]), .B(n13), .Y(n43) );
  ENOX1 U87 ( .A(n2), .B(n38), .C(N46), .D(n45), .Y(N55) );
  INVX1 U88 ( .A(ntrancnt[1]), .Y(n13) );
endmodule


module phyidd_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module phyidd_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n17), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n10), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(A[0]), .Y(n18) );
  INVX1 U2 ( .A(B[2]), .Y(n14) );
  INVX1 U3 ( .A(B[3]), .Y(n15) );
  INVX1 U4 ( .A(B[4]), .Y(n13) );
  INVX1 U5 ( .A(B[5]), .Y(n11) );
  INVX1 U6 ( .A(B[1]), .Y(n17) );
  NAND21X1 U7 ( .B(n16), .A(n18), .Y(carry[1]) );
  INVX1 U8 ( .A(B[6]), .Y(n12) );
  INVX1 U9 ( .A(B[7]), .Y(n10) );
  INVX1 U10 ( .A(B[0]), .Y(n16) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module phyidd_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n18), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n10), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(B[2]), .Y(n14) );
  INVX1 U2 ( .A(B[3]), .Y(n15) );
  INVX1 U3 ( .A(B[4]), .Y(n13) );
  INVX1 U4 ( .A(B[5]), .Y(n11) );
  INVX1 U5 ( .A(B[1]), .Y(n18) );
  NAND21X1 U6 ( .B(n17), .A(n16), .Y(carry[1]) );
  INVX1 U7 ( .A(A[0]), .Y(n16) );
  INVX1 U8 ( .A(B[6]), .Y(n12) );
  INVX1 U9 ( .A(B[7]), .Y(n10) );
  INVX1 U10 ( .A(B[0]), .Y(n17) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_a0 ( i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, 
        r_rxdb_opt, r_ords_ena, r_pshords, r_rgdcrc, prx_cccnt, prx_rst, 
        prx_setsta, prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, 
        prx_fifopsh, prx_fifowdat, pff_txreq, pid_gobusy, pid_goidle, 
        pid_ccidle, pcc_rxgood, prx_crcstart, prx_crcshfi4, prx_crcsidat, 
        prx_rxcode, prx_adpn, prx_rcvdords, prx_eoprcvd, prx_fsm, clk, srstz, 
        test_si, test_so, test_se );
  input [1:0] r_rxdb_opt;
  input [6:0] r_ords_ena;
  output [1:0] prx_cccnt;
  output [1:0] prx_rst;
  output [6:0] prx_setsta;
  output [7:0] prx_fifowdat;
  output [3:0] prx_crcsidat;
  output [4:0] prx_rxcode;
  output [5:0] prx_adpn;
  output [2:0] prx_rcvdords;
  output [3:0] prx_fsm;
  input i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_pshords,
         r_rgdcrc, pff_txreq, pid_gobusy, pid_goidle, pid_ccidle, pcc_rxgood,
         clk, srstz, test_si, test_se;
  output prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, prx_fifopsh,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd, test_so;
  wire   N31, N32, N33, db_gohi, db_golo, cctrans, shrtrans, N58, N59, N60,
         N61, N70, N71, N72, N73, N74, N75, N76, N96, N153, N154, N155, N156,
         N157, ps_ords_ena, cs_ords_ena, N236, N239, N246, N247, N248, N249,
         N250, N275, N276, N277, N278, N279, net10639, net10645, net10650,
         net10655, net10660, net10665, net10670, n214, n284, n187, n188, n189,
         n190, n191, n192, n271, n17, n74, n79, n80, n84, n87, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n125, n126, n127, n128,
         n131, n132, n134, n138, n139, n140, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n154, n156, n157, n159, n160, n162,
         n164, n165, n166, n167, n170, n171, n172, n173, n174, n176, n213,
         n215, n1, n3, n4, n5, n6, n7, n8, n9, n11, n15, n18, n20, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n81, n82,
         n83, n85, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n129, n130, n133, n135, n136,
         n137, n141, n142, n153, n155, n158, n161, n163, n168, n169, n175,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283;
  wire   [5:0] cccnt;
  wire   [2:0] ps_dat5b;
  wire   [2:0] bcnt;
  wire   [7:3] ordsbuf;
  wire   [5:2] add_83_carry;

  HAD1X1 add_83_U1_1_1 ( .A(cccnt[1]), .B(cccnt[0]), .CO(add_83_carry[2]), 
        .SO(N58) );
  HAD1X1 add_83_U1_1_2 ( .A(cccnt[2]), .B(add_83_carry[2]), .CO(
        add_83_carry[3]), .SO(N59) );
  HAD1X1 add_83_U1_1_3 ( .A(cccnt[3]), .B(add_83_carry[3]), .CO(
        add_83_carry[4]), .SO(N60) );
  HAD1X1 add_83_U1_1_4 ( .A(cccnt[4]), .B(add_83_carry[4]), .CO(
        add_83_carry[5]), .SO(N61) );
  phyrx_db u0_phyrx_db ( .clk(clk), .srstz(srstz), .x_cc(i_cc), .ptx_txact(n4), 
        .r_rxdb_opt(r_rxdb_opt), .gohi(db_gohi), .golo(db_golo), .gotrans(
        prx_trans), .test_si(n271), .test_so(test_so), .test_se(test_se) );
  phyrx_adp u0_phyrx_adp ( .clk(clk), .srstz(srstz), .gohi(db_gohi), .golo(
        db_golo), .gobusy(pid_gobusy), .goidle(pid_goidle), .i_ccidle(
        pid_ccidle), .k0_det(n17), .r_adprx_en(r_adprx_en), .r_adp2nd(r_adp2nd), .adp_val(prx_adpn), .d_cc(prx_d_cc), .cctrans(cctrans), .test_si(shrtrans), 
        .test_so(n271), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 clk_gate_cccnt_reg ( .CLK(clk), .EN(N70), 
        .ENCLK(net10639), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 clk_gate_cs_dat5b_reg ( .CLK(clk), .EN(N153), 
        .ENCLK(net10645), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 clk_gate_bcnt_reg ( .CLK(clk), .EN(N236), 
        .ENCLK(net10650), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 clk_gate_cs_dat4b_reg ( .CLK(clk), .EN(n213), 
        .ENCLK(net10655), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 clk_gate_ordsbuf_reg ( .CLK(clk), .EN(n215), 
        .ENCLK(net10660), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 clk_gate_ordsbuf_reg_0 ( .CLK(clk), .EN(N250), .ENCLK(net10665), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 clk_gate_cs_bmni_reg ( .CLK(clk), .EN(N275), 
        .ENCLK(net10670), .TE(test_se) );
  SDFFQX1 ordsbuf_reg_4_ ( .D(prx_fifowdat[4]), .SIN(ordsbuf[3]), .SMC(test_se), .C(net10660), .Q(ordsbuf[4]) );
  SDFFQX1 ordsbuf_reg_7_ ( .D(prx_fifowdat[7]), .SIN(ordsbuf[6]), .SMC(test_se), .C(net10660), .Q(ordsbuf[7]) );
  SDFFQX1 ordsbuf_reg_6_ ( .D(prx_fifowdat[6]), .SIN(ordsbuf[5]), .SMC(test_se), .C(net10660), .Q(ordsbuf[6]) );
  SDFFQX1 cs_dat4b_reg_2_ ( .D(prx_fifowdat[6]), .SIN(prx_fifowdat[1]), .SMC(
        test_se), .C(net10655), .Q(prx_fifowdat[2]) );
  SDFFQX1 ordsbuf_reg_5_ ( .D(prx_fifowdat[5]), .SIN(ordsbuf[4]), .SMC(test_se), .C(net10660), .Q(ordsbuf[5]) );
  SDFFQX1 ordsbuf_reg_3_ ( .D(N249), .SIN(prx_rcvdords[2]), .SMC(test_se), .C(
        net10665), .Q(ordsbuf[3]) );
  SDFFQX1 cs_dat4b_reg_1_ ( .D(prx_fifowdat[5]), .SIN(prx_fifowdat[0]), .SMC(
        test_se), .C(net10655), .Q(prx_fifowdat[1]) );
  SDFFQX1 cs_dat4b_reg_0_ ( .D(prx_fifowdat[4]), .SIN(n3), .SMC(test_se), .C(
        net10655), .Q(prx_fifowdat[0]) );
  SDFFQX1 cs_dat4b_reg_3_ ( .D(prx_crcsidat[3]), .SIN(prx_fifowdat[2]), .SMC(
        test_se), .C(net10655), .Q(prx_rxcode[3]) );
  SDFFQX1 cs_dat4b_reg_4_ ( .D(N96), .SIN(prx_rxcode[3]), .SMC(test_se), .C(
        net10655), .Q(prx_rxcode[4]) );
  SDFFQX1 bcnt_reg_0_ ( .D(n256), .SIN(test_si), .SMC(test_se), .C(net10650), 
        .Q(bcnt[0]) );
  SDFFQX1 bcnt_reg_1_ ( .D(n262), .SIN(bcnt[0]), .SMC(test_se), .C(net10650), 
        .Q(bcnt[1]) );
  SDFFQX1 bcnt_reg_2_ ( .D(N239), .SIN(bcnt[1]), .SMC(test_se), .C(net10650), 
        .Q(bcnt[2]) );
  SDFFQX1 cs_bmni_reg_2_ ( .D(N278), .SIN(prx_fsm[1]), .SMC(test_se), .C(
        net10670), .Q(prx_fsm[2]) );
  SDFFQX1 cs_bmni_reg_1_ ( .D(N277), .SIN(prx_fsm[0]), .SMC(test_se), .C(
        net10670), .Q(prx_fsm[1]) );
  SDFFQX1 cs_bmni_reg_0_ ( .D(N276), .SIN(cccnt[5]), .SMC(test_se), .C(
        net10670), .Q(prx_fsm[0]) );
  SDFFQX1 cs_bmni_reg_3_ ( .D(N279), .SIN(prx_fsm[2]), .SMC(test_se), .C(
        net10670), .Q(prx_fsm[3]) );
  SDFFQX1 cs_dat5b_reg_0_ ( .D(N154), .SIN(prx_rxcode[4]), .SMC(test_se), .C(
        net10645), .Q(ps_dat5b[0]) );
  SDFFQX1 cs_dat5b_reg_1_ ( .D(N155), .SIN(ps_dat5b[0]), .SMC(test_se), .C(
        net10645), .Q(ps_dat5b[1]) );
  SDFFQX1 cs_dat5b_reg_2_ ( .D(N156), .SIN(ps_dat5b[1]), .SMC(test_se), .C(
        net10645), .Q(ps_dat5b[2]) );
  SDFFQX1 cs_dat5b_reg_3_ ( .D(N157), .SIN(ps_dat5b[2]), .SMC(test_se), .C(
        net10645), .Q(prx_bmc) );
  SDFFQX1 cccnt_reg_4_ ( .D(N75), .SIN(cccnt[3]), .SMC(test_se), .C(net10639), 
        .Q(cccnt[4]) );
  SDFFQX1 cccnt_reg_3_ ( .D(N74), .SIN(cccnt[2]), .SMC(test_se), .C(net10639), 
        .Q(cccnt[3]) );
  SDFFQX1 cccnt_reg_1_ ( .D(N72), .SIN(cccnt[0]), .SMC(test_se), .C(net10639), 
        .Q(cccnt[1]) );
  SDFFQX1 cccnt_reg_2_ ( .D(N73), .SIN(cccnt[1]), .SMC(test_se), .C(net10639), 
        .Q(cccnt[2]) );
  SDFFQX1 cccnt_reg_0_ ( .D(N71), .SIN(bcnt[2]), .SMC(test_se), .C(net10639), 
        .Q(cccnt[0]) );
  SDFFQX1 shrtrans_reg ( .D(n214), .SIN(ordsbuf[7]), .SMC(test_se), .C(clk), 
        .Q(shrtrans) );
  SDFFQX1 cccnt_reg_5_ ( .D(N76), .SIN(cccnt[4]), .SMC(test_se), .C(net10639), 
        .Q(cccnt[5]) );
  SDFFQX1 ordsbuf_reg_1_ ( .D(N247), .SIN(prx_rcvdords[0]), .SMC(test_se), .C(
        net10665), .Q(prx_rcvdords[1]) );
  SDFFQX1 ordsbuf_reg_2_ ( .D(N248), .SIN(prx_rcvdords[1]), .SMC(test_se), .C(
        net10665), .Q(prx_rcvdords[2]) );
  SDFFQX1 ordsbuf_reg_0_ ( .D(N246), .SIN(prx_bmc), .SMC(test_se), .C(net10665), .Q(prx_rcvdords[0]) );
  NOR21XL U223 ( .B(r_ords_ena[0]), .A(n282), .Y(n192) );
  MUX4X1 U220 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[4]), .D2(r_ords_ena[5]), 
        .D3(r_ords_ena[6]), .S0(N31), .S1(N32), .Y(n187) );
  MUX2X1 U219 ( .D0(r_ords_ena[1]), .D1(r_ords_ena[2]), .S(N31), .Y(n188) );
  NOR21XL U218 ( .B(r_ords_ena[0]), .A(n257), .Y(n189) );
  MUX3X1 U217 ( .D0(n189), .D1(n188), .D2(n187), .S0(N32), .S1(N33), .Y(
        ps_ords_ena) );
  MUX4XL U44 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[4]), .D2(r_ords_ena[5]), 
        .D3(r_ords_ena[6]), .S0(prx_rcvdords[0]), .S1(prx_rcvdords[1]), .Y(
        n190) );
  MUX2XL U43 ( .D0(r_ords_ena[1]), .D1(r_ords_ena[2]), .S(prx_rcvdords[0]), 
        .Y(n191) );
  MUX3XL U42 ( .D0(n192), .D1(n191), .D2(n190), .S0(prx_rcvdords[1]), .S1(
        prx_rcvdords[2]), .Y(cs_ords_ena) );
  INVX3 U3 ( .A(prx_fifowdat[5]), .Y(n18) );
  NAND31X2 U4 ( .C(n50), .A(n49), .B(n48), .Y(prx_fifowdat[5]) );
  NAND21X2 U5 ( .B(ps_dat5b[1]), .A(n223), .Y(n55) );
  INVX1 U6 ( .A(n49), .Y(n42) );
  AOI21BBXL U7 ( .B(n55), .C(n116), .A(n54), .Y(n56) );
  AO21X1 U8 ( .B(prx_fsm[1]), .C(n121), .A(n120), .Y(n123) );
  NAND21X1 U9 ( .B(n116), .A(n223), .Y(n53) );
  NOR2X1 U10 ( .A(n117), .B(n225), .Y(n7) );
  NAND31X1 U11 ( .C(n42), .A(n41), .B(n40), .Y(n43) );
  NAND21X1 U12 ( .B(n223), .A(prx_bmc), .Y(n136) );
  NAND21X1 U13 ( .B(n59), .A(n33), .Y(n35) );
  MUX2X1 U14 ( .D0(ps_dat5b[1]), .D1(n114), .S(prx_bmc), .Y(n115) );
  NAND21X1 U15 ( .B(n59), .A(n58), .Y(n60) );
  NAND21X1 U16 ( .B(n57), .A(n56), .Y(n58) );
  NAND21XL U17 ( .B(n46), .A(n45), .Y(prx_fifowdat[4]) );
  NAND3X1 U18 ( .A(ps_dat5b[2]), .B(n39), .C(ps_dat5b[0]), .Y(n1) );
  NAND21X2 U19 ( .B(n61), .A(n60), .Y(prx_fifowdat[6]) );
  NAND21X1 U20 ( .B(n46), .A(n45), .Y(n284) );
  MUX2IX1 U21 ( .D0(n44), .D1(n43), .S(ps_dat5b[0]), .Y(n45) );
  INVX1 U22 ( .A(n111), .Y(n3) );
  BUFX3 U23 ( .A(ptx_txact), .Y(n4) );
  BUFX3 U24 ( .A(prx_fifowdat[0]), .Y(prx_rxcode[0]) );
  BUFX3 U25 ( .A(prx_fifowdat[2]), .Y(prx_rxcode[2]) );
  BUFX3 U26 ( .A(prx_fifowdat[1]), .Y(prx_rxcode[1]) );
  NOR21X1 U27 ( .B(ps_dat5b[0]), .A(n55), .Y(n50) );
  OR2X1 U28 ( .A(n36), .B(n6), .Y(N96) );
  AND2XL U29 ( .A(n79), .B(n7), .Y(n5) );
  AND2XL U30 ( .A(n185), .B(n15), .Y(n186) );
  NAND21XL U31 ( .B(n86), .A(n89), .Y(n88) );
  MUX2BXL U32 ( .D0(n35), .D1(n1), .S(n223), .Y(n6) );
  AO21XL U33 ( .B(n9), .C(n118), .A(n5), .Y(prx_crcshfi4) );
  AND4XL U34 ( .A(n227), .B(n136), .C(n135), .D(n133), .Y(prx_setsta[0]) );
  INVXL U35 ( .A(prx_rcvdords[0]), .Y(n282) );
  NOR42XL U36 ( .C(ordsbuf[7]), .D(ordsbuf[5]), .A(n276), .B(ordsbuf[4]), .Y(
        n170) );
  NAND3XL U37 ( .A(n259), .B(n274), .C(prx_rcvdords[1]), .Y(n104) );
  NAND42X1 U38 ( .C(n279), .D(n161), .A(ordsbuf[3]), .B(n165), .Y(n163) );
  INVXL U39 ( .A(prx_rcvdords[1]), .Y(n281) );
  INVXL U40 ( .A(prx_rcvdords[2]), .Y(n280) );
  NAND21X1 U41 ( .B(n167), .A(n201), .Y(n159) );
  INVX1 U45 ( .A(n155), .Y(n201) );
  NAND21X1 U46 ( .B(n224), .A(n89), .Y(N153) );
  INVX1 U47 ( .A(n85), .Y(n89) );
  NAND21X1 U48 ( .B(n232), .A(n264), .Y(n85) );
  INVX1 U49 ( .A(pid_goidle), .Y(n265) );
  INVX1 U50 ( .A(srstz), .Y(n22) );
  INVX1 U51 ( .A(n245), .Y(n227) );
  INVX1 U52 ( .A(n168), .Y(n204) );
  NAND21X1 U53 ( .B(n15), .A(n204), .Y(n155) );
  OA22X1 U54 ( .A(n272), .B(n167), .C(n155), .D(n153), .Y(n158) );
  INVX1 U55 ( .A(n172), .Y(n153) );
  NOR2X1 U56 ( .A(n146), .B(n147), .Y(n126) );
  AO21X1 U57 ( .B(n211), .C(n210), .A(n209), .Y(N32) );
  INVX1 U58 ( .A(n127), .Y(n210) );
  NAND21X1 U59 ( .B(n148), .A(n106), .Y(n209) );
  INVX1 U60 ( .A(N31), .Y(n257) );
  INVX1 U61 ( .A(n118), .Y(n70) );
  NAND2X1 U62 ( .A(N33), .B(N32), .Y(n74) );
  OAI21X1 U63 ( .B(n162), .C(n272), .A(n167), .Y(n172) );
  INVX1 U64 ( .A(n167), .Y(n269) );
  INVX1 U65 ( .A(n206), .Y(n197) );
  NAND21X1 U66 ( .B(n22), .A(n108), .Y(n232) );
  INVX1 U67 ( .A(n251), .Y(n253) );
  INVX1 U68 ( .A(n88), .Y(n224) );
  INVX1 U69 ( .A(n134), .Y(n274) );
  INVX1 U70 ( .A(n244), .Y(n235) );
  INVX1 U71 ( .A(pid_gobusy), .Y(n264) );
  INVX1 U72 ( .A(n212), .Y(n255) );
  AND2X1 U73 ( .A(n255), .B(prx_fifowdat[3]), .Y(N249) );
  INVX1 U74 ( .A(n129), .Y(n86) );
  INVX2 U75 ( .A(n62), .Y(n185) );
  NAND32X1 U76 ( .B(n24), .C(n25), .A(n90), .Y(n219) );
  INVX1 U77 ( .A(n96), .Y(n24) );
  INVX1 U78 ( .A(n142), .Y(prx_cccnt[0]) );
  NAND21X1 U79 ( .B(n121), .A(n77), .Y(n245) );
  NAND32X1 U80 ( .B(n73), .C(n121), .A(n71), .Y(n212) );
  NAND32X1 U81 ( .B(n73), .C(n122), .A(n121), .Y(n75) );
  INVX1 U82 ( .A(n169), .Y(prx_fifowdat[3]) );
  NAND31X1 U83 ( .C(pff_txreq), .A(n94), .B(n93), .Y(n107) );
  NAND21X1 U84 ( .B(n142), .A(n4), .Y(n93) );
  AO21X1 U85 ( .B(n222), .C(n216), .A(n22), .Y(N71) );
  AO21X1 U86 ( .B(N59), .C(n222), .A(n22), .Y(N73) );
  AO21X1 U87 ( .B(N60), .C(n222), .A(n22), .Y(N74) );
  AO21X1 U88 ( .B(N58), .C(n222), .A(n22), .Y(N72) );
  AO21X1 U89 ( .B(N61), .C(n222), .A(n22), .Y(N75) );
  INVX1 U90 ( .A(n217), .Y(n222) );
  NAND32X1 U91 ( .B(n22), .C(n107), .A(n217), .Y(N70) );
  NAND31XL U92 ( .C(prx_fifowdat[6]), .A(prx_fifowdat[7]), .B(prx_fifowdat[5]), 
        .Y(n168) );
  NAND31X1 U93 ( .C(n200), .A(n199), .B(n98), .Y(n105) );
  NOR2X1 U94 ( .A(n159), .B(n134), .Y(n200) );
  NAND21X1 U95 ( .B(n267), .A(n198), .Y(n199) );
  NAND21X1 U96 ( .B(n197), .A(n196), .Y(n198) );
  OAI21X1 U97 ( .B(n160), .C(n269), .A(n195), .Y(n202) );
  NOR2X1 U98 ( .A(n162), .B(n134), .Y(n160) );
  NOR2X1 U99 ( .A(n105), .B(n145), .Y(n127) );
  NAND4X1 U100 ( .A(n261), .B(n126), .C(n127), .D(n138), .Y(n106) );
  INVX1 U101 ( .A(n148), .Y(n261) );
  OAI21X1 U102 ( .B(n134), .C(n139), .A(n140), .Y(n138) );
  AOI32X1 U103 ( .A(n275), .B(n281), .C(n259), .D(n143), .E(n201), .Y(n140) );
  NAND4X1 U104 ( .A(n97), .B(n98), .C(n99), .D(n100), .Y(n79) );
  AOI211X1 U105 ( .C(n263), .D(n275), .A(n101), .B(n102), .Y(n100) );
  AOI21X1 U106 ( .B(n103), .C(n104), .A(n105), .Y(n101) );
  INVX1 U107 ( .A(n106), .Y(n263) );
  OAI211X1 U108 ( .C(n267), .D(n180), .A(n179), .B(n178), .Y(n147) );
  INVX1 U109 ( .A(n102), .Y(n178) );
  NAND32X1 U110 ( .B(n167), .C(n272), .A(n204), .Y(n179) );
  AOI32X1 U111 ( .A(n172), .B(n195), .C(n15), .D(n170), .E(n181), .Y(n180) );
  OAI211X1 U112 ( .C(n272), .D(n159), .A(n173), .B(n103), .Y(n146) );
  NAND43X1 U113 ( .B(n169), .C(n158), .D(prx_rxcode[0]), .A(n176), .Y(n173) );
  NOR2X1 U114 ( .A(n267), .B(n278), .Y(n176) );
  INVX1 U115 ( .A(n208), .Y(n211) );
  OAI211X1 U116 ( .C(n128), .D(n105), .A(n106), .B(n211), .Y(N31) );
  AOI21BX1 U117 ( .C(n146), .B(n147), .A(n145), .Y(n128) );
  OAI21X1 U118 ( .B(n125), .C(n208), .A(n207), .Y(N33) );
  NAND21X1 U119 ( .B(n126), .A(n127), .Y(n125) );
  INVX1 U120 ( .A(n209), .Y(n207) );
  NOR2X1 U121 ( .A(n257), .B(n74), .Y(prx_rst[0]) );
  NOR2X1 U122 ( .A(N31), .B(n74), .Y(prx_rst[1]) );
  INVX1 U123 ( .A(ps_ords_ena), .Y(n237) );
  INVXL U124 ( .A(N96), .Y(n69) );
  INVX1 U125 ( .A(n124), .Y(prx_setsta[6]) );
  NAND32X1 U126 ( .B(n137), .C(n141), .A(prx_eoprcvd), .Y(n124) );
  AND3X1 U127 ( .A(prx_eoprcvd), .B(pcc_rxgood), .C(n137), .Y(prx_setsta[3])
         );
  OA21X1 U128 ( .B(n231), .C(n242), .A(n235), .Y(N279) );
  INVX1 U129 ( .A(n230), .Y(n231) );
  INVX1 U130 ( .A(n112), .Y(prx_eoprcvd) );
  NAND32X1 U131 ( .B(n111), .C(n110), .A(n109), .Y(n112) );
  INVX1 U132 ( .A(cs_ords_ena), .Y(n110) );
  INVX1 U133 ( .A(n108), .Y(n109) );
  OAI211X1 U134 ( .C(n144), .D(n139), .A(n149), .B(n99), .Y(n148) );
  OAI211X1 U135 ( .C(n152), .D(n193), .A(prx_fifowdat[7]), .B(n186), .Y(n149)
         );
  INVX1 U136 ( .A(n139), .Y(n193) );
  NOR2X1 U137 ( .A(n268), .B(n144), .Y(n152) );
  AOI31X1 U138 ( .A(n247), .B(n246), .C(n245), .D(n244), .Y(N277) );
  INVX1 U139 ( .A(n243), .Y(n246) );
  INVX1 U140 ( .A(n242), .Y(n247) );
  AOI21X1 U141 ( .B(n241), .C(n240), .A(n244), .Y(N278) );
  AO21X1 U142 ( .B(n79), .C(ps_ords_ena), .A(n239), .Y(n241) );
  NAND21X1 U143 ( .B(n225), .A(n74), .Y(n239) );
  GEN2XL U144 ( .D(n238), .E(n237), .C(n236), .B(n235), .A(n234), .Y(N276) );
  NOR5X1 U145 ( .A(n264), .B(n233), .C(n232), .D(pid_goidle), .E(n4), .Y(n234)
         );
  INVX1 U146 ( .A(n239), .Y(n238) );
  OAI22AX1 U147 ( .D(N32), .C(n225), .A(n267), .B(n212), .Y(N247) );
  OAI22AX1 U148 ( .D(N33), .C(n225), .A(n278), .B(n212), .Y(N248) );
  INVX1 U149 ( .A(n113), .Y(n114) );
  OAI22X1 U150 ( .A(n257), .B(n225), .C(n279), .D(n212), .Y(N246) );
  NAND21X1 U151 ( .B(n194), .A(n274), .Y(n206) );
  NAND2X1 U152 ( .A(n131), .B(n283), .Y(n167) );
  INVX1 U153 ( .A(n177), .Y(n183) );
  NAND21X1 U154 ( .B(n279), .A(prx_fifowdat[3]), .Y(n177) );
  INVX1 U155 ( .A(n170), .Y(n272) );
  OAI21X1 U156 ( .B(n268), .C(n134), .A(n139), .Y(n143) );
  NOR2X1 U157 ( .A(n283), .B(n131), .Y(n162) );
  INVX1 U158 ( .A(n194), .Y(n181) );
  NOR32XL U159 ( .B(n171), .C(n279), .A(n164), .Y(n102) );
  NOR32XL U160 ( .B(n150), .C(n283), .A(n280), .Y(n156) );
  NAND21X1 U161 ( .B(n184), .A(n156), .Y(n139) );
  NAND3X1 U162 ( .A(n277), .B(n276), .C(n157), .Y(n134) );
  INVX1 U163 ( .A(n161), .Y(n260) );
  NAND3X1 U164 ( .A(n259), .B(n281), .C(n273), .Y(n98) );
  OAI21BBX1 U165 ( .A(n227), .B(n135), .C(n233), .Y(n83) );
  INVX1 U166 ( .A(n233), .Y(prx_idle) );
  NAND4X1 U167 ( .A(n150), .B(n279), .C(n260), .D(n151), .Y(n99) );
  NOR3XL U168 ( .A(n280), .B(n144), .C(n278), .Y(n151) );
  INVX1 U169 ( .A(n249), .Y(n256) );
  INVX1 U170 ( .A(n164), .Y(n273) );
  NAND42X1 U171 ( .C(n232), .D(pid_goidle), .A(n81), .B(n78), .Y(N275) );
  NAND31X1 U172 ( .C(n233), .A(n266), .B(pid_gobusy), .Y(n78) );
  NAND21X1 U173 ( .B(n244), .A(n76), .Y(n81) );
  NAND42X1 U174 ( .C(n243), .D(n236), .A(n229), .B(n225), .Y(n76) );
  NAND4X1 U175 ( .A(n278), .B(n279), .C(n131), .D(n132), .Y(n97) );
  NOR21XL U176 ( .B(n260), .A(n134), .Y(n132) );
  INVX1 U177 ( .A(n144), .Y(n275) );
  INVX1 U178 ( .A(pcc_rxgood), .Y(n141) );
  INVX1 U179 ( .A(n229), .Y(n119) );
  INVX1 U180 ( .A(n4), .Y(n266) );
  NAND32X1 U181 ( .B(n73), .C(n111), .A(n122), .Y(n230) );
  NAND21X1 U182 ( .B(n255), .A(n240), .Y(n243) );
  NAND2X1 U183 ( .A(n226), .B(n230), .Y(n236) );
  INVX1 U184 ( .A(n65), .Y(n66) );
  NAND21X1 U185 ( .B(n51), .A(n47), .Y(n48) );
  NAND21X1 U186 ( .B(prx_bmc), .A(ps_dat5b[0]), .Y(n47) );
  INVX1 U187 ( .A(shrtrans), .Y(n30) );
  INVX1 U188 ( .A(n219), .Y(n32) );
  INVX1 U189 ( .A(n218), .Y(n31) );
  NAND21X1 U190 ( .B(n136), .A(n113), .Y(n40) );
  NOR21XL U191 ( .B(ps_dat5b[0]), .A(n51), .Y(n61) );
  NOR21XL U192 ( .B(n59), .A(n51), .Y(n46) );
  NOR32XL U193 ( .B(n116), .C(prx_bmc), .A(n55), .Y(n44) );
  OR3XL U194 ( .A(bcnt[1]), .B(n250), .C(bcnt[0]), .Y(n68) );
  OAI21BBX1 U195 ( .A(r_pshords), .B(N250), .C(n8), .Y(prx_fifopsh) );
  NAND3X1 U196 ( .A(n123), .B(n122), .C(n9), .Y(n8) );
  NOR2XL U197 ( .A(n117), .B(n111), .Y(n9) );
  GEN2XL U198 ( .D(shrtrans), .E(n216), .C(n29), .B(n28), .A(n27), .Y(n218) );
  AND2X1 U199 ( .A(n65), .B(n91), .Y(n27) );
  INVX1 U200 ( .A(n25), .Y(n28) );
  NAND21X1 U201 ( .B(n29), .A(cccnt[0]), .Y(n96) );
  AO21X1 U202 ( .B(cccnt[2]), .C(cccnt[1]), .A(cccnt[5]), .Y(n25) );
  NAND21X1 U203 ( .B(n26), .A(cccnt[4]), .Y(n65) );
  INVX1 U204 ( .A(cccnt[5]), .Y(n91) );
  INVX1 U205 ( .A(cccnt[3]), .Y(n26) );
  INVX1 U206 ( .A(cccnt[0]), .Y(n216) );
  INVX1 U207 ( .A(cccnt[2]), .Y(n29) );
  NAND43X1 U208 ( .B(n92), .C(n91), .D(n96), .A(n90), .Y(n142) );
  INVX1 U209 ( .A(cccnt[1]), .Y(n92) );
  INVX1 U210 ( .A(n23), .Y(n90) );
  NAND21X1 U211 ( .B(cccnt[4]), .A(n26), .Y(n23) );
  NAND21X1 U212 ( .B(ps_dat5b[1]), .A(ps_dat5b[2]), .Y(n113) );
  NAND21X1 U213 ( .B(ps_dat5b[0]), .A(n37), .Y(n33) );
  INVX1 U214 ( .A(ps_dat5b[1]), .Y(n37) );
  INVX1 U215 ( .A(ps_dat5b[2]), .Y(n116) );
  INVX1 U216 ( .A(prx_bmc), .Y(n59) );
  INVX1 U221 ( .A(n34), .Y(n39) );
  NAND21X1 U222 ( .B(n37), .A(prx_bmc), .Y(n34) );
  INVX1 U224 ( .A(prx_fsm[3]), .Y(n111) );
  INVX1 U225 ( .A(prx_fsm[0]), .Y(n121) );
  INVX1 U226 ( .A(n64), .Y(n77) );
  NAND21X1 U227 ( .B(prx_fsm[1]), .A(n71), .Y(n64) );
  INVX1 U228 ( .A(n63), .Y(n71) );
  NAND21X1 U229 ( .B(prx_fsm[2]), .A(n111), .Y(n63) );
  INVX1 U230 ( .A(bcnt[2]), .Y(n250) );
  OR2X1 U231 ( .A(prx_fsm[3]), .B(n75), .Y(n225) );
  INVX1 U232 ( .A(n72), .Y(n120) );
  NAND21X1 U233 ( .B(prx_fsm[1]), .A(prx_fsm[0]), .Y(n72) );
  INVX1 U234 ( .A(prx_fsm[2]), .Y(n122) );
  INVX1 U235 ( .A(prx_fsm[1]), .Y(n73) );
  MUX2IX1 U236 ( .D0(prx_rxcode[4]), .D1(prx_rxcode[3]), .S(prx_fsm[3]), .Y(
        n169) );
  OAI31XL U237 ( .A(n87), .B(n91), .C(n96), .D(n95), .Y(n217) );
  NAND3X1 U238 ( .A(cccnt[3]), .B(cccnt[1]), .C(cccnt[4]), .Y(n87) );
  INVX1 U239 ( .A(n107), .Y(n95) );
  OAI21X1 U240 ( .B(n84), .C(n217), .A(srstz), .Y(N76) );
  XNOR2XL U241 ( .A(cccnt[5]), .B(add_83_carry[5]), .Y(n84) );
  MUX2XL U242 ( .D0(N96), .D1(prx_crcsidat[3]), .S(prx_fsm[3]), .Y(
        prx_fifowdat[7]) );
  INVX1 U243 ( .A(n175), .Y(n195) );
  NAND43X1 U244 ( .B(prx_fifowdat[2]), .C(n169), .D(n168), .A(prx_fifowdat[0]), 
        .Y(n175) );
  NOR2XL U245 ( .A(n130), .B(n11), .Y(prx_crcsidat[3]) );
  AOI21X1 U246 ( .B(ps_dat5b[1]), .C(n116), .A(n115), .Y(n11) );
  OAI221X1 U247 ( .A(prx_fifowdat[1]), .B(n182), .C(n164), .D(n159), .E(n104), 
        .Y(n145) );
  OAI21X1 U248 ( .B(n162), .C(n164), .A(n167), .Y(n166) );
  AOI32X1 U249 ( .A(n269), .B(n274), .C(n204), .D(n203), .E(n267), .Y(n205) );
  INVX1 U250 ( .A(n202), .Y(n203) );
  AND2XL U251 ( .A(n7), .B(ps_ords_ena), .Y(prx_setsta[1]) );
  AND2XL U252 ( .A(n7), .B(n237), .Y(prx_setsta[2]) );
  OAI211X1 U253 ( .C(prx_fsm[0]), .D(n230), .A(n229), .B(n228), .Y(n242) );
  OA22X1 U254 ( .A(n227), .B(n226), .C(n239), .D(n237), .Y(n228) );
  AND2X1 U255 ( .A(prx_eoprcvd), .B(n141), .Y(prx_setsta[4]) );
  NOR21XL U256 ( .B(n150), .A(prx_rcvdords[2]), .Y(n131) );
  NAND32X1 U257 ( .B(prx_fifowdat[2]), .C(n167), .A(n183), .Y(n194) );
  NAND32X1 U258 ( .B(n278), .C(prx_fifowdat[1]), .A(n183), .Y(n184) );
  INVX1 U259 ( .A(n154), .Y(n268) );
  GEN2XL U260 ( .D(prx_rcvdords[2]), .E(n150), .C(n283), .B(n258), .A(n156), 
        .Y(n154) );
  INVX1 U261 ( .A(n184), .Y(n258) );
  NOR3XL U262 ( .A(n282), .B(prx_rcvdords[1]), .C(n270), .Y(n150) );
  INVX1 U263 ( .A(ordsbuf[3]), .Y(n270) );
  NOR43XL U264 ( .B(prx_rcvdords[2]), .C(n260), .D(n174), .A(n281), .Y(n171)
         );
  NOR3XL U265 ( .A(n270), .B(prx_rcvdords[0]), .C(prx_fifowdat[2]), .Y(n174)
         );
  INVX1 U266 ( .A(n163), .Y(n259) );
  NOR3XL U267 ( .A(n282), .B(prx_rcvdords[2]), .C(prx_fifowdat[2]), .Y(n165)
         );
  NAND32X1 U268 ( .B(n267), .C(r_exist1st), .A(prx_fifowdat[3]), .Y(n161) );
  INVX1 U269 ( .A(prx_fifowdat[0]), .Y(n279) );
  INVX1 U270 ( .A(prx_fifowdat[1]), .Y(n267) );
  INVX1 U271 ( .A(prx_fifowdat[2]), .Y(n278) );
  AND2X1 U272 ( .A(ordsbuf[7]), .B(ordsbuf[4]), .Y(n157) );
  NOR4XL U273 ( .A(n80), .B(cccnt[2]), .C(cccnt[5]), .D(cccnt[3]), .Y(
        prx_cccnt[1]) );
  NAND3X1 U274 ( .A(cccnt[0]), .B(cccnt[1]), .C(cccnt[4]), .Y(n80) );
  INVX1 U275 ( .A(r_ordrs4), .Y(n283) );
  NAND3X1 U276 ( .A(n171), .B(prx_fifowdat[0]), .C(n170), .Y(n103) );
  INVX1 U277 ( .A(ordsbuf[6]), .Y(n276) );
  INVX1 U278 ( .A(ordsbuf[5]), .Y(n277) );
  NAND21X1 U279 ( .B(bcnt[0]), .A(n253), .Y(n249) );
  MUX2X1 U280 ( .D0(n254), .D1(n256), .S(bcnt[1]), .Y(n262) );
  AND2X1 U281 ( .A(bcnt[0]), .B(n253), .Y(n254) );
  NAND3X1 U282 ( .A(n157), .B(n276), .C(ordsbuf[5]), .Y(n164) );
  NAND3X1 U283 ( .A(n157), .B(n277), .C(ordsbuf[6]), .Y(n144) );
  INVX1 U284 ( .A(r_rgdcrc), .Y(n137) );
  OAI22X1 U285 ( .A(n252), .B(n251), .C(n250), .D(n249), .Y(N239) );
  MUX2BXL U286 ( .D0(n250), .D1(n248), .S(bcnt[1]), .Y(n252) );
  AND2X1 U287 ( .A(bcnt[0]), .B(n250), .Y(n248) );
  AND2X1 U288 ( .A(n224), .B(prx_bmc), .Y(N156) );
  AND2X1 U289 ( .A(n224), .B(ps_dat5b[2]), .Y(N155) );
  AND2X1 U290 ( .A(n224), .B(ps_dat5b[1]), .Y(N154) );
  NAND21X1 U291 ( .B(n75), .A(prx_fsm[3]), .Y(n229) );
  AND3X1 U292 ( .A(pid_goidle), .B(cs_ords_ena), .C(prx_fsm[3]), .Y(
        prx_setsta[5]) );
  AND2X1 U293 ( .A(n221), .B(srstz), .Y(n214) );
  AND3X1 U294 ( .A(n30), .B(n219), .C(n218), .Y(n220) );
  NAND21X1 U295 ( .B(prx_fsm[0]), .A(n77), .Y(n233) );
  NAND21X1 U296 ( .B(prx_fsm[2]), .A(n120), .Y(n226) );
  OR2X1 U297 ( .A(bcnt[2]), .B(bcnt[1]), .Y(n135) );
  NAND43X1 U298 ( .B(prx_fsm[0]), .C(prx_fsm[2]), .D(n3), .A(prx_fsm[1]), .Y(
        n240) );
  INVX1 U299 ( .A(n20), .Y(prx_crcsidat[2]) );
  INVXL U300 ( .A(prx_fifowdat[6]), .Y(n20) );
  INVX1 U301 ( .A(n18), .Y(prx_crcsidat[1]) );
  INVX1 U302 ( .A(n15), .Y(prx_crcsidat[0]) );
  INVXL U303 ( .A(prx_fifowdat[4]), .Y(n15) );
  NAND21X2 U304 ( .B(n39), .A(n38), .Y(n49) );
  NOR21XL U305 ( .B(n37), .A(n52), .Y(n36) );
  NOR21X1 U306 ( .B(ps_dat5b[0]), .A(n52), .Y(n57) );
  XOR2X1 U307 ( .A(n130), .B(ps_dat5b[2]), .Y(n52) );
  INVX1 U308 ( .A(n82), .Y(n215) );
  NAND21X1 U309 ( .B(n212), .A(n213), .Y(n82) );
  INVXL U310 ( .A(n67), .Y(n17) );
  OAI211X1 U311 ( .C(n284), .D(n185), .A(n227), .B(N96), .Y(n67) );
  AND2X2 U312 ( .A(n53), .B(ps_dat5b[1]), .Y(n54) );
  INVX2 U313 ( .A(n53), .Y(n38) );
  NAND43X2 U314 ( .B(n32), .C(n31), .D(n30), .A(cctrans), .Y(n130) );
  OAI221XL U315 ( .A(prx_fifowdat[1]), .B(n206), .C(prx_fifowdat[4]), .D(n205), 
        .E(n97), .Y(n208) );
  NAND21XL U316 ( .B(n202), .A(prx_fifowdat[4]), .Y(n196) );
  AOI32XL U317 ( .A(n166), .B(n195), .C(prx_fifowdat[4]), .D(n273), .E(n181), 
        .Y(n182) );
  NAND21X2 U318 ( .B(n18), .A(prx_fifowdat[6]), .Y(n62) );
  NAND43X1 U319 ( .B(n69), .C(n20), .D(prx_fifowdat[5]), .A(n15), .Y(n118) );
  AND2XL U320 ( .A(n224), .B(n223), .Y(N157) );
  NAND31XL U321 ( .C(ps_dat5b[2]), .A(ps_dat5b[1]), .B(n223), .Y(n41) );
  NAND32XL U322 ( .B(n213), .C(n22), .A(n251), .Y(N236) );
  NAND43X1 U323 ( .B(n22), .C(n213), .D(n83), .A(n129), .Y(n251) );
  AO21XL U324 ( .B(n119), .C(n213), .A(n5), .Y(prx_crcstart) );
  AO21XL U325 ( .B(n213), .C(n227), .A(prx_setsta[6]), .Y(prx_fiforst) );
  INVX1 U326 ( .A(n117), .Y(n213) );
  NAND43X1 U327 ( .B(n70), .C(n117), .D(n22), .A(n265), .Y(n244) );
  NAND21XL U328 ( .B(n117), .A(n70), .Y(n108) );
  OA21XL U329 ( .B(prx_bmc), .C(n130), .A(n129), .Y(n133) );
  NAND32X1 U330 ( .B(n116), .C(n37), .A(n130), .Y(n51) );
  INVX3 U331 ( .A(n130), .Y(n223) );
  NAND21X1 U332 ( .B(n7), .A(n82), .Y(N250) );
  MUX2XL U333 ( .D0(shrtrans), .D1(n220), .S(cctrans), .Y(n221) );
  NAND21XL U334 ( .B(n4), .A(cctrans), .Y(n94) );
  GEN2XL U335 ( .D(n66), .E(cccnt[2]), .C(cccnt[5]), .B(cctrans), .A(n223), 
        .Y(n129) );
  AO21X4 U336 ( .B(n68), .C(n67), .A(n86), .Y(n117) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_adp ( clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, 
        r_adprx_en, r_adp2nd, adp_val, d_cc, cctrans, test_si, test_so, 
        test_se );
  output [5:0] adp_val;
  input clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, r_adprx_en,
         r_adp2nd, test_si, test_se;
  output d_cc, cctrans, test_so;
  wire   dcnt_n_2_, dcnt_n_1_, dcnt_n_0_, N49, N50, N51, N52, N53, N54, N55,
         N97, N98, N99, N100, N101, N102, N103, N104, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N169, N170, N172, N173, net10687, net10693, net10698, net10703,
         n115, n36, n37, n38, n39, n40, n44, n46, n47, n48, n56, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n81, n82, n84, n85,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n41, n42, n43, n45, n49, n50, n51, n52, n53, n54,
         n55, n57, n58, n71, n73, n74, n75, n76, n77, n78, n79, n80, n83, n86,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7;
  wire   [7:0] dcnt_h;
  wire   [5:0] adp_v0;
  wire   [5:0] dcnt_e;

  SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 clk_gate_adp_n_reg ( .CLK(clk), .EN(N49), 
        .ENCLK(net10687), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 clk_gate_dcnt_e_reg ( .CLK(clk), .EN(N130), 
        .ENCLK(net10693), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 clk_gate_dcnt_h_reg ( .CLK(clk), .EN(N137), 
        .ENCLK(net10698), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 clk_gate_dcnt_n_reg ( .CLK(clk), .EN(N169), 
        .ENCLK(net10703), .TE(test_se) );
  phyrx_adp_DW01_inc_0 add_385 ( .A(dcnt_h), .SUM({N104, N103, N102, N101, 
        N100, N99, N98, N97}) );
  phyrx_adp_DW_div_tc_6 div_338 ( .a({n4, dcnt_h}), .b({1'b0, 1'b1, 1'b1, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, adp_v0}), .remainder({SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7}), .divide_by_0() );
  SDFFQX1 dcnt_h_reg_6_ ( .D(N144), .SIN(dcnt_h[5]), .SMC(test_se), .C(
        net10698), .Q(dcnt_h[6]) );
  SDFFQX1 dcnt_h_reg_4_ ( .D(N142), .SIN(dcnt_h[3]), .SMC(test_se), .C(
        net10698), .Q(dcnt_h[4]) );
  SDFFQX1 dcnt_h_reg_5_ ( .D(N143), .SIN(dcnt_h[4]), .SMC(test_se), .C(
        net10698), .Q(dcnt_h[5]) );
  SDFFQX1 dcnt_h_reg_1_ ( .D(N139), .SIN(dcnt_h[0]), .SMC(test_se), .C(
        net10698), .Q(dcnt_h[1]) );
  SDFFQX1 dcnt_h_reg_2_ ( .D(N140), .SIN(dcnt_h[1]), .SMC(test_se), .C(
        net10698), .Q(dcnt_h[2]) );
  SDFFQX1 dcnt_h_reg_3_ ( .D(N141), .SIN(dcnt_h[2]), .SMC(test_se), .C(
        net10698), .Q(dcnt_h[3]) );
  SDFFQX1 dcnt_h_reg_0_ ( .D(N138), .SIN(dcnt_e[5]), .SMC(test_se), .C(
        net10698), .Q(dcnt_h[0]) );
  SDFFQX1 dcnt_h_reg_7_ ( .D(N145), .SIN(dcnt_h[6]), .SMC(test_se), .C(
        net10698), .Q(dcnt_h[7]) );
  SDFFQX1 adp_n_reg_5_ ( .D(N55), .SIN(adp_val[4]), .SMC(test_se), .C(net10687), .Q(adp_val[5]) );
  SDFFQX1 adp_n_reg_0_ ( .D(N50), .SIN(test_si), .SMC(test_se), .C(net10687), 
        .Q(adp_val[0]) );
  SDFFQX1 adp_n_reg_4_ ( .D(N54), .SIN(adp_val[3]), .SMC(test_se), .C(net10687), .Q(adp_val[4]) );
  SDFFQX1 cs_d_cc_reg ( .D(n115), .SIN(adp_val[5]), .SMC(test_se), .C(clk), 
        .Q(d_cc) );
  SDFFQX1 adp_n_reg_1_ ( .D(N51), .SIN(adp_val[0]), .SMC(test_se), .C(net10687), .Q(adp_val[1]) );
  SDFFQX1 dcnt_n_reg_3_ ( .D(N173), .SIN(dcnt_n_2_), .SMC(test_se), .C(
        net10703), .Q(test_so) );
  SDFFQX1 dcnt_e_reg_1_ ( .D(N132), .SIN(dcnt_e[0]), .SMC(test_se), .C(
        net10693), .Q(dcnt_e[1]) );
  SDFFQX1 adp_n_reg_3_ ( .D(N53), .SIN(adp_val[2]), .SMC(test_se), .C(net10687), .Q(adp_val[3]) );
  SDFFQX1 adp_n_reg_2_ ( .D(N52), .SIN(adp_val[1]), .SMC(test_se), .C(net10687), .Q(adp_val[2]) );
  SDFFQX1 dcnt_e_reg_2_ ( .D(N133), .SIN(dcnt_e[1]), .SMC(test_se), .C(
        net10693), .Q(dcnt_e[2]) );
  SDFFQX1 dcnt_e_reg_5_ ( .D(N136), .SIN(dcnt_e[4]), .SMC(test_se), .C(
        net10693), .Q(dcnt_e[5]) );
  SDFFQX1 dcnt_e_reg_4_ ( .D(N135), .SIN(dcnt_e[3]), .SMC(test_se), .C(
        net10693), .Q(dcnt_e[4]) );
  SDFFQX1 dcnt_n_reg_2_ ( .D(N172), .SIN(dcnt_n_1_), .SMC(test_se), .C(
        net10703), .Q(dcnt_n_2_) );
  SDFFQX1 dcnt_n_reg_1_ ( .D(n134), .SIN(dcnt_n_0_), .SMC(test_se), .C(
        net10703), .Q(dcnt_n_1_) );
  SDFFQX1 dcnt_e_reg_0_ ( .D(N131), .SIN(d_cc), .SMC(test_se), .C(net10693), 
        .Q(dcnt_e[0]) );
  SDFFQX1 dcnt_e_reg_3_ ( .D(N134), .SIN(dcnt_e[2]), .SMC(test_se), .C(
        net10693), .Q(dcnt_e[3]) );
  SDFFQX1 dcnt_n_reg_0_ ( .D(N170), .SIN(n4), .SMC(test_se), .C(net10703), .Q(
        dcnt_n_0_) );
  INVXL U5 ( .A(golo), .Y(n24) );
  INVXL U6 ( .A(gohi), .Y(n25) );
  MUX2X1 U7 ( .D0(n25), .D1(n24), .S(d_cc), .Y(n55) );
  NAND21X1 U8 ( .B(n31), .A(n30), .Y(n105) );
  INVX1 U9 ( .A(dcnt_h[7]), .Y(n3) );
  INVX1 U10 ( .A(n3), .Y(n4) );
  AND2XL U11 ( .A(adp_val[4]), .B(gohi), .Y(n23) );
  XNOR2XL U12 ( .A(n113), .B(adp_val[0]), .Y(n9) );
  OR3XL U13 ( .A(dcnt_e[2]), .B(dcnt_e[1]), .C(dcnt_e[3]), .Y(n34) );
  NOR3XL U14 ( .A(goidle), .B(gobusy), .C(n13), .Y(n72) );
  INVXL U15 ( .A(n58), .Y(n35) );
  NAND32XL U16 ( .B(n108), .C(n42), .A(n71), .Y(n83) );
  AND3XL U17 ( .A(dcnt_e[3]), .B(dcnt_e[4]), .C(n74), .Y(n76) );
  XOR2XL U18 ( .A(test_so), .B(adp_val[3]), .Y(n14) );
  XOR2XL U19 ( .A(adp_val[2]), .B(dcnt_n_2_), .Y(n15) );
  INVXL U20 ( .A(dcnt_e[0]), .Y(n108) );
  NAND2X1 U21 ( .A(n75), .B(n17), .Y(n27) );
  NAND43X1 U22 ( .B(adp_val[0]), .C(adp_val[1]), .D(adp_val[2]), .A(n16), .Y(
        n17) );
  NAND31XL U23 ( .C(n108), .A(dcnt_e[2]), .B(dcnt_e[1]), .Y(n41) );
  INVXL U24 ( .A(adp_val[3]), .Y(n16) );
  AND2XL U25 ( .A(dcnt_e[5]), .B(n42), .Y(n43) );
  NAND21XL U26 ( .B(n45), .A(dcnt_e[0]), .Y(n51) );
  OAI22AXL U27 ( .D(srstz), .C(n104), .A(dcnt_n_0_), .B(n111), .Y(N170) );
  OR4XL U28 ( .A(n19), .B(n18), .C(n27), .D(n5), .Y(n104) );
  OR4XL U29 ( .A(test_so), .B(dcnt_n_2_), .C(dcnt_n_1_), .D(dcnt_n_0_), .Y(n5)
         );
  OR2XL U30 ( .A(dcnt_e[5]), .B(n83), .Y(n78) );
  AOI211XL U31 ( .C(n113), .D(n112), .A(n111), .B(n110), .Y(n134) );
  INVXL U32 ( .A(dcnt_n_1_), .Y(n112) );
  OR4XL U33 ( .A(n7), .B(n27), .C(n13), .D(n11), .Y(n111) );
  NAND21XL U34 ( .B(dcnt_e[5]), .A(n10), .Y(n80) );
  NOR2XL U35 ( .A(n135), .B(dcnt_e[2]), .Y(n88) );
  NOR2XL U36 ( .A(dcnt_e[1]), .B(dcnt_e[0]), .Y(n100) );
  NOR2XL U37 ( .A(n82), .B(dcnt_e[4]), .Y(n81) );
  NAND2XL U38 ( .A(dcnt_n_0_), .B(dcnt_n_1_), .Y(n47) );
  INVXL U39 ( .A(dcnt_e[3]), .Y(n136) );
  INVXL U40 ( .A(dcnt_n_2_), .Y(n132) );
  INVXL U41 ( .A(dcnt_e[5]), .Y(n116) );
  INVX1 U42 ( .A(n13), .Y(n12) );
  INVX1 U43 ( .A(k0_det), .Y(n133) );
  INVX1 U44 ( .A(srstz), .Y(n13) );
  INVX1 U45 ( .A(n72), .Y(n119) );
  OAI211X1 U46 ( .C(n40), .D(n39), .A(n38), .B(n37), .Y(n85) );
  NAND2X1 U47 ( .A(n40), .B(n97), .Y(n95) );
  OR2X1 U48 ( .A(n95), .B(n93), .Y(n92) );
  OAI21X1 U49 ( .B(n96), .C(n126), .A(n91), .Y(n36) );
  OAI2B11X1 U50 ( .D(n97), .C(n36), .A(n98), .B(n95), .Y(n39) );
  NAND32X1 U51 ( .B(n40), .C(n97), .A(n36), .Y(n98) );
  OAI211X1 U52 ( .C(n93), .D(n36), .A(n94), .B(n92), .Y(n38) );
  NAND3X1 U53 ( .A(n95), .B(n36), .C(n93), .Y(n94) );
  INVX1 U54 ( .A(n96), .Y(n125) );
  INVX1 U55 ( .A(n107), .Y(n124) );
  NAND21X1 U56 ( .B(n10), .A(n58), .Y(n75) );
  INVX1 U57 ( .A(n34), .Y(n71) );
  AND2X1 U58 ( .A(n7), .B(n26), .Y(n29) );
  INVX1 U59 ( .A(n27), .Y(n28) );
  NOR32XL U60 ( .B(n91), .C(n125), .A(adp_v0[0]), .Y(n40) );
  XOR2X1 U61 ( .A(n89), .B(n90), .Y(n37) );
  OAI21BBX1 U62 ( .A(n91), .B(adp_v0[3]), .C(n125), .Y(n90) );
  NAND2X1 U63 ( .A(n36), .B(n92), .Y(n89) );
  OAI21X1 U64 ( .B(n99), .C(n126), .A(adp_v0[5]), .Y(n91) );
  NOR3XL U65 ( .A(adp_v0[1]), .B(adp_v0[3]), .C(adp_v0[2]), .Y(n99) );
  INVX1 U66 ( .A(adp_v0[4]), .Y(n126) );
  NAND2X1 U67 ( .A(n84), .B(n124), .Y(N134) );
  AOI32X1 U68 ( .A(n85), .B(n101), .C(n86), .D(n87), .E(n109), .Y(n84) );
  INVX1 U69 ( .A(n78), .Y(n101) );
  OAI21X1 U70 ( .B(n88), .C(n136), .A(n82), .Y(n87) );
  OA21X1 U71 ( .B(adp_v0[2]), .C(n96), .A(n91), .Y(n93) );
  OAI21X1 U72 ( .B(adp_v0[1]), .C(n96), .A(n91), .Y(n97) );
  NOR2X1 U73 ( .A(n126), .B(adp_v0[5]), .Y(n96) );
  NOR21XL U74 ( .B(n117), .A(n39), .Y(N51) );
  NOR21XL U75 ( .B(n117), .A(n37), .Y(N53) );
  NOR21XL U76 ( .B(n117), .A(n38), .Y(N52) );
  NOR21XL U77 ( .B(n117), .A(n40), .Y(N50) );
  AND2X1 U78 ( .A(n36), .B(n117), .Y(N54) );
  AO21X1 U79 ( .B(n109), .C(n102), .A(n119), .Y(n107) );
  AO21X1 U80 ( .B(n109), .C(n108), .A(n107), .Y(N131) );
  INVX1 U81 ( .A(n77), .Y(n86) );
  OAI31XL U82 ( .A(n81), .B(n116), .C(n103), .D(n124), .Y(N136) );
  INVX1 U83 ( .A(n103), .Y(n109) );
  INVX1 U84 ( .A(n121), .Y(n123) );
  NAND32X1 U85 ( .B(n120), .C(n119), .A(n118), .Y(n121) );
  NOR3XL U86 ( .A(n120), .B(n118), .C(n119), .Y(n6) );
  OAI221X1 U87 ( .A(n54), .B(n77), .C(n133), .D(n102), .E(n72), .Y(N130) );
  INVX1 U88 ( .A(n80), .Y(n54) );
  NAND32X1 U89 ( .B(n35), .C(n34), .A(n33), .Y(n45) );
  INVX1 U90 ( .A(n53), .Y(n33) );
  NAND43X1 U91 ( .B(n114), .C(n20), .D(n7), .A(n12), .Y(N169) );
  INVX1 U92 ( .A(n104), .Y(n20) );
  NAND21X1 U93 ( .B(n117), .A(n12), .Y(N49) );
  AND2X1 U94 ( .A(n117), .B(n116), .Y(N55) );
  NOR21XL U95 ( .B(n114), .A(n48), .Y(N172) );
  XNOR2XL U96 ( .A(n47), .B(n132), .Y(n48) );
  INVX1 U97 ( .A(n111), .Y(n114) );
  INVX1 U98 ( .A(n69), .Y(n131) );
  INVX1 U99 ( .A(n67), .Y(n130) );
  INVX1 U100 ( .A(n65), .Y(n129) );
  INVX1 U101 ( .A(n63), .Y(n128) );
  INVX1 U102 ( .A(n61), .Y(n127) );
  NAND2X1 U103 ( .A(n88), .B(n136), .Y(n82) );
  INVX1 U104 ( .A(n100), .Y(n135) );
  MUX2X1 U105 ( .D0(n23), .D1(n22), .S(d_cc), .Y(n31) );
  XOR2X1 U106 ( .A(n42), .B(dcnt_e[5]), .Y(n58) );
  NAND21X1 U107 ( .B(dcnt_e[0]), .A(n71), .Y(n49) );
  NOR41XL U108 ( .D(n8), .A(n15), .B(n14), .C(n9), .Y(n7) );
  XNOR2XL U109 ( .A(adp_val[1]), .B(dcnt_n_1_), .Y(n8) );
  NOR2X1 U110 ( .A(dcnt_e[4]), .B(n49), .Y(n10) );
  INVX1 U111 ( .A(dcnt_e[4]), .Y(n42) );
  INVX1 U112 ( .A(dcnt_n_0_), .Y(n113) );
  XOR2X1 U113 ( .A(n21), .B(d_cc), .Y(n26) );
  INVX1 U114 ( .A(n41), .Y(n74) );
  INVX1 U115 ( .A(adp_val[4]), .Y(n21) );
  AO21X1 U116 ( .B(r_adprx_en), .C(k0_det), .A(n53), .Y(n77) );
  OAI211X1 U117 ( .C(r_adp2nd), .D(n83), .A(n80), .B(n79), .Y(n103) );
  AND2X1 U118 ( .A(n86), .B(n78), .Y(n79) );
  GEN2XL U119 ( .D(n82), .E(dcnt_e[4]), .C(n81), .B(n109), .A(n107), .Y(N135)
         );
  GEN2XL U120 ( .D(n135), .E(dcnt_e[2]), .C(n88), .B(n109), .A(n107), .Y(N133)
         );
  GEN2XL U121 ( .D(dcnt_e[1]), .E(dcnt_e[0]), .C(n100), .B(n109), .A(n107), 
        .Y(N132) );
  NAND43X1 U122 ( .B(n74), .C(n52), .D(dcnt_e[3]), .A(n50), .Y(n120) );
  NOR32XL U123 ( .B(n49), .C(n45), .A(n43), .Y(n50) );
  AO22AXL U124 ( .A(N100), .B(n6), .C(n123), .D(n66), .Y(N141) );
  AOI21X1 U125 ( .B(dcnt_h[3]), .C(n130), .A(n65), .Y(n66) );
  AO22AXL U126 ( .A(N99), .B(n6), .C(n123), .D(n68), .Y(N140) );
  AOI21X1 U127 ( .B(dcnt_h[2]), .C(n131), .A(n67), .Y(n68) );
  AO22AXL U128 ( .A(N98), .B(n6), .C(n123), .D(n70), .Y(N139) );
  AOI21X1 U129 ( .B(dcnt_h[1]), .C(dcnt_h[0]), .A(n69), .Y(n70) );
  AO22AXL U130 ( .A(N102), .B(n6), .C(n123), .D(n62), .Y(N143) );
  AOI21X1 U131 ( .B(dcnt_h[5]), .C(n128), .A(n61), .Y(n62) );
  AO22AXL U132 ( .A(N101), .B(n6), .C(n123), .D(n64), .Y(N142) );
  AOI21X1 U133 ( .B(dcnt_h[4]), .C(n129), .A(n63), .Y(n64) );
  AO22AXL U134 ( .A(N103), .B(n6), .C(n123), .D(n60), .Y(N144) );
  AOI21X1 U135 ( .B(dcnt_h[6]), .C(n127), .A(n59), .Y(n60) );
  AO22AXL U136 ( .A(N104), .B(n6), .C(n123), .D(n56), .Y(N145) );
  XNOR2XL U137 ( .A(dcnt_h[7]), .B(n59), .Y(n56) );
  AO22X1 U138 ( .A(N97), .B(n6), .C(n123), .D(n122), .Y(N138) );
  INVX1 U139 ( .A(dcnt_h[0]), .Y(n122) );
  OAI31XL U140 ( .A(i_ccidle), .B(n32), .C(n78), .D(n133), .Y(n52) );
  NAND42X1 U141 ( .C(n52), .D(n119), .A(n51), .B(n120), .Y(N137) );
  INVX1 U142 ( .A(n26), .Y(n18) );
  MUX2XL U143 ( .D0(n25), .D1(n24), .S(adp_val[4]), .Y(n19) );
  INVX1 U144 ( .A(n73), .Y(n117) );
  NAND5XL U145 ( .A(n12), .B(dcnt_e[0]), .C(n71), .D(n58), .E(n57), .Y(n73) );
  AND2X1 U146 ( .A(n106), .B(n12), .Y(n115) );
  NOR4XL U147 ( .A(test_so), .B(dcnt_n_0_), .C(dcnt_n_1_), .D(dcnt_n_2_), .Y(
        n11) );
  NOR21XL U148 ( .B(n114), .A(n44), .Y(N173) );
  XNOR2XL U149 ( .A(test_so), .B(n46), .Y(n44) );
  NOR2X1 U150 ( .A(n132), .B(n47), .Y(n46) );
  NOR2X1 U151 ( .A(n131), .B(dcnt_h[2]), .Y(n67) );
  NOR2X1 U152 ( .A(n130), .B(dcnt_h[3]), .Y(n65) );
  NOR2X1 U153 ( .A(n129), .B(dcnt_h[4]), .Y(n63) );
  NOR2X1 U154 ( .A(n128), .B(dcnt_h[5]), .Y(n61) );
  NOR2X1 U155 ( .A(dcnt_h[1]), .B(dcnt_h[0]), .Y(n69) );
  INVX1 U156 ( .A(n47), .Y(n110) );
  NOR2X1 U157 ( .A(n127), .B(dcnt_h[6]), .Y(n59) );
  INVX1 U158 ( .A(d_cc), .Y(n118) );
  INVX1 U159 ( .A(r_adprx_en), .Y(n102) );
  XOR2XL U160 ( .A(n105), .B(d_cc), .Y(n106) );
  OA21X1 U161 ( .B(n76), .C(n75), .A(n105), .Y(cctrans) );
  NAND21XL U162 ( .B(i_ccidle), .A(n105), .Y(n53) );
  INVXL U163 ( .A(n105), .Y(n32) );
  MUX2BX2 U164 ( .D0(n55), .D1(n29), .S(n28), .Y(n30) );
  INVXL U165 ( .A(n55), .Y(n57) );
  AND2XL U166 ( .A(golo), .B(n21), .Y(n22) );
endmodule


module phyrx_adp_DW_div_tc_6 ( a, b, quotient, remainder, divide_by_0 );
  input [8:0] a;
  input [3:0] b;
  output [8:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   u_div_SumTmp_1__0_, u_div_SumTmp_1__2_, u_div_SumTmp_2__0_,
         u_div_SumTmp_3__0_, u_div_SumTmp_4__0_, u_div_SumTmp_5__0_,
         u_div_CryTmp_0__2_, u_div_CryTmp_0__3_, u_div_CryTmp_0__4_,
         u_div_CryTmp_1__4_, u_div_CryTmp_2__4_, u_div_CryTmp_3__4_,
         u_div_CryTmp_4__4_, u_div_CryTmp_5__4_, u_div_PartRem_1__2_,
         u_div_PartRem_1__3_, u_div_PartRem_2__3_, u_div_PartRem_3__3_,
         u_div_PartRem_4__3_, u_div_PartRem_5__3_, u_div_PartRem_7__0_,
         u_div_PartRem_7__1_, n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12,
         n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32;
  wire   [5:1] u_div_QIncCry;
  wire   [5:0] u_div_QInv;
  wire   [6:1] u_div_AIncCry;
  wire   [6:0] u_div_AInv;

  HAD1X1 u_div_u_ha_AInc_6 ( .A(u_div_AInv[6]), .B(u_div_AIncCry[6]), .CO(
        u_div_PartRem_7__1_), .SO(u_div_PartRem_7__0_) );
  HAD1X1 u_div_u_ha_AInc_5 ( .A(u_div_AInv[5]), .B(u_div_AIncCry[5]), .CO(
        u_div_AIncCry[6]), .SO(u_div_SumTmp_5__0_) );
  HAD1X1 u_div_u_ha_AInc_4 ( .A(u_div_AInv[4]), .B(u_div_AIncCry[4]), .CO(
        u_div_AIncCry[5]), .SO(u_div_SumTmp_4__0_) );
  HAD1X1 u_div_u_ha_AInc_3 ( .A(u_div_AInv[3]), .B(u_div_AIncCry[3]), .CO(
        u_div_AIncCry[4]), .SO(u_div_SumTmp_3__0_) );
  HAD1X1 u_div_u_ha_AInc_2 ( .A(u_div_AInv[2]), .B(u_div_AIncCry[2]), .CO(
        u_div_AIncCry[3]), .SO(u_div_SumTmp_2__0_) );
  HAD1X1 u_div_u_ha_AInc_1 ( .A(u_div_AInv[1]), .B(u_div_AIncCry[1]), .CO(
        u_div_AIncCry[2]), .SO(u_div_SumTmp_1__0_) );
  HAD1X1 u_div_u_ha_QInc_4 ( .A(u_div_QInv[4]), .B(u_div_QIncCry[4]), .CO(
        u_div_QIncCry[5]), .SO(quotient[4]) );
  HAD1X1 u_div_u_ha_QInc_3 ( .A(u_div_QInv[3]), .B(u_div_QIncCry[3]), .CO(
        u_div_QIncCry[4]), .SO(quotient[3]) );
  HAD1X1 u_div_u_ha_QInc_2 ( .A(u_div_QInv[2]), .B(u_div_QIncCry[2]), .CO(
        u_div_QIncCry[3]), .SO(quotient[2]) );
  HAD1X1 u_div_u_ha_QInc_1 ( .A(u_div_QInv[1]), .B(u_div_QIncCry[1]), .CO(
        u_div_QIncCry[2]), .SO(quotient[1]) );
  HAD1X1 u_div_u_ha_QInc_0 ( .A(u_div_QInv[0]), .B(a[7]), .CO(u_div_QIncCry[1]), .SO(quotient[0]) );
  XOR2X1 u_div_u_ha_QInc_5 ( .A(u_div_QInv[5]), .B(u_div_QIncCry[5]), .Y(
        quotient[5]) );
  AND2X1 u_div_u_ha_AInc_0 ( .A(u_div_AInv[0]), .B(a[8]), .Y(u_div_AIncCry[1])
         );
  INVX1 U1 ( .A(n18), .Y(n28) );
  INVX1 U2 ( .A(n19), .Y(n27) );
  INVX1 U3 ( .A(n20), .Y(n25) );
  XOR2X1 U4 ( .A(n26), .B(n25), .Y(u_div_SumTmp_1__2_) );
  NAND21X1 U5 ( .B(u_div_PartRem_3__3_), .A(n2), .Y(u_div_CryTmp_2__4_) );
  MUX2IX1 U6 ( .D0(n18), .D1(n6), .S(u_div_CryTmp_3__4_), .Y(
        u_div_PartRem_3__3_) );
  NAND2X1 U7 ( .A(n27), .B(n12), .Y(n2) );
  XNOR2XL U8 ( .A(n11), .B(n28), .Y(n6) );
  MUX2AXL U9 ( .D0(n10), .D1(n10), .S(u_div_CryTmp_4__4_), .Y(n18) );
  MUX2AXL U10 ( .D0(n11), .D1(n11), .S(u_div_CryTmp_3__4_), .Y(n19) );
  NAND21X1 U11 ( .B(u_div_PartRem_2__3_), .A(n4), .Y(u_div_CryTmp_1__4_) );
  MUX2IX1 U12 ( .D0(n19), .D1(n7), .S(u_div_CryTmp_2__4_), .Y(
        u_div_PartRem_2__3_) );
  NAND2X1 U13 ( .A(n25), .B(n26), .Y(n4) );
  XNOR2XL U14 ( .A(n12), .B(n27), .Y(n7) );
  NAND21X1 U15 ( .B(u_div_PartRem_4__3_), .A(n1), .Y(u_div_CryTmp_3__4_) );
  MUX2IX1 U16 ( .D0(n17), .D1(n5), .S(u_div_CryTmp_4__4_), .Y(
        u_div_PartRem_4__3_) );
  NAND2X1 U17 ( .A(n28), .B(n11), .Y(n1) );
  XNOR2XL U18 ( .A(n10), .B(n31), .Y(n5) );
  MUX2AXL U19 ( .D0(n12), .D1(n12), .S(u_div_CryTmp_2__4_), .Y(n20) );
  MUX2AXL U20 ( .D0(n21), .D1(n21), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__2_) );
  INVX1 U21 ( .A(u_div_CryTmp_0__3_), .Y(n23) );
  NOR21XL U22 ( .B(u_div_CryTmp_0__2_), .A(n24), .Y(u_div_CryTmp_0__3_) );
  MUX2IX1 U23 ( .D0(n32), .D1(n32), .S(u_div_CryTmp_1__4_), .Y(
        u_div_CryTmp_0__2_) );
  INVX1 U24 ( .A(u_div_PartRem_1__2_), .Y(n24) );
  INVX1 U25 ( .A(n17), .Y(n31) );
  INVX1 U26 ( .A(n21), .Y(n26) );
  MUX2AXL U27 ( .D0(u_div_PartRem_7__0_), .D1(u_div_PartRem_7__0_), .S(
        u_div_CryTmp_5__4_), .Y(n17) );
  AND2X1 U28 ( .A(u_div_PartRem_7__1_), .B(u_div_PartRem_7__0_), .Y(
        u_div_CryTmp_5__4_) );
  NAND21X1 U29 ( .B(u_div_PartRem_5__3_), .A(n3), .Y(u_div_CryTmp_4__4_) );
  MUX2IX1 U30 ( .D0(n29), .D1(n8), .S(u_div_CryTmp_5__4_), .Y(
        u_div_PartRem_5__3_) );
  NAND2X1 U31 ( .A(n31), .B(n10), .Y(n3) );
  INVX1 U32 ( .A(u_div_PartRem_7__1_), .Y(n29) );
  MUX2IX1 U33 ( .D0(u_div_SumTmp_2__0_), .D1(u_div_SumTmp_2__0_), .S(
        u_div_CryTmp_2__4_), .Y(n21) );
  MUX2X1 U34 ( .D0(u_div_SumTmp_5__0_), .D1(u_div_SumTmp_5__0_), .S(
        u_div_CryTmp_5__4_), .Y(n10) );
  MUX2X1 U35 ( .D0(u_div_SumTmp_4__0_), .D1(u_div_SumTmp_4__0_), .S(
        u_div_CryTmp_4__4_), .Y(n11) );
  MUX2X1 U36 ( .D0(u_div_SumTmp_3__0_), .D1(u_div_SumTmp_3__0_), .S(
        u_div_CryTmp_3__4_), .Y(n12) );
  XNOR2XL U37 ( .A(u_div_PartRem_7__0_), .B(u_div_PartRem_7__1_), .Y(n8) );
  INVX1 U38 ( .A(u_div_SumTmp_1__0_), .Y(n32) );
  XOR2X1 U39 ( .A(a[8]), .B(a[6]), .Y(u_div_AInv[6]) );
  XOR2X1 U40 ( .A(a[7]), .B(u_div_CryTmp_4__4_), .Y(u_div_QInv[4]) );
  XOR2X1 U41 ( .A(a[7]), .B(u_div_CryTmp_0__4_), .Y(u_div_QInv[0]) );
  NAND21X1 U42 ( .B(u_div_PartRem_1__3_), .A(n23), .Y(u_div_CryTmp_0__4_) );
  MUX2AXL U43 ( .D0(n20), .D1(u_div_SumTmp_1__2_), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__3_) );
  XOR2X1 U44 ( .A(a[8]), .B(a[2]), .Y(u_div_AInv[2]) );
  XOR2X1 U45 ( .A(a[8]), .B(a[3]), .Y(u_div_AInv[3]) );
  XOR2X1 U46 ( .A(a[8]), .B(a[4]), .Y(u_div_AInv[4]) );
  XOR2X1 U47 ( .A(a[8]), .B(a[5]), .Y(u_div_AInv[5]) );
  XOR2X1 U48 ( .A(a[7]), .B(u_div_CryTmp_1__4_), .Y(u_div_QInv[1]) );
  XOR2X1 U49 ( .A(a[7]), .B(u_div_CryTmp_2__4_), .Y(u_div_QInv[2]) );
  XOR2X1 U50 ( .A(a[7]), .B(u_div_CryTmp_3__4_), .Y(u_div_QInv[3]) );
  XOR2X1 U51 ( .A(a[8]), .B(a[1]), .Y(u_div_AInv[1]) );
  XOR2X1 U52 ( .A(a[8]), .B(a[0]), .Y(u_div_AInv[0]) );
  XNOR2XL U53 ( .A(a[7]), .B(n30), .Y(u_div_QInv[5]) );
  INVX1 U54 ( .A(u_div_CryTmp_5__4_), .Y(n30) );
endmodule


module phyrx_adp_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_db ( clk, srstz, x_cc, ptx_txact, r_rxdb_opt, gohi, golo, gotrans, 
        test_si, test_so, test_se );
  input [1:0] r_rxdb_opt;
  input clk, srstz, x_cc, ptx_txact, test_si, test_se;
  output gohi, golo, gotrans, test_so;
  wire   cc_buf_6_, cc_buf_5_, cc_buf_4_, cc_buf_3_, cc_buf_0_, N11, N12, N13,
         N14, N15, N16, N17, N18, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46;

  SDFFQX1 cc_buf_reg_3_ ( .D(N14), .SIN(n17), .SMC(test_se), .C(clk), .Q(
        cc_buf_3_) );
  SDFFQX1 cc_buf_reg_7_ ( .D(N18), .SIN(cc_buf_6_), .SMC(test_se), .C(clk), 
        .Q(test_so) );
  SDFFQX1 cc_buf_reg_5_ ( .D(N16), .SIN(cc_buf_4_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_5_) );
  SDFFQX1 cc_buf_reg_6_ ( .D(N17), .SIN(cc_buf_5_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_6_) );
  SDFFQXX2 cc_buf_reg_2_ ( .D(N13), .SIN(n2), .SMC(test_se), .C(clk), .Q(n17), 
        .XQ(n1) );
  SDFFQX1 cc_buf_reg_4_ ( .D(N15), .SIN(cc_buf_3_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_4_) );
  SDFFQXX2 cc_buf_reg_1_ ( .D(N12), .SIN(cc_buf_0_), .SMC(test_se), .C(clk), 
        .Q(n2), .XQ(n3) );
  SDFFQX1 cc_buf_reg_0_ ( .D(N11), .SIN(test_si), .SMC(test_se), .C(clk), .Q(
        cc_buf_0_) );
  MUX2X1 U3 ( .D0(n46), .D1(n45), .S(r_rxdb_opt[0]), .Y(gohi) );
  NAND2X1 U4 ( .A(n5), .B(n6), .Y(n25) );
  NAND2X1 U5 ( .A(n4), .B(cc_buf_0_), .Y(n6) );
  INVX2 U6 ( .A(n24), .Y(n4) );
  INVX1 U7 ( .A(cc_buf_3_), .Y(n10) );
  NAND2X1 U8 ( .A(n24), .B(n23), .Y(n5) );
  INVX1 U9 ( .A(n29), .Y(n28) );
  NAND21X1 U10 ( .B(n30), .A(n29), .Y(n32) );
  NAND2X2 U11 ( .A(n7), .B(n8), .Y(n24) );
  NAND2X1 U12 ( .A(n2), .B(n17), .Y(n8) );
  NAND2X1 U13 ( .A(n3), .B(n1), .Y(n7) );
  NAND21X1 U14 ( .B(n31), .A(n18), .Y(n41) );
  XNOR2X1 U15 ( .A(n35), .B(n13), .Y(n43) );
  INVXL U16 ( .A(cc_buf_6_), .Y(n16) );
  INVX1 U17 ( .A(n35), .Y(n12) );
  NAND2X1 U18 ( .A(n33), .B(n32), .Y(n13) );
  NAND2X1 U19 ( .A(n30), .B(n28), .Y(n33) );
  NAND21XL U20 ( .B(n14), .A(n27), .Y(n42) );
  AO21XL U21 ( .B(cc_buf_5_), .C(cc_buf_4_), .A(n9), .Y(n29) );
  INVXL U22 ( .A(test_so), .Y(n15) );
  XOR3XL U23 ( .A(n25), .B(cc_buf_6_), .C(test_so), .Y(n34) );
  NOR2XL U24 ( .A(n26), .B(n10), .Y(n9) );
  INVXL U25 ( .A(n41), .Y(n44) );
  AOI21XL U26 ( .B(n26), .C(n10), .A(n9), .Y(n11) );
  INVXL U27 ( .A(cc_buf_0_), .Y(n23) );
  INVXL U28 ( .A(n21), .Y(gotrans) );
  AND2XL U29 ( .A(cc_buf_6_), .B(n19), .Y(N18) );
  AND2XL U30 ( .A(cc_buf_5_), .B(n19), .Y(N17) );
  AND2XL U31 ( .A(cc_buf_4_), .B(n19), .Y(N16) );
  AND2XL U32 ( .A(cc_buf_3_), .B(n19), .Y(N15) );
  INVX1 U33 ( .A(n20), .Y(n19) );
  INVX1 U34 ( .A(srstz), .Y(n20) );
  AOI21AX1 U35 ( .B(n12), .C(n33), .A(n32), .Y(n18) );
  INVX1 U36 ( .A(n42), .Y(n31) );
  NOR21XL U37 ( .B(x_cc), .A(n20), .Y(N11) );
  NAND21X1 U38 ( .B(n34), .A(n11), .Y(n35) );
  NAND21X1 U39 ( .B(n11), .A(n34), .Y(n36) );
  AO21XL U40 ( .B(n3), .C(n23), .A(n40), .Y(n21) );
  INVX1 U41 ( .A(n22), .Y(n40) );
  MAJ3X1 U42 ( .A(n25), .B(n16), .C(n15), .Y(n14) );
  XNOR2XL U43 ( .A(cc_buf_4_), .B(cc_buf_5_), .Y(n26) );
  ENOXL U44 ( .A(n24), .B(n23), .C(n2), .D(n17), .Y(n27) );
  AND2XL U45 ( .A(cc_buf_0_), .B(n19), .Y(N12) );
  XOR2X1 U46 ( .A(n27), .B(n14), .Y(n30) );
  NAND31X1 U47 ( .C(n43), .A(n36), .B(n35), .Y(n37) );
  NAND21X2 U48 ( .B(n41), .A(n37), .Y(n38) );
  OAI22X1 U49 ( .A(n44), .B(n43), .C(n18), .D(n42), .Y(n45) );
  AND2X1 U50 ( .A(n17), .B(n19), .Y(N14) );
  AND3XL U51 ( .A(n17), .B(cc_buf_3_), .C(n40), .Y(n46) );
  NAND42XL U52 ( .C(cc_buf_3_), .D(n17), .A(n22), .B(n21), .Y(n39) );
  NOR32XL U53 ( .B(n2), .C(n19), .A(ptx_txact), .Y(N13) );
  NAND21XL U54 ( .B(n23), .A(n2), .Y(n22) );
  MUX2IX4 U55 ( .D0(n39), .D1(n38), .S(r_rxdb_opt[1]), .Y(golo) );
endmodule


module i2cslv_a0 ( i_sda, i_scl, o_sda, i_deva, i_inc, i_fwnak, i_fwack, o_we, 
        o_re, o_r_early, o_idle, o_dec, o_busev, o_ofs, o_lt_ofs, o_wdat, 
        o_lt_buf, o_dbgpo, i_rdat, i_rd_mem, i_clk, i_rstz, i_prefetch, 
        test_si, test_se );
  input [7:1] i_deva;
  output [3:0] o_busev;
  output [7:0] o_ofs;
  output [7:0] o_lt_ofs;
  output [7:0] o_wdat;
  output [7:0] o_lt_buf;
  output [7:0] o_dbgpo;
  input [7:0] i_rdat;
  input i_sda, i_scl, i_inc, i_fwnak, i_fwack, i_rd_mem, i_clk, i_rstz,
         i_prefetch, test_si, test_se;
  output o_sda, o_we, o_re, o_r_early, o_idle, o_dec;
  wire   i2c_scl, sdafall, cs_rwb, N74, N75, N76, N77, N78, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, ps_rwbuf_0_, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, net10720, net10726, net10731, net10736,
         net10741, n118, n119, n120, n121, n11, n12, n13, n14, n15, n61, n64,
         n79, n83, n88, n99, n100, n116, n124, n127, n130, n135, n1, n2, n3,
         n4, n5, n6, n8, n9, n10, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n62, n63, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n80, n81, n82, n84, n85,
         n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n117, n122, n123, n125, n126, n128, n129, n131,
         n132, n133, n134, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164;
  wire   [1:0] cs_sta;

  INVX1 U6 ( .A(n15), .Y(n12) );
  INVX1 U7 ( .A(n15), .Y(n13) );
  INVX1 U8 ( .A(n15), .Y(n14) );
  INVX1 U10 ( .A(n15), .Y(n11) );
  INVX1 U11 ( .A(i_rstz), .Y(n15) );
  i2cdbnc_a0_1 db_scl ( .i_clk(i_clk), .i_rstz(n11), .i_i2c(i_scl), .r_opt({
        1'b1, 1'b0}), .o_i2c(i2c_scl), .rise(o_dbgpo[6]), .fall(o_dbgpo[7]), 
        .test_si(cs_sta[1]), .test_se(test_se) );
  i2cdbnc_a0_0 db_sda ( .i_clk(i_clk), .i_rstz(n11), .i_i2c(i_sda), .r_opt({
        1'b0, 1'b0}), .o_i2c(ps_rwbuf_0_), .rise(o_dbgpo[5]), .fall(sdafall), 
        .test_si(i2c_scl), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 clk_gate_cs_bit_reg ( .CLK(i_clk), .EN(N74), 
        .ENCLK(net10720), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 clk_gate_adcnt_reg ( .CLK(i_clk), .EN(N114), 
        .ENCLK(net10726), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 clk_gate_rwbuf_reg ( .CLK(i_clk), .EN(N144), 
        .ENCLK(net10731), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 clk_gate_lt_buf_reg ( .CLK(i_clk), .EN(N179), .ENCLK(net10736), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 clk_gate_lt_ofs_reg ( .CLK(i_clk), .EN(
        o_busev[0]), .ENCLK(net10741), .TE(test_se) );
  SDFFSQX1 sdat_reg ( .D(n118), .SIN(o_wdat[7]), .SMC(test_se), .C(i_clk), 
        .XS(n12), .Q(o_sda) );
  SDFFQX1 lt_ofs_reg_7_ ( .D(o_wdat[7]), .SIN(o_lt_ofs[6]), .SMC(test_se), .C(
        net10741), .Q(o_lt_ofs[7]) );
  SDFFQX1 lt_ofs_reg_6_ ( .D(o_wdat[6]), .SIN(o_lt_ofs[5]), .SMC(test_se), .C(
        net10741), .Q(o_lt_ofs[6]) );
  SDFFQX1 lt_ofs_reg_0_ ( .D(o_wdat[0]), .SIN(o_lt_buf[7]), .SMC(test_se), .C(
        net10741), .Q(o_lt_ofs[0]) );
  SDFFQX1 lt_ofs_reg_1_ ( .D(o_wdat[1]), .SIN(o_lt_ofs[0]), .SMC(test_se), .C(
        net10741), .Q(o_lt_ofs[1]) );
  SDFFQX1 lt_buf_reg_7_ ( .D(N187), .SIN(o_lt_buf[6]), .SMC(test_se), .C(
        net10736), .Q(o_lt_buf[7]) );
  SDFFQX1 lt_buf_reg_6_ ( .D(N186), .SIN(o_lt_buf[5]), .SMC(test_se), .C(
        net10736), .Q(o_lt_buf[6]) );
  SDFFQX1 lt_buf_reg_3_ ( .D(N183), .SIN(o_lt_buf[2]), .SMC(test_se), .C(
        net10736), .Q(o_lt_buf[3]) );
  SDFFQX1 lt_buf_reg_1_ ( .D(N181), .SIN(o_lt_buf[0]), .SMC(test_se), .C(
        net10736), .Q(o_lt_buf[1]) );
  SDFFQX1 lt_buf_reg_0_ ( .D(N180), .SIN(ps_rwbuf_0_), .SMC(test_se), .C(
        net10736), .Q(o_lt_buf[0]) );
  SDFFQX1 lt_ofs_reg_5_ ( .D(o_wdat[5]), .SIN(o_lt_ofs[4]), .SMC(test_se), .C(
        net10741), .Q(o_lt_ofs[5]) );
  SDFFQX1 lt_ofs_reg_4_ ( .D(o_wdat[4]), .SIN(o_lt_ofs[3]), .SMC(test_se), .C(
        net10741), .Q(o_lt_ofs[4]) );
  SDFFQX1 lt_ofs_reg_3_ ( .D(o_wdat[3]), .SIN(o_lt_ofs[2]), .SMC(test_se), .C(
        net10741), .Q(o_lt_ofs[3]) );
  SDFFQX1 lt_buf_reg_5_ ( .D(N185), .SIN(o_lt_buf[4]), .SMC(test_se), .C(
        net10736), .Q(o_lt_buf[5]) );
  SDFFQX1 lt_buf_reg_4_ ( .D(N184), .SIN(o_lt_buf[3]), .SMC(test_se), .C(
        net10736), .Q(o_lt_buf[4]) );
  SDFFQX1 lt_buf_reg_2_ ( .D(N182), .SIN(o_lt_buf[1]), .SMC(test_se), .C(
        net10736), .Q(o_lt_buf[2]) );
  SDFFQX1 lt_ofs_reg_2_ ( .D(o_wdat[2]), .SIN(o_lt_ofs[1]), .SMC(test_se), .C(
        net10741), .Q(o_lt_ofs[2]) );
  SDFFRQX1 adcnt_reg_1_ ( .D(N107), .SIN(o_ofs[0]), .SMC(test_se), .C(net10726), .XR(n13), .Q(o_ofs[1]) );
  SDFFRQX1 adcnt_reg_3_ ( .D(N109), .SIN(o_ofs[2]), .SMC(test_se), .C(net10726), .XR(n13), .Q(o_ofs[3]) );
  SDFFRQX1 adcnt_reg_5_ ( .D(N111), .SIN(o_ofs[4]), .SMC(test_se), .C(net10726), .XR(n13), .Q(o_ofs[5]) );
  SDFFRQX1 adcnt_reg_6_ ( .D(N112), .SIN(o_ofs[5]), .SMC(test_se), .C(net10726), .XR(n14), .Q(o_ofs[6]) );
  SDFFRQX1 adcnt_reg_2_ ( .D(N108), .SIN(o_ofs[1]), .SMC(test_se), .C(net10726), .XR(n13), .Q(o_ofs[2]) );
  SDFFRQX1 adcnt_reg_0_ ( .D(N106), .SIN(test_si), .SMC(test_se), .C(net10726), 
        .XR(n13), .Q(o_ofs[0]) );
  SDFFRQX1 adcnt_reg_4_ ( .D(N110), .SIN(o_ofs[3]), .SMC(test_se), .C(net10726), .XR(n13), .Q(o_ofs[4]) );
  SDFFRQX1 cs_rwb_reg ( .D(n119), .SIN(o_dbgpo[3]), .SMC(test_se), .C(i_clk), 
        .XR(n13), .Q(cs_rwb) );
  SDFFRQX1 adcnt_reg_7_ ( .D(N113), .SIN(o_ofs[6]), .SMC(test_se), .C(net10726), .XR(n13), .Q(o_ofs[7]) );
  SDFFSQX1 rwbuf_reg_6_ ( .D(N142), .SIN(o_wdat[5]), .SMC(test_se), .C(
        net10731), .XS(n12), .Q(o_wdat[6]) );
  SDFFSQX1 rwbuf_reg_4_ ( .D(N140), .SIN(o_wdat[3]), .SMC(test_se), .C(
        net10731), .XS(n12), .Q(o_wdat[4]) );
  SDFFSQX1 rwbuf_reg_5_ ( .D(N141), .SIN(o_wdat[4]), .SMC(test_se), .C(
        net10731), .XS(n12), .Q(o_wdat[5]) );
  SDFFSQX1 rwbuf_reg_1_ ( .D(N137), .SIN(o_wdat[0]), .SMC(test_se), .C(
        net10731), .XS(n13), .Q(o_wdat[1]) );
  SDFFSQX1 rwbuf_reg_3_ ( .D(N139), .SIN(o_wdat[2]), .SMC(test_se), .C(
        net10731), .XS(n12), .Q(o_wdat[3]) );
  SDFFSQX1 rwbuf_reg_7_ ( .D(N143), .SIN(o_wdat[6]), .SMC(test_se), .C(
        net10731), .XS(n11), .Q(o_wdat[7]) );
  SDFFSQX1 rwbuf_reg_0_ ( .D(N136), .SIN(o_lt_ofs[7]), .SMC(test_se), .C(
        net10731), .XS(n11), .Q(o_wdat[0]) );
  SDFFSQX1 cs_bit_reg_0_ ( .D(N75), .SIN(o_ofs[7]), .SMC(test_se), .C(net10720), .XS(n12), .Q(o_dbgpo[0]) );
  SDFFSQX1 cs_bit_reg_2_ ( .D(N77), .SIN(o_dbgpo[1]), .SMC(test_se), .C(
        net10720), .XS(n12), .Q(o_dbgpo[2]) );
  SDFFSQX1 rwbuf_reg_2_ ( .D(N138), .SIN(o_wdat[1]), .SMC(test_se), .C(
        net10731), .XS(n12), .Q(o_wdat[2]) );
  SDFFSQX1 cs_bit_reg_1_ ( .D(N76), .SIN(o_dbgpo[0]), .SMC(test_se), .C(
        net10720), .XS(n12), .Q(o_dbgpo[1]) );
  SDFFSQX1 cs_bit_reg_3_ ( .D(N78), .SIN(o_dbgpo[2]), .SMC(test_se), .C(
        net10720), .XS(n12), .Q(o_dbgpo[3]) );
  SDFFRQX1 cs_sta_reg_1_ ( .D(n121), .SIN(cs_sta[0]), .SMC(test_se), .C(i_clk), 
        .XR(n14), .Q(cs_sta[1]) );
  SDFFRQX1 cs_sta_reg_0_ ( .D(n120), .SIN(cs_rwb), .SMC(test_se), .C(i_clk), 
        .XR(n13), .Q(cs_sta[0]) );
  OA21X1 U3 ( .B(n151), .C(n150), .A(n149), .Y(n152) );
  INVX1 U4 ( .A(n140), .Y(n41) );
  INVX1 U5 ( .A(n82), .Y(n148) );
  INVX1 U9 ( .A(n90), .Y(n89) );
  INVX1 U12 ( .A(n25), .Y(o_busev[0]) );
  INVX1 U13 ( .A(o_dbgpo[7]), .Y(n160) );
  AOI21X1 U14 ( .B(n112), .C(n104), .A(n111), .Y(n1) );
  AOI21X1 U15 ( .B(n112), .C(n109), .A(n111), .Y(n2) );
  AOI21X1 U16 ( .B(n112), .C(n125), .A(n111), .Y(n3) );
  NAND21X1 U17 ( .B(n144), .A(n158), .Y(n91) );
  AOI21X1 U18 ( .B(n112), .C(n101), .A(n111), .Y(n4) );
  OR2X1 U19 ( .A(n158), .B(n64), .Y(N74) );
  INVX1 U20 ( .A(n73), .Y(n26) );
  AND2X1 U21 ( .A(n111), .B(n144), .Y(o_dec) );
  BUFX3 U22 ( .A(o_busev[3]), .Y(o_dbgpo[4]) );
  NAND5XL U23 ( .A(o_busev[1]), .B(n58), .C(n56), .D(n59), .E(n18), .Y(n140)
         );
  AND4X1 U24 ( .A(n53), .B(n57), .C(n55), .D(n54), .Y(n18) );
  INVX1 U25 ( .A(o_dbgpo[6]), .Y(n69) );
  INVX1 U26 ( .A(n17), .Y(o_busev[1]) );
  NAND32X1 U27 ( .B(n145), .C(n69), .A(n111), .Y(n17) );
  AND3X1 U28 ( .A(o_dbgpo[6]), .B(n112), .C(n46), .Y(o_re) );
  MUX2X1 U29 ( .D0(n43), .D1(n131), .S(i_prefetch), .Y(o_r_early) );
  MUX2X1 U30 ( .D0(n45), .D1(n143), .S(i_prefetch), .Y(n46) );
  INVX1 U31 ( .A(n42), .Y(n131) );
  NAND21X1 U32 ( .B(n44), .A(n41), .Y(n42) );
  NAND21X1 U33 ( .B(n95), .A(n144), .Y(n82) );
  AND4X1 U34 ( .A(o_dbgpo[6]), .B(n111), .C(n40), .D(n148), .Y(n43) );
  INVX1 U35 ( .A(n68), .Y(n40) );
  INVX1 U36 ( .A(n96), .Y(n144) );
  INVX1 U37 ( .A(n146), .Y(n111) );
  INVX1 U38 ( .A(n48), .Y(n51) );
  AND2X1 U39 ( .A(n148), .B(n44), .Y(n45) );
  INVX1 U40 ( .A(n142), .Y(o_we) );
  INVX1 U41 ( .A(n126), .Y(n112) );
  INVX1 U42 ( .A(n93), .Y(n30) );
  MUX2AXL U43 ( .D0(n5), .D1(n100), .S(n148), .Y(n149) );
  AOI21X1 U44 ( .B(n151), .C(n147), .A(n146), .Y(n5) );
  NAND32X1 U45 ( .B(n69), .C(n97), .A(n96), .Y(n90) );
  INVX1 U46 ( .A(i_rd_mem), .Y(n159) );
  ENOX1 U47 ( .A(n139), .B(n90), .C(n97), .D(i_rdat[7]), .Y(N143) );
  OA21X1 U48 ( .B(n89), .C(n97), .A(n88), .Y(N144) );
  NAND32X1 U49 ( .B(n145), .C(n117), .A(o_dbgpo[7]), .Y(n25) );
  NAND21X1 U50 ( .B(i_prefetch), .A(n68), .Y(n147) );
  INVX1 U51 ( .A(n127), .Y(n104) );
  INVX1 U52 ( .A(n79), .Y(o_busev[2]) );
  INVX1 U53 ( .A(n61), .Y(o_busev[3]) );
  OR4X1 U54 ( .A(n69), .B(o_dbgpo[7]), .C(n146), .D(n147), .Y(n72) );
  NAND2X1 U55 ( .A(n61), .B(n79), .Y(n64) );
  INVX1 U56 ( .A(n76), .Y(n86) );
  GEN2XL U57 ( .D(n153), .E(o_dbgpo[7]), .C(n75), .B(n144), .A(n74), .Y(n76)
         );
  NAND21X1 U58 ( .B(n64), .A(n73), .Y(n74) );
  INVX1 U59 ( .A(n72), .Y(n75) );
  INVX1 U60 ( .A(n130), .Y(n109) );
  INVX1 U61 ( .A(n135), .Y(n125) );
  INVX1 U62 ( .A(n145), .Y(n151) );
  INVX1 U63 ( .A(n53), .Y(n65) );
  INVX1 U64 ( .A(n54), .Y(n63) );
  INVX1 U65 ( .A(n55), .Y(n62) );
  NAND21X1 U66 ( .B(n146), .A(o_dbgpo[7]), .Y(n73) );
  GEN2XL U67 ( .D(n144), .E(n95), .C(n29), .B(n28), .A(n27), .Y(N114) );
  AND2X1 U68 ( .A(n112), .B(o_dbgpo[7]), .Y(n28) );
  NAND21X1 U69 ( .B(n26), .A(n25), .Y(n27) );
  MUX2X1 U70 ( .D0(n143), .D1(n24), .S(i_prefetch), .Y(n29) );
  NAND21X1 U71 ( .B(n41), .A(n142), .Y(N179) );
  OR2X1 U72 ( .A(n94), .B(n6), .Y(N76) );
  AOI21X1 U73 ( .B(n93), .C(n92), .A(n91), .Y(n6) );
  INVX1 U74 ( .A(n47), .Y(n158) );
  NAND32X1 U75 ( .B(n160), .C(o_idle), .A(n88), .Y(n47) );
  OAI22X1 U76 ( .A(n142), .B(n133), .C(n140), .D(n132), .Y(N181) );
  OAI22X1 U77 ( .A(n142), .B(n134), .C(n140), .D(n133), .Y(N182) );
  OAI22X1 U78 ( .A(n142), .B(n136), .C(n140), .D(n134), .Y(N183) );
  OAI22X1 U79 ( .A(n142), .B(n137), .C(n140), .D(n136), .Y(N184) );
  OAI22X1 U80 ( .A(n142), .B(n138), .C(n140), .D(n137), .Y(N185) );
  OAI22X1 U81 ( .A(n142), .B(n139), .C(n140), .D(n138), .Y(N186) );
  OAI22X1 U82 ( .A(n142), .B(n141), .C(n140), .D(n139), .Y(N187) );
  INVX1 U83 ( .A(n49), .Y(n94) );
  NAND21X1 U84 ( .B(n61), .A(n79), .Y(n49) );
  INVX1 U85 ( .A(i_inc), .Y(n101) );
  INVX1 U86 ( .A(n117), .Y(n129) );
  NAND43X1 U87 ( .B(o_dbgpo[3]), .C(o_dbgpo[2]), .D(o_dbgpo[1]), .A(o_dbgpo[0]), .Y(n145) );
  NAND43X1 U88 ( .B(n39), .C(n38), .D(n37), .A(n36), .Y(n68) );
  XOR2X1 U89 ( .A(i_deva[1]), .B(o_wdat[1]), .Y(n39) );
  NOR32XL U90 ( .B(n35), .C(n34), .A(n33), .Y(n36) );
  XOR2X1 U91 ( .A(i_deva[3]), .B(o_wdat[3]), .Y(n38) );
  NAND21X1 U92 ( .B(o_dbgpo[3]), .A(n51), .Y(n96) );
  NAND21X1 U93 ( .B(cs_sta[0]), .A(n153), .Y(n146) );
  NAND21X1 U94 ( .B(o_dbgpo[0]), .A(n21), .Y(n92) );
  XOR2X1 U95 ( .A(n134), .B(i_deva[3]), .Y(n54) );
  XOR2X1 U96 ( .A(n138), .B(i_deva[6]), .Y(n55) );
  XOR2X1 U97 ( .A(n132), .B(i_deva[1]), .Y(n53) );
  OR2X1 U98 ( .A(o_dbgpo[2]), .B(n92), .Y(n48) );
  NAND21X1 U99 ( .B(n32), .A(n31), .Y(n33) );
  XNOR2XL U100 ( .A(i_deva[7]), .B(o_wdat[7]), .Y(n31) );
  XOR2X1 U101 ( .A(i_deva[5]), .B(o_wdat[5]), .Y(n32) );
  XOR2X1 U102 ( .A(n139), .B(i_deva[7]), .Y(n56) );
  XOR2X1 U103 ( .A(n136), .B(i_deva[4]), .Y(n59) );
  XOR2X1 U104 ( .A(n137), .B(i_deva[5]), .Y(n58) );
  XOR2X1 U105 ( .A(n133), .B(i_deva[2]), .Y(n57) );
  XOR2X1 U106 ( .A(n139), .B(i_deva[6]), .Y(n35) );
  XOR2X1 U107 ( .A(n137), .B(i_deva[4]), .Y(n34) );
  XOR2X1 U108 ( .A(o_wdat[2]), .B(i_deva[2]), .Y(n37) );
  INVX1 U109 ( .A(cs_sta[1]), .Y(n153) );
  INVX1 U110 ( .A(o_dbgpo[1]), .Y(n21) );
  INVX1 U111 ( .A(n23), .Y(n143) );
  NAND21X1 U112 ( .B(n145), .A(cs_rwb), .Y(n23) );
  INVX1 U113 ( .A(o_wdat[6]), .Y(n139) );
  INVX1 U114 ( .A(o_wdat[4]), .Y(n137) );
  INVX1 U115 ( .A(o_wdat[2]), .Y(n134) );
  INVX1 U116 ( .A(o_wdat[5]), .Y(n138) );
  INVX1 U117 ( .A(o_wdat[1]), .Y(n133) );
  INVX1 U118 ( .A(o_wdat[3]), .Y(n136) );
  INVX1 U119 ( .A(o_wdat[0]), .Y(n132) );
  NAND43X1 U120 ( .B(cs_rwb), .C(n126), .D(n145), .A(o_dbgpo[7]), .Y(n142) );
  NAND21X1 U121 ( .B(cs_sta[0]), .A(cs_sta[1]), .Y(n126) );
  INVX1 U122 ( .A(cs_rwb), .Y(n95) );
  INVX1 U123 ( .A(ps_rwbuf_0_), .Y(n44) );
  NAND21X1 U124 ( .B(n66), .A(o_dbgpo[1]), .Y(n93) );
  AND3X1 U125 ( .A(o_dbgpo[3]), .B(o_dbgpo[2]), .C(n30), .Y(o_idle) );
  INVX1 U126 ( .A(o_dbgpo[0]), .Y(n66) );
  AOI22X1 U127 ( .A(i_rd_mem), .B(i_rdat[7]), .C(n159), .D(o_wdat[7]), .Y(n100) );
  AOI221XL U128 ( .A(ps_rwbuf_0_), .B(n144), .C(n99), .D(n145), .E(n143), .Y(
        n154) );
  NAND2X1 U129 ( .A(n100), .B(cs_rwb), .Y(n99) );
  MUX2X1 U130 ( .D0(n157), .D1(n156), .S(n160), .Y(n118) );
  MUX3X1 U131 ( .D0(o_sda), .D1(i_rdat[7]), .D2(i_fwnak), .S0(n155), .S1(n83), 
        .Y(n156) );
  OAI211X1 U132 ( .C(n154), .D(n153), .A(n88), .B(n152), .Y(n157) );
  XOR2X1 U133 ( .A(i_fwnak), .B(i_fwack), .Y(n83) );
  NAND21X1 U134 ( .B(n155), .A(n22), .Y(n97) );
  NAND43X1 U135 ( .B(n116), .C(o_dbgpo[3]), .D(o_dbgpo[2]), .A(n21), .Y(n22)
         );
  NAND3X1 U136 ( .A(cs_rwb), .B(n88), .C(i_rd_mem), .Y(n116) );
  AO22X1 U137 ( .A(n89), .B(o_wdat[3]), .C(i_rdat[4]), .D(n97), .Y(N140) );
  AO22X1 U138 ( .A(n89), .B(o_wdat[2]), .C(i_rdat[3]), .D(n97), .Y(N139) );
  AO22X1 U139 ( .A(n89), .B(o_wdat[1]), .C(i_rdat[2]), .D(n97), .Y(N138) );
  AO22X1 U140 ( .A(n89), .B(o_wdat[0]), .C(i_rdat[1]), .D(n97), .Y(N137) );
  AO22X1 U141 ( .A(n89), .B(o_wdat[5]), .C(i_rdat[6]), .D(n97), .Y(N142) );
  INVX1 U142 ( .A(n20), .Y(n155) );
  NAND6XL U143 ( .A(o_dbgpo[3]), .B(cs_rwb), .C(n88), .D(n51), .E(n19), .F(
        i_rd_mem), .Y(n20) );
  INVX1 U144 ( .A(i2c_scl), .Y(n19) );
  OAI21BBX1 U145 ( .A(i_rdat[0]), .B(n97), .C(n8), .Y(N136) );
  NAND4X1 U146 ( .A(o_dbgpo[6]), .B(ps_rwbuf_0_), .C(n96), .D(n95), .Y(n8) );
  NOR32XL U147 ( .B(o_ofs[2]), .C(n135), .A(n162), .Y(n130) );
  NOR32XL U148 ( .B(o_ofs[0]), .C(i_inc), .A(n161), .Y(n135) );
  NOR32XL U149 ( .B(o_ofs[4]), .C(n130), .A(n163), .Y(n127) );
  NAND3X1 U150 ( .A(i2c_scl), .B(n160), .C(sdafall), .Y(n79) );
  AO21X1 U151 ( .B(n129), .C(o_wdat[6]), .A(n105), .Y(N112) );
  OAI32X1 U152 ( .A(n126), .B(n104), .C(o_ofs[6]), .D(n1), .E(n103), .Y(n105)
         );
  INVX1 U153 ( .A(o_ofs[6]), .Y(n103) );
  NAND3X1 U154 ( .A(i2c_scl), .B(n160), .C(o_dbgpo[5]), .Y(n61) );
  OAI222XL U155 ( .A(n164), .B(n1), .C(n80), .D(n126), .E(n141), .F(n117), .Y(
        N113) );
  MUX2BXL U156 ( .D0(o_ofs[6]), .D1(n78), .S(n164), .Y(n80) );
  INVX1 U157 ( .A(o_ofs[7]), .Y(n164) );
  AND2X1 U158 ( .A(o_ofs[6]), .B(n127), .Y(n78) );
  INVX1 U159 ( .A(o_ofs[1]), .Y(n161) );
  NAND21X1 U160 ( .B(cs_sta[1]), .A(cs_sta[0]), .Y(n117) );
  AO21X1 U161 ( .B(n70), .C(n72), .A(n64), .Y(n81) );
  NAND5XL U162 ( .A(n124), .B(o_dbgpo[1]), .C(i_prefetch), .D(n67), .E(n66), 
        .Y(n70) );
  NAND43X1 U163 ( .B(n65), .C(n63), .D(n62), .A(n60), .Y(n67) );
  AND4X1 U164 ( .A(n59), .B(n58), .C(n57), .D(n56), .Y(n60) );
  MUX2X1 U165 ( .D0(n77), .D1(cs_sta[0]), .S(n86), .Y(n120) );
  NAND21X1 U166 ( .B(n71), .A(n81), .Y(n77) );
  AND4X1 U167 ( .A(n144), .B(n150), .C(n95), .D(n52), .Y(n71) );
  INVX1 U168 ( .A(n64), .Y(n52) );
  MUX2X1 U169 ( .D0(n87), .D1(cs_sta[1]), .S(n86), .Y(n121) );
  NAND21X1 U170 ( .B(n85), .A(n84), .Y(n87) );
  AO21X1 U171 ( .B(n82), .C(n150), .A(n64), .Y(n84) );
  INVX1 U172 ( .A(n81), .Y(n85) );
  NAND2X1 U173 ( .A(cs_sta[0]), .B(cs_sta[1]), .Y(n88) );
  OAI222XL U174 ( .A(n163), .B(n2), .C(n107), .D(n126), .E(n138), .F(n117), 
        .Y(N111) );
  MUX2BXL U175 ( .D0(o_ofs[4]), .D1(n106), .S(n163), .Y(n107) );
  AND2X1 U176 ( .A(o_ofs[4]), .B(n130), .Y(n106) );
  AO21X1 U177 ( .B(n129), .C(o_wdat[4]), .A(n110), .Y(N110) );
  OAI32X1 U178 ( .A(n126), .B(n109), .C(o_ofs[4]), .D(n2), .E(n108), .Y(n110)
         );
  INVX1 U179 ( .A(o_ofs[4]), .Y(n108) );
  AO21X1 U180 ( .B(n129), .C(o_wdat[2]), .A(n128), .Y(N108) );
  OAI32X1 U181 ( .A(n126), .B(n125), .C(o_ofs[2]), .D(n3), .E(n123), .Y(n128)
         );
  INVX1 U182 ( .A(o_ofs[2]), .Y(n123) );
  INVX1 U183 ( .A(o_ofs[3]), .Y(n162) );
  GEN2XL U184 ( .D(o_dbgpo[3]), .E(n48), .C(n144), .B(n158), .A(n64), .Y(N78)
         );
  GEN2XL U185 ( .D(o_dbgpo[2]), .E(n92), .C(n51), .B(n50), .A(n94), .Y(N77) );
  INVX1 U186 ( .A(n91), .Y(n50) );
  MUX2BXL U187 ( .D0(ps_rwbuf_0_), .D1(n9), .S(n10), .Y(n119) );
  NAND2X1 U188 ( .A(cs_rwb), .B(n79), .Y(n9) );
  NAND2X1 U189 ( .A(n79), .B(o_busev[1]), .Y(n10) );
  AO21X1 U190 ( .B(o_wdat[0]), .C(o_we), .A(n131), .Y(N180) );
  OAI222XL U191 ( .A(n162), .B(n3), .C(n114), .D(n126), .E(n136), .F(n117), 
        .Y(N109) );
  MUX2BXL U192 ( .D0(o_ofs[2]), .D1(n113), .S(n162), .Y(n114) );
  AND2X1 U193 ( .A(o_ofs[2]), .B(n135), .Y(n113) );
  OAI222XL U194 ( .A(n161), .B(n4), .C(n122), .D(n126), .E(n133), .F(n117), 
        .Y(N107) );
  MUX2BXL U195 ( .D0(o_ofs[0]), .D1(n115), .S(n161), .Y(n122) );
  AND2X1 U196 ( .A(o_ofs[0]), .B(i_inc), .Y(n115) );
  AO21X1 U197 ( .B(n129), .C(o_wdat[0]), .A(n102), .Y(N106) );
  OAI32X1 U198 ( .A(n126), .B(n101), .C(o_ofs[0]), .D(n4), .E(n98), .Y(n102)
         );
  INVX1 U199 ( .A(o_ofs[0]), .Y(n98) );
  INVX1 U200 ( .A(o_ofs[5]), .Y(n163) );
  OAI21AX1 U201 ( .B(o_dbgpo[0]), .C(n91), .A(n64), .Y(N75) );
  NOR2X1 U202 ( .A(o_dbgpo[3]), .B(o_dbgpo[2]), .Y(n124) );
  AND4X1 U203 ( .A(o_dbgpo[1]), .B(cs_rwb), .C(n124), .D(n66), .Y(n24) );
  INVX1 U204 ( .A(cs_sta[0]), .Y(n150) );
  INVX1 U205 ( .A(o_wdat[7]), .Y(n141) );
  AO22XL U206 ( .A(n89), .B(o_wdat[4]), .C(i_rdat[5]), .D(n97), .Y(N141) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2cdbnc_a0_0 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall, test_si, 
        test_se );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c, test_si, test_se;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n7, n5, n6, n8, n1, n2;

  SDFFSQX1 d_i2c_reg_2_ ( .D(N19), .SIN(N19), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(d_i2c_2_) );
  SDFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .SIN(test_si), .SMC(test_se), .C(i_clk), 
        .XS(i_rstz), .Q(N18) );
  SDFFSQX1 d_i2c_reg_1_ ( .D(N18), .SIN(N18), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(N19) );
  SDFFSQXX1 r_i2c_reg ( .D(n7), .SIN(d_i2c_2_), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(o_i2c), .XQ(n1) );
  OAI21X1 U3 ( .B(fall), .C(n1), .A(n5), .Y(n7) );
  OAI211X1 U4 ( .C(r_opt[0]), .D(d_i2c_2_), .A(n1), .B(n6), .Y(n5) );
  AND2X1 U5 ( .A(N18), .B(N19), .Y(n6) );
  INVX1 U6 ( .A(n5), .Y(rise) );
  AOI211X1 U7 ( .C(n2), .D(d_i2c_2_), .A(n1), .B(n8), .Y(fall) );
  INVX1 U8 ( .A(r_opt[1]), .Y(n2) );
  OR2X1 U9 ( .A(N19), .B(N18), .Y(n8) );
endmodule


module i2cdbnc_a0_1 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall, test_si, 
        test_se );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c, test_si, test_se;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n6, n1, n2, n3, n4;

  SDFFSQX1 d_i2c_reg_1_ ( .D(N18), .SIN(N18), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(N19) );
  SDFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .SIN(test_si), .SMC(test_se), .C(i_clk), 
        .XS(i_rstz), .Q(N18) );
  SDFFSQX1 d_i2c_reg_2_ ( .D(N19), .SIN(N19), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(d_i2c_2_) );
  SDFFSQXX1 r_i2c_reg ( .D(n6), .SIN(d_i2c_2_), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(o_i2c), .XQ(n3) );
  INVX1 U3 ( .A(n4), .Y(fall) );
  NOR43XL U4 ( .B(N18), .C(N19), .D(n3), .A(n2), .Y(rise) );
  NOR2X1 U5 ( .A(r_opt[0]), .B(d_i2c_2_), .Y(n2) );
  NAND42X1 U6 ( .C(N19), .D(N18), .A(n1), .B(o_i2c), .Y(n4) );
  NAND21X1 U7 ( .B(r_opt[1]), .A(d_i2c_2_), .Y(n1) );
  AO21X1 U8 ( .B(o_i2c), .C(n4), .A(rise), .Y(n6) );
endmodule


module regbank_a0 ( srci, dm_fault, cc1_di, cc2_di, di_rd_det, di_stbovp, 
        i_tmrf, i_vcbyval, dnchk_en, r_pwrv_upd, aswkup, ps_pwrdn, r_sleep, 
        r_pwrdn, r_ocdrv_enz, r_osc_stop, r_osc_lo, r_osc_gate, r_fw_pwrv, 
        r_cvcwr, r_cvofs, r_otpi_gate, r_pwrctl, r_pwr_i, r_cvctl, r_srcctl, 
        r_dpdmctl, r_ccrx, r_cctrx, r_ccctl, r_fcpwr, r_fcpre, fcp_r_dat, 
        fcp_r_sta, fcp_r_msk, fcp_r_ctl, fcp_r_crc, fcp_r_acc, fcp_r_tui, 
        r_accctl, r_bclk_sel, r_dacwr, r_dac_en, r_sar_en, r_adofs, r_isofs, 
        x_daclsb, r_comp_opt, dac_r_ctl, dac_r_comp, dac_r_cmpsta, dac_r_vs, 
        REVID, atpg_en, sfr_r, sfr_w, set_hold, bkpt_hold, cpurst, sfr_addr, 
        sfr_wdat, sfr_rdat, ff_p0, di_p0, ictlr_idle, ictlr_inc, r_inst_ofs, 
        r_psrd, r_pswr, r_fortxdat, r_fortxrdy, r_fortxen, r_ana_tm, r_gpio_tm, 
        r_gpio_ie, r_gpio_oe, r_gpio_pu, r_gpio_pd, r_gpio_s0, r_gpio_s1, 
        r_gpio_s2, r_gpio_s3, r_regtrm, i_pc, i_goidle, i_gobusy, i_i2c_idle, 
        bus_idle, i2c_stretch, i_i2c_rwbuf, i_i2c_ltbuf, i_i2c_ofs, o_intr, 
        r_auto_gdcrc, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, r_unlock, 
        r_first, r_last, r_fiforst, r_set_cpmsgid, r_txendk, r_txnumk, 
        r_txshrt, r_auto_discard, r_hold_mcu, r_txauto, r_rxords_ena, r_spec, 
        r_dat_spec, r_dat_portrole, r_dat_datarole, r_discard, r_pshords, 
        r_pg0_sel, r_strtch, r_i2c_attr, r_i2c_ninc, r_hwi2c_en, r_i2c_fwnak, 
        r_i2c_fwack, r_i2c_deva, i2c_ev, prl_c0set, prl_cany0, prl_discard, 
        prl_GCTxDone, prl_cpmsgid, pff_ack, prx_rst, pff_obsd, pff_full, 
        pff_empty, ptx_ack, pff_ptr, prx_adpn, pff_rdat, pff_rxpart, 
        prx_rcvinf, ptx_fsm, prx_fsm, prl_fsm, prx_setsta, clk_1500k, clk_500k, 
        clk_500, clk, xrstz, xclk, dbgpo, srstz, prstz, test_si2, test_si1, 
        test_so2, test_so1, test_se );
  input [5:0] srci;
  output [11:0] r_fw_pwrv;
  output [1:0] r_cvcwr;
  input [15:0] r_cvofs;
  output [7:4] r_pwrctl;
  output [7:0] r_pwr_i;
  output [7:0] r_cvctl;
  output [7:0] r_srcctl;
  output [7:0] r_dpdmctl;
  output [7:0] r_ccrx;
  output [7:0] r_cctrx;
  output [7:0] r_ccctl;
  output [6:0] r_fcpwr;
  input [7:0] fcp_r_dat;
  input [7:0] fcp_r_sta;
  input [7:0] fcp_r_msk;
  input [7:0] fcp_r_ctl;
  input [7:0] fcp_r_crc;
  input [7:0] fcp_r_acc;
  input [7:0] fcp_r_tui;
  input [7:0] r_accctl;
  output [14:0] r_dacwr;
  input [7:0] r_dac_en;
  input [7:0] r_sar_en;
  input [7:0] r_adofs;
  input [7:0] r_isofs;
  input [5:0] x_daclsb;
  output [7:0] r_comp_opt;
  input [7:0] dac_r_ctl;
  input [7:0] dac_r_comp;
  input [7:0] dac_r_cmpsta;
  input [63:0] dac_r_vs;
  input [6:0] REVID;
  input [7:0] sfr_addr;
  input [7:0] sfr_wdat;
  output [7:0] sfr_rdat;
  input [7:0] ff_p0;
  input [7:0] di_p0;
  output [14:0] r_inst_ofs;
  output [3:0] r_ana_tm;
  output [1:0] r_gpio_ie;
  output [6:0] r_gpio_oe;
  output [6:0] r_gpio_pu;
  output [6:0] r_gpio_pd;
  output [2:0] r_gpio_s0;
  output [2:0] r_gpio_s1;
  output [2:0] r_gpio_s2;
  output [2:0] r_gpio_s3;
  output [55:0] r_regtrm;
  input [15:0] i_pc;
  input [7:0] i_i2c_rwbuf;
  input [7:0] i_i2c_ltbuf;
  input [7:0] i_i2c_ofs;
  output [4:0] o_intr;
  output [1:0] r_auto_gdcrc;
  output [4:0] r_txnumk;
  output [6:0] r_txauto;
  output [6:0] r_rxords_ena;
  output [1:0] r_spec;
  output [1:0] r_dat_spec;
  output [3:0] r_pg0_sel;
  output [7:1] r_i2c_deva;
  input [7:0] i2c_ev;
  input [2:0] prl_cpmsgid;
  input [1:0] pff_ack;
  input [1:0] prx_rst;
  input [5:0] pff_ptr;
  input [5:0] prx_adpn;
  input [7:0] pff_rdat;
  input [15:0] pff_rxpart;
  input [4:0] prx_rcvinf;
  input [2:0] ptx_fsm;
  input [3:0] prx_fsm;
  input [3:0] prl_fsm;
  input [6:0] prx_setsta;
  output [31:0] dbgpo;
  input dm_fault, cc1_di, cc2_di, di_rd_det, di_stbovp, i_tmrf, i_vcbyval,
         dnchk_en, atpg_en, sfr_r, sfr_w, set_hold, bkpt_hold, cpurst,
         ictlr_idle, ictlr_inc, i_goidle, i_gobusy, i_i2c_idle, prl_c0set,
         prl_cany0, prl_discard, prl_GCTxDone, pff_obsd, pff_full, pff_empty,
         ptx_ack, clk_1500k, clk_500k, clk_500, clk, xrstz, xclk, test_si2,
         test_si1, test_se;
  output r_pwrv_upd, aswkup, ps_pwrdn, r_sleep, r_pwrdn, r_ocdrv_enz,
         r_osc_stop, r_osc_lo, r_osc_gate, r_otpi_gate, r_fcpre, r_bclk_sel,
         r_psrd, r_pswr, r_fortxdat, r_fortxrdy, r_fortxen, r_gpio_tm,
         bus_idle, i2c_stretch, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop,
         r_unlock, r_first, r_last, r_fiforst, r_set_cpmsgid, r_txendk,
         r_txshrt, r_auto_discard, r_hold_mcu, r_dat_portrole, r_dat_datarole,
         r_discard, r_pshords, r_strtch, r_i2c_attr, r_i2c_ninc, r_hwi2c_en,
         r_i2c_fwnak, r_i2c_fwack, srstz, prstz, test_so2, test_so1;
  wire   we_246, we_245, we_232, we_231, we_230, we_228, we_227, we_222,
         we_217, we_215, we_214, we_213, we_211, we_209, we_203, we_191,
         we_187, we_182, we_181, we_176, we_175, we_172, we_171, we_148,
         we_143, regF4_7_, regF4_3, regE3_0, regD4_6_, regD4_5_, regD4_4_,
         regD4_3_, regD4_2_, regD4_1_, regD4_0_, regD3_7_, regD3_3, reg25_0_,
         reg19_7_, reg12_1, reg11_7_, reg11_4, regAD_7, N23, N24, N25, N26,
         N27, N29, N30, N31, N32, N33, N34, N35, N36, upd01, phyrst, upd12,
         upd18, upd19, upd20, upd21, lt_reg26_0, i2c_mode_upd, i2c_mode_wdat,
         upd31, N81, as_p0_chg, dmf_wkup, p0_chg_clr, di_stbovp_clr,
         di_rd_det_clr, dm_fault_clr, pwrdn_rstz, osc_low_clr, osc_low_rstz,
         r_pos_gate, osc_gate_n_2_, osc_gate_n_1_, osc_gate_n_0_, m_ovp,
         m_ovp_sta, setAE_7, m_scp, m_scp_sta, s_ovp, s_ovp_sta, s_scp,
         s_scp_sta, net10758, n1209, n1210, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n26, n71, n74,
         n75, n79, n80, n81, n83, n85, n95, n100, n101, n102, n103, n105, n106,
         n107, n109, n111, n112, n113, n114, n116, n117, n118, n119, n120,
         n121, n122, n124, n125, n126, n128, n129, n132, n133, n134, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n164, n165, n167, n168, n169, n170, n171, n172, n173, n174, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n1,
         n2, n3, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72,
         n73, n76, n77, n78, n82, n84, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n96, n97, n98, n99, n104, n108, n110, n115, n123, n127, n130,
         n131, n135, n136, n137, n138, n139, n163, n166, n175, n176, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151,
         SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153,
         SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155,
         SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157,
         SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159,
         SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161,
         SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163,
         SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165,
         SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167,
         SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169,
         SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171,
         SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173,
         SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175,
         SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177,
         SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179,
         SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181,
         SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183,
         SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185,
         SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187,
         SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189,
         SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191,
         SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193,
         SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195,
         SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197,
         SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199,
         SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201,
         SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203,
         SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205,
         SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207,
         SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209,
         SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211,
         SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213,
         SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215,
         SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217,
         SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219,
         SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221,
         SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223,
         SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225,
         SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227,
         SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229,
         SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231,
         SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233,
         SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235,
         SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237,
         SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239,
         SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241,
         SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243,
         SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245,
         SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247,
         SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249,
         SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251,
         SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253,
         SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255,
         SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257,
         SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259,
         SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261,
         SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263,
         SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265,
         SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267,
         SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269,
         SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271,
         SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273,
         SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275,
         SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277,
         SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279,
         SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281,
         SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283,
         SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285,
         SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287,
         SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289,
         SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291,
         SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293,
         SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295,
         SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297,
         SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299,
         SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301,
         SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303,
         SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305,
         SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307,
         SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309,
         SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311,
         SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313,
         SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315,
         SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317,
         SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319,
         SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321,
         SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323,
         SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325,
         SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327,
         SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329,
         SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331,
         SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333,
         SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335,
         SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337,
         SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339,
         SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341,
         SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343,
         SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345,
         SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347,
         SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349,
         SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351,
         SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353,
         SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355,
         SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357,
         SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359,
         SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361,
         SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363,
         SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365,
         SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367,
         SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369,
         SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371,
         SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373,
         SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375,
         SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377,
         SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379,
         SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381,
         SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383,
         SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385,
         SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387,
         SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389,
         SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391,
         SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393,
         SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395,
         SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397,
         SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399,
         SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401,
         SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403,
         SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405,
         SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407,
         SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409,
         SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411,
         SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413,
         SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415,
         SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417,
         SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419,
         SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421,
         SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423,
         SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425,
         SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427,
         SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429,
         SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431,
         SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433,
         SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435,
         SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437,
         SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439,
         SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441,
         SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443,
         SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445,
         SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447,
         SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449,
         SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451,
         SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453,
         SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455,
         SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457,
         SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459,
         SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461,
         SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463,
         SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465,
         SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467,
         SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469,
         SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471,
         SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473,
         SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475,
         SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477,
         SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479,
         SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481,
         SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483,
         SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485,
         SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487,
         SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489,
         SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491,
         SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493,
         SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495,
         SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497,
         SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499,
         SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501,
         SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503,
         SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505,
         SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507,
         SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509,
         SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511,
         SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513,
         SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515,
         SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517,
         SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519,
         SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521,
         SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523,
         SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525,
         SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527,
         SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529,
         SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531,
         SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533,
         SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535,
         SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537,
         SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539,
         SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541,
         SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543,
         SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545,
         SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547,
         SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549,
         SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551,
         SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553,
         SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555,
         SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557,
         SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559,
         SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561,
         SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563,
         SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565,
         SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567,
         SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569,
         SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571,
         SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573,
         SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575,
         SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577,
         SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579,
         SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581,
         SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583,
         SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585,
         SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587,
         SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589,
         SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591,
         SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593,
         SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595,
         SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597,
         SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599,
         SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601,
         SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603,
         SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605,
         SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607,
         SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609,
         SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611,
         SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613,
         SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615,
         SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617,
         SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619,
         SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621,
         SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623,
         SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625,
         SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627,
         SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629,
         SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631,
         SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633,
         SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635,
         SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637,
         SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639,
         SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641,
         SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643,
         SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645,
         SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647,
         SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649,
         SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651,
         SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653,
         SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655,
         SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657,
         SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659,
         SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661,
         SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663,
         SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665,
         SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667,
         SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669,
         SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671,
         SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673,
         SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675,
         SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677,
         SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679,
         SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681,
         SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683,
         SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685,
         SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687,
         SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689,
         SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691,
         SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693,
         SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695,
         SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697,
         SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699,
         SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701,
         SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703,
         SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705,
         SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707,
         SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709,
         SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711,
         SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713,
         SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715,
         SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717,
         SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719,
         SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721,
         SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723,
         SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725,
         SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727,
         SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729,
         SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731,
         SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733,
         SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735,
         SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737,
         SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739,
         SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741,
         SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743,
         SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745,
         SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747,
         SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749,
         SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751,
         SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753,
         SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755,
         SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757,
         SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759,
         SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761,
         SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763,
         SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765,
         SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767,
         SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769,
         SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771,
         SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773,
         SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775,
         SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777,
         SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779,
         SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781,
         SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783,
         SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785,
         SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787,
         SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789,
         SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791,
         SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793,
         SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795,
         SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797,
         SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799,
         SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801,
         SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803,
         SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805,
         SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807,
         SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809,
         SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811,
         SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813,
         SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815,
         SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817,
         SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819,
         SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821,
         SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823,
         SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825,
         SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827,
         SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829,
         SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831,
         SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833,
         SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835,
         SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837,
         SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839,
         SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841,
         SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843,
         SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845,
         SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847,
         SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849,
         SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851,
         SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853,
         SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855,
         SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857,
         SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859,
         SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861,
         SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863,
         SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865,
         SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867,
         SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869,
         SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871,
         SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873,
         SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875,
         SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877,
         SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879,
         SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881,
         SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883,
         SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885,
         SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887,
         SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889,
         SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891,
         SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893,
         SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895,
         SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897,
         SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899,
         SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901,
         SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903,
         SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905,
         SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907,
         SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909,
         SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911,
         SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913,
         SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915,
         SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917,
         SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919,
         SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921,
         SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923,
         SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925,
         SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927,
         SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929,
         SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931,
         SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933,
         SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935,
         SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937,
         SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939,
         SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941,
         SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943,
         SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945,
         SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947,
         SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949,
         SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951,
         SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953,
         SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955,
         SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957,
         SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959,
         SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961,
         SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963,
         SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965,
         SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967,
         SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969,
         SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971,
         SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973,
         SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975,
         SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977,
         SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979,
         SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981,
         SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983,
         SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985,
         SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987,
         SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989,
         SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991,
         SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993,
         SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995,
         SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997,
         SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999,
         SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001,
         SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003,
         SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005,
         SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007,
         SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009,
         SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011,
         SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013,
         SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015,
         SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017;
  wire   [167:162] we;
  wire   [3:2] regE3;
  wire   [7:0] regDF;
  wire   [7:0] regDE;
  wire   [7:0] reg31;
  wire   [7:0] reg30;
  wire   [7:0] reg28;
  wire   [7:0] reg27;
  wire   [7:1] reg21;
  wire   [4:0] reg20;
  wire   [7:3] reg12;
  wire   [7:0] reg06;
  wire   [7:0] reg05;
  wire   [7:0] regAF;
  wire   [7:0] regAE;
  wire   [5:0] regAD;
  wire   [7:0] regAC;
  wire   [7:0] regAB;
  wire   [7:0] reg94;
  wire   [7:0] irqAE;
  wire   [7:0] irqDF;
  wire   [7:0] irq28;
  wire   [7:0] irq04;
  wire   [7:0] irq03;
  wire   [1:0] drstz;
  wire   [4:0] rstcnt;
  wire   [1:0] r_phyrst;
  wire   [7:0] wd01;
  wire   [7:0] clr03;
  wire   [7:0] set03;
  wire   [7:0] clr04;
  wire   [7:0] set04;
  wire   [7:0] wd12;
  wire   [14:0] inst_ofs_plus;
  wire   [7:0] wd18;
  wire   [7:0] wd19;
  wire   [7:0] wd20;
  wire   [7:0] wd21;
  wire   [7:0] clr28;
  wire   [2:0] oscdwn_shft;
  wire   [7:0] d_p0;
  wire   [7:0] setDF;
  wire   [7:0] clrDF;
  wire   [7:0] clrAE;
  wire   [5:0] setAE;
  wire   [3:0] lt_regE4_3_0;
  wire   [4:2] add_179_carry;

  AND2X1 U0_MASK_0 ( .A(oscdwn_shft[2]), .B(as_p0_chg), .Y(p0_chg_clr) );
  AND2X1 U0_MASK_1 ( .A(test_so2), .B(di_stbovp), .Y(di_stbovp_clr) );
  AND2X1 U0_MASK_2 ( .A(regD4_6_), .B(di_rd_det), .Y(di_rd_det_clr) );
  AND2X1 U0_MASK_3 ( .A(r_srcctl[7]), .B(dmf_wkup), .Y(dm_fault_clr) );
  AND2X1 U0_MASK_4 ( .A(regD4_5_), .B(aswkup), .Y(osc_low_clr) );
  HAD1X1 add_179_U1_1_1 ( .A(N26), .B(N27), .CO(add_179_carry[2]), .SO(N29) );
  HAD1X1 add_179_U1_1_2 ( .A(N25), .B(add_179_carry[2]), .CO(add_179_carry[3]), 
        .SO(N30) );
  HAD1X1 add_179_U1_1_3 ( .A(N24), .B(add_179_carry[3]), .CO(add_179_carry[4]), 
        .SO(N31) );
  glreg_a0_79 u0_reg00 ( .clk(clk), .arstz(n58), .we(we_176), .wdat({n254, 
        n246, n238, n231, n225, n218, n208, n203}), .rdat({r_txendk, r_txauto}), .test_si(n311), .test_se(test_se) );
  glreg_a0_78 u0_reg01 ( .clk(clk), .arstz(n40), .we(upd01), .wdat(wd01), 
        .rdat({r_last, r_first, r_unlock, r_txnumk}), .test_si(r_txendk), 
        .test_se(test_se) );
  glsta_a0_6 u0_reg03 ( .clk(clk), .arstz(n49), .rst0(n18), .set2({set03[7:4], 
        n71, set03[2:0]}), .clr1(clr03), .rdat(dbgpo[7:0]), .irq(irq03), 
        .test_si(r_last), .test_se(test_se) );
  glsta_a0_5 u0_reg04 ( .clk(clk), .arstz(n41), .rst0(n19), .set2(set04), 
        .clr1(clr04), .rdat(dbgpo[15:8]), .irq(irq04), .test_si(dbgpo[7]), 
        .test_se(test_se) );
  glreg_a0_77 u0_reg05 ( .clk(clk), .arstz(n46), .we(we_181), .wdat({n255, 
        sfr_wdat[6], n237, n231, n226, n219, n208, n202}), .rdat(reg05), 
        .test_si(dbgpo[15]), .test_se(test_se) );
  glreg_a0_76 u0_reg06 ( .clk(clk), .arstz(n50), .we(we_182), .wdat({n255, 
        n243, n237, n231, n225, n218, n208, n203}), .rdat(reg06), .test_si(
        reg05[7]), .test_se(test_se) );
  glreg_a0_75 u0_reg11 ( .clk(clk), .arstz(n51), .we(we_187), .wdat({n255, 
        sfr_wdat[6], n237, n231, n226, n219, n209, n203}), .rdat({reg11_7_, 
        r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0]}), .test_si(r_dpdmctl[7]), .test_se(test_se) );
  glreg_a0_74 u0_reg12 ( .clk(clk), .arstz(n52), .we(upd12), .wdat(wd12), 
        .rdat({reg12, r_txshrt, reg12_1, r_pshords}), .test_si(reg11_7_), 
        .test_se(test_se) );
  glreg_WIDTH5_2 u0_reg14 ( .clk(clk), .arstz(n90), .we(r_set_cpmsgid), .wdat(
        {n255, n244, n238, n231, n226}), .rdat({r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1]}), .test_si(reg12[7]), 
        .test_se(test_se) );
  glreg_a0_73 u0_reg15 ( .clk(clk), .arstz(n54), .we(we_191), .wdat({n255, 
        n243, n238, n232, n226, n219, n210, n204}), .rdat(dbgpo[31:24]), 
        .test_si(r_auto_gdcrc[0]), .test_se(test_se) );
  glreg_a0_72 u0_reg18 ( .clk(clk), .arstz(n55), .we(upd18), .wdat(wd18), 
        .rdat(r_inst_ofs[7:0]), .test_si(dbgpo[31]), .test_se(test_se) );
  glreg_a0_71 u0_reg19 ( .clk(clk), .arstz(n56), .we(upd19), .wdat(wd19), 
        .rdat({reg19_7_, r_inst_ofs[14:8]}), .test_si(r_inst_ofs[7]), 
        .test_se(test_se) );
  glreg_a0_70 u0_reg20 ( .clk(clk), .arstz(n61), .we(upd20), .wdat(wd20), 
        .rdat({r_dat_spec, r_dat_datarole, reg20}), .test_si(n11), .test_se(
        test_se) );
  glreg_a0_69 u0_reg21 ( .clk(clk), .arstz(n67), .we(upd21), .wdat(wd21), 
        .rdat({reg21, r_dat_portrole}), .test_si(r_dat_spec[1]), .test_se(
        test_se) );
  glreg_6_00000018 u0_reg25 ( .clk(clk), .arstz(n84), .we(n199), .wdat({n238, 
        sfr_wdat[4], n225, n220, n209, n203}), .rdat({r_i2c_attr, r_pg0_sel, 
        reg25_0_}), .test_si(reg21[7]), .test_se(test_se) );
  glreg_WIDTH1_6 u0_reg26 ( .clk(clk), .arstz(n98), .we(n198), .wdat(n202), 
        .rdat(lt_reg26_0), .test_si(r_i2c_attr), .test_se(test_se) );
  glreg_1_1 u1_reg26 ( .clk(clk), .arstz(n98), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat(r_hwi2c_en), .test_si(n306), .test_se(test_se)
         );
  glreg_7_70 u2_reg26 ( .clk(clk), .arstz(n82), .we(n198), .wdat({n254, n246, 
        n237, n231, n226, n219, n209}), .rdat(r_i2c_deva), .test_si(n303), 
        .test_se(test_se) );
  glreg_a0_68 u0_reg27 ( .clk(clk), .arstz(n78), .we(we_203), .wdat({n255, 
        n243, n238, n231, n226, n219, n209, n203}), .rdat(reg27), .test_si(
        lt_reg26_0), .test_se(test_se) );
  glsta_a0_4 u0_reg28 ( .clk(clk), .arstz(n77), .rst0(1'b0), .set2(i2c_ev), 
        .clr1(clr28), .rdat(reg28), .irq(irq28), .test_si(reg27[7]), .test_se(
        test_se) );
  glreg_a0_67 u0_reg31 ( .clk(clk), .arstz(n76), .we(upd31), .wdat(i_pc[15:8]), 
        .rdat(reg31), .test_si(reg28[7]), .test_se(test_se) );
  glreg_8_00000001 u0_regD1 ( .clk(clk), .arstz(n39), .we(we_209), .wdat({n255, 
        n243, n238, n231, n226, n219, n209, n202}), .rdat({r_exist1st, 
        r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, r_gpio_oe[6], r_gpio_pu[6], 
        r_gpio_pd[6]}), .test_si(regAF[7]), .test_se(test_se) );
  glreg_8_00000011 u0_regD3 ( .clk(clk), .arstz(n37), .we(we_211), .wdat({n255, 
        n243, n238, n234, n226, n219, n209, n202}), .rdat({regD3_7_, 
        r_gpio_oe[5], r_gpio_pu[5], r_gpio_pd[5], regD3_3, r_gpio_oe[4], 
        r_gpio_pu[4], r_gpio_pd[4]}), .test_si(r_exist1st), .test_se(test_se)
         );
  glreg_WIDTH3 u4_regD4 ( .clk(clk), .arstz(n98), .we(n360), .wdat({n255, n243, 
        n238}), .rdat({test_so2, regD4_6_, regD4_5_}), .test_si(regD4_4_), 
        .test_se(test_se) );
  glreg_WIDTH2_2 u3_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n360), .wdat({
        n234, n225}), .rdat({regD4_4_, regD4_3_}), .test_si(regD4_2_), 
        .test_se(test_se) );
  glreg_WIDTH1_5 u2_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n360), .wdat(
        n218), .rdat(regD4_2_), .test_si(r_i2c_deva[7]), .test_se(test_se) );
  glreg_WIDTH1_4 u1_regD4 ( .clk(clk), .arstz(osc_low_rstz), .we(n9), .wdat(
        n208), .rdat(regD4_1_), .test_si(r_hwi2c_en), .test_se(test_se) );
  glreg_WIDTH1_3 u0_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n360), .wdat(
        n202), .rdat(regD4_0_), .test_si(regD3_7_), .test_se(test_se) );
  glreg_8_000000f0 u0_regD5 ( .clk(clk), .arstz(n33), .we(we_213), .wdat({n254, 
        n246, n237, n234, n226, n219, n209, n203}), .rdat({r_gpio_pu[3:0], 
        r_gpio_pd[3:0]}), .test_si(regD4_0_), .test_se(test_se) );
  glreg_8_00000098 u0_regD6 ( .clk(clk), .arstz(n34), .we(we_214), .wdat({n254, 
        n243, n238, n234, n225, n219, n209, n203}), .rdat({r_gpio_oe[1], 
        r_gpio_s1, r_gpio_oe[0], r_gpio_s0}), .test_si(r_gpio_pu[3]), 
        .test_se(test_se) );
  glreg_8_00000032 u0_regD7 ( .clk(clk), .arstz(n35), .we(we_215), .wdat({n255, 
        n243, n237, n234, n227, n219, n208, n203}), .rdat({r_gpio_oe[3], 
        r_gpio_s3, r_gpio_oe[2], r_gpio_s2}), .test_si(r_gpio_oe[1]), 
        .test_se(test_se) );
  glreg_a0_66 u0_regD9 ( .clk(clk), .arstz(n72), .we(we_217), .wdat({n256, 
        n243, n238, n231, n227, n220, n209, n203}), .rdat({r_ana_tm, 
        r_fortxdat, r_fortxrdy, r_fortxen, r_sleep}), .test_si(r_gpio_oe[3]), 
        .test_se(test_se) );
  glreg_a0_65 u0_regDE ( .clk(clk), .arstz(n70), .we(we_222), .wdat({n256, 
        n243, n239, n232, n227, n220, n209, n203}), .rdat(regDE), .test_si(
        r_ana_tm[3]), .test_se(test_se) );
  glsta_a0_3 u0_regDF ( .clk(clk), .arstz(n73), .rst0(1'b0), .set2(setDF), 
        .clr1(clrDF), .rdat(regDF), .irq(irqDF), .test_si(regDE[7]), .test_se(
        test_se) );
  glreg_a0_64 u0_reg8F ( .clk(clk), .arstz(n68), .we(we_143), .wdat({n256, 
        n244, n239, n232, n227, n220, n210, n204}), .rdat(r_dpdmctl), 
        .test_si(reg06[7]), .test_se(test_se) );
  glreg_WIDTH4 u0_reg94 ( .clk(clk), .arstz(n93), .we(we_148), .wdat({n244, 
        n239, n232, n227}), .rdat(reg94[6:3]), .test_si(reg31[7]), .test_se(
        test_se) );
  glreg_a0_63 u0_regA1 ( .clk(clk), .arstz(n66), .we(we[162]), .wdat({n256, 
        n244, n239, n232, n227, n220, n210, n204}), .rdat(r_regtrm[7:0]), 
        .test_si(reg94[6]), .test_se(test_se) );
  glreg_a0_62 u0_regA2 ( .clk(clk), .arstz(n69), .we(we[162]), .wdat({n256, 
        n244, n239, n232, n227, n220, n210, n204}), .rdat(r_regtrm[15:8]), 
        .test_si(r_regtrm[7]), .test_se(test_se) );
  glreg_a0_61 u0_regA3 ( .clk(clk), .arstz(n64), .we(we[163]), .wdat({n256, 
        n244, n239, n232, n227, n220, n210, n204}), .rdat(r_regtrm[23:16]), 
        .test_si(r_regtrm[15]), .test_se(test_se) );
  glreg_a0_60 u0_regA4 ( .clk(clk), .arstz(n63), .we(we[164]), .wdat({n256, 
        n244, n239, n232, n227, n220, n210, n204}), .rdat(r_regtrm[31:24]), 
        .test_si(r_regtrm[23]), .test_se(test_se) );
  glreg_a0_59 u0_regA5 ( .clk(clk), .arstz(n62), .we(we[165]), .wdat({n256, 
        n244, n239, n232, n227, n220, n210, n204}), .rdat(r_regtrm[39:32]), 
        .test_si(r_regtrm[31]), .test_se(test_se) );
  glreg_a0_58 u0_regA6 ( .clk(clk), .arstz(n65), .we(we[166]), .wdat({n256, 
        n244, n239, n232, n228, n220, n210, n204}), .rdat(r_regtrm[47:40]), 
        .test_si(r_regtrm[39]), .test_se(test_se) );
  glreg_a0_57 u0_regA7 ( .clk(clk), .arstz(n60), .we(we[167]), .wdat({n257, 
        n244, n240, n233, n228, n221, n210, n204}), .rdat(r_regtrm[55:48]), 
        .test_si(r_regtrm[47]), .test_se(test_se) );
  glreg_a0_56 u0_regAB ( .clk(clk), .arstz(n59), .we(we_171), .wdat({n257, 
        n245, n240, n233, n228, n221, n210, n204}), .rdat(regAB), .test_si(
        r_regtrm[55]), .test_se(test_se) );
  glreg_8_00000028 u0_regAC ( .clk(clk), .arstz(n36), .we(we_172), .wdat({n257, 
        n245, n237, n233, n225, n221, n211, n205}), .rdat(regAC), .test_si(
        regAB[7]), .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_2 u2_ovp_db ( .o_dbc(reg94[2]), .o_chg(), .i_org(
        srci[2]), .clk(clk_500), .rstz(n89), .test_si(n304), .test_so(n303), 
        .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_1 u1_ocp_db ( .o_dbc(reg94[1]), .o_chg(), .i_org(
        srci[1]), .clk(clk_500), .rstz(n88), .test_si(n308), .test_so(n307), 
        .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_0 u1_uvp_db ( .o_dbc(reg94[0]), .o_chg(), .i_org(
        srci[0]), .clk(clk_500), .rstz(n87), .test_si(n305), .test_so(n304), 
        .test_se(test_se) );
  dbnc_a0_2 u1_ovp_db ( .o_dbc(m_ovp), .o_chg(m_ovp_sta), .i_org(srci[2]), 
        .clk(clk_500k), .rstz(n86), .test_si(n307), .test_so(n306), .test_se(
        test_se) );
  dbnc_WIDTH3_TIMEOUT5_4 u0_otpi_db ( .o_dbc(regAD[3]), .o_chg(setAE[3]), 
        .i_org(srci[5]), .clk(clk_1500k), .rstz(n91), .test_si(n314), 
        .test_so(n313), .test_se(test_se) );
  dbnc_WIDTH3_TIMEOUT5_3 u0_ocp_db ( .o_dbc(regAD[1]), .o_chg(setAE[1]), 
        .i_org(srci[1]), .clk(clk_1500k), .rstz(n92), .test_si(n315), 
        .test_so(n314), .test_se(test_se) );
  dbnc_WIDTH3_TIMEOUT5_2 u0_uvp_db ( .o_dbc(regAD[0]), .o_chg(setAE[0]), 
        .i_org(srci[0]), .clk(clk_1500k), .rstz(n90), .test_si(n310), 
        .test_so(n309), .test_se(test_se) );
  dbnc_WIDTH3_TIMEOUT5_1 u1_scp_db ( .o_dbc(m_scp), .o_chg(m_scp_sta), .i_org(
        srci[3]), .clk(clk_1500k), .rstz(n92), .test_si(r_fw_pwrv[3]), 
        .test_so(n305), .test_se(test_se) );
  dbnc_WIDTH3_TIMEOUT5_0 u0_dmf_db ( .o_dbc(regAD_7), .o_chg(setAE_7), .i_org(
        dm_fault), .clk(clk_1500k), .rstz(n91), .test_si(n316), .test_so(n315), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_13 u0_otps_db ( .o_dbc(reg94[7]), .o_chg(), .i_org(
        srci[5]), .clk(clk), .rstz(n94), .test_si(n313), .test_so(n312), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_12 u0_cc1_db ( .o_dbc(regF4_3), .o_chg(), .i_org(cc1_di), .clk(clk), .rstz(n96), .test_si(rstcnt[4]), .test_so(n317), .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_11 u0_cc2_db ( .o_dbc(regF4_7_), .o_chg(), .i_org(
        cc2_di), .clk(clk), .rstz(n94), .test_si(n317), .test_so(n316), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_10 u0_ovp_db ( .o_dbc(s_ovp), .o_chg(s_ovp_sta), 
        .i_org(srci[2]), .clk(clk), .rstz(n96), .test_si(n312), .test_so(n311), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_9 u0_scp_db ( .o_dbc(s_scp), .o_chg(s_scp_sta), .i_org(
        srci[3]), .clk(clk), .rstz(n97), .test_si(r_cctrx[7]), .test_so(n310), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_8 u0_v5oc_db ( .o_dbc(regAD[5]), .o_chg(setAE[5]), 
        .i_org(srci[4]), .clk(clk), .rstz(n97), .test_si(n309), .test_so(n308), 
        .test_se(test_se) );
  glsta_a0_2 u0_regAE ( .clk(clk), .arstz(n57), .rst0(1'b0), .set2({setAE_7, 
        1'b0, setAE}), .clr1(clrAE), .rdat(regAE), .irq(irqAE), .test_si(
        regAC[7]), .test_se(test_se) );
  glreg_a0_55 u0_regAF ( .clk(clk), .arstz(n48), .we(we_175), .wdat({n257, 
        n245, n240, n233, n228, n221, n211, n205}), .rdat(regAF), .test_si(
        regAE[7]), .test_se(test_se) );
  glreg_a0_54 u0_regE3 ( .clk(clk), .arstz(n47), .we(we_227), .wdat({n257, 
        n245, n240, n233, n228, n221, n211, n205}), .rdat({r_srcctl[7:4], 
        regE3, r_srcctl[1], regE3_0}), .test_si(regDF[7]), .test_se(test_se)
         );
  glreg_4_00000004 u1_regE4 ( .clk(clk), .arstz(n93), .we(r_pwrv_upd), .wdat(
        lt_regE4_3_0), .rdat(r_fw_pwrv[3:0]), .test_si(regD4_1_), .test_se(
        test_se) );
  glreg_8_00000004 u0_regE4 ( .clk(clk), .arstz(n38), .we(we_228), .wdat({n257, 
        n245, n240, n233, n228, n218, n211, n205}), .rdat({r_pwrctl, 
        lt_regE4_3_0}), .test_si(r_srcctl[7]), .test_se(test_se) );
  glreg_8_0000001f u0_regE5 ( .clk(clk), .arstz(n32), .we(r_pwrv_upd), .wdat({
        n257, n245, n240, n234, n225, n218, n208, n202}), .rdat(
        r_fw_pwrv[11:4]), .test_si(r_pwrctl[7]), .test_se(test_se) );
  glreg_a0_53 u0_regE6 ( .clk(clk), .arstz(n45), .we(we_230), .wdat({n257, 
        n245, n240, n233, n228, n221, n211, n205}), .rdat(r_ccrx), .test_si(
        r_fw_pwrv[11]), .test_se(test_se) );
  glreg_a0_52 u0_regE7 ( .clk(clk), .arstz(n44), .we(we_231), .wdat({n257, 
        n245, n240, n233, n228, n221, n211, n205}), .rdat(r_ccctl), .test_si(
        r_ccrx[7]), .test_se(test_se) );
  glreg_a0_51 u0_regE8 ( .clk(clk), .arstz(n53), .we(we_232), .wdat({n257, 
        n245, n240, n233, n228, n221, n211, n205}), .rdat(r_comp_opt), 
        .test_si(r_ccctl[7]), .test_se(test_se) );
  glreg_a0_50 u0_regF5 ( .clk(clk), .arstz(n43), .we(we_245), .wdat({n254, 
        n245, n237, n233, n225, n221, n211, n205}), .rdat(r_cvctl), .test_si(
        r_comp_opt[7]), .test_se(test_se) );
  glreg_a0_49 u0_regF6 ( .clk(clk), .arstz(n42), .we(we_246), .wdat({n256, 
        n246, n239, n231, n226, n218, n208, n202}), .rdat(r_cctrx), .test_si(
        r_cvctl[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_regbank_a0 clk_gate_rstcnt_reg ( .CLK(clk), .EN(N23), 
        .ENCLK(net10758), .TE(test_se) );
  regbank_a0_DW01_add_0 add_527 ( .A(regAC), .B(regAB), .CI(1'b0), .SUM(
        r_pwr_i), .CO() );
  regbank_a0_DW01_inc_0 add_303 ( .A({1'b0, r_inst_ofs}), .SUM({
        SYNOPSYS_UNCONNECTED_1, inst_ofs_plus}) );
  regbank_a0_DW_rightsh_1 srl_132 ( .A({dac_r_vs, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, r_cctrx, r_cvctl, regF4_7_, x_daclsb[5:3], regF4_3, 
        x_daclsb[2:0], r_sar_en, r_dac_en, dac_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_comp_opt, r_ccctl, r_ccrx, r_fw_pwrv[11:4], r_pwrctl, r_fw_pwrv[3:0], 
        r_srcctl[7:4], regE3, r_srcctl[1], regE3_0, dac_r_cmpsta, dac_r_comp, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, regDF, regDE, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_ana_tm, r_fortxdat, 
        r_fortxrdy, r_fortxen, r_sleep, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, r_gpio_oe[3], r_gpio_s3, r_gpio_oe[2], r_gpio_s2, 
        r_gpio_oe[1], r_gpio_s1, r_gpio_oe[0], r_gpio_s0, r_gpio_pu[3:0], 
        r_gpio_pd[3:0], test_so2, regD4_6_, regD4_5_, regD4_4_, regD4_3_, 
        regD4_2_, regD4_1_, regD4_0_, regD3_7_, r_gpio_oe[5], r_gpio_pu[5], 
        r_gpio_pd[5], regD3_3, r_gpio_oe[4], r_gpio_pu[4], r_gpio_pd[4], 
        i_i2c_rwbuf, r_exist1st, r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, 
        r_gpio_oe[6], r_gpio_pu[6], r_gpio_pd[6], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, reg31, reg30, i_i2c_ltbuf, reg28, reg27, r_i2c_deva, 
        r_hwi2c_en, 1'b0, 1'b0, r_i2c_attr, r_pg0_sel, reg25_0_, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, prx_rcvinf[4], REVID, 
        prx_rcvinf[3], ptx_fsm, prx_fsm, reg21, r_dat_portrole, r_dat_spec, 
        r_dat_datarole, reg20, n12, r_inst_ofs, i_i2c_ofs, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, dbgpo[31:24], r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1], prl_cpmsgid, n14, 
        prx_rcvinf[2:0], prl_fsm, reg12, r_txshrt, reg12_1, r_pshords, 
        reg11_7_, r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0], 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, pff_empty, 
        pff_full, pff_ptr, reg06, reg05, dbgpo[15:0], pff_rdat, r_last, 
        r_first, r_unlock, r_txnumk, r_txendk, r_txauto, regAF, regAE, regAD_7, 
        1'b0, regAD, regAC, regAB, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_regtrm, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, fcp_r_crc, fcp_r_dat, fcp_r_msk, fcp_r_sta, 
        fcp_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, fcp_r_acc, r_accctl, fcp_r_tui, reg94, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, r_isofs, r_adofs, r_dpdmctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_cvofs, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .DATA_TC(1'b0), .SH({sfr_addr[6:1], n176, 
        1'b0, 1'b0, 1'b0}), .B({SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, 
        SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, 
        SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, 
        SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, 
        SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, 
        SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, 
        SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, 
        SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, 
        SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, 
        SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, 
        SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, 
        SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, 
        SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, 
        SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, 
        SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, 
        SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, 
        SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, 
        SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, 
        SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, 
        SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, 
        SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, 
        SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, 
        SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, 
        SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, 
        SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, 
        SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, 
        SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, 
        SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, 
        SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, 
        SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, 
        SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, 
        SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, 
        SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, 
        SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, 
        SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, 
        SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, 
        SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, 
        SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, 
        SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, 
        SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, 
        SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, 
        SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, 
        SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, 
        SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, 
        SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, 
        SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, 
        SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, 
        SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, 
        SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, 
        SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, 
        SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, 
        SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, 
        SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, 
        SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, 
        SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, 
        SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, 
        SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, 
        SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, 
        SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, 
        SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, 
        SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, 
        SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, 
        SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, 
        SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, 
        SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, 
        SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, 
        SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, 
        SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, 
        SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, 
        SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, 
        SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, 
        SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, 
        SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, 
        SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, 
        SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, 
        SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, 
        SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, 
        SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, 
        SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, 
        SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, 
        SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, 
        SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, 
        SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, 
        SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, 
        SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, 
        SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, 
        SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, 
        SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, 
        SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, 
        SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, 
        SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, 
        SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, 
        SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, 
        SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, 
        SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, 
        SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, 
        SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, 
        SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, 
        SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, 
        SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, 
        SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, 
        SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, 
        SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, 
        SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, 
        SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, 
        SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, 
        SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, 
        SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, 
        SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, 
        SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, 
        SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, 
        SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, 
        SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, 
        SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, 
        SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, 
        SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, 
        SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, 
        SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, 
        SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, 
        SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, 
        SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, 
        SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, 
        SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, 
        SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, 
        SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, 
        SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, 
        SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, 
        SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, 
        SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, 
        SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, 
        SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, 
        SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, 
        SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, 
        SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, 
        SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, 
        SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, 
        SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, 
        SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, 
        SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, 
        SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, 
        SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, 
        SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, 
        SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, 
        SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, 
        SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, 
        SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, 
        SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, 
        SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, 
        SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, 
        SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, 
        SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, 
        SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, 
        SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, 
        SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, 
        SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, 
        SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, 
        SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, 
        SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, 
        SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, 
        SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, 
        SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, 
        SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, 
        SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, 
        SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, 
        SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, 
        SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, 
        SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, 
        SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, 
        SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, 
        SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, 
        SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, 
        SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, 
        SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, 
        SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, 
        SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, 
        SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, 
        SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, 
        SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, 
        SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, 
        SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, 
        SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, 
        SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, 
        SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, 
        SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, 
        SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, 
        SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, 
        SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, 
        SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, 
        SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, 
        SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, 
        SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, 
        SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, 
        SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, 
        SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, 
        SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, 
        SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, 
        SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, 
        SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, 
        SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, 
        SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, 
        SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, 
        SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, 
        SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, 
        SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, 
        SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, 
        SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, 
        SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, 
        SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, 
        SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, 
        SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, 
        SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, 
        SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, 
        SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, 
        SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, 
        SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, 
        SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, 
        SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, 
        SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, 
        SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, 
        SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, 
        SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, 
        SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, 
        SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, 
        SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, 
        SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, 
        SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, 
        SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, 
        SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, 
        SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, 
        SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, 
        SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, 
        SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, 
        SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, 
        SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, 
        SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, 
        SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, 
        SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, 
        SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, 
        SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, 
        SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, 
        SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, 
        SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, 
        SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, 
        SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, 
        SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, 
        SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, 
        SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, 
        SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, 
        SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, 
        SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, 
        SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, 
        SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, 
        SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, 
        SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, 
        SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, 
        SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, 
        SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, 
        SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, 
        SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, 
        SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, 
        SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, 
        SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, 
        SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, 
        SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, 
        SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, 
        SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, 
        SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, 
        SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, 
        SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, 
        SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, 
        SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, 
        SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, 
        SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, 
        SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, 
        SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, 
        SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, 
        SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, 
        SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, 
        SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, 
        SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017, sfr_rdat}) );
  SDFFRQX1 r_phyrst_reg_0_ ( .D(n1210), .SIN(oscdwn_shft[2]), .SMC(test_se), 
        .C(clk), .XR(n2), .Q(r_phyrst[0]) );
  SDFFRQX1 rstcnt_reg_0_ ( .D(N36), .SIN(r_phyrst[1]), .SMC(test_se), .C(
        net10758), .XR(n3), .Q(rstcnt[0]) );
  SDFFRQX1 d_p0_reg_7_ ( .D(ff_p0[7]), .SIN(d_p0[6]), .SMC(test_se), .C(clk), 
        .XR(n381), .Q(d_p0[7]) );
  SDFFRQX1 d_p0_reg_6_ ( .D(ff_p0[6]), .SIN(d_p0[5]), .SMC(test_se), .C(clk), 
        .XR(n381), .Q(d_p0[6]) );
  SDFFRQX1 d_p0_reg_5_ ( .D(ff_p0[5]), .SIN(d_p0[4]), .SMC(test_se), .C(clk), 
        .XR(n381), .Q(d_p0[5]) );
  SDFFRQX1 d_p0_reg_4_ ( .D(ff_p0[4]), .SIN(d_p0[3]), .SMC(test_se), .C(clk), 
        .XR(n381), .Q(d_p0[4]) );
  SDFFRQX1 d_p0_reg_3_ ( .D(ff_p0[3]), .SIN(d_p0[2]), .SMC(test_se), .C(clk), 
        .XR(n381), .Q(d_p0[3]) );
  SDFFRQX1 d_p0_reg_2_ ( .D(ff_p0[2]), .SIN(d_p0[1]), .SMC(test_se), .C(clk), 
        .XR(n381), .Q(d_p0[2]) );
  SDFFRQX1 d_p0_reg_1_ ( .D(ff_p0[1]), .SIN(d_p0[0]), .SMC(test_se), .C(clk), 
        .XR(n381), .Q(d_p0[1]) );
  SDFFRQX1 d_p0_reg_0_ ( .D(ff_p0[0]), .SIN(test_si2), .SMC(test_se), .C(clk), 
        .XR(n381), .Q(d_p0[0]) );
  SDFFRQX1 r_phyrst_reg_1_ ( .D(n1209), .SIN(r_phyrst[0]), .SMC(test_se), .C(
        clk), .XR(n2), .Q(r_phyrst[1]) );
  SDFFQX1 oscdwn_shft_reg_2_ ( .D(n355), .SIN(oscdwn_shft[1]), .SMC(test_se), 
        .C(clk), .Q(oscdwn_shft[2]) );
  SDFFQX1 oscdwn_shft_reg_1_ ( .D(oscdwn_shft[0]), .SIN(oscdwn_shft[0]), .SMC(
        test_se), .C(clk), .Q(oscdwn_shft[1]) );
  SDFFRQX1 drstz_reg_1_ ( .D(drstz[0]), .SIN(drstz[0]), .SMC(test_se), .C(clk), 
        .XR(n3), .Q(drstz[1]) );
  SDFFNRQX1 osc_gate_n_reg_1_ ( .D(osc_gate_n_0_), .SIN(osc_gate_n_0_), .SMC(
        test_se), .XC(xclk), .XR(n2), .Q(osc_gate_n_1_) );
  SDFFRQX1 rstcnt_reg_3_ ( .D(N33), .SIN(rstcnt[2]), .SMC(test_se), .C(
        net10758), .XR(n2), .Q(rstcnt[3]) );
  SDFFRQX1 rstcnt_reg_1_ ( .D(N35), .SIN(rstcnt[0]), .SMC(test_se), .C(
        net10758), .XR(n3), .Q(rstcnt[1]) );
  SDFFRQX1 rstcnt_reg_2_ ( .D(N34), .SIN(rstcnt[1]), .SMC(test_se), .C(
        net10758), .XR(n2), .Q(rstcnt[2]) );
  SDFFRQX1 rstcnt_reg_4_ ( .D(N32), .SIN(rstcnt[3]), .SMC(test_se), .C(
        net10758), .XR(n3), .Q(rstcnt[4]) );
  SDFFNRQX1 osc_gate_n_reg_3_ ( .D(osc_gate_n_2_), .SIN(osc_gate_n_2_), .SMC(
        test_se), .XC(xclk), .XR(n3), .Q(test_so1) );
  SDFFNRQX1 osc_gate_n_reg_0_ ( .D(r_pos_gate), .SIN(test_si1), .SMC(test_se), 
        .XC(xclk), .XR(n3), .Q(osc_gate_n_0_) );
  SDFFNRQX1 osc_gate_n_reg_2_ ( .D(osc_gate_n_1_), .SIN(osc_gate_n_1_), .SMC(
        test_se), .XC(xclk), .XR(n2), .Q(osc_gate_n_2_) );
  OAI21X1 U406 ( .B(n197), .C(n384), .A(n264), .Y(srstz) );
  SDFFQX1 oscdwn_shft_reg_0_ ( .D(N81), .SIN(drstz[1]), .SMC(test_se), .C(clk), 
        .Q(oscdwn_shft[0]) );
  SDFFRQX1 drstz_reg_0_ ( .D(1'b1), .SIN(d_p0[7]), .SMC(test_se), .C(clk), 
        .XR(n2), .Q(drstz[0]) );
  INVX2 U7 ( .A(n321), .Y(n351) );
  INVX1 U8 ( .A(n201), .Y(n176) );
  INVX1 U9 ( .A(sfr_w), .Y(n301) );
  NAND21X1 U11 ( .B(n200), .A(n269), .Y(n321) );
  INVX1 U12 ( .A(n268), .Y(n269) );
  MUX2X1 U13 ( .D0(pff_rxpart[6]), .D1(n246), .S(n298), .Y(wd20[6]) );
  MUX2X1 U14 ( .D0(pff_rxpart[5]), .D1(n240), .S(n298), .Y(wd20[5]) );
  INVXL U15 ( .A(xrstz), .Y(n1) );
  INVXL U16 ( .A(n1), .Y(n2) );
  INVXL U17 ( .A(n1), .Y(n3) );
  INVXL U18 ( .A(n284), .Y(n9) );
  INVX1 U19 ( .A(reg19_7_), .Y(n10) );
  INVX1 U20 ( .A(n10), .Y(n11) );
  INVX1 U21 ( .A(n10), .Y(n12) );
  INVX1 U22 ( .A(prl_cany0), .Y(n13) );
  INVX1 U23 ( .A(n13), .Y(n14) );
  INVX1 U24 ( .A(n358), .Y(n15) );
  INVX1 U25 ( .A(n362), .Y(n16) );
  BUFX3 U26 ( .A(n103), .Y(n17) );
  NOR2X1 U27 ( .A(n141), .B(prl_c0set), .Y(phyrst) );
  INVX1 U28 ( .A(phyrst), .Y(n18) );
  INVX1 U29 ( .A(phyrst), .Y(n19) );
  NOR21XL U30 ( .B(pff_ack[0]), .A(prl_cany0), .Y(set04[4]) );
  BUFX3 U31 ( .A(pff_ptr[4]), .Y(dbgpo[20]) );
  BUFX3 U32 ( .A(pff_ptr[0]), .Y(dbgpo[16]) );
  BUFX3 U33 ( .A(pff_ptr[5]), .Y(dbgpo[21]) );
  BUFX3 U34 ( .A(pff_ptr[2]), .Y(dbgpo[18]) );
  BUFX3 U35 ( .A(pff_ptr[3]), .Y(dbgpo[19]) );
  BUFX3 U36 ( .A(pff_ptr[1]), .Y(dbgpo[17]) );
  INVXL U37 ( .A(n201), .Y(n200) );
  NAND21XL U38 ( .B(n95), .A(n351), .Y(n359) );
  AND2XL U39 ( .A(n344), .B(n351), .Y(r_dacwr[11]) );
  NOR21XL U40 ( .B(n351), .A(n132), .Y(r_fcpwr[1]) );
  AND2XL U41 ( .A(n272), .B(n351), .Y(we_172) );
  AND2XL U42 ( .A(n350), .B(n351), .Y(we_148) );
  NAND32XL U43 ( .B(n325), .C(n278), .A(n201), .Y(n79) );
  NAND21XL U44 ( .B(n335), .A(n176), .Y(n270) );
  AND4XL U45 ( .A(n327), .B(n335), .C(n326), .D(n201), .Y(we_176) );
  NAND21XL U46 ( .B(n265), .A(sfr_addr[2]), .Y(n335) );
  NAND21XL U47 ( .B(n265), .A(sfr_addr[1]), .Y(n326) );
  NAND21XL U48 ( .B(n265), .A(sfr_addr[3]), .Y(n289) );
  MUX2XL U49 ( .D0(i_pc[1]), .D1(prx_adpn[1]), .S(n12), .Y(reg30[1]) );
  AND3X1 U50 ( .A(n9), .B(n224), .C(n355), .Y(ps_pwrdn) );
  ENOXL U51 ( .A(n216), .B(n111), .C(r_txnumk[1]), .D(n111), .Y(wd01[1]) );
  ENOXL U52 ( .A(n223), .B(n16), .C(r_txnumk[2]), .D(n111), .Y(wd01[2]) );
  MUX2XL U53 ( .D0(r_txnumk[3]), .D1(n229), .S(n362), .Y(wd01[3]) );
  INVX1 U54 ( .A(n258), .Y(n254) );
  INVX1 U55 ( .A(n213), .Y(n208) );
  INVX1 U56 ( .A(n251), .Y(n245) );
  INVX1 U57 ( .A(n261), .Y(n257) );
  INVX1 U58 ( .A(n260), .Y(n256) );
  INVX1 U59 ( .A(n215), .Y(n210) );
  INVX1 U60 ( .A(n250), .Y(n244) );
  INVX1 U61 ( .A(n214), .Y(n209) );
  INVX1 U62 ( .A(n249), .Y(n243) );
  INVX1 U63 ( .A(n259), .Y(n255) );
  INVX1 U64 ( .A(n212), .Y(n211) );
  INVX1 U65 ( .A(n230), .Y(n224) );
  INVX1 U66 ( .A(n230), .Y(n225) );
  BUFX3 U67 ( .A(n217), .Y(n213) );
  BUFX3 U68 ( .A(n253), .Y(n248) );
  BUFX3 U69 ( .A(n263), .Y(n258) );
  NAND2X1 U70 ( .A(n206), .B(n222), .Y(n129) );
  NOR3XL U71 ( .A(n133), .B(n236), .C(n222), .Y(r_discard) );
  AND2X1 U72 ( .A(n323), .B(n237), .Y(clr04[5]) );
  AND2X1 U73 ( .A(n323), .B(n208), .Y(clr04[1]) );
  AND2X1 U74 ( .A(n323), .B(n234), .Y(clr04[4]) );
  AND2X1 U75 ( .A(n323), .B(n202), .Y(clr04[0]) );
  AND2X1 U76 ( .A(n323), .B(n246), .Y(clr04[6]) );
  AND2X1 U77 ( .A(n323), .B(n218), .Y(clr04[2]) );
  AND2X1 U78 ( .A(n323), .B(n254), .Y(clr04[7]) );
  AND2X1 U79 ( .A(n323), .B(n224), .Y(clr04[3]) );
  INVX1 U80 ( .A(n223), .Y(n218) );
  INVX1 U81 ( .A(n207), .Y(n202) );
  INVX1 U82 ( .A(n242), .Y(n237) );
  BUFX3 U83 ( .A(n217), .Y(n212) );
  BUFX3 U84 ( .A(n247), .Y(n250) );
  BUFX3 U85 ( .A(n263), .Y(n259) );
  BUFX3 U86 ( .A(n251), .Y(n249) );
  BUFX3 U87 ( .A(n253), .Y(n251) );
  BUFX3 U88 ( .A(n259), .Y(n260) );
  BUFX3 U89 ( .A(n212), .Y(n214) );
  INVX1 U90 ( .A(n235), .Y(n234) );
  INVX1 U91 ( .A(n236), .Y(n233) );
  INVX1 U92 ( .A(n242), .Y(n239) );
  INVX1 U93 ( .A(n230), .Y(n227) );
  INVX1 U94 ( .A(n223), .Y(n220) );
  INVX1 U95 ( .A(n236), .Y(n232) );
  INVX1 U96 ( .A(n207), .Y(n204) );
  INVX1 U97 ( .A(n223), .Y(n219) );
  INVX1 U98 ( .A(n230), .Y(n226) );
  INVX1 U99 ( .A(n242), .Y(n238) );
  INVX1 U100 ( .A(n207), .Y(n203) );
  INVX1 U101 ( .A(n236), .Y(n231) );
  INVX1 U102 ( .A(n223), .Y(n221) );
  INVX1 U103 ( .A(n242), .Y(n240) );
  INVX1 U104 ( .A(n230), .Y(n228) );
  INVX1 U105 ( .A(n207), .Y(n205) );
  BUFX3 U106 ( .A(n259), .Y(n261) );
  BUFX3 U107 ( .A(n212), .Y(n215) );
  BUFX3 U108 ( .A(n247), .Y(n252) );
  BUFX3 U109 ( .A(n259), .Y(n262) );
  BUFX3 U110 ( .A(n212), .Y(n216) );
  INVX1 U111 ( .A(n230), .Y(n229) );
  INVX1 U112 ( .A(n247), .Y(n246) );
  INVX1 U113 ( .A(n104), .Y(n92) );
  INVX1 U114 ( .A(n123), .Y(n91) );
  INVX1 U115 ( .A(n136), .Y(n90) );
  INVX1 U116 ( .A(n104), .Y(n93) );
  INVX1 U117 ( .A(n138), .Y(n39) );
  INVX1 U118 ( .A(n99), .Y(n97) );
  INVX1 U119 ( .A(n138), .Y(n57) );
  INVX1 U120 ( .A(n115), .Y(n73) );
  INVX1 U121 ( .A(n115), .Y(n77) );
  INVX1 U122 ( .A(n139), .Y(n41) );
  INVX1 U123 ( .A(n138), .Y(n49) );
  INVX1 U124 ( .A(n131), .Y(n42) );
  INVX1 U125 ( .A(n131), .Y(n43) );
  INVX1 U126 ( .A(n142), .Y(n53) );
  INVX1 U127 ( .A(n131), .Y(n44) );
  INVX1 U128 ( .A(n108), .Y(n45) );
  INVX1 U129 ( .A(n110), .Y(n47) );
  INVX1 U130 ( .A(n135), .Y(n48) );
  INVX1 U131 ( .A(n99), .Y(n96) );
  INVX1 U132 ( .A(n104), .Y(n94) );
  INVX1 U133 ( .A(n136), .Y(n59) );
  INVX1 U134 ( .A(n139), .Y(n60) );
  INVX1 U135 ( .A(n127), .Y(n65) );
  INVX1 U136 ( .A(n130), .Y(n62) );
  INVX1 U137 ( .A(n127), .Y(n63) );
  INVX1 U138 ( .A(n127), .Y(n64) );
  INVX1 U139 ( .A(n123), .Y(n69) );
  INVX1 U140 ( .A(n130), .Y(n66) );
  INVX1 U141 ( .A(n138), .Y(n68) );
  INVX1 U142 ( .A(n123), .Y(n70) );
  INVX1 U143 ( .A(n123), .Y(n72) );
  INVX1 U144 ( .A(n115), .Y(n76) );
  INVX1 U145 ( .A(n110), .Y(n78) );
  INVX1 U146 ( .A(n99), .Y(n67) );
  INVX1 U147 ( .A(n135), .Y(n61) );
  INVX1 U148 ( .A(n130), .Y(n56) );
  INVX1 U149 ( .A(n130), .Y(n55) );
  INVX1 U150 ( .A(n130), .Y(n54) );
  INVX1 U151 ( .A(n123), .Y(n52) );
  INVX1 U152 ( .A(n115), .Y(n51) );
  INVX1 U153 ( .A(n131), .Y(n50) );
  INVX1 U154 ( .A(n139), .Y(n46) );
  INVX1 U155 ( .A(n127), .Y(n40) );
  INVX1 U156 ( .A(n104), .Y(n58) );
  INVX1 U157 ( .A(n110), .Y(n82) );
  INVX1 U158 ( .A(n110), .Y(n84) );
  INVX1 U159 ( .A(n108), .Y(n86) );
  INVX1 U160 ( .A(n108), .Y(n87) );
  INVX1 U161 ( .A(n108), .Y(n88) );
  INVX1 U162 ( .A(n104), .Y(n89) );
  INVX1 U163 ( .A(n99), .Y(n98) );
  INVX1 U164 ( .A(sfr_wdat[3]), .Y(n230) );
  INVX1 U165 ( .A(sfr_wdat[7]), .Y(n263) );
  INVX1 U166 ( .A(sfr_wdat[5]), .Y(n241) );
  INVX1 U167 ( .A(sfr_wdat[1]), .Y(n217) );
  INVX1 U168 ( .A(sfr_wdat[4]), .Y(n236) );
  INVX1 U169 ( .A(sfr_wdat[2]), .Y(n222) );
  INVX1 U170 ( .A(sfr_wdat[0]), .Y(n206) );
  INVX1 U171 ( .A(n300), .Y(n318) );
  NAND5XL U172 ( .A(n246), .B(n254), .C(n224), .D(n207), .E(n356), .Y(n133) );
  INVX1 U173 ( .A(n128), .Y(n356) );
  NOR2X1 U174 ( .A(n248), .B(n364), .Y(r_i2c_fwnak) );
  NOR2X1 U175 ( .A(n259), .B(n364), .Y(r_i2c_fwack) );
  NAND21X1 U176 ( .B(n117), .A(n175), .Y(n105) );
  INVX1 U177 ( .A(n75), .Y(n353) );
  INVX1 U178 ( .A(n322), .Y(n323) );
  AND2X1 U179 ( .A(n293), .B(n237), .Y(clr28[5]) );
  AND2X1 U180 ( .A(n293), .B(n208), .Y(clr28[1]) );
  AND2X1 U181 ( .A(n293), .B(n234), .Y(clr28[4]) );
  AND2X1 U182 ( .A(n293), .B(n202), .Y(clr28[0]) );
  AND2X1 U183 ( .A(n293), .B(n246), .Y(clr28[6]) );
  AND2X1 U184 ( .A(n293), .B(n218), .Y(clr28[2]) );
  AND2X1 U185 ( .A(n293), .B(n254), .Y(clr28[7]) );
  AND2X1 U186 ( .A(n293), .B(n224), .Y(clr28[3]) );
  INVX1 U187 ( .A(n359), .Y(n357) );
  NOR2X1 U188 ( .A(n242), .B(n177), .Y(clr03[5]) );
  NOR2X1 U189 ( .A(n214), .B(n177), .Y(clr03[1]) );
  NOR2X1 U190 ( .A(n235), .B(n177), .Y(clr03[4]) );
  NOR2X1 U191 ( .A(n207), .B(n177), .Y(clr03[0]) );
  NOR2X1 U192 ( .A(n251), .B(n177), .Y(clr03[6]) );
  NOR2X1 U193 ( .A(n223), .B(n177), .Y(clr03[2]) );
  NOR2X1 U194 ( .A(n260), .B(n177), .Y(clr03[7]) );
  INVX1 U195 ( .A(n111), .Y(n362) );
  NOR21XL U196 ( .B(n224), .A(n174), .Y(clrAE[3]) );
  NOR21XL U197 ( .B(n224), .A(n177), .Y(clr03[3]) );
  INVX1 U198 ( .A(n363), .Y(n198) );
  NOR2X1 U199 ( .A(n241), .B(n174), .Y(clrAE[5]) );
  NOR2X1 U200 ( .A(n213), .B(n174), .Y(clrAE[1]) );
  INVX1 U201 ( .A(sfr_wdat[0]), .Y(n207) );
  NOR2X1 U202 ( .A(n235), .B(n174), .Y(clrAE[4]) );
  NOR2X1 U203 ( .A(n207), .B(n174), .Y(clrAE[0]) );
  INVX1 U204 ( .A(n364), .Y(n199) );
  NOR2X1 U205 ( .A(n250), .B(n174), .Y(clrAE[6]) );
  NOR2X1 U206 ( .A(n223), .B(n174), .Y(clrAE[2]) );
  NOR2X1 U207 ( .A(n259), .B(n174), .Y(clrAE[7]) );
  NOR2X1 U208 ( .A(n75), .B(n100), .Y(we[165]) );
  INVX1 U209 ( .A(n101), .Y(n342) );
  NOR21XL U210 ( .B(n351), .A(n100), .Y(we[164]) );
  INVX1 U211 ( .A(sfr_wdat[2]), .Y(n223) );
  NOR2X1 U212 ( .A(n100), .B(n101), .Y(we[162]) );
  INVX1 U213 ( .A(sfr_wdat[5]), .Y(n242) );
  AND2X1 U214 ( .A(n302), .B(n327), .Y(we_181) );
  AND2X1 U215 ( .A(n283), .B(n347), .Y(we_215) );
  AND2X1 U216 ( .A(n283), .B(n302), .Y(we_213) );
  INVX1 U217 ( .A(sfr_wdat[4]), .Y(n235) );
  BUFX3 U218 ( .A(n253), .Y(n247) );
  INVX1 U219 ( .A(sfr_wdat[6]), .Y(n253) );
  INVX1 U220 ( .A(n175), .Y(n163) );
  INVX1 U221 ( .A(n175), .Y(n166) );
  INVX1 U222 ( .A(n136), .Y(n33) );
  INVX1 U223 ( .A(n136), .Y(n35) );
  INVX1 U224 ( .A(n136), .Y(n34) );
  INVX1 U225 ( .A(n135), .Y(n36) );
  INVX1 U226 ( .A(n135), .Y(n37) );
  INVX1 U227 ( .A(n135), .Y(n38) );
  INVX1 U228 ( .A(n137), .Y(n131) );
  INVX1 U229 ( .A(n137), .Y(n108) );
  INVX1 U230 ( .A(n137), .Y(n127) );
  INVX1 U231 ( .A(n26), .Y(n104) );
  INVX1 U232 ( .A(n26), .Y(n123) );
  INVX1 U233 ( .A(n137), .Y(n115) );
  INVX1 U234 ( .A(n137), .Y(n99) );
  INVX1 U235 ( .A(n137), .Y(n110) );
  INVX1 U236 ( .A(n26), .Y(n130) );
  INVX1 U237 ( .A(sfr_addr[0]), .Y(n201) );
  NAND21X1 U238 ( .B(n276), .A(n277), .Y(n300) );
  NOR2X1 U239 ( .A(n75), .B(n134), .Y(r_dacwr[5]) );
  AND2X1 U240 ( .A(n344), .B(n346), .Y(r_dacwr[8]) );
  INVX1 U241 ( .A(n85), .Y(n346) );
  NAND21X1 U242 ( .B(n336), .A(n294), .Y(n101) );
  NOR2X1 U243 ( .A(n101), .B(n134), .Y(r_dacwr[2]) );
  NOR21XL U244 ( .B(n351), .A(n134), .Y(r_dacwr[4]) );
  NOR2X1 U245 ( .A(n83), .B(n134), .Y(r_dacwr[3]) );
  NOR2X1 U246 ( .A(n85), .B(n134), .Y(r_dacwr[1]) );
  NOR2X1 U247 ( .A(n79), .B(n134), .Y(r_dacwr[0]) );
  NOR2X1 U248 ( .A(n81), .B(n134), .Y(r_dacwr[7]) );
  NOR2X1 U249 ( .A(n74), .B(n134), .Y(r_dacwr[6]) );
  NAND21X1 U250 ( .B(n331), .A(n366), .Y(r_fiforst) );
  INVX1 U251 ( .A(prl_c0set), .Y(n366) );
  NOR6XL U252 ( .A(n129), .B(n225), .C(n128), .D(n254), .E(sfr_wdat[4]), .F(
        n246), .Y(n331) );
  NAND43X1 U253 ( .B(n337), .C(n330), .D(n208), .A(n241), .Y(n128) );
  NAND21X1 U254 ( .B(n200), .A(n325), .Y(n336) );
  INVX1 U255 ( .A(n330), .Y(n347) );
  INVX1 U256 ( .A(n121), .Y(r_fifopsh) );
  NOR2X1 U257 ( .A(n74), .B(n132), .Y(r_fcpwr[3]) );
  INVX1 U258 ( .A(n81), .Y(n339) );
  INVX1 U259 ( .A(n320), .Y(n332) );
  NAND21X1 U260 ( .B(n319), .A(n318), .Y(n320) );
  NAND21X1 U261 ( .B(n85), .A(n338), .Y(n364) );
  NAND21X1 U262 ( .B(n75), .A(n299), .Y(n103) );
  NAND21X1 U263 ( .B(n324), .A(n325), .Y(n177) );
  NAND21X1 U264 ( .B(n101), .A(n338), .Y(n363) );
  INVX1 U265 ( .A(n292), .Y(n293) );
  AND2X1 U266 ( .A(n350), .B(n353), .Y(r_fcpwr[4]) );
  NAND21X1 U267 ( .B(n83), .A(n299), .Y(n117) );
  NOR2X1 U268 ( .A(n75), .B(n80), .Y(r_pwrv_upd) );
  INVX1 U269 ( .A(n297), .Y(n298) );
  NAND21X1 U270 ( .B(n74), .A(n272), .Y(n174) );
  OR2X1 U271 ( .A(n325), .B(n324), .Y(n111) );
  NOR2X1 U272 ( .A(n80), .B(n101), .Y(r_dacwr[12]) );
  NOR2X1 U273 ( .A(n74), .B(n95), .Y(r_set_cpmsgid) );
  NOR21XL U274 ( .B(n224), .A(n173), .Y(clrDF[3]) );
  AND2X1 U275 ( .A(n344), .B(n353), .Y(we_245) );
  NOR2X1 U276 ( .A(n241), .B(n173), .Y(clrDF[5]) );
  NOR2X1 U277 ( .A(n212), .B(n173), .Y(clrDF[1]) );
  NOR2X1 U278 ( .A(n235), .B(n173), .Y(clrDF[4]) );
  NOR2X1 U279 ( .A(n206), .B(n173), .Y(clrDF[0]) );
  NOR2X1 U280 ( .A(n249), .B(n173), .Y(clrDF[6]) );
  NOR2X1 U281 ( .A(n222), .B(n173), .Y(clrDF[2]) );
  NOR2X1 U282 ( .A(n258), .B(n173), .Y(clrDF[7]) );
  NOR2X1 U283 ( .A(n81), .B(n132), .Y(r_fcpwr[5]) );
  NOR2X1 U284 ( .A(n75), .B(n132), .Y(r_fcpwr[2]) );
  AO21X1 U285 ( .B(n299), .C(n342), .A(n163), .Y(upd18) );
  INVX1 U286 ( .A(n83), .Y(n343) );
  INVX1 U287 ( .A(n74), .Y(n349) );
  AND3X1 U288 ( .A(n280), .B(n349), .C(n279), .Y(we_222) );
  AND3X1 U289 ( .A(n280), .B(n279), .C(n346), .Y(we_217) );
  INVX1 U290 ( .A(n337), .Y(n327) );
  INVX1 U291 ( .A(n79), .Y(n345) );
  NOR21XL U292 ( .B(n351), .A(n80), .Y(we_228) );
  AND2X1 U293 ( .A(n287), .B(n325), .Y(we_211) );
  AND2X1 U294 ( .A(n350), .B(n349), .Y(r_fcpwr[6]) );
  AND2X1 U295 ( .A(n350), .B(n346), .Y(r_dacwr[14]) );
  AND2X1 U296 ( .A(n350), .B(n345), .Y(r_dacwr[13]) );
  AND2X1 U297 ( .A(n344), .B(n343), .Y(r_dacwr[10]) );
  AND2X1 U298 ( .A(n344), .B(n342), .Y(r_dacwr[9]) );
  AND2X1 U299 ( .A(n344), .B(n349), .Y(we_246) );
  AND2X1 U300 ( .A(n272), .B(n339), .Y(we_175) );
  AND2X1 U301 ( .A(n272), .B(n343), .Y(we_171) );
  AND2X1 U302 ( .A(n338), .B(n343), .Y(we_203) );
  NOR2X1 U303 ( .A(n83), .B(n95), .Y(we_187) );
  NOR2X1 U304 ( .A(n83), .B(n132), .Y(r_fcpwr[0]) );
  NOR2X1 U305 ( .A(n83), .B(n100), .Y(we[163]) );
  NOR2X1 U306 ( .A(n80), .B(n81), .Y(we_231) );
  NOR2X1 U307 ( .A(n80), .B(n83), .Y(we_227) );
  INVX1 U308 ( .A(n285), .Y(n283) );
  AND2X1 U309 ( .A(n283), .B(n20), .Y(we_214) );
  AND2X1 U310 ( .A(n20), .B(n327), .Y(we_182) );
  NOR2X1 U311 ( .A(n81), .B(n95), .Y(we_191) );
  NOR2X1 U312 ( .A(n74), .B(n80), .Y(we_230) );
  NOR2X1 U313 ( .A(n81), .B(n100), .Y(we[167]) );
  NOR2X1 U314 ( .A(n74), .B(n100), .Y(we[166]) );
  NAND21X1 U315 ( .B(n319), .A(n354), .Y(n100) );
  INVX1 U316 ( .A(n273), .Y(n354) );
  INVX1 U317 ( .A(n348), .Y(n279) );
  INVX1 U318 ( .A(n282), .Y(n302) );
  NAND21X1 U319 ( .B(n325), .A(n281), .Y(n282) );
  INVX1 U320 ( .A(N30), .Y(n379) );
  INVX1 U321 ( .A(ictlr_inc), .Y(n175) );
  INVX1 U322 ( .A(n139), .Y(n32) );
  INVX1 U323 ( .A(atpg_en), .Y(n264) );
  INVX1 U324 ( .A(n139), .Y(n137) );
  INVX1 U325 ( .A(n26), .Y(n136) );
  INVX1 U326 ( .A(n26), .Y(n135) );
  INVX1 U327 ( .A(n284), .Y(n360) );
  NAND32X1 U328 ( .B(n300), .C(n295), .A(n351), .Y(n284) );
  INVX1 U329 ( .A(n289), .Y(n276) );
  INVX1 U330 ( .A(n288), .Y(n277) );
  NAND32X1 U331 ( .B(n201), .C(n278), .A(n326), .Y(n85) );
  NAND21XL U332 ( .B(n301), .A(n347), .Y(n81) );
  NAND21XL U333 ( .B(n301), .A(n20), .Y(n74) );
  NAND32X1 U334 ( .B(n201), .C(n326), .A(n294), .Y(n83) );
  INVX1 U335 ( .A(n278), .Y(n294) );
  INVX1 U336 ( .A(n335), .Y(n333) );
  NAND21X1 U337 ( .B(n348), .A(n341), .Y(n134) );
  NAND21X1 U338 ( .B(n289), .A(n277), .Y(n348) );
  NAND32XL U339 ( .B(n319), .C(n301), .A(n318), .Y(n337) );
  NAND21X1 U340 ( .B(n326), .A(n281), .Y(n330) );
  NOR2X1 U341 ( .A(n335), .B(n336), .Y(n20) );
  INVX1 U342 ( .A(n267), .Y(n344) );
  NAND21X1 U343 ( .B(n300), .A(n341), .Y(n267) );
  INVX1 U344 ( .A(n270), .Y(n281) );
  NAND32X1 U345 ( .B(n337), .C(n336), .A(n335), .Y(n121) );
  INVX1 U346 ( .A(n326), .Y(n325) );
  INVX1 U347 ( .A(n102), .Y(n319) );
  INVX1 U348 ( .A(n290), .Y(n338) );
  NAND32X1 U349 ( .B(n289), .C(n295), .A(n288), .Y(n290) );
  NAND21X1 U350 ( .B(n348), .A(n352), .Y(n132) );
  NAND32X1 U351 ( .B(n337), .C(n201), .A(n335), .Y(n324) );
  ENOX1 U352 ( .A(n103), .B(n262), .C(pff_rxpart[15]), .D(n103), .Y(wd21[7])
         );
  NAND32X1 U353 ( .B(n81), .C(n295), .A(n279), .Y(n173) );
  INVX1 U354 ( .A(n275), .Y(n350) );
  NAND21X1 U355 ( .B(n300), .A(n352), .Y(n275) );
  MUX2X1 U356 ( .D0(pff_rxpart[1]), .D1(n211), .S(n298), .Y(wd20[1]) );
  AND3X1 U357 ( .A(n354), .B(n353), .C(n352), .Y(r_cvcwr[1]) );
  NAND4X1 U358 ( .A(n117), .B(n118), .C(n119), .D(n175), .Y(upd19) );
  NAND32XL U359 ( .B(n301), .C(n300), .A(n280), .Y(n285) );
  INVX1 U360 ( .A(n286), .Y(n287) );
  NAND32X1 U361 ( .B(n201), .C(n285), .A(n335), .Y(n286) );
  AND4X1 U362 ( .A(n276), .B(n339), .C(n352), .D(n288), .Y(we_143) );
  AND4X1 U363 ( .A(n341), .B(n276), .C(n288), .D(n345), .Y(we_232) );
  AND3XL U364 ( .A(n354), .B(n351), .C(n352), .Y(r_cvcwr[0]) );
  AND2X1 U365 ( .A(n287), .B(n326), .Y(we_209) );
  NAND21X1 U366 ( .B(n348), .A(n102), .Y(n95) );
  NAND21X1 U367 ( .B(n273), .A(n341), .Y(n80) );
  INVX1 U368 ( .A(n296), .Y(n299) );
  NAND21X1 U369 ( .B(n295), .A(n354), .Y(n296) );
  INVX1 U370 ( .A(n271), .Y(n272) );
  NAND32X1 U371 ( .B(n289), .C(n319), .A(n288), .Y(n271) );
  INVX1 U372 ( .A(n295), .Y(n280) );
  NAND21X1 U373 ( .B(n277), .A(n289), .Y(n273) );
  INVX1 U374 ( .A(n116), .Y(n71) );
  XOR2X1 U375 ( .A(N31), .B(N32), .Y(N33) );
  XNOR2XL U376 ( .A(n379), .B(N29), .Y(N35) );
  XNOR2XL U377 ( .A(N31), .B(n379), .Y(N34) );
  INVX1 U378 ( .A(n26), .Y(n138) );
  INVX1 U379 ( .A(n26), .Y(n139) );
  BUFX3 U380 ( .A(pff_empty), .Y(dbgpo[23]) );
  BUFX3 U381 ( .A(pff_full), .Y(dbgpo[22]) );
  NAND21XL U382 ( .B(n265), .A(sfr_addr[4]), .Y(n288) );
  INVX1 U383 ( .A(n266), .Y(n341) );
  INVX1 U384 ( .A(n334), .Y(r_fifopop) );
  NAND43X1 U385 ( .B(n365), .C(n333), .D(n336), .A(n332), .Y(n334) );
  INVX1 U386 ( .A(n172), .Y(bus_idle) );
  INVX1 U387 ( .A(n291), .Y(n340) );
  NAND21X1 U388 ( .B(n365), .A(n338), .Y(n291) );
  NAND42X1 U389 ( .C(n133), .D(n218), .A(n165), .B(n235), .Y(n119) );
  NAND2X1 U390 ( .A(n380), .B(n119), .Y(n141) );
  NOR32XL U391 ( .B(n350), .C(n347), .A(n365), .Y(r_fcpre) );
  NAND2X1 U392 ( .A(n107), .B(n357), .Y(n106) );
  INVX1 U393 ( .A(n274), .Y(n352) );
  MUX2X1 U394 ( .D0(n228), .D1(pff_rxpart[11]), .S(n103), .Y(wd21[3]) );
  OAI22X1 U395 ( .A(n175), .B(n10), .C(n262), .D(n105), .Y(wd19[7]) );
  AO22AXL U396 ( .A(inst_ofs_plus[11]), .B(n163), .C(n224), .D(n105), .Y(
        wd19[3]) );
  ENOX1 U397 ( .A(n17), .B(n235), .C(pff_rxpart[12]), .D(n103), .Y(wd21[4]) );
  ENOX1 U398 ( .A(n17), .B(n223), .C(pff_rxpart[10]), .D(n103), .Y(wd21[2]) );
  ENOX1 U399 ( .A(n17), .B(n215), .C(pff_rxpart[9]), .D(n103), .Y(wd21[1]) );
  ENOX1 U400 ( .A(n17), .B(n242), .C(pff_rxpart[13]), .D(n103), .Y(wd21[5]) );
  ENOX1 U401 ( .A(n17), .B(n252), .C(pff_rxpart[14]), .D(n103), .Y(wd21[6]) );
  NAND2X1 U402 ( .A(n114), .B(n17), .Y(upd21) );
  NAND4X1 U403 ( .A(n202), .B(n218), .C(n192), .D(n193), .Y(n118) );
  NOR4XL U404 ( .A(n254), .B(n224), .C(n247), .D(n235), .Y(n193) );
  NOR21XL U405 ( .B(n165), .A(n128), .Y(n192) );
  OA21X1 U407 ( .B(prx_rst[0]), .C(prx_rst[1]), .A(set03[1]), .Y(set03[7]) );
  NAND43X1 U408 ( .B(set_hold), .C(cpurst), .D(n357), .A(n107), .Y(upd12) );
  MUX2X1 U409 ( .D0(pff_rxpart[0]), .D1(n205), .S(n298), .Y(wd20[0]) );
  MUX2X1 U410 ( .D0(pff_rxpart[2]), .D1(n221), .S(n298), .Y(wd20[2]) );
  MUX2X1 U411 ( .D0(pff_rxpart[7]), .D1(sfr_wdat[7]), .S(n298), .Y(wd20[7]) );
  MUX2X1 U412 ( .D0(pff_rxpart[3]), .D1(n229), .S(n298), .Y(wd20[3]) );
  MUX2X1 U413 ( .D0(pff_rxpart[4]), .D1(n234), .S(n298), .Y(wd20[4]) );
  NAND21X1 U414 ( .B(n298), .A(n114), .Y(upd20) );
  OAI32X1 U415 ( .A(n369), .B(r_fifopsh), .C(n362), .D(n261), .E(n111), .Y(
        wd01[7]) );
  ENOX1 U416 ( .A(n242), .B(n105), .C(inst_ofs_plus[13]), .D(n166), .Y(wd19[5]) );
  ENOX1 U417 ( .A(n235), .B(n105), .C(inst_ofs_plus[12]), .D(n166), .Y(wd19[4]) );
  ENOX1 U418 ( .A(n216), .B(n105), .C(inst_ofs_plus[9]), .D(n166), .Y(wd19[1])
         );
  ENOX1 U419 ( .A(n222), .B(n105), .C(inst_ofs_plus[10]), .D(n166), .Y(wd19[2]) );
  ENOX1 U420 ( .A(n206), .B(n105), .C(inst_ofs_plus[8]), .D(n166), .Y(wd19[0])
         );
  OAI211X1 U421 ( .C(n369), .D(n121), .A(n16), .B(n112), .Y(upd01) );
  AND3X1 U422 ( .A(n20), .B(n10), .C(n340), .Y(upd31) );
  MUX2X1 U423 ( .D0(n225), .D1(inst_ofs_plus[3]), .S(n163), .Y(wd18[3]) );
  ENOX1 U424 ( .A(n163), .B(n223), .C(inst_ofs_plus[2]), .D(ictlr_inc), .Y(
        wd18[2]) );
  ENOX1 U425 ( .A(n163), .B(n235), .C(inst_ofs_plus[4]), .D(ictlr_inc), .Y(
        wd18[4]) );
  ENOX1 U426 ( .A(n163), .B(n242), .C(inst_ofs_plus[5]), .D(n166), .Y(wd18[5])
         );
  ENOX1 U427 ( .A(n163), .B(n215), .C(inst_ofs_plus[1]), .D(ictlr_inc), .Y(
        wd18[1]) );
  ENOX1 U428 ( .A(n163), .B(n261), .C(inst_ofs_plus[7]), .D(n166), .Y(wd18[7])
         );
  ENOX1 U429 ( .A(n163), .B(n252), .C(inst_ofs_plus[6]), .D(n166), .Y(wd18[6])
         );
  NAND2X1 U430 ( .A(prx_setsta[3]), .B(n13), .Y(n116) );
  AND2X1 U431 ( .A(prx_setsta[6]), .B(n13), .Y(set03[6]) );
  XNOR2XL U432 ( .A(N24), .B(n383), .Y(N25) );
  XNOR2XL U433 ( .A(N25), .B(n382), .Y(N26) );
  AND2X1 U434 ( .A(i_goidle), .B(n13), .Y(set04[1]) );
  XNOR2XL U435 ( .A(n385), .B(add_179_carry[4]), .Y(N32) );
  XNOR2XL U436 ( .A(N27), .B(N29), .Y(N36) );
  NOR2X1 U437 ( .A(n13), .B(i_goidle), .Y(n167) );
  NAND2X1 U438 ( .A(n126), .B(n361), .Y(N81) );
  INVX1 U439 ( .A(n142), .Y(n381) );
  XNOR2XL U440 ( .A(di_p0[3]), .B(n372), .Y(n185) );
  XNOR2XL U441 ( .A(di_p0[5]), .B(n371), .Y(n187) );
  XNOR2XL U442 ( .A(di_p0[7]), .B(n370), .Y(n189) );
  XNOR2XL U443 ( .A(di_p0[4]), .B(n377), .Y(n188) );
  XNOR2XL U444 ( .A(di_p0[6]), .B(n375), .Y(n190) );
  XNOR2XL U445 ( .A(di_p0[2]), .B(n376), .Y(n186) );
  NAND2X1 U446 ( .A(n264), .B(aswkup), .Y(pwrdn_rstz) );
  AND2X1 U447 ( .A(dnchk_en), .B(dm_fault), .Y(dmf_wkup) );
  INVX1 U448 ( .A(n142), .Y(n26) );
  MUX2X1 U449 ( .D0(i_pc[0]), .D1(prx_adpn[0]), .S(n12), .Y(reg30[0]) );
  MUX2X1 U450 ( .D0(i_pc[3]), .D1(prx_adpn[3]), .S(n11), .Y(reg30[3]) );
  AND2X1 U451 ( .A(i_pc[6]), .B(n10), .Y(reg30[6]) );
  AND2X1 U452 ( .A(i_pc[7]), .B(n10), .Y(reg30[7]) );
  MUX2X1 U453 ( .D0(s_scp), .D1(m_scp), .S(reg94[5]), .Y(regAD[4]) );
  MUX2X1 U454 ( .D0(i_pc[2]), .D1(prx_adpn[2]), .S(reg19_7_), .Y(reg30[2]) );
  MUX2X1 U455 ( .D0(i_pc[5]), .D1(prx_adpn[5]), .S(n12), .Y(reg30[5]) );
  MUX2X1 U456 ( .D0(s_ovp), .D1(m_ovp), .S(reg94[4]), .Y(regAD[2]) );
  INVX1 U457 ( .A(n140), .Y(n355) );
  OAI211X1 U458 ( .C(ictlr_idle), .D(n329), .A(oscdwn_shft[1]), .B(bus_idle), 
        .Y(n140) );
  AND2X1 U459 ( .A(n126), .B(regD4_1_), .Y(n329) );
  MUX2X1 U460 ( .D0(i_pc[4]), .D1(prx_adpn[4]), .S(n11), .Y(reg30[4]) );
  OR4X1 U461 ( .A(osc_gate_n_1_), .B(osc_gate_n_0_), .C(test_so1), .D(
        osc_gate_n_2_), .Y(r_osc_gate) );
  AOI211X1 U462 ( .C(n383), .D(n382), .A(rstcnt[3]), .B(n385), .Y(n197) );
  INVX1 U463 ( .A(rstcnt[4]), .Y(n385) );
  INVX1 U464 ( .A(rstcnt[2]), .Y(n383) );
  INVX1 U465 ( .A(rstcnt[1]), .Y(n382) );
  NAND42X1 U466 ( .C(n14), .D(n328), .A(i_i2c_idle), .B(n196), .Y(n172) );
  INVX1 U467 ( .A(prx_rcvinf[4]), .Y(n328) );
  NOR3XL U468 ( .A(ptx_fsm[0]), .B(ptx_fsm[2]), .C(ptx_fsm[1]), .Y(n196) );
  INVX1 U469 ( .A(sfr_r), .Y(n365) );
  NOR21XL U470 ( .B(pff_ack[1]), .A(prl_cany0), .Y(set04[5]) );
  NAND4X1 U471 ( .A(n155), .B(n156), .C(n157), .D(n158), .Y(o_intr[1]) );
  AOI22X1 U472 ( .A(reg06[0]), .B(irq04[0]), .C(reg06[1]), .D(irq04[1]), .Y(
        n158) );
  AOI22X1 U473 ( .A(reg06[6]), .B(irq04[6]), .C(reg06[7]), .D(irq04[7]), .Y(
        n155) );
  AOI22X1 U474 ( .A(reg06[4]), .B(irq04[4]), .C(reg06[5]), .D(irq04[5]), .Y(
        n156) );
  INVX1 U475 ( .A(drstz[1]), .Y(n384) );
  AND3X1 U476 ( .A(n347), .B(n11), .C(n340), .Y(r_psrd) );
  NOR2X1 U477 ( .A(regD4_2_), .B(regD4_0_), .Y(n126) );
  NAND32X1 U478 ( .B(bkpt_hold), .C(reg12[3]), .A(n126), .Y(r_hold_mcu) );
  AND3X1 U479 ( .A(n339), .B(n12), .C(n338), .Y(r_pswr) );
  AND2X1 U480 ( .A(regD4_2_), .B(oscdwn_shft[2]), .Y(r_pos_gate) );
  ENOX1 U481 ( .A(n207), .B(n363), .C(n363), .D(lt_reg26_0), .Y(i2c_mode_wdat)
         );
  AOI21X1 U482 ( .B(n171), .C(n363), .A(n172), .Y(i2c_mode_upd) );
  XNOR2XL U483 ( .A(r_hwi2c_en), .B(lt_reg26_0), .Y(n171) );
  OAI32X1 U484 ( .A(n378), .B(r_phyrst[1]), .C(n367), .D(r_phyrst[0]), .E(n164), .Y(n1210) );
  INVX1 U485 ( .A(n167), .Y(n367) );
  AOI21X1 U486 ( .B(reg11_7_), .C(set03[7]), .A(n141), .Y(n164) );
  OAI21BX1 U487 ( .C(reg12[3]), .B(n107), .A(n109), .Y(wd12[3]) );
  AOI32X1 U488 ( .A(set_hold), .B(n107), .C(n359), .D(n224), .E(n358), .Y(n109) );
  INVX1 U489 ( .A(n106), .Y(n358) );
  ENOX1 U490 ( .A(n17), .B(n207), .C(pff_rxpart[8]), .D(n103), .Y(wd21[0]) );
  NOR21XL U491 ( .B(n112), .A(n113), .Y(wd01[6]) );
  AOI22X1 U492 ( .A(n362), .B(n246), .C(r_first), .D(n111), .Y(n113) );
  NAND2X1 U493 ( .A(n21), .B(n107), .Y(wd12[4]) );
  MUX2IX1 U494 ( .D0(reg12[4]), .D1(n234), .S(n357), .Y(n21) );
  NAND4X1 U495 ( .A(n159), .B(n160), .C(n161), .D(n162), .Y(o_intr[0]) );
  AOI22X1 U496 ( .A(reg05[4]), .B(irq03[4]), .C(reg05[5]), .D(irq03[5]), .Y(
        n160) );
  AOI22X1 U497 ( .A(reg05[2]), .B(irq03[2]), .C(reg05[3]), .D(irq03[3]), .Y(
        n161) );
  OAI21X1 U498 ( .B(r_fifopsh), .C(r_fifopop), .A(r_first), .Y(n112) );
  AOI22X1 U499 ( .A(reg05[0]), .B(irq03[0]), .C(reg05[1]), .D(irq03[1]), .Y(
        n162) );
  AOI22X1 U500 ( .A(reg05[6]), .B(irq03[6]), .C(reg05[7]), .D(irq03[7]), .Y(
        n159) );
  NOR21XL U501 ( .B(prx_setsta[1]), .A(n14), .Y(set03[1]) );
  NOR21XL U502 ( .B(prx_setsta[2]), .A(prl_cany0), .Y(set03[2]) );
  OAI21X1 U503 ( .B(n191), .C(n172), .A(n118), .Y(N23) );
  NOR21XL U504 ( .B(n120), .A(rstcnt[4]), .Y(n191) );
  ENOX1 U505 ( .A(n252), .B(n105), .C(inst_ofs_plus[14]), .D(n166), .Y(wd19[6]) );
  ENOX1 U506 ( .A(n223), .B(n106), .C(r_txshrt), .D(n106), .Y(wd12[2]) );
  ENOX1 U507 ( .A(n242), .B(n106), .C(reg12[5]), .D(n106), .Y(wd12[5]) );
  ENOX1 U508 ( .A(n235), .B(n16), .C(r_txnumk[4]), .D(n111), .Y(wd01[4]) );
  ENOX1 U509 ( .A(n242), .B(n16), .C(r_unlock), .D(n111), .Y(wd01[5]) );
  ENOX1 U510 ( .A(n206), .B(n106), .C(r_pshords), .D(n106), .Y(wd12[0]) );
  ENOX1 U511 ( .A(n216), .B(n15), .C(reg12_1), .D(n106), .Y(wd12[1]) );
  ENOX1 U512 ( .A(n252), .B(n15), .C(reg12[6]), .D(n106), .Y(wd12[6]) );
  ENOX1 U513 ( .A(n262), .B(n15), .C(reg12[7]), .D(n106), .Y(wd12[7]) );
  AO22AXL U514 ( .A(r_txnumk[0]), .B(n111), .C(sfr_wdat[0]), .D(n111), .Y(
        wd01[0]) );
  NAND3X1 U515 ( .A(n168), .B(n169), .C(n170), .Y(i2c_stretch) );
  AOI22X1 U516 ( .A(reg28[2]), .B(reg27[2]), .C(reg28[3]), .D(reg27[3]), .Y(
        n168) );
  AOI22X1 U517 ( .A(reg28[0]), .B(reg27[0]), .C(reg28[1]), .D(reg27[1]), .Y(
        n169) );
  AOI222XL U518 ( .A(reg28[7]), .B(reg27[7]), .C(reg28[4]), .D(reg27[4]), .E(
        reg28[6]), .F(reg27[6]), .Y(n170) );
  ENOX1 U519 ( .A(n163), .B(n207), .C(inst_ofs_plus[0]), .D(n166), .Y(wd18[0])
         );
  NOR21XL U520 ( .B(pff_obsd), .A(n14), .Y(set04[3]) );
  NOR21XL U521 ( .B(oscdwn_shft[2]), .A(n361), .Y(r_osc_lo) );
  AOI22X1 U522 ( .A(reg06[2]), .B(irq04[2]), .C(reg06[3]), .D(irq04[3]), .Y(
        n157) );
  INVX1 U523 ( .A(regD4_1_), .Y(n361) );
  AND2X1 U524 ( .A(regD4_0_), .B(oscdwn_shft[2]), .Y(r_osc_stop) );
  NOR21XL U525 ( .B(prx_setsta[4]), .A(prl_cany0), .Y(set03[4]) );
  AOI21BBXL U526 ( .B(r_auto_gdcrc[1]), .C(n116), .A(set03[6]), .Y(n114) );
  AO21X1 U527 ( .B(n124), .C(n125), .A(reg11_4), .Y(r_rxords_ena[4]) );
  NOR3XL U528 ( .A(r_rxords_ena[0]), .B(r_rxords_ena[2]), .C(r_rxords_ena[1]), 
        .Y(n124) );
  NOR3XL U529 ( .A(r_rxords_ena[3]), .B(r_rxords_ena[6]), .C(r_rxords_ena[5]), 
        .Y(n125) );
  OAI31XL U530 ( .A(n197), .B(r_phyrst[1]), .C(n384), .D(n264), .Y(prstz) );
  NOR21XL U531 ( .B(prl_GCTxDone), .A(n14), .Y(set04[6]) );
  NOR21XL U532 ( .B(prx_setsta[5]), .A(prl_cany0), .Y(set03[5]) );
  AOI22X1 U533 ( .A(reg27[6]), .B(irq28[6]), .C(reg27[7]), .D(irq28[7]), .Y(
        n151) );
  NAND4X1 U534 ( .A(n151), .B(n152), .C(n153), .D(n154), .Y(o_intr[2]) );
  AOI22X1 U535 ( .A(reg27[4]), .B(irq28[4]), .C(reg27[5]), .D(irq28[5]), .Y(
        n152) );
  AOI22X1 U536 ( .A(reg27[0]), .B(irq28[0]), .C(reg27[1]), .D(irq28[1]), .Y(
        n154) );
  NOR21XL U537 ( .B(ptx_ack), .A(prl_cany0), .Y(set04[0]) );
  NOR21XL U538 ( .B(i_gobusy), .A(prl_cany0), .Y(set04[2]) );
  XNOR2XL U539 ( .A(n385), .B(rstcnt[3]), .Y(N24) );
  XOR2X1 U540 ( .A(N26), .B(rstcnt[0]), .Y(N27) );
  AOI221XL U541 ( .A(regAF[4]), .B(regAE[4]), .C(regAF[2]), .D(regAE[2]), .E(
        n368), .Y(r_srcctl[0]) );
  INVX1 U542 ( .A(regE3_0), .Y(n368) );
  AOI22X1 U543 ( .A(reg27[2]), .B(irq28[2]), .C(reg27[3]), .D(irq28[3]), .Y(
        n153) );
  AND2X1 U544 ( .A(reg94[7]), .B(reg94[6]), .Y(r_otpi_gate) );
  AO22AXL U545 ( .A(reg94[4]), .B(m_ovp_sta), .C(s_ovp_sta), .D(reg94[4]), .Y(
        setAE[2]) );
  AO22AXL U546 ( .A(reg94[5]), .B(m_scp_sta), .C(s_scp_sta), .D(reg94[5]), .Y(
        setAE[4]) );
  AND2X1 U547 ( .A(regD4_4_), .B(oscdwn_shft[2]), .Y(r_ocdrv_enz) );
  NOR21XL U548 ( .B(prl_discard), .A(prl_cany0), .Y(set04[7]) );
  AND2X1 U549 ( .A(regD4_3_), .B(oscdwn_shft[2]), .Y(r_pwrdn) );
  NAND4X1 U550 ( .A(n143), .B(n144), .C(n145), .D(n146), .Y(o_intr[4]) );
  AOI22X1 U551 ( .A(regAF[6]), .B(irqAE[6]), .C(regAF[7]), .D(irqAE[7]), .Y(
        n143) );
  AOI22X1 U552 ( .A(regAF[0]), .B(irqAE[0]), .C(regAF[1]), .D(irqAE[1]), .Y(
        n146) );
  AOI22X1 U553 ( .A(irqAE[2]), .B(regAF[2]), .C(regAF[3]), .D(irqAE[3]), .Y(
        n145) );
  OAI32X1 U554 ( .A(n378), .B(r_phyrst[1]), .C(n167), .D(r_phyrst[0]), .E(n380), .Y(n1209) );
  AOI22X1 U555 ( .A(irqAE[4]), .B(regAF[4]), .C(irqAE[5]), .D(regAF[5]), .Y(
        n144) );
  INVX1 U556 ( .A(reg25_0_), .Y(r_i2c_ninc) );
  NOR21XL U557 ( .B(prx_setsta[0]), .A(prl_cany0), .Y(set03[0]) );
  XNOR2XL U558 ( .A(d_p0[0]), .B(n374), .Y(setDF[0]) );
  XNOR2XL U559 ( .A(d_p0[1]), .B(n373), .Y(setDF[1]) );
  XNOR2XL U560 ( .A(d_p0[2]), .B(n376), .Y(setDF[2]) );
  XNOR2XL U561 ( .A(d_p0[3]), .B(n372), .Y(setDF[3]) );
  XNOR2XL U562 ( .A(d_p0[4]), .B(n377), .Y(setDF[4]) );
  NAND2X1 U563 ( .A(rstcnt[4]), .B(n120), .Y(n107) );
  NOR42XL U564 ( .C(n194), .D(r_inst_ofs[10]), .A(r_inst_ofs[8]), .B(n195), 
        .Y(n165) );
  NAND4X1 U565 ( .A(r_inst_ofs[14]), .B(r_inst_ofs[13]), .C(r_inst_ofs[12]), 
        .D(r_inst_ofs[11]), .Y(n195) );
  NOR2X1 U566 ( .A(n12), .B(r_inst_ofs[9]), .Y(n194) );
  AOI22X1 U567 ( .A(regDE[0]), .B(irqDF[0]), .C(regDE[1]), .D(irqDF[1]), .Y(
        n150) );
  NOR4XL U568 ( .A(rstcnt[0]), .B(rstcnt[1]), .C(rstcnt[2]), .D(rstcnt[3]), 
        .Y(n120) );
  AOI22X1 U569 ( .A(regDE[2]), .B(irqDF[2]), .C(regDE[3]), .D(irqDF[3]), .Y(
        n149) );
  XNOR2XL U570 ( .A(d_p0[6]), .B(n375), .Y(setDF[6]) );
  XNOR2XL U571 ( .A(d_p0[7]), .B(n370), .Y(setDF[7]) );
  XNOR2XL U572 ( .A(d_p0[5]), .B(n371), .Y(setDF[5]) );
  INVX1 U573 ( .A(ff_p0[1]), .Y(n373) );
  INVX1 U574 ( .A(ff_p0[6]), .Y(n375) );
  INVX1 U575 ( .A(ff_p0[0]), .Y(n374) );
  INVX1 U576 ( .A(ff_p0[3]), .Y(n372) );
  INVX1 U577 ( .A(ff_p0[2]), .Y(n376) );
  INVX1 U578 ( .A(ff_p0[5]), .Y(n371) );
  INVX1 U579 ( .A(ff_p0[4]), .Y(n377) );
  INVX1 U580 ( .A(ff_p0[7]), .Y(n370) );
  NAND4X1 U581 ( .A(n147), .B(n148), .C(n149), .D(n150), .Y(o_intr[3]) );
  AOI22X1 U582 ( .A(regDE[6]), .B(irqDF[6]), .C(regDE[7]), .D(irqDF[7]), .Y(
        n147) );
  AOI22X1 U583 ( .A(regDE[4]), .B(irqDF[4]), .C(regDE[5]), .D(irqDF[5]), .Y(
        n148) );
  INVX1 U584 ( .A(r_phyrst[1]), .Y(n380) );
  INVX1 U585 ( .A(r_last), .Y(n369) );
  INVX1 U586 ( .A(r_phyrst[0]), .Y(n378) );
  INVX1 U587 ( .A(regD3_3), .Y(r_gpio_ie[0]) );
  NAND42X1 U588 ( .C(di_stbovp_clr), .D(di_rd_det_clr), .A(n381), .B(n178), 
        .Y(aswkup) );
  NOR3XL U589 ( .A(dm_fault_clr), .B(p0_chg_clr), .C(i_tmrf), .Y(n178) );
  INVX1 U590 ( .A(regD3_7_), .Y(r_gpio_ie[1]) );
  NAND2X1 U591 ( .A(n3), .B(srstz), .Y(n142) );
  OAI21X1 U592 ( .B(osc_low_clr), .C(n142), .A(n264), .Y(osc_low_rstz) );
  AOI22X1 U593 ( .A(regDE[1]), .B(n183), .C(regDE[0]), .D(n184), .Y(n182) );
  XNOR2XL U594 ( .A(di_p0[0]), .B(n374), .Y(n184) );
  XNOR2XL U595 ( .A(di_p0[1]), .B(n373), .Y(n183) );
  AOI22X1 U596 ( .A(regAF[5]), .B(regAE[5]), .C(regAD[5]), .D(i_vcbyval), .Y(
        n122) );
  AND2X1 U597 ( .A(regE3[3]), .B(n122), .Y(r_srcctl[3]) );
  AND2X1 U598 ( .A(regE3[2]), .B(n122), .Y(r_srcctl[2]) );
  NAND4X1 U599 ( .A(n179), .B(n180), .C(n181), .D(n182), .Y(as_p0_chg) );
  AOI22X1 U600 ( .A(regDE[7]), .B(n189), .C(regDE[6]), .D(n190), .Y(n179) );
  AOI22X1 U601 ( .A(regDE[5]), .B(n187), .C(regDE[4]), .D(n188), .Y(n180) );
  AOI22X1 U602 ( .A(regDE[3]), .B(n185), .C(regDE[2]), .D(n186), .Y(n181) );
  INVX1 U603 ( .A(sfr_addr[7]), .Y(n265) );
  NAND21XL U604 ( .B(n268), .A(n176), .Y(n75) );
  NAND32X1 U605 ( .B(n335), .C(n301), .A(n326), .Y(n268) );
  NAND21XL U606 ( .B(n321), .A(n332), .Y(n322) );
  NAND21XL U607 ( .B(n321), .A(n299), .Y(n297) );
  NAND21XL U608 ( .B(n321), .A(n338), .Y(n292) );
  NAND21XL U609 ( .B(n333), .A(sfr_w), .Y(n278) );
  NOR2XL U610 ( .A(n31), .B(sfr_addr[6]), .Y(n102) );
  NAND21XL U611 ( .B(sfr_addr[6]), .A(n31), .Y(n274) );
  NAND21XL U612 ( .B(n31), .A(sfr_addr[6]), .Y(n266) );
  INVXL U613 ( .A(sfr_addr[5]), .Y(n31) );
  NAND21XL U614 ( .B(sfr_addr[5]), .A(sfr_addr[6]), .Y(n295) );
endmodule


module regbank_a0_DW_rightsh_1 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n59, n61,
         n63, n64, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n90, n91, n93, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n106, n107, n108, n109,
         n110, n111, n112, n113, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n195, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n308, n309, n312, n313,
         n314, n316, n317, n318, n319, n320, n497, n503, n509, n510, n515,
         n516, n521, n527, n528, n533, n534, n539, n540, n545, n546, n551,
         n552, n557, n558, n563, n564, n575, n576, n581, n582, n585, n586,
         n589, n590, n597, n598, n601, n602, n605, n609, n610, n617, n618,
         n621, n622, n625, n626, n629, n630, n633, n634, n637, n638, n641,
         n642, n645, n646, n649, n650, n653, n654, n657, n658, n661, n662,
         n665, n666, n669, n670, n673, n674, n677, n678, n681, n684, n687,
         n690, n693, n696, n699, n702, n705, n706, n709, n710, n713, n714,
         n717, n718, n721, n722, n725, n726, n729, n730, n733, n734, n737,
         n740, n743, n746, n749, n752, n755, n758, n761, n762, n765, n766,
         n769, n770, n773, n774, n777, n778, n781, n782, n785, n786, n789,
         n790, n795, n796, n801, n802, n807, n808, n813, n814, n819, n825,
         n826, n831, n832, n837, n838, n843, n844, n855, n856, n861, n862,
         n867, n868, n873, n879, n880, n885, n886, n891, n892, n897, n898,
         n903, n904, n910, n915, n916, n927, n928, n933, n934, n937, n938,
         n941, n942, n945, n946, n949, n950, n953, n954, n957, n961, n962,
         n965, n966, n969, n970, n973, n974, n977, n978, n981, n982, n985,
         n986, n989, n993, n994, n997, n998, n1009, n1010, n1015, n1016, n1021,
         n1022, n1027, n1028, n1034, n1039, n1040, n1045, n1046, n1049, n1050,
         n1053, n1054, n1057, n1058, n1061, n1062, n1065, n1066, n1069, n1070,
         n1073, n1074, n1077, n1078, n1081, n1082, n1085, n1086, n1093, n1094,
         n1097, n1098, n1101, n1102, n1105, n1106, n1109, n1110, n1113, n1114,
         n1117, n1118, n1121, n1122, n1125, n1126, n1129, n1130, n1133, n1134,
         n1137, n1138, n1141, n1142, n1145, n1146, n1149, n1153, n1154, n1157,
         n1158, n1161, n1162, n1166, n1169, n1170, n1173, n1177, n1178, n1181,
         n1182, n1185, n1186, n1189, n1190, n1193, n1194, n1197, n1198, n1201,
         n1202, n1205, n1206, n1209, n1210, n1213, n1214, n1217, n1218, n1221,
         n1222, n1225, n1226, n1230, n1233, n1234, n1237, n1238, n1241, n1244,
         n1247, n1250, n1253, n1256, n1259, n1262, n1269, n1272, n1275, n1278,
         n1281, n1284, n1287, n1290, n1293, n1296, n1299, n1302, n1305, n1308,
         n1311, n1312, n1315, n1316, n1319, n1320, n1323, n1324, n1327, n1328,
         n1331, n1335, n1336, n1339, n1340, n1343, n1344, n1347, n1348, n1351,
         n1352, n1355, n1356, n1359, n1360, n1363, n1367, n1368, n1371, n1372,
         n1377, n1378, n1395, n1396, n1401, n1402, n1407, n1413, n1414, n1419,
         n1420, n1425, n1426, n1431, n1432, n1437, n1438, n1443, n1449, n1450,
         n1461, n1462, n1467, n1468, n1471, n1472, n1475, n1476, n1479, n1480,
         n1483, n1487, n1488, n1491, n1495, n1499, n1500, n1503, n1504, n1507,
         n1508, n1511, n1512, n1515, n1516, n1519, n1520, n1523, n1524, n1527,
         n1528, n1531, n1532, n1535, n1536, n1539, n1540, n1543, n1544, n1547,
         n1548, n1551, n1552, n1555, n1556, n1559, n1560, n1563, n1564, n1584,
         n1588, n1592, n1593, n1594, n1596, n1597, n1598, n1599, n1600, n1602,
         n1608, n1610, n1611, n1613, n1614, n1616, n1618, n1620, n1622, n1624,
         n1626, n1628, n1629, n1630, n1631, n1632, n1634, n1636, n1639, n1640,
         n1641, n1642, n1644, n1645, n1646, n1647, n1648, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1668, n1671, n1672, n1674, n1677, n1678, n1682, n1686, n1688, n1693,
         n1694, n1696, n1698, n1712, n1716, n1719, n1720, n1721, n1722, n1724,
         n1725, n1726, n1727, n1728, n1730, n1736, n1738, n1739, n1741, n1742,
         n1744, n1746, n1748, n1750, n1751, n1752, n1754, n1756, n1757, n1758,
         n1759, n1760, n1762, n1764, n1767, n1768, n1769, n1770, n1772, n1773,
         n1774, n1775, n1776, n1780, n1781, n1785, n1796, n1800, n1802, n1805,
         n1806, n1810, n1814, n1815, n1816, n1821, n1822, n1823, n1824, n1826,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998;

  MUX2IX4 U14 ( .D0(n27), .D1(n43), .S(n3852), .Y(n11) );
  MUX2IX4 U22 ( .D0(n19), .D1(n35), .S(n3853), .Y(n3) );
  MUX2IX4 U30 ( .D0(n75), .D1(n107), .S(n3855), .Y(n43) );
  MUX2IX4 U51 ( .D0(n54), .D1(n86), .S(n3857), .Y(n22) );
  MUX2IX4 U53 ( .D0(n52), .D1(n84), .S(n3857), .Y(n20) );
  MUX2IX4 U83 ( .D0(n150), .D1(n214), .S(n3861), .Y(n86) );
  AO22X1 U515 ( .A(n3851), .B(A[254]), .C(n3952), .D(A[766]), .Y(n497) );
  AO22X1 U525 ( .A(n3974), .B(A[253]), .C(n3988), .D(A[765]), .Y(n503) );
  AO22X1 U534 ( .A(n3851), .B(A[508]), .C(n3988), .D(A[1020]), .Y(n510) );
  AO22X1 U540 ( .A(n516), .B(n3762), .C(n515), .D(n3911), .Y(n1826) );
  AO22X1 U544 ( .A(n3851), .B(A[507]), .C(n3956), .D(A[1019]), .Y(n516) );
  AO22X1 U555 ( .A(n3974), .B(A[250]), .C(n3988), .D(A[762]), .Y(n521) );
  AO22X1 U560 ( .A(n528), .B(n3793), .C(n527), .D(n3911), .Y(n1824) );
  AO22X1 U564 ( .A(n3975), .B(A[505]), .C(n3953), .D(A[1017]), .Y(n528) );
  AO22X1 U570 ( .A(n534), .B(n3762), .C(n533), .D(n3798), .Y(n1823) );
  AO22X1 U574 ( .A(n3971), .B(A[504]), .C(n3953), .D(A[1016]), .Y(n534) );
  AO22X1 U580 ( .A(n540), .B(n3687), .C(n539), .D(n3911), .Y(n1822) );
  AO22X1 U584 ( .A(n3974), .B(A[503]), .C(n3953), .D(A[1015]), .Y(n540) );
  AO22X1 U590 ( .A(n546), .B(n3900), .C(n545), .D(n3911), .Y(n1821) );
  AO22X1 U594 ( .A(n3972), .B(A[502]), .C(n3953), .D(A[1014]), .Y(n546) );
  AO22X1 U604 ( .A(n3981), .B(A[501]), .C(n3953), .D(A[1013]), .Y(n552) );
  AO22X1 U605 ( .A(n3981), .B(A[245]), .C(n3953), .D(A[757]), .Y(n551) );
  AO22X1 U614 ( .A(n3972), .B(A[500]), .C(n3954), .D(A[1012]), .Y(n558) );
  AO22X1 U615 ( .A(n3977), .B(A[244]), .C(n3953), .D(A[756]), .Y(n557) );
  AO22X1 U624 ( .A(n3981), .B(A[499]), .C(n3954), .D(A[1011]), .Y(n564) );
  AO22X1 U625 ( .A(n3981), .B(A[243]), .C(n3954), .D(A[755]), .Y(n563) );
  AO22X1 U640 ( .A(n576), .B(n3687), .C(n575), .D(n3914), .Y(n1816) );
  AO22X1 U644 ( .A(n3981), .B(A[497]), .C(n3954), .D(A[1009]), .Y(n576) );
  AO22X1 U650 ( .A(n582), .B(n3900), .C(n581), .D(n3914), .Y(n1815) );
  AO22X1 U654 ( .A(n3974), .B(A[496]), .C(n3957), .D(A[1008]), .Y(n582) );
  NOR2X1 U664 ( .A(n3947), .B(A[239]), .Y(n585) );
  NOR2X1 U672 ( .A(n3947), .B(A[238]), .Y(n589) );
  NOR2X1 U688 ( .A(n3946), .B(A[236]), .Y(n597) );
  NOR2X1 U696 ( .A(n3946), .B(A[235]), .Y(n601) );
  NOR2X1 U712 ( .A(n3946), .B(A[233]), .Y(n609) );
  NOR2X1 U728 ( .A(n3946), .B(A[231]), .Y(n617) );
  NOR2X1 U736 ( .A(n3946), .B(A[230]), .Y(n621) );
  NOR2X1 U744 ( .A(n3944), .B(A[229]), .Y(n625) );
  NOR2X1 U752 ( .A(n3944), .B(A[228]), .Y(n629) );
  NOR2X1 U760 ( .A(n3946), .B(A[227]), .Y(n633) );
  NOR2X1 U776 ( .A(n3944), .B(A[225]), .Y(n641) );
  NOR2X1 U784 ( .A(n3944), .B(A[224]), .Y(n645) );
  NOR2X1 U792 ( .A(n3944), .B(A[223]), .Y(n649) );
  NOR2X1 U800 ( .A(n3944), .B(A[222]), .Y(n653) );
  NOR2X1 U808 ( .A(n3945), .B(A[221]), .Y(n657) );
  NOR2X1 U816 ( .A(n3944), .B(A[220]), .Y(n661) );
  NOR2X1 U824 ( .A(n3945), .B(A[219]), .Y(n665) );
  NOR2X1 U832 ( .A(n3944), .B(A[218]), .Y(n669) );
  NOR2X1 U840 ( .A(n3944), .B(A[217]), .Y(n673) );
  NOR2X1 U848 ( .A(n3944), .B(A[216]), .Y(n677) );
  NOR2X1 U1031 ( .A(n3945), .B(A[447]), .Y(n762) );
  NOR2X1 U1039 ( .A(n3945), .B(A[446]), .Y(n766) );
  NOR2X1 U1047 ( .A(n3945), .B(A[445]), .Y(n770) );
  NOR2X1 U1063 ( .A(n3946), .B(A[443]), .Y(n778) );
  NOR2X1 U1071 ( .A(n3945), .B(A[442]), .Y(n782) );
  NOR2X1 U1079 ( .A(n3945), .B(A[441]), .Y(n786) );
  NOR2X1 U1087 ( .A(n3946), .B(A[440]), .Y(n790) );
  AO22X1 U1092 ( .A(n796), .B(n3892), .C(n795), .D(n3915), .Y(n1758) );
  AO22X1 U1096 ( .A(n3982), .B(A[439]), .C(n3952), .D(A[951]), .Y(n796) );
  AO22X1 U1097 ( .A(n3982), .B(A[183]), .C(n3961), .D(A[695]), .Y(n795) );
  AO22X1 U1102 ( .A(n802), .B(n3899), .C(n801), .D(n3914), .Y(n1757) );
  AO22X1 U1106 ( .A(n3981), .B(A[438]), .C(n3961), .D(A[950]), .Y(n802) );
  AO22X1 U1107 ( .A(n3981), .B(A[182]), .C(n3961), .D(A[694]), .Y(n801) );
  AO22X1 U1116 ( .A(n3982), .B(A[437]), .C(n3961), .D(A[949]), .Y(n808) );
  AO22X1 U1117 ( .A(n3982), .B(A[181]), .C(n3990), .D(A[693]), .Y(n807) );
  AO22X1 U1126 ( .A(n3974), .B(A[436]), .C(n3835), .D(A[948]), .Y(n814) );
  AO22X1 U1137 ( .A(n3983), .B(A[179]), .C(n3958), .D(A[691]), .Y(n819) );
  AO22X1 U1147 ( .A(n3973), .B(A[178]), .C(n3958), .D(A[690]), .Y(n825) );
  AO22X1 U1152 ( .A(n832), .B(n3892), .C(n831), .D(n3910), .Y(n1752) );
  AO22X1 U1156 ( .A(n3983), .B(A[433]), .C(n3958), .D(A[945]), .Y(n832) );
  AO22X1 U1157 ( .A(n3983), .B(A[177]), .C(n3958), .D(A[689]), .Y(n831) );
  AO22X1 U1162 ( .A(n838), .B(n3899), .C(n837), .D(n3915), .Y(n1751) );
  AO22X1 U1166 ( .A(n3973), .B(A[432]), .C(n3958), .D(A[944]), .Y(n838) );
  AO22X1 U1167 ( .A(n3973), .B(A[176]), .C(n3958), .D(A[688]), .Y(n837) );
  AO22X1 U1172 ( .A(n844), .B(n3890), .C(n843), .D(n3910), .Y(n1750) );
  AO22X1 U1176 ( .A(n3983), .B(A[431]), .C(n3958), .D(A[943]), .Y(n844) );
  AO22X1 U1177 ( .A(n3983), .B(A[175]), .C(n3958), .D(A[687]), .Y(n843) );
  AO22X1 U1192 ( .A(n856), .B(n3898), .C(n855), .D(n3910), .Y(n1748) );
  AO22X1 U1196 ( .A(n3965), .B(A[429]), .C(n3957), .D(A[941]), .Y(n856) );
  AO22X1 U1206 ( .A(n3974), .B(A[428]), .C(n3957), .D(A[940]), .Y(n862) );
  AO22X1 U1207 ( .A(n3974), .B(A[172]), .C(n3957), .D(A[684]), .Y(n861) );
  AO22X1 U1212 ( .A(n868), .B(n3899), .C(n867), .D(n3909), .Y(n1746) );
  AO22X1 U1216 ( .A(n3984), .B(A[427]), .C(n3957), .D(A[939]), .Y(n868) );
  AO22X1 U1217 ( .A(n3984), .B(A[171]), .C(n3957), .D(A[683]), .Y(n867) );
  AO22X1 U1232 ( .A(n880), .B(n3898), .C(n879), .D(n3909), .Y(n1744) );
  AO22X1 U1236 ( .A(n3984), .B(A[425]), .C(n3960), .D(A[937]), .Y(n880) );
  AO22X1 U1237 ( .A(n3984), .B(A[169]), .C(n3956), .D(A[681]), .Y(n879) );
  AO22X1 U1246 ( .A(n3974), .B(A[424]), .C(n3988), .D(A[936]), .Y(n886) );
  AO22X1 U1247 ( .A(n3974), .B(A[168]), .C(n3988), .D(A[680]), .Y(n885) );
  AO22X1 U1252 ( .A(n892), .B(n3884), .C(n891), .D(n3909), .Y(n1742) );
  AO22X1 U1256 ( .A(n3984), .B(A[423]), .C(n3960), .D(A[935]), .Y(n892) );
  AO22X1 U1257 ( .A(n3985), .B(A[167]), .C(n3960), .D(A[679]), .Y(n891) );
  AO22X1 U1262 ( .A(n898), .B(n3899), .C(n897), .D(n3916), .Y(n1741) );
  AO22X1 U1266 ( .A(n3975), .B(A[422]), .C(n3956), .D(A[934]), .Y(n898) );
  AO22X1 U1267 ( .A(n3975), .B(A[166]), .C(n3960), .D(A[678]), .Y(n897) );
  AO22X1 U1277 ( .A(n3985), .B(A[165]), .C(n3955), .D(A[677]), .Y(n903) );
  AO22X1 U1286 ( .A(n3975), .B(A[420]), .C(n3955), .D(A[932]), .Y(n910) );
  AO22X1 U1292 ( .A(n916), .B(n3898), .C(n915), .D(n3909), .Y(n1738) );
  AO22X1 U1296 ( .A(n3985), .B(A[419]), .C(n3955), .D(A[931]), .Y(n916) );
  AO22X1 U1297 ( .A(n3985), .B(A[163]), .C(n3955), .D(A[675]), .Y(n915) );
  AO22X1 U1312 ( .A(n928), .B(n3899), .C(n927), .D(n3909), .Y(n1736) );
  AO22X1 U1316 ( .A(n3985), .B(A[417]), .C(n3955), .D(A[929]), .Y(n928) );
  AO22X1 U1317 ( .A(n3964), .B(A[161]), .C(n3955), .D(A[673]), .Y(n927) );
  AO22X1 U1326 ( .A(n3976), .B(A[416]), .C(n3955), .D(A[928]), .Y(n934) );
  AO22X1 U1327 ( .A(n3976), .B(A[160]), .C(n3954), .D(A[672]), .Y(n933) );
  NOR21X1 U1360 ( .B(n3934), .A(A[668]), .Y(n949) );
  AO22X1 U1474 ( .A(n3976), .B(A[398]), .C(n3963), .D(A[910]), .Y(n1010) );
  AO22X1 U1475 ( .A(n3976), .B(A[142]), .C(n3963), .D(A[654]), .Y(n1009) );
  AO22X1 U1480 ( .A(n1016), .B(n3898), .C(n1015), .D(n3912), .Y(n1716) );
  AO22X1 U1484 ( .A(n3973), .B(A[397]), .C(n3963), .D(A[909]), .Y(n1016) );
  AO22X1 U1485 ( .A(n3968), .B(A[141]), .C(n3962), .D(A[653]), .Y(n1015) );
  AO22X1 U1494 ( .A(n3976), .B(A[396]), .C(n3962), .D(A[908]), .Y(n1022) );
  AO22X1 U1495 ( .A(n3977), .B(A[140]), .C(n3962), .D(A[652]), .Y(n1021) );
  AO22X1 U1504 ( .A(n3985), .B(A[395]), .C(n3962), .D(A[907]), .Y(n1028) );
  AO22X1 U1505 ( .A(n3984), .B(A[139]), .C(n3962), .D(A[651]), .Y(n1027) );
  AO22X1 U1514 ( .A(n3977), .B(A[394]), .C(n3962), .D(A[906]), .Y(n1034) );
  AO22X1 U1520 ( .A(n1040), .B(n3897), .C(n1039), .D(n3914), .Y(n1712) );
  AO22X1 U1524 ( .A(n3985), .B(A[393]), .C(n3962), .D(A[905]), .Y(n1040) );
  AO22X1 U1525 ( .A(n3977), .B(A[137]), .C(n3962), .D(A[649]), .Y(n1039) );
  AO22X1 U1534 ( .A(n3977), .B(A[392]), .C(n3962), .D(A[904]), .Y(n1046) );
  AO22X1 U1535 ( .A(n3977), .B(A[136]), .C(n3961), .D(A[648]), .Y(n1045) );
  NOR2X1 U1543 ( .A(n3952), .B(A[391]), .Y(n1050) );
  NOR2X1 U1551 ( .A(n3952), .B(A[390]), .Y(n1054) );
  NOR2X1 U1559 ( .A(n3951), .B(A[389]), .Y(n1058) );
  NOR2X1 U1567 ( .A(n3951), .B(A[388]), .Y(n1062) );
  NOR2X1 U1575 ( .A(n3951), .B(A[387]), .Y(n1066) );
  NOR2X1 U1583 ( .A(n3951), .B(A[386]), .Y(n1070) );
  NOR2X1 U1592 ( .A(n3950), .B(A[129]), .Y(n1073) );
  NOR2X1 U1599 ( .A(n3950), .B(A[384]), .Y(n1078) );
  NOR2X1 U1607 ( .A(n3950), .B(A[383]), .Y(n1082) );
  NOR2X1 U1615 ( .A(n3950), .B(A[382]), .Y(n1086) );
  NOR2X1 U1631 ( .A(n3950), .B(A[380]), .Y(n1094) );
  NOR2X1 U1639 ( .A(n3950), .B(A[379]), .Y(n1098) );
  NOR2X1 U1647 ( .A(n3949), .B(A[378]), .Y(n1102) );
  NOR2X1 U1655 ( .A(n3947), .B(A[377]), .Y(n1106) );
  NOR2X1 U1663 ( .A(n3949), .B(A[376]), .Y(n1110) );
  NOR2X1 U1671 ( .A(n3949), .B(A[375]), .Y(n1114) );
  NOR2X1 U1679 ( .A(n3949), .B(A[374]), .Y(n1118) );
  NOR2X1 U1687 ( .A(n3949), .B(A[373]), .Y(n1122) );
  NOR2X1 U1703 ( .A(n3948), .B(A[371]), .Y(n1130) );
  NOR2X1 U1711 ( .A(n3948), .B(A[370]), .Y(n1134) );
  NOR2X1 U1719 ( .A(n3948), .B(A[369]), .Y(n1138) );
  NOR2X1 U1727 ( .A(n3948), .B(A[368]), .Y(n1142) );
  NOR2X1 U1735 ( .A(n3948), .B(A[367]), .Y(n1146) );
  NOR2X1 U1751 ( .A(n3948), .B(A[365]), .Y(n1154) );
  NOR2X1 U1767 ( .A(n3947), .B(A[363]), .Y(n1162) );
  NOR2X1 U1775 ( .A(n3947), .B(A[362]), .Y(n1166) );
  NOR2X1 U1783 ( .A(n3947), .B(A[361]), .Y(n1170) );
  NOR2X1 U1799 ( .A(n3947), .B(A[359]), .Y(n1178) );
  NOR2X1 U1807 ( .A(n3951), .B(A[358]), .Y(n1182) );
  NOR2X1 U1815 ( .A(n3947), .B(A[357]), .Y(n1186) );
  NOR2X1 U1823 ( .A(n3947), .B(A[356]), .Y(n1190) );
  NOR2X1 U1831 ( .A(n3948), .B(A[355]), .Y(n1194) );
  NOR2X1 U1839 ( .A(n3948), .B(A[354]), .Y(n1198) );
  NOR2X1 U1847 ( .A(n3948), .B(A[353]), .Y(n1202) );
  NOR2X1 U1855 ( .A(n3949), .B(A[352]), .Y(n1206) );
  NOR2X1 U1863 ( .A(n3949), .B(A[351]), .Y(n1210) );
  NOR2X1 U1871 ( .A(n3949), .B(A[350]), .Y(n1214) );
  NOR2X1 U1879 ( .A(n3949), .B(A[349]), .Y(n1218) );
  NOR2X1 U1887 ( .A(n3950), .B(A[348]), .Y(n1222) );
  NOR2X1 U1895 ( .A(n3950), .B(A[347]), .Y(n1226) );
  NOR2X1 U1911 ( .A(n3952), .B(A[345]), .Y(n1234) );
  NOR2X1 U1919 ( .A(n3952), .B(A[344]), .Y(n1238) );
  NAND21X1 U1924 ( .B(n3793), .A(n1241), .Y(n1662) );
  NAND21X1 U1931 ( .B(n3793), .A(n1244), .Y(n1661) );
  NAND21X1 U1938 ( .B(n3896), .A(n1247), .Y(n1660) );
  NAND21X1 U1945 ( .B(n3896), .A(n1250), .Y(n1659) );
  NOR21X1 U1948 ( .B(n3939), .A(A[596]), .Y(n1250) );
  NAND21X1 U1952 ( .B(n3896), .A(n1253), .Y(n1658) );
  NAND21X1 U1966 ( .B(n3896), .A(n1259), .Y(n1656) );
  NAND21X1 U1973 ( .B(n3896), .A(n1262), .Y(n1655) );
  NAND21X1 U1980 ( .B(n3896), .A(n3933), .Y(n1654) );
  NAND21X1 U1986 ( .B(n3896), .A(n3933), .Y(n1653) );
  NAND21X1 U1992 ( .B(n3896), .A(n1269), .Y(n1652) );
  NOR21X1 U2002 ( .B(n3938), .A(A[588]), .Y(n1272) );
  NAND21X1 U2006 ( .B(n3897), .A(n1275), .Y(n1650) );
  NAND21X1 U2020 ( .B(n3897), .A(n1281), .Y(n1648) );
  NAND21X1 U2027 ( .B(n3897), .A(n1284), .Y(n1647) );
  NOR21X1 U2134 ( .B(n3940), .A(A[570]), .Y(n1331) );
  AO22X1 U2218 ( .A(n1378), .B(n3762), .C(n1377), .D(n3911), .Y(n1622) );
  AO22X1 U2222 ( .A(n3977), .B(A[303]), .C(n3961), .D(A[815]), .Y(n1378) );
  AO22X1 U2223 ( .A(n3978), .B(A[47]), .C(n3961), .D(A[559]), .Y(n1377) );
  AO22X1 U2252 ( .A(n3969), .B(A[300]), .C(n3960), .D(A[812]), .Y(n1396) );
  AO22X1 U2258 ( .A(n1402), .B(n3793), .C(n1401), .D(n3914), .Y(n1618) );
  AO22X1 U2262 ( .A(n3978), .B(A[299]), .C(n3956), .D(A[811]), .Y(n1402) );
  AO22X1 U2263 ( .A(n3978), .B(A[43]), .C(n3956), .D(A[555]), .Y(n1401) );
  AO22X1 U2273 ( .A(n3969), .B(A[42]), .C(n3988), .D(A[554]), .Y(n1407) );
  AO22X1 U2278 ( .A(n1414), .B(n3687), .C(n1413), .D(n3915), .Y(n1616) );
  AO22X1 U2282 ( .A(n3978), .B(A[297]), .C(n3988), .D(A[809]), .Y(n1414) );
  AO22X1 U2283 ( .A(n3979), .B(A[41]), .C(n3960), .D(A[553]), .Y(n1413) );
  AO22X1 U2292 ( .A(n3969), .B(A[296]), .C(n3988), .D(A[808]), .Y(n1420) );
  AO22X1 U2293 ( .A(n3965), .B(A[40]), .C(n3959), .D(A[552]), .Y(n1419) );
  AO22X1 U2298 ( .A(n1426), .B(n3900), .C(n1425), .D(n3915), .Y(n1614) );
  AO22X1 U2302 ( .A(n3979), .B(A[295]), .C(n3959), .D(A[807]), .Y(n1426) );
  AO22X1 U2303 ( .A(n3979), .B(A[39]), .C(n3959), .D(A[551]), .Y(n1425) );
  AO22X1 U2308 ( .A(n1432), .B(n3900), .C(n1431), .D(n3917), .Y(n1613) );
  AO22X1 U2312 ( .A(n3970), .B(A[294]), .C(n3959), .D(A[806]), .Y(n1432) );
  AO22X1 U2322 ( .A(n3979), .B(A[293]), .C(n3959), .D(A[805]), .Y(n1438) );
  AO22X1 U2323 ( .A(n3979), .B(A[37]), .C(n3959), .D(A[549]), .Y(n1437) );
  AO22X1 U2338 ( .A(n1450), .B(n3901), .C(n1449), .D(n3914), .Y(n1610) );
  AO22X1 U2358 ( .A(n1462), .B(n3900), .C(n1461), .D(n3914), .Y(n1608) );
  AO22X1 U2362 ( .A(n3980), .B(A[289]), .C(n3963), .D(A[801]), .Y(n1462) );
  AO22X1 U2363 ( .A(n3980), .B(A[33]), .C(n3942), .D(A[545]), .Y(n1461) );
  AO22X1 U2372 ( .A(n3851), .B(A[288]), .C(n3940), .D(A[800]), .Y(n1468) );
  AO22X1 U2373 ( .A(n3851), .B(A[32]), .C(n3958), .D(A[544]), .Y(n1467) );
  INVX1 U2611 ( .A(n3968), .Y(n3927) );
  INVX2 U2612 ( .A(n3991), .Y(n3968) );
  BUFX6 U2613 ( .A(n3931), .Y(n3648) );
  MUX2X1 U2614 ( .D0(n669), .D1(n670), .S(n3890), .Y(n3805) );
  MUX2XL U2615 ( .D0(n1102), .D1(n1101), .S(n3917), .Y(n3839) );
  MUX2X1 U2616 ( .D0(n1133), .D1(n1134), .S(n3882), .Y(n3803) );
  EORXL U2617 ( .A(n873), .B(n3916), .C(n3814), .D(n3912), .Y(n3844) );
  MUX2X1 U2618 ( .D0(n725), .D1(n726), .S(n3889), .Y(n3840) );
  MUX2IX1 U2619 ( .D0(n3843), .D1(n3845), .S(n3878), .Y(n123) );
  NOR21XL U2620 ( .B(n3935), .A(A[661]), .Y(n977) );
  NOR21XL U2621 ( .B(n3942), .A(A[537]), .Y(n1495) );
  NOR21XL U2622 ( .B(n3942), .A(A[604]), .Y(n1221) );
  NOR21XL U2623 ( .B(n3941), .A(A[540]), .Y(n1483) );
  MUX2IXL U2624 ( .D0(A[476]), .D1(A[988]), .S(n3989), .Y(n662) );
  MUX2IX1 U2625 ( .D0(n3671), .D1(n3651), .S(n3874), .Y(n165) );
  MUX2IX1 U2626 ( .D0(n3678), .D1(n3749), .S(n3877), .Y(n133) );
  INVX2 U2627 ( .A(n3880), .Y(n3867) );
  MUX2IX1 U2628 ( .D0(n148), .D1(n212), .S(n3861), .Y(n84) );
  MUX2IX1 U2629 ( .D0(n68), .D1(n100), .S(n3856), .Y(n36) );
  MUX2X1 U2630 ( .D0(n3688), .D1(n3689), .S(n3857), .Y(n28) );
  MUX2IX1 U2631 ( .D0(n70), .D1(n102), .S(n3856), .Y(n38) );
  MUX2IX1 U2632 ( .D0(n134), .D1(n198), .S(n3863), .Y(n70) );
  MUX2IX1 U2633 ( .D0(n18), .D1(n34), .S(n3853), .Y(n2) );
  EORX1 U2634 ( .A(n3955), .B(A[930]), .C(n3955), .D(n3821), .Y(n3849) );
  NOR21XL U2635 ( .B(n3943), .A(A[610]), .Y(n1197) );
  NOR21XL U2636 ( .B(n3933), .A(A[961]), .Y(n755) );
  NOR21XL U2637 ( .B(n3930), .A(A[660]), .Y(n981) );
  NOR21XL U2638 ( .B(n3937), .A(A[834]), .Y(n1302) );
  NOR21XL U2639 ( .B(n3937), .A(A[836]), .Y(n1296) );
  NOR21XL U2640 ( .B(n3686), .A(A[964]), .Y(n746) );
  MUX2X1 U2641 ( .D0(n1611), .D1(n1739), .S(n3876), .Y(n149) );
  ENOX1 U2642 ( .A(n3763), .B(n3762), .C(n910), .D(n3897), .Y(n1739) );
  MUX2IX1 U2643 ( .D0(n3747), .D1(n3669), .S(n3869), .Y(n213) );
  MUX2X1 U2644 ( .D0(n1189), .D1(n1190), .S(n3885), .Y(n3747) );
  NOR21XL U2645 ( .B(n3993), .A(A[612]), .Y(n1189) );
  NOR21XL U2646 ( .B(n3943), .A(A[524]), .Y(n1547) );
  MUX2IX1 U2647 ( .D0(n3748), .D1(n3654), .S(n3868), .Y(n221) );
  NOR2X1 U2648 ( .A(n3948), .B(A[364]), .Y(n1158) );
  MUX2IX1 U2649 ( .D0(n3673), .D1(n3652), .S(n3875), .Y(n157) );
  MUX2IX1 U2650 ( .D0(n309), .D1(n3656), .S(n3872), .Y(n189) );
  NOR21XL U2651 ( .B(n3935), .A(A[972]), .Y(n718) );
  NOR21XL U2652 ( .B(n3933), .A(A[960]), .Y(n758) );
  NOR21XL U2653 ( .B(n3937), .A(A[616]), .Y(n1173) );
  MUX2X1 U2654 ( .D0(n1613), .D1(n1741), .S(n3875), .Y(n151) );
  MUX2IX1 U2655 ( .D0(n139), .D1(n203), .S(n3862), .Y(n75) );
  MUX2IX1 U2656 ( .D0(n3838), .D1(n3837), .S(n3877), .Y(n139) );
  MUX2IX1 U2657 ( .D0(n171), .D1(n235), .S(n3859), .Y(n107) );
  MUX2IX1 U2658 ( .D0(n67), .D1(n99), .S(n3856), .Y(n35) );
  MUX2IX1 U2659 ( .D0(n59), .D1(n91), .S(n3857), .Y(n27) );
  MUX2IX1 U2660 ( .D0(n123), .D1(n187), .S(n3864), .Y(n59) );
  NOR21XL U2661 ( .B(n3935), .A(A[973]), .Y(n714) );
  NOR21XL U2662 ( .B(n3935), .A(A[717]), .Y(n713) );
  EORX1 U2663 ( .A(n503), .B(n3798), .C(n3795), .D(n3909), .Y(n3794) );
  OR2X1 U2664 ( .A(n3950), .B(A[381]), .Y(n3810) );
  MUX2X1 U2665 ( .D0(n1628), .D1(n1756), .S(n3874), .Y(n166) );
  NOR21XL U2666 ( .B(n3940), .A(A[565]), .Y(n1351) );
  MUX2X1 U2667 ( .D0(n1596), .D1(n1724), .S(n3877), .Y(n134) );
  MUX2IX1 U2668 ( .D0(n3792), .D1(n3806), .S(n3876), .Y(n150) );
  MUX2IX1 U2669 ( .D0(n3705), .D1(n3657), .S(n3869), .Y(n214) );
  MUX2IX1 U2670 ( .D0(n66), .D1(n98), .S(n3856), .Y(n34) );
  MUX2IX1 U2671 ( .D0(n50), .D1(n82), .S(n3856), .Y(n18) );
  MUX2BXL U2672 ( .D0(n3711), .D1(n178), .S(n3865), .Y(n50) );
  MUX2IX1 U2673 ( .D0(n146), .D1(n210), .S(n3862), .Y(n82) );
  MUX2IX1 U2674 ( .D0(n74), .D1(n106), .S(n3855), .Y(n42) );
  MUX2IX1 U2675 ( .D0(n138), .D1(n202), .S(n3862), .Y(n74) );
  MUX2X1 U2676 ( .D0(n1600), .D1(n1728), .S(n3877), .Y(n138) );
  MUX2BXL U2677 ( .D0(n3702), .D1(n90), .S(n3857), .Y(n26) );
  MUX2IX1 U2678 ( .D0(n173), .D1(n237), .S(n3859), .Y(n109) );
  MUX2IX1 U2679 ( .D0(n3751), .D1(n3660), .S(n3867), .Y(n237) );
  MUX2IX1 U2680 ( .D0(n3750), .D1(n3667), .S(n3873), .Y(n173) );
  MUX2IX1 U2681 ( .D0(n141), .D1(n205), .S(n3862), .Y(n77) );
  MUX2IX1 U2682 ( .D0(n3655), .D1(n3752), .S(n3870), .Y(n205) );
  MUX2IX1 U2683 ( .D0(n69), .D1(n101), .S(n3856), .Y(n37) );
  MUX2IX1 U2684 ( .D0(n133), .D1(n197), .S(n3863), .Y(n69) );
  MUX2IX1 U2685 ( .D0(n53), .D1(n85), .S(n3857), .Y(n21) );
  MUX2IX1 U2686 ( .D0(n117), .D1(n181), .S(n3864), .Y(n53) );
  MUX2IX1 U2687 ( .D0(n213), .D1(n149), .S(n3866), .Y(n85) );
  MUX2IX1 U2688 ( .D0(n3649), .D1(n3679), .S(n3872), .Y(n181) );
  MUX2IX1 U2689 ( .D0(n61), .D1(n93), .S(n3856), .Y(n29) );
  MUX2IX1 U2690 ( .D0(n125), .D1(n189), .S(n3864), .Y(n61) );
  MUX2IX1 U2691 ( .D0(n157), .D1(n221), .S(n3860), .Y(n93) );
  MUX2IX1 U2692 ( .D0(n3658), .D1(n3833), .S(n3878), .Y(n125) );
  MUX2AXL U2693 ( .D0(n3692), .D1(n1719), .S(n3878), .Y(n129) );
  MUX2IX1 U2694 ( .D0(n3653), .D1(n3681), .S(n3876), .Y(n145) );
  MUX2IX1 U2695 ( .D0(n3650), .D1(n3680), .S(n3875), .Y(n153) );
  MUX2IX1 U2696 ( .D0(n3707), .D1(n3659), .S(n3878), .Y(n121) );
  MUX2AXL U2697 ( .D0(n3706), .D1(n1823), .S(n3867), .Y(n233) );
  INVX1 U2698 ( .A(n3880), .Y(n3877) );
  INVX1 U2699 ( .A(n3866), .Y(n3859) );
  MUX2IX1 U2700 ( .D0(n5), .D1(n13), .S(SH[3]), .Y(B[4]) );
  MUX2IX1 U2701 ( .D0(n29), .D1(n45), .S(n3852), .Y(n13) );
  MUX2IX1 U2702 ( .D0(n21), .D1(n37), .S(n3853), .Y(n5) );
  MUX2IX1 U2703 ( .D0(n77), .D1(n109), .S(n3855), .Y(n45) );
  MUX2IX1 U2704 ( .D0(n28), .D1(n44), .S(n3852), .Y(n12) );
  MUX2IX1 U2705 ( .D0(n20), .D1(n36), .S(n3853), .Y(n4) );
  MUX2IX1 U2706 ( .D0(n22), .D1(n38), .S(n3853), .Y(n6) );
  MUX2IX1 U2707 ( .D0(n30), .D1(n46), .S(n3852), .Y(n14) );
  MUX2IX1 U2708 ( .D0(n4), .D1(n12), .S(SH[3]), .Y(B[3]) );
  INVX1 U2709 ( .A(n3992), .Y(n3969) );
  INVX1 U2710 ( .A(SH[8]), .Y(n3922) );
  INVXL U2711 ( .A(n3996), .Y(n3994) );
  INVX1 U2712 ( .A(n3994), .Y(n3970) );
  INVX1 U2713 ( .A(SH[9]), .Y(n3998) );
  INVXL U2714 ( .A(n3997), .Y(n3990) );
  INVX1 U2715 ( .A(n3924), .Y(n3918) );
  INVXL U2716 ( .A(n3998), .Y(n3986) );
  INVX1 U2717 ( .A(SH[9]), .Y(n3996) );
  INVX1 U2718 ( .A(n3997), .Y(n3993) );
  INVX1 U2719 ( .A(n3922), .Y(n3812) );
  INVX1 U2720 ( .A(n3916), .Y(n3897) );
  INVX1 U2721 ( .A(n3916), .Y(n3896) );
  AND2X1 U2722 ( .A(n1296), .B(n3894), .Y(n3649) );
  AOI22X1 U2723 ( .A(n1420), .B(n3901), .C(n1419), .D(n3917), .Y(n3650) );
  AOI22X1 U2724 ( .A(n814), .B(n3890), .C(n813), .D(n3914), .Y(n3651) );
  AOI22X1 U2725 ( .A(n862), .B(n3898), .C(n861), .D(n3915), .Y(n3652) );
  AOI22X1 U2726 ( .A(n1468), .B(n3687), .C(n1467), .D(n3911), .Y(n3653) );
  MUX2X1 U2727 ( .D0(n597), .D1(n598), .S(n3891), .Y(n3654) );
  MUX2X1 U2728 ( .D0(n1221), .D1(n1222), .S(n3887), .Y(n3655) );
  MUX2X1 U2729 ( .D0(n717), .D1(n718), .S(n3889), .Y(n3656) );
  MUX2X1 U2730 ( .D0(n625), .D1(n626), .S(n3892), .Y(n3657) );
  MUX2X1 U2731 ( .D0(n1547), .D1(n1548), .S(n3893), .Y(n3658) );
  AOI22X1 U2732 ( .A(n1046), .B(n3899), .C(n1045), .D(n3913), .Y(n3659) );
  AOI22X1 U2733 ( .A(n510), .B(n3687), .C(n509), .D(n3798), .Y(n3660) );
  MUX2X1 U2734 ( .D0(n637), .D1(n638), .S(n3891), .Y(n3661) );
  MUX2X1 U2735 ( .D0(n1209), .D1(n1210), .S(n3887), .Y(n3662) );
  MUX2X1 U2736 ( .D0(n1213), .D1(n1214), .S(n3887), .Y(n3663) );
  MUX2X1 U2737 ( .D0(n765), .D1(n766), .S(n3800), .Y(n3664) );
  MUX2X1 U2738 ( .D0(n761), .D1(n762), .S(n3801), .Y(n3665) );
  MUX2X1 U2739 ( .D0(n1149), .D1(n3964), .S(n3882), .Y(n3666) );
  MUX2X1 U2740 ( .D0(n773), .D1(n774), .S(n3800), .Y(n3667) );
  MUX2X1 U2741 ( .D0(n3788), .D1(n1230), .S(n3888), .Y(n3668) );
  MUX2X1 U2742 ( .D0(n629), .D1(n630), .S(n3891), .Y(n3669) );
  MUX2X1 U2743 ( .D0(n949), .D1(n950), .S(n3887), .Y(n3670) );
  MUX2X1 U2744 ( .D0(n1355), .D1(n1356), .S(n3801), .Y(n3671) );
  MUX2X1 U2745 ( .D0(n781), .D1(n782), .S(n3801), .Y(n3672) );
  AOI22X1 U2746 ( .A(n1396), .B(n3900), .C(n1395), .D(n3913), .Y(n3673) );
  AND2X1 U2747 ( .A(n681), .B(n3895), .Y(n3674) );
  AOI22X1 U2748 ( .A(n564), .B(n3901), .C(n563), .D(n3909), .Y(n3675) );
  AOI22X1 U2749 ( .A(n1010), .B(n3897), .C(n1009), .D(n3912), .Y(n3676) );
  AOI22X1 U2750 ( .A(n1028), .B(n3897), .C(n1027), .D(n3911), .Y(n3677) );
  MUX2X1 U2751 ( .D0(n1515), .D1(n1516), .S(n3893), .Y(n3678) );
  AND2X1 U2752 ( .A(n746), .B(n3895), .Y(n3679) );
  AOI22X1 U2753 ( .A(n886), .B(n3899), .C(n885), .D(n3916), .Y(n3680) );
  AOI22X1 U2754 ( .A(n934), .B(n3898), .C(n933), .D(n3917), .Y(n3681) );
  MUX2X1 U2755 ( .D0(n1479), .D1(n1480), .S(n3890), .Y(n3682) );
  AND2X1 U2756 ( .A(n687), .B(n3895), .Y(n3683) );
  AND2X1 U2757 ( .A(n690), .B(n3895), .Y(n3684) );
  MUX2IX1 U2758 ( .D0(A[914]), .D1(A[402]), .S(n3851), .Y(n3685) );
  INVX1 U2759 ( .A(n3967), .Y(n3686) );
  NOR21XL U2760 ( .B(n3686), .A(A[620]), .Y(n1157) );
  AOI22BXL U2761 ( .B(n3686), .A(A[162]), .D(n3972), .C(A[674]), .Y(n3850) );
  NOR21XL U2762 ( .B(n3990), .A(A[628]), .Y(n1125) );
  NOR21XL U2763 ( .B(n3990), .A(A[622]), .Y(n1149) );
  NOR21XL U2764 ( .B(n3835), .A(A[621]), .Y(n1153) );
  INVX1 U2765 ( .A(n3987), .Y(n3967) );
  INVX1 U2766 ( .A(n3982), .Y(n3988) );
  INVX1 U2767 ( .A(n3902), .Y(n3687) );
  INVX1 U2768 ( .A(n3900), .Y(n3917) );
  INVX1 U2769 ( .A(n3994), .Y(n3965) );
  MUX2X1 U2770 ( .D0(n126), .D1(n190), .S(n3864), .Y(n3691) );
  INVX1 U2771 ( .A(n3966), .Y(n3955) );
  INVX1 U2772 ( .A(n3880), .Y(n3878) );
  INVX1 U2773 ( .A(n3989), .Y(n3976) );
  MUX2IX1 U2774 ( .D0(n165), .D1(n229), .S(n3860), .Y(n101) );
  MUX2X1 U2775 ( .D0(n3690), .D1(n3691), .S(n3858), .Y(n30) );
  MUX2X1 U2776 ( .D0(n1688), .D1(n1816), .S(n3868), .Y(n226) );
  MUX2IX1 U2777 ( .D0(A[412]), .D1(A[924]), .S(n3926), .Y(n950) );
  AOI22X1 U2778 ( .A(n3970), .B(A[292]), .C(n3959), .D(A[804]), .Y(n3760) );
  MUX2XL U2779 ( .D0(n945), .D1(n946), .S(n3887), .Y(n3717) );
  MUX2XL U2780 ( .D0(n124), .D1(n188), .S(n3864), .Y(n3688) );
  MUX2X1 U2781 ( .D0(n156), .D1(n220), .S(n3861), .Y(n3689) );
  INVX1 U2782 ( .A(n3904), .Y(n3893) );
  INVX1 U2783 ( .A(n3966), .Y(n3948) );
  INVXL U2784 ( .A(n3998), .Y(n3959) );
  INVXL U2785 ( .A(n3902), .Y(n3901) );
  INVX1 U2786 ( .A(n3998), .Y(n3953) );
  INVX1 U2787 ( .A(n3970), .Y(n3952) );
  INVXL U2788 ( .A(n3866), .Y(n3863) );
  INVX1 U2789 ( .A(n3866), .Y(n3862) );
  INVX1 U2790 ( .A(n3964), .Y(n3961) );
  INVX1 U2791 ( .A(n3964), .Y(n3963) );
  MUX2IX1 U2792 ( .D0(n3784), .D1(n3791), .S(n3868), .Y(n229) );
  MUX2XL U2793 ( .D0(n1539), .D1(n1540), .S(n3893), .Y(n3703) );
  MUX2IX1 U2794 ( .D0(n142), .D1(n206), .S(n3862), .Y(n78) );
  MUX2XL U2795 ( .D0(n122), .D1(n186), .S(n3864), .Y(n3702) );
  MUX2XL U2796 ( .D0(n1531), .D1(n1532), .S(n3893), .Y(n3692) );
  MUX2IXL U2797 ( .D0(n1519), .D1(n1520), .S(n3893), .Y(n1594) );
  MUX2IXL U2798 ( .D0(A[275]), .D1(A[787]), .S(n3932), .Y(n1520) );
  MUX2IX1 U2799 ( .D0(A[413]), .D1(A[925]), .S(n3927), .Y(n946) );
  AO22XL U2800 ( .A(n3970), .B(A[38]), .C(n3959), .D(A[550]), .Y(n1431) );
  OAI22AX1 U2801 ( .D(n3716), .C(n3919), .A(n3847), .B(n3917), .Y(n1620) );
  INVX1 U2802 ( .A(n3902), .Y(n3900) );
  INVX1 U2803 ( .A(n3858), .Y(n3856) );
  INVXL U2804 ( .A(n3866), .Y(n3864) );
  INVX1 U2805 ( .A(n3858), .Y(n3857) );
  MUX2IX1 U2806 ( .D0(n3756), .D1(n3670), .S(n3876), .Y(n141) );
  MUX2IX1 U2807 ( .D0(n163), .D1(n227), .S(n3860), .Y(n99) );
  MUX2X1 U2808 ( .D0(n1636), .D1(n1764), .S(n3873), .Y(n174) );
  MUX2X1 U2809 ( .D0(n1185), .D1(n1186), .S(n3885), .Y(n3705) );
  MUX2X1 U2810 ( .D0(n153), .D1(n217), .S(n3861), .Y(n3699) );
  MUX2IX1 U2811 ( .D0(n3825), .D1(n3840), .S(n3872), .Y(n187) );
  MUX2IX1 U2812 ( .D0(n118), .D1(n182), .S(n3864), .Y(n54) );
  MUX2X1 U2813 ( .D0(n1618), .D1(n1746), .S(n3875), .Y(n156) );
  MUX2X1 U2814 ( .D0(n1693), .D1(n1821), .S(n3867), .Y(n231) );
  AO22XL U2815 ( .A(n3979), .B(A[291]), .C(n3959), .D(A[803]), .Y(n1450) );
  AO22XL U2816 ( .A(n3980), .B(A[35]), .C(n3992), .D(A[547]), .Y(n1449) );
  AO22XL U2817 ( .A(n3970), .B(A[36]), .C(n3959), .D(A[548]), .Y(n1443) );
  MUX2IX1 U2818 ( .D0(n3803), .D1(n3830), .S(n3868), .Y(n227) );
  MUX2IXL U2819 ( .D0(n119), .D1(n183), .S(n3864), .Y(n55) );
  MUX2IX1 U2820 ( .D0(n3682), .D1(n3717), .S(n3876), .Y(n142) );
  MUX2X1 U2821 ( .D0(n1696), .D1(n1824), .S(n3867), .Y(n234) );
  MUX2IX1 U2822 ( .D0(n155), .D1(n219), .S(n3861), .Y(n91) );
  MUX2IX1 U2823 ( .D0(n3726), .D1(n3722), .S(n3870), .Y(n202) );
  MUX2XL U2824 ( .D0(n121), .D1(n185), .S(n3864), .Y(n3698) );
  MUX2X1 U2825 ( .D0(n158), .D1(n222), .S(n3860), .Y(n3690) );
  NAND2XL U2826 ( .A(n1302), .B(n3894), .Y(n1641) );
  MUX2IX4 U2827 ( .D0(n3), .D1(n11), .S(SH[3]), .Y(B[2]) );
  OR2X1 U2828 ( .A(n3946), .B(A[237]), .Y(n3786) );
  AND2XL U2829 ( .A(n3909), .B(n1278), .Y(n3825) );
  NOR21XL U2830 ( .B(n3993), .A(A[530]), .Y(n1523) );
  MUX2IX1 U2831 ( .D0(A[285]), .D1(A[797]), .S(n3992), .Y(n1480) );
  AO22AXL U2832 ( .A(n1443), .B(n3914), .C(n3687), .D(n3760), .Y(n1611) );
  INVXL U2833 ( .A(n1660), .Y(n318) );
  AO22XL U2834 ( .A(n3851), .B(A[251]), .C(n3986), .D(A[763]), .Y(n515) );
  NOR21XL U2835 ( .B(n3939), .A(A[594]), .Y(n1256) );
  MUX2XL U2836 ( .D0(n161), .D1(n225), .S(n3860), .Y(n3695) );
  MUX2IXL U2837 ( .D0(n162), .D1(n226), .S(n3860), .Y(n98) );
  MUX2IXL U2838 ( .D0(n164), .D1(n228), .S(n3860), .Y(n100) );
  MUX2IXL U2839 ( .D0(n166), .D1(n230), .S(n3860), .Y(n102) );
  INVX1 U2840 ( .A(n3854), .Y(n3852) );
  INVX1 U2841 ( .A(n3965), .Y(n3949) );
  INVXL U2842 ( .A(n3866), .Y(n3860) );
  AND2XL U2843 ( .A(n3741), .B(n3879), .Y(n3711) );
  MUX2AXL U2844 ( .D0(n130), .D1(n3704), .S(n3863), .Y(n66) );
  MUX2XL U2845 ( .D0(n129), .D1(n193), .S(n3863), .Y(n3694) );
  INVXL U2846 ( .A(n1483), .Y(n3737) );
  MUX2IXL U2847 ( .D0(n3737), .D1(n3832), .S(n3800), .Y(n3756) );
  MUX2XL U2848 ( .D0(A[493]), .D1(A[1005]), .S(n3930), .Y(n3787) );
  MUX2AX1 U2849 ( .D0(A[188]), .D1(n3804), .S(n3928), .Y(n773) );
  MUX2IXL U2850 ( .D0(A[477]), .D1(A[989]), .S(n3835), .Y(n658) );
  NOR21XL U2851 ( .B(n3937), .A(A[837]), .Y(n1293) );
  INVXL U2852 ( .A(n3904), .Y(n3894) );
  INVXL U2853 ( .A(n3966), .Y(n3941) );
  INVXL U2854 ( .A(n3967), .Y(n3934) );
  INVXL U2855 ( .A(n3812), .Y(n3906) );
  INVXL U2856 ( .A(n3880), .Y(n3879) );
  MUX2IXL U2857 ( .D0(n160), .D1(n224), .S(n3860), .Y(n96) );
  MUX2IX1 U2858 ( .D0(n26), .D1(n42), .S(n3852), .Y(n10) );
  INVXL U2859 ( .A(SH[7]), .Y(n3881) );
  NAND2XL U2860 ( .A(n3718), .B(n3879), .Y(n119) );
  MUX2XL U2861 ( .D0(n314), .D1(n3714), .S(n3871), .Y(n3704) );
  MUX2X1 U2862 ( .D0(n1602), .D1(n1730), .S(n3877), .Y(n140) );
  MUX2XL U2863 ( .D0(n1632), .D1(n1760), .S(n3874), .Y(n170) );
  MUX2IXL U2864 ( .D0(n320), .D1(n3674), .S(n3871), .Y(n200) );
  INVXL U2865 ( .A(n1651), .Y(n309) );
  MUX2IX1 U2866 ( .D0(n170), .D1(n234), .S(n3859), .Y(n106) );
  MUX2AXL U2867 ( .D0(n3693), .D1(n1751), .S(n3874), .Y(n161) );
  MUX2XL U2868 ( .D0(n1640), .D1(n1768), .S(n3873), .Y(n178) );
  MUX2BXL U2869 ( .D0(n1671), .D1(n3696), .S(n3870), .Y(n209) );
  MUX2XL U2870 ( .D0(n1616), .D1(n1744), .S(n3875), .Y(n154) );
  MUX2X1 U2871 ( .D0(n1657), .D1(n1785), .S(n3871), .Y(n195) );
  AO22X1 U2872 ( .A(n3978), .B(A[45]), .C(n3956), .D(A[557]), .Y(n3716) );
  MUX2IX1 U2873 ( .D0(n3834), .D1(n3844), .S(n3875), .Y(n155) );
  NOR21XL U2874 ( .B(n3942), .A(A[532]), .Y(n1515) );
  MUX2IXL U2875 ( .D0(n1335), .D1(n1336), .S(n3800), .Y(n1632) );
  MUX2IXL U2876 ( .D0(A[316]), .D1(A[828]), .S(n3927), .Y(n1324) );
  NOR21XL U2877 ( .B(n3935), .A(A[716]), .Y(n717) );
  MUX2IXL U2878 ( .D0(A[484]), .D1(A[996]), .S(n3932), .Y(n630) );
  MUX2XL U2879 ( .D0(n1073), .D1(n1074), .S(n3884), .Y(n3741) );
  AO22XL U2880 ( .A(n3982), .B(A[241]), .C(n3954), .D(A[753]), .Y(n575) );
  AO22XL U2881 ( .A(n3851), .B(A[249]), .C(n3956), .D(A[761]), .Y(n527) );
  MUX2XL U2882 ( .D0(n1169), .D1(n1170), .S(n3801), .Y(n3720) );
  INVXL U2883 ( .A(n3986), .Y(n3978) );
  INVXL U2884 ( .A(n3793), .Y(n3798) );
  INVXL U2885 ( .A(n3970), .Y(n3950) );
  INVXL U2886 ( .A(n3982), .Y(n3936) );
  INVXL U2887 ( .A(n3997), .Y(n3962) );
  INVXL U2888 ( .A(n3982), .Y(n3945) );
  INVXL U2889 ( .A(n3965), .Y(n3951) );
  INVX1 U2890 ( .A(n3987), .Y(n3982) );
  INVXL U2891 ( .A(n3986), .Y(n3985) );
  MUX2IX1 U2892 ( .D0(n63), .D1(n95), .S(n3856), .Y(n31) );
  MUX2IX1 U2893 ( .D0(n64), .D1(n96), .S(n3856), .Y(n32) );
  MUX2IX1 U2894 ( .D0(n80), .D1(n112), .S(n3855), .Y(n48) );
  NAND2X1 U2895 ( .A(n3775), .B(n3879), .Y(n117) );
  MUX2IX1 U2896 ( .D0(n72), .D1(n104), .S(n3855), .Y(n40) );
  MUX2IX1 U2897 ( .D0(n168), .D1(n232), .S(n3859), .Y(n104) );
  NAND2XL U2898 ( .A(n3776), .B(n3879), .Y(n118) );
  MUX2IX1 U2899 ( .D0(n3738), .D1(n3773), .S(n3867), .Y(n239) );
  MUX2IX1 U2900 ( .D0(n175), .D1(n239), .S(n3859), .Y(n111) );
  MUX2X1 U2901 ( .D0(n1597), .D1(n1725), .S(n3877), .Y(n135) );
  MUX2IX1 U2902 ( .D0(n176), .D1(n240), .S(n3859), .Y(n112) );
  MUX2IX1 U2903 ( .D0(n55), .D1(n87), .S(n3857), .Y(n23) );
  MUX2X1 U2904 ( .D0(n1323), .D1(n1324), .S(n3888), .Y(n3750) );
  MUX2X1 U2905 ( .D0(n1624), .D1(n1752), .S(n3874), .Y(n162) );
  MUX2IX1 U2906 ( .D0(n131), .D1(n195), .S(n3863), .Y(n67) );
  MUX2X1 U2907 ( .D0(n1093), .D1(n1094), .S(n3883), .Y(n3751) );
  MUX2X1 U2908 ( .D0(n645), .D1(n646), .S(n3890), .Y(n3696) );
  MUX2X1 U2909 ( .D0(n1614), .D1(n1742), .S(n3875), .Y(n152) );
  MUX2X1 U2910 ( .D0(n1653), .D1(n1781), .S(n3871), .Y(n191) );
  MUX2X1 U2911 ( .D0(n1698), .D1(n1826), .S(n3867), .Y(n236) );
  MUX2X1 U2912 ( .D0(n1594), .D1(n1722), .S(n3877), .Y(n132) );
  MUX2X1 U2913 ( .D0(n1598), .D1(n1726), .S(n3877), .Y(n136) );
  MUX2X1 U2914 ( .D0(n605), .D1(n3790), .S(n3793), .Y(n3709) );
  AND2XL U2915 ( .A(n693), .B(n3793), .Y(n3715) );
  AND2XL U2916 ( .A(n684), .B(n3762), .Y(n3712) );
  MUX2IXL U2917 ( .D0(n3783), .D1(n3785), .S(n3868), .Y(n222) );
  MUX2IXL U2918 ( .D0(n318), .D1(n3683), .S(n3871), .Y(n198) );
  MUX2XL U2919 ( .D0(n1644), .D1(n1772), .S(n3872), .Y(n182) );
  MUX2X1 U2920 ( .D0(n1599), .D1(n1727), .S(n3877), .Y(n137) );
  MUX2XL U2921 ( .D0(n1652), .D1(n1780), .S(n3872), .Y(n190) );
  AND2XL U2922 ( .A(n702), .B(n3762), .Y(n3713) );
  MUX2IXL U2923 ( .D0(n317), .D1(n3684), .S(n3871), .Y(n197) );
  MUX2IX1 U2924 ( .D0(A[490]), .D1(A[1002]), .S(n3945), .Y(n3790) );
  AO22XL U2925 ( .A(n3985), .B(A[421]), .C(n3960), .D(A[933]), .Y(n904) );
  NOR21XL U2926 ( .B(n3941), .A(A[564]), .Y(n1355) );
  NOR2XL U2927 ( .A(n3945), .B(A[444]), .Y(n774) );
  NOR2XL U2928 ( .A(n3952), .B(A[346]), .Y(n1230) );
  NOR2XL U2929 ( .A(n3952), .B(A[385]), .Y(n1074) );
  NOR21XL U2930 ( .B(n3941), .A(A[562]), .Y(n1363) );
  MUX2IX1 U2931 ( .D0(n3848), .D1(n3816), .S(n3881), .Y(n147) );
  AOI22X1 U2932 ( .A(n3969), .B(A[46]), .C(n3961), .D(A[558]), .Y(n3766) );
  MUX2IXL U2933 ( .D0(n1217), .D1(n1218), .S(n3887), .Y(n1668) );
  NOR21XL U2934 ( .B(n3942), .A(A[605]), .Y(n1217) );
  MUX2IXL U2935 ( .D0(n713), .D1(n714), .S(n3801), .Y(n1780) );
  MUX2IXL U2936 ( .D0(n977), .D1(n978), .S(n3886), .Y(n1724) );
  MUX2IXL U2937 ( .D0(A[405]), .D1(A[917]), .S(n3926), .Y(n978) );
  NOR21XL U2938 ( .B(n3939), .A(A[597]), .Y(n1247) );
  NOR21XL U2939 ( .B(n3938), .A(A[589]), .Y(n1269) );
  NOR21XL U2940 ( .B(n3936), .A(A[629]), .Y(n1121) );
  NOR2XL U2941 ( .A(n3952), .B(A[135]), .Y(n1049) );
  NOR2XL U2942 ( .A(n3951), .B(A[134]), .Y(n1053) );
  NOR2XL U2943 ( .A(n3951), .B(A[131]), .Y(n1065) );
  NOR2XL U2944 ( .A(n3950), .B(A[128]), .Y(n1077) );
  MUX2XL U2945 ( .D0(n1057), .D1(n1058), .S(n3884), .Y(n3776) );
  NOR2XL U2946 ( .A(n3951), .B(A[133]), .Y(n1057) );
  NOR21XL U2947 ( .B(n3943), .A(A[525]), .Y(n1543) );
  NOR21XL U2948 ( .B(n3941), .A(A[541]), .Y(n1479) );
  INVX1 U2949 ( .A(n3903), .Y(n3898) );
  INVXL U2950 ( .A(n3996), .Y(n3954) );
  INVXL U2951 ( .A(n3971), .Y(n3944) );
  INVXL U2952 ( .A(n3967), .Y(n3946) );
  INVXL U2953 ( .A(n3982), .Y(n3947) );
  INVXL U2954 ( .A(n3970), .Y(n3957) );
  INVXL U2955 ( .A(n3975), .Y(n3938) );
  INVXL U2956 ( .A(n3972), .Y(n3943) );
  INVXL U2957 ( .A(n3967), .Y(n3937) );
  INVXL U2958 ( .A(n3812), .Y(n3907) );
  INVXL U2959 ( .A(n3866), .Y(n3861) );
  INVXL U2960 ( .A(n3987), .Y(n3981) );
  INVX1 U2961 ( .A(n3920), .Y(n3908) );
  INVXL U2962 ( .A(n3866), .Y(n3865) );
  INVX1 U2963 ( .A(n3921), .Y(n3905) );
  MUX2IXL U2964 ( .D0(n127), .D1(n191), .S(n3863), .Y(n63) );
  MUX2XL U2965 ( .D0(n1593), .D1(n1721), .S(n3877), .Y(n131) );
  MUX2IXL U2966 ( .D0(n1523), .D1(n1524), .S(n3900), .Y(n1593) );
  NAND2XL U2967 ( .A(n696), .B(n3895), .Y(n1785) );
  MUX2XL U2968 ( .D0(n1551), .D1(n1552), .S(n3894), .Y(n3746) );
  MUX2IX1 U2969 ( .D0(n76), .D1(n108), .S(n3855), .Y(n44) );
  MUX2IXL U2970 ( .D0(n140), .D1(n204), .S(n3862), .Y(n76) );
  MUX2IXL U2971 ( .D0(n172), .D1(n236), .S(n3859), .Y(n108) );
  MUX2IXL U2972 ( .D0(n3727), .D1(n3723), .S(n3870), .Y(n204) );
  MUX2XL U2973 ( .D0(n1371), .D1(n1372), .S(n3800), .Y(n3693) );
  MUX2XL U2974 ( .D0(n1631), .D1(n1759), .S(n3874), .Y(n169) );
  MUX2X1 U2975 ( .D0(n3694), .D1(n3695), .S(n3856), .Y(n33) );
  MUX2IXL U2976 ( .D0(n159), .D1(n223), .S(n3860), .Y(n95) );
  MUX2IXL U2977 ( .D0(n3666), .D1(n3732), .S(n3868), .Y(n223) );
  MUX2IXL U2978 ( .D0(n3764), .D1(n3757), .S(n3875), .Y(n159) );
  MUX2XL U2979 ( .D0(n1674), .D1(n1802), .S(n3869), .Y(n212) );
  MUX2IXL U2980 ( .D0(n144), .D1(n208), .S(n3862), .Y(n80) );
  MUX2IXL U2981 ( .D0(n3662), .D1(n3721), .S(n3870), .Y(n208) );
  MUX2IXL U2982 ( .D0(n3744), .D1(n3719), .S(n3876), .Y(n144) );
  MUX2IXL U2983 ( .D0(n143), .D1(n207), .S(n3862), .Y(n79) );
  MUX2IXL U2984 ( .D0(n3663), .D1(n3733), .S(n3870), .Y(n207) );
  MUX2IXL U2985 ( .D0(n132), .D1(n3697), .S(n3863), .Y(n68) );
  MUX2IXL U2986 ( .D0(n316), .D1(n3715), .S(n3871), .Y(n3697) );
  MUX2IXL U2987 ( .D0(n145), .D1(n209), .S(n3862), .Y(n81) );
  NAND2XL U2988 ( .A(n3743), .B(n3879), .Y(n113) );
  MUX2X1 U2989 ( .D0(n3698), .D1(n3699), .S(n3857), .Y(n25) );
  MUX2IXL U2990 ( .D0(n151), .D1(n215), .S(n3861), .Y(n87) );
  MUX2IXL U2991 ( .D0(n308), .D1(n3728), .S(n3872), .Y(n188) );
  MUX2X1 U2992 ( .D0(n3700), .D1(n3701), .S(n3855), .Y(n41) );
  MUX2XL U2993 ( .D0(n137), .D1(n201), .S(n3862), .Y(n3700) );
  MUX2X1 U2994 ( .D0(n169), .D1(n233), .S(n3859), .Y(n3701) );
  MUX2IXL U2995 ( .D0(n136), .D1(n200), .S(n3863), .Y(n72) );
  MUX2IXL U2996 ( .D0(n135), .D1(n199), .S(n3863), .Y(n71) );
  MUX2IXL U2997 ( .D0(n167), .D1(n231), .S(n3859), .Y(n103) );
  MUX2IXL U2998 ( .D0(n319), .D1(n3712), .S(n3871), .Y(n199) );
  MUX2IXL U2999 ( .D0(n128), .D1(n192), .S(n3863), .Y(n64) );
  MUX2IXL U3000 ( .D0(n312), .D1(n3745), .S(n3871), .Y(n192) );
  MUX2IXL U3001 ( .D0(n3725), .D1(n3770), .S(n3878), .Y(n128) );
  NAND2XL U3002 ( .A(n3740), .B(n3879), .Y(n116) );
  MUX2IX2 U3003 ( .D0(n116), .D1(n180), .S(n3865), .Y(n52) );
  MUX2IXL U3004 ( .D0(n3724), .D1(n3665), .S(n3873), .Y(n176) );
  MUX2IXL U3005 ( .D0(n3730), .D1(n3767), .S(n3867), .Y(n240) );
  MUX2IXL U3006 ( .D0(n3734), .D1(n3664), .S(n3873), .Y(n175) );
  NAND21XL U3007 ( .B(n3897), .A(n1272), .Y(n1651) );
  MUX2X1 U3008 ( .D0(n1641), .D1(n1769), .S(n3873), .Y(n179) );
  MUX2XL U3009 ( .D0(n981), .D1(n982), .S(n3886), .Y(n3749) );
  MUX2XL U3010 ( .D0(n1157), .D1(n1158), .S(n3882), .Y(n3748) );
  MUX2XL U3011 ( .D0(n1109), .D1(n1110), .S(n3883), .Y(n3706) );
  MUX2XL U3012 ( .D0(n1563), .D1(n1564), .S(n3888), .Y(n3707) );
  NAND2XL U3013 ( .A(n752), .B(n3895), .Y(n1769) );
  NAND2XL U3014 ( .A(n743), .B(n3895), .Y(n1772) );
  MUX2X1 U3015 ( .D0(n661), .D1(n662), .S(n3890), .Y(n3752) );
  MUX2XL U3016 ( .D0(n1647), .D1(n1775), .S(n3872), .Y(n185) );
  MUX2XL U3017 ( .D0(n1645), .D1(n1773), .S(n3872), .Y(n183) );
  MUX2AXL U3018 ( .D0(n3708), .D1(n1815), .S(n3868), .Y(n225) );
  MUX2XL U3019 ( .D0(n1141), .D1(n1142), .S(n3882), .Y(n3708) );
  MUX2XL U3020 ( .D0(n1610), .D1(n1738), .S(n3876), .Y(n148) );
  MUX2XL U3021 ( .D0(n1622), .D1(n1750), .S(n3875), .Y(n160) );
  NAND2XL U3022 ( .A(n1293), .B(n3894), .Y(n1644) );
  MUX2XL U3023 ( .D0(n1129), .D1(n1130), .S(n3883), .Y(n3710) );
  MUX2XL U3024 ( .D0(n1584), .D1(n1712), .S(n3878), .Y(n122) );
  MUX2XL U3025 ( .D0(n1648), .D1(n1776), .S(n3872), .Y(n186) );
  MUX2XL U3026 ( .D0(n1592), .D1(n1720), .S(n3878), .Y(n130) );
  MUX2XL U3027 ( .D0(n1678), .D1(n1806), .S(n3869), .Y(n216) );
  MUX2IXL U3028 ( .D0(n56), .D1(n88), .S(n3857), .Y(n24) );
  MUX2IXL U3029 ( .D0(n120), .D1(n184), .S(n3864), .Y(n56) );
  MUX2IXL U3030 ( .D0(n152), .D1(n216), .S(n3861), .Y(n88) );
  NAND2XL U3031 ( .A(n3742), .B(n3879), .Y(n120) );
  MUX2XL U3032 ( .D0(n1646), .D1(n1774), .S(n3872), .Y(n184) );
  MUX2XL U3033 ( .D0(n1608), .D1(n1736), .S(n3876), .Y(n146) );
  AND2XL U3034 ( .A(n699), .B(n3762), .Y(n3714) );
  MUX2IXL U3035 ( .D0(n3786), .D1(n3787), .S(n3893), .Y(n3785) );
  MUX2IXL U3036 ( .D0(A[492]), .D1(A[1004]), .S(n3648), .Y(n598) );
  MUX2IXL U3037 ( .D0(n1205), .D1(n1206), .S(n3887), .Y(n1671) );
  MUX2IXL U3038 ( .D0(n585), .D1(n586), .S(n3893), .Y(n1814) );
  MUX2IXL U3039 ( .D0(A[495]), .D1(A[1007]), .S(n3835), .Y(n586) );
  MUX2IXL U3040 ( .D0(A[191]), .D1(A[703]), .S(n3929), .Y(n761) );
  MUX2IXL U3041 ( .D0(A[317]), .D1(A[829]), .S(n3927), .Y(n1320) );
  MUX2IXL U3042 ( .D0(n621), .D1(n622), .S(n3891), .Y(n1805) );
  MUX2IXL U3043 ( .D0(n709), .D1(n710), .S(n3801), .Y(n1781) );
  MUX2IXL U3044 ( .D0(n733), .D1(n734), .S(n3801), .Y(n1775) );
  MUX2IXL U3045 ( .D0(A[120]), .D1(A[632]), .S(n3925), .Y(n1109) );
  AOI22XL U3046 ( .A(n1438), .B(n3901), .C(n1437), .D(n3916), .Y(n3792) );
  MUX2IXL U3047 ( .D0(n1339), .D1(n1340), .S(n3889), .Y(n1631) );
  MUX2IXL U3048 ( .D0(n965), .D1(n966), .S(n3886), .Y(n1727) );
  MUX2IXL U3049 ( .D0(A[408]), .D1(A[920]), .S(n3926), .Y(n966) );
  MUX2IXL U3050 ( .D0(n973), .D1(n974), .S(n3886), .Y(n1725) );
  MUX2IXL U3051 ( .D0(n969), .D1(n970), .S(n3886), .Y(n1726) );
  MUX2IXL U3052 ( .D0(A[407]), .D1(A[919]), .S(n3929), .Y(n970) );
  MUX2IXL U3053 ( .D0(A[184]), .D1(A[696]), .S(n3927), .Y(n789) );
  MUX2IXL U3054 ( .D0(n777), .D1(n778), .S(n3889), .Y(n1762) );
  MUX2IX1 U3055 ( .D0(A[308]), .D1(A[820]), .S(n3929), .Y(n1356) );
  MUX2IXL U3056 ( .D0(n997), .D1(n998), .S(n3885), .Y(n1719) );
  MUX2IXL U3057 ( .D0(A[400]), .D1(A[912]), .S(n3925), .Y(n998) );
  MUX2IXL U3058 ( .D0(n601), .D1(n602), .S(n3892), .Y(n1810) );
  MUX2IXL U3059 ( .D0(A[491]), .D1(A[1003]), .S(n3648), .Y(n602) );
  MUX2IXL U3060 ( .D0(n633), .D1(n634), .S(n3892), .Y(n1802) );
  AOI22BXL U3061 ( .B(n3765), .A(n3687), .D(n3766), .C(n3913), .Y(n3764) );
  MUX2IXL U3062 ( .D0(A[480]), .D1(A[992]), .S(n3933), .Y(n646) );
  MUX2IXL U3063 ( .D0(A[123]), .D1(A[635]), .S(n3925), .Y(n1097) );
  MUX2IXL U3064 ( .D0(A[309]), .D1(A[821]), .S(n3928), .Y(n1352) );
  MUX2IXL U3065 ( .D0(A[266]), .D1(A[778]), .S(n3930), .Y(n1556) );
  MUX2IXL U3066 ( .D0(n1487), .D1(n1488), .S(n3890), .Y(n1602) );
  MUX2IXL U3067 ( .D0(A[283]), .D1(A[795]), .S(n3933), .Y(n1488) );
  MUX2IXL U3068 ( .D0(A[190]), .D1(A[702]), .S(n3929), .Y(n765) );
  MUX2IXL U3069 ( .D0(A[269]), .D1(A[781]), .S(n3930), .Y(n1544) );
  AOI22AXL U3070 ( .A(n497), .B(n3910), .D(n3774), .C(n3762), .Y(n3773) );
  MUX2XL U3071 ( .D0(n1053), .D1(n1054), .S(n3884), .Y(n3718) );
  MUX2XL U3072 ( .D0(n3755), .D1(n1491), .S(n3912), .Y(n3838) );
  NOR2XL U3073 ( .A(n3946), .B(A[234]), .Y(n605) );
  NOR21XL U3074 ( .B(n3939), .A(A[600]), .Y(n1237) );
  MUX2XL U3075 ( .D0(n937), .D1(n938), .S(n3887), .Y(n3719) );
  MUX2XL U3076 ( .D0(n649), .D1(n650), .S(n3891), .Y(n3721) );
  MUX2XL U3077 ( .D0(n673), .D1(n674), .S(n3891), .Y(n3722) );
  MUX2XL U3078 ( .D0(n665), .D1(n666), .S(n3801), .Y(n3723) );
  MUX2XL U3079 ( .D0(n1311), .D1(n1312), .S(n3888), .Y(n3724) );
  MUX2XL U3080 ( .D0(n1535), .D1(n1536), .S(n3894), .Y(n3725) );
  MUX2XL U3081 ( .D0(n1233), .D1(n1234), .S(n3888), .Y(n3726) );
  MUX2XL U3082 ( .D0(n1225), .D1(n1226), .S(n3888), .Y(n3727) );
  MUX2XL U3083 ( .D0(n721), .D1(n722), .S(n3889), .Y(n3728) );
  MUX2XL U3084 ( .D0(n677), .D1(n678), .S(n3890), .Y(n3729) );
  MUX2XL U3085 ( .D0(n1081), .D1(n1082), .S(n3884), .Y(n3730) );
  MUX2X1 U3086 ( .D0(n609), .D1(n610), .S(n3793), .Y(n3731) );
  MUX2XL U3087 ( .D0(n1061), .D1(n1062), .S(n3884), .Y(n3775) );
  NOR2XL U3088 ( .A(n3951), .B(A[132]), .Y(n1061) );
  MUX2XL U3089 ( .D0(n1069), .D1(n1070), .S(n3884), .Y(n3802) );
  NOR2XL U3090 ( .A(n3951), .B(A[130]), .Y(n1069) );
  MUX2XL U3091 ( .D0(n589), .D1(n590), .S(n3892), .Y(n3732) );
  MUX2XL U3092 ( .D0(n653), .D1(n654), .S(n3891), .Y(n3733) );
  MUX2XL U3093 ( .D0(n1315), .D1(n1316), .S(n3888), .Y(n3734) );
  MUX2XL U3094 ( .D0(n941), .D1(n942), .S(n3887), .Y(n3735) );
  MUX2XL U3095 ( .D0(n1475), .D1(n1476), .S(n3889), .Y(n3736) );
  MUX2BXL U3096 ( .D0(n1173), .D1(n3781), .S(n3885), .Y(n3780) );
  AO22XL U3097 ( .A(n3971), .B(A[252]), .C(n3953), .D(A[764]), .Y(n509) );
  AO22AXL U3098 ( .A(n819), .B(n3910), .C(n3899), .D(n3761), .Y(n1754) );
  AO22XL U3099 ( .A(n3981), .B(A[240]), .C(n3954), .D(A[752]), .Y(n581) );
  AO22XL U3100 ( .A(n3972), .B(A[246]), .C(n3953), .D(A[758]), .Y(n545) );
  MUX2XL U3101 ( .D0(n1085), .D1(n1086), .S(n3884), .Y(n3738) );
  MUX2XL U3102 ( .D0(n1125), .D1(n1126), .S(n3883), .Y(n3784) );
  NOR2XL U3103 ( .A(n3949), .B(A[372]), .Y(n1126) );
  MUX2IXL U3104 ( .D0(n3739), .D1(n1495), .S(n3909), .Y(n1600) );
  MUX2IXL U3105 ( .D0(A[281]), .D1(A[793]), .S(n3933), .Y(n3739) );
  MUX2IXL U3106 ( .D0(A[268]), .D1(A[780]), .S(n3930), .Y(n1548) );
  INVXL U3107 ( .A(n3916), .Y(n3762) );
  MUX2IXL U3108 ( .D0(n641), .D1(n642), .S(n3891), .Y(n1800) );
  MUX2IXL U3109 ( .D0(A[481]), .D1(A[993]), .S(n3933), .Y(n642) );
  MUX2IXL U3110 ( .D0(n993), .D1(n994), .S(n3886), .Y(n1720) );
  MUX2IXL U3111 ( .D0(A[401]), .D1(A[913]), .S(n3925), .Y(n994) );
  MUX2IXL U3112 ( .D0(n1177), .D1(n1178), .S(n3885), .Y(n1678) );
  AOI22BXL U3113 ( .B(n3771), .A(n3898), .D(n3772), .C(n3912), .Y(n3770) );
  MUX2IXL U3114 ( .D0(A[264]), .D1(A[776]), .S(n3930), .Y(n1564) );
  MUX2IXL U3115 ( .D0(A[265]), .D1(A[777]), .S(n3835), .Y(n1560) );
  AOI22BXL U3116 ( .B(n3768), .A(n3762), .D(n3769), .C(n3914), .Y(n3767) );
  MUX2XL U3117 ( .D0(n1065), .D1(n1066), .S(n3884), .Y(n3740) );
  MUX2XL U3118 ( .D0(n1049), .D1(n1050), .S(n3885), .Y(n3742) );
  MUX2XL U3119 ( .D0(n1077), .D1(n1078), .S(n3884), .Y(n3743) );
  MUX2XL U3120 ( .D0(n1471), .D1(n1472), .S(n3890), .Y(n3744) );
  MUX2XL U3121 ( .D0(n705), .D1(n706), .S(n3890), .Y(n3745) );
  INVXL U3122 ( .A(n1656), .Y(n314) );
  AO22XL U3123 ( .A(n3981), .B(A[247]), .C(n3954), .D(A[759]), .Y(n539) );
  AO22XL U3124 ( .A(n3971), .B(A[248]), .C(n3953), .D(A[760]), .Y(n533) );
  INVXL U3125 ( .A(n3986), .Y(n3979) );
  INVXL U3126 ( .A(n3986), .Y(n3980) );
  INVX1 U3127 ( .A(n3687), .Y(n3913) );
  INVX1 U3128 ( .A(n3901), .Y(n3817) );
  INVX1 U3129 ( .A(n3854), .Y(n3853) );
  INVXL U3130 ( .A(n3968), .Y(n3931) );
  INVX1 U3131 ( .A(n3908), .Y(n3885) );
  INVX1 U3132 ( .A(n3907), .Y(n3886) );
  INVXL U3133 ( .A(n3966), .Y(n3940) );
  INVX1 U3134 ( .A(n3964), .Y(n3930) );
  INVX1 U3135 ( .A(n3907), .Y(n3888) );
  INVX1 U3136 ( .A(n3907), .Y(n3887) );
  INVX1 U3137 ( .A(n3906), .Y(n3800) );
  INVX1 U3138 ( .A(n3906), .Y(n3801) );
  INVX1 U3139 ( .A(n3906), .Y(n3889) );
  INVX1 U3140 ( .A(n3908), .Y(n3883) );
  INVX1 U3141 ( .A(n3908), .Y(n3884) );
  INVXL U3142 ( .A(n3904), .Y(n3895) );
  INVXL U3143 ( .A(n3968), .Y(n3929) );
  INVX1 U3144 ( .A(n3967), .Y(n3932) );
  INVX1 U3145 ( .A(n3964), .Y(n3928) );
  INVXL U3146 ( .A(n3968), .Y(n3925) );
  INVXL U3147 ( .A(n3968), .Y(n3926) );
  INVXL U3148 ( .A(n3967), .Y(n3933) );
  INVXL U3149 ( .A(n3998), .Y(n3958) );
  INVXL U3150 ( .A(n3903), .Y(n3899) );
  INVXL U3151 ( .A(n3968), .Y(n3956) );
  INVXL U3152 ( .A(n3966), .Y(n3939) );
  INVX1 U3153 ( .A(n3967), .Y(n3935) );
  INVX1 U3154 ( .A(n3967), .Y(n3960) );
  INVX1 U3155 ( .A(SH[4]), .Y(n3854) );
  INVX1 U3156 ( .A(n3905), .Y(n3892) );
  INVX1 U3157 ( .A(n3905), .Y(n3890) );
  INVX1 U3158 ( .A(n3881), .Y(n3869) );
  INVX1 U3159 ( .A(n3881), .Y(n3868) );
  INVX1 U3160 ( .A(n3881), .Y(n3876) );
  INVX1 U3161 ( .A(n3905), .Y(n3891) );
  INVX1 U3162 ( .A(n3924), .Y(n3882) );
  INVX1 U3163 ( .A(n3880), .Y(n3870) );
  INVX1 U3164 ( .A(n3881), .Y(n3871) );
  INVX1 U3165 ( .A(n3880), .Y(n3872) );
  INVX1 U3166 ( .A(n3881), .Y(n3873) );
  INVX1 U3167 ( .A(n3881), .Y(n3874) );
  INVX1 U3168 ( .A(n3881), .Y(n3875) );
  INVX1 U3169 ( .A(n3812), .Y(n3902) );
  INVX1 U3170 ( .A(n3924), .Y(n3793) );
  INVX1 U3171 ( .A(n3919), .Y(n3912) );
  INVXL U3172 ( .A(n3989), .Y(n3977) );
  INVXL U3173 ( .A(n3986), .Y(n3984) );
  INVXL U3174 ( .A(n3990), .Y(n3973) );
  INVXL U3175 ( .A(n3989), .Y(n3975) );
  INVX1 U3176 ( .A(n3921), .Y(n3916) );
  MUX2IX1 U3177 ( .D0(n32), .D1(n48), .S(n3852), .Y(n16) );
  MUX2IX1 U3178 ( .D0(n31), .D1(n47), .S(n3852), .Y(n15) );
  MUX2IX1 U3179 ( .D0(n2), .D1(n10), .S(SH[3]), .Y(B[1]) );
  INVX2 U3180 ( .A(n3995), .Y(n3964) );
  INVX1 U3181 ( .A(n3858), .Y(n3855) );
  INVX1 U3182 ( .A(SH[6]), .Y(n3866) );
  INVX1 U3183 ( .A(SH[5]), .Y(n3858) );
  INVX1 U3184 ( .A(SH[7]), .Y(n3880) );
  MUX2X1 U3185 ( .D0(n1620), .D1(n1748), .S(n3875), .Y(n158) );
  MUX2X1 U3186 ( .D0(n1629), .D1(n1757), .S(n3874), .Y(n167) );
  MUX2IXL U3187 ( .D0(n1347), .D1(n1348), .S(n3801), .Y(n1629) );
  NOR21XL U3188 ( .B(n3936), .A(A[980]), .Y(n690) );
  MUX2X1 U3189 ( .D0(n1588), .D1(n1716), .S(n3878), .Y(n126) );
  MUX2IXL U3190 ( .D0(n1543), .D1(n1544), .S(n3894), .Y(n1588) );
  MUX2IXL U3191 ( .D0(n1137), .D1(n1138), .S(n3882), .Y(n1688) );
  MUX2X1 U3192 ( .D0(n1686), .D1(n1814), .S(n3868), .Y(n224) );
  MUX2IXL U3193 ( .D0(n1145), .D1(n1146), .S(n3882), .Y(n1686) );
  MUX2IXL U3194 ( .D0(n1193), .D1(n1194), .S(n3885), .Y(n1674) );
  MUX2X1 U3195 ( .D0(n1682), .D1(n1810), .S(n3869), .Y(n220) );
  MUX2IXL U3196 ( .D0(n1161), .D1(n1162), .S(n3882), .Y(n1682) );
  MUX2IX1 U3197 ( .D0(n3710), .D1(n3675), .S(n3868), .Y(n228) );
  MUX2X1 U3198 ( .D0(n1677), .D1(n1805), .S(n3869), .Y(n215) );
  MUX2IXL U3199 ( .D0(n1181), .D1(n1182), .S(n3885), .Y(n1677) );
  MUX2IXL U3200 ( .D0(n617), .D1(n618), .S(n3892), .Y(n1806) );
  MUX2IX1 U3201 ( .D0(n3780), .D1(n3777), .S(n3869), .Y(n217) );
  MUX2IX1 U3202 ( .D0(n154), .D1(n218), .S(n3861), .Y(n90) );
  MUX2IX1 U3203 ( .D0(n3720), .D1(n3731), .S(n3869), .Y(n218) );
  MUX2IXL U3204 ( .D0(n1499), .D1(n1500), .S(n3892), .Y(n1599) );
  MUX2IX1 U3205 ( .D0(n51), .D1(n83), .S(n3857), .Y(n19) );
  MUX2IX1 U3206 ( .D0(n115), .D1(n179), .S(n3865), .Y(n51) );
  MUX2IX1 U3207 ( .D0(n147), .D1(n211), .S(n3861), .Y(n83) );
  MUX2IX1 U3208 ( .D0(n1511), .D1(n1512), .S(n3893), .Y(n1596) );
  MUX2IXL U3209 ( .D0(n961), .D1(n962), .S(n3886), .Y(n1728) );
  MUX2IX1 U3210 ( .D0(n3836), .D1(n3672), .S(n3873), .Y(n171) );
  MUX2IXL U3211 ( .D0(n985), .D1(n986), .S(n3886), .Y(n1722) );
  MUX2X1 U3212 ( .D0(n1634), .D1(n1762), .S(n3873), .Y(n172) );
  MUX2IXL U3213 ( .D0(n1327), .D1(n1328), .S(n3888), .Y(n1634) );
  MUX2IXL U3214 ( .D0(n953), .D1(n954), .S(n3887), .Y(n1730) );
  MUX2IXL U3215 ( .D0(n1507), .D1(n1508), .S(n3892), .Y(n1597) );
  MUX2IXL U3216 ( .D0(n1503), .D1(n1504), .S(n3893), .Y(n1598) );
  MUX2X1 U3217 ( .D0(n1694), .D1(n1822), .S(n3867), .Y(n232) );
  MUX2IXL U3218 ( .D0(n1113), .D1(n1114), .S(n3883), .Y(n1694) );
  MUX2IX1 U3219 ( .D0(n49), .D1(n81), .S(SH[5]), .Y(n17) );
  MUX2IX1 U3220 ( .D0(n113), .D1(n177), .S(n3865), .Y(n49) );
  MUX2X1 U3221 ( .D0(n1639), .D1(n1767), .S(n3873), .Y(n177) );
  NAND2XL U3222 ( .A(n1308), .B(n3894), .Y(n1639) );
  MUX2X1 U3223 ( .D0(n1672), .D1(n1800), .S(n3870), .Y(n210) );
  MUX2IXL U3224 ( .D0(n1201), .D1(n1202), .S(n3885), .Y(n1672) );
  NAND2XL U3225 ( .A(n1305), .B(n3895), .Y(n1640) );
  MUX2X1 U3226 ( .D0(n1668), .D1(n1796), .S(n3870), .Y(n206) );
  MUX2IXL U3227 ( .D0(n657), .D1(n658), .S(n3891), .Y(n1796) );
  NAND2XL U3228 ( .A(n1287), .B(n3894), .Y(n1646) );
  NAND2XL U3229 ( .A(n1290), .B(n3895), .Y(n1645) );
  MUX2X1 U3230 ( .D0(n1642), .D1(n1770), .S(n3873), .Y(n180) );
  NAND2XL U3231 ( .A(n1299), .B(n3894), .Y(n1642) );
  MUX2IX1 U3232 ( .D0(n3668), .D1(n3805), .S(n3870), .Y(n203) );
  MUX2IXL U3233 ( .D0(n729), .D1(n730), .S(n3889), .Y(n1776) );
  INVX1 U3234 ( .A(n1654), .Y(n312) );
  NOR21XL U3235 ( .B(n3934), .A(A[969]), .Y(n730) );
  MUX2IXL U3236 ( .D0(n789), .D1(n790), .S(n3800), .Y(n1759) );
  MUX2IX1 U3237 ( .D0(n1351), .D1(n1352), .S(n3800), .Y(n1628) );
  MUX2X1 U3238 ( .D0(n1630), .D1(n1758), .S(n3874), .Y(n168) );
  MUX2IXL U3239 ( .D0(n1343), .D1(n1344), .S(n3800), .Y(n1630) );
  MUX2IXL U3240 ( .D0(n785), .D1(n786), .S(n3800), .Y(n1760) );
  MUX2X1 U3241 ( .D0(n1626), .D1(n1754), .S(n3874), .Y(n164) );
  MUX2IXL U3242 ( .D0(n1359), .D1(n1360), .S(n3889), .Y(n1626) );
  MUX2IX1 U3243 ( .D0(n313), .D1(n3713), .S(n3871), .Y(n193) );
  MUX2IX1 U3244 ( .D0(n3782), .D1(n3729), .S(n3870), .Y(n201) );
  MUX2IX1 U3245 ( .D0(n71), .D1(n103), .S(n3855), .Y(n39) );
  MUX2IXL U3246 ( .D0(n1527), .D1(n1528), .S(n3894), .Y(n1592) );
  MUX2IX1 U3247 ( .D0(n3709), .D1(n3842), .S(n3881), .Y(n219) );
  MUX2IX1 U3248 ( .D0(n78), .D1(n110), .S(n3855), .Y(n46) );
  MUX2IXL U3249 ( .D0(n1117), .D1(n1118), .S(n3883), .Y(n1693) );
  MUX2IX1 U3250 ( .D0(n1319), .D1(n1320), .S(n3888), .Y(n1636) );
  MUX2IXL U3251 ( .D0(n3736), .D1(n3735), .S(n3876), .Y(n143) );
  NOR21XL U3252 ( .B(n3936), .A(A[978]), .Y(n696) );
  NAND2XL U3253 ( .A(n749), .B(n3896), .Y(n1770) );
  NOR21XL U3254 ( .B(n3989), .A(A[963]), .Y(n749) );
  NAND2XL U3255 ( .A(n740), .B(n3793), .Y(n1773) );
  NOR21XL U3256 ( .B(n3686), .A(A[966]), .Y(n740) );
  NAND2XL U3257 ( .A(n737), .B(n3895), .Y(n1774) );
  NOR21XL U3258 ( .B(n3686), .A(A[967]), .Y(n737) );
  NOR21XL U3259 ( .B(n3992), .A(A[965]), .Y(n743) );
  NAND2XL U3260 ( .A(n755), .B(n3793), .Y(n1768) );
  MUX2IXL U3261 ( .D0(n1367), .D1(n1368), .S(n3889), .Y(n1624) );
  MUX2IXL U3262 ( .D0(n1559), .D1(n1560), .S(n3882), .Y(n1584) );
  MUX2IXL U3263 ( .D0(n1097), .D1(n1098), .S(n3883), .Y(n1698) );
  MUX2IXL U3264 ( .D0(n1105), .D1(n1106), .S(n3883), .Y(n1696) );
  NOR21XL U3265 ( .B(n3989), .A(A[962]), .Y(n752) );
  NOR21XL U3266 ( .B(n3936), .A(A[981]), .Y(n687) );
  NOR21XL U3267 ( .B(n3936), .A(A[977]), .Y(n699) );
  NOR21XL U3268 ( .B(n3936), .A(A[979]), .Y(n693) );
  NOR21XL U3269 ( .B(n3926), .A(A[976]), .Y(n702) );
  NOR21XL U3270 ( .B(n3936), .A(A[982]), .Y(n684) );
  NOR21XL U3271 ( .B(n3937), .A(A[983]), .Y(n681) );
  MUX2IX1 U3272 ( .D0(n7), .D1(n15), .S(SH[3]), .Y(B[6]) );
  MUX2IX1 U3273 ( .D0(n23), .D1(n39), .S(n3852), .Y(n7) );
  MUX2IX1 U3274 ( .D0(n1), .D1(n9), .S(SH[3]), .Y(B[0]) );
  MUX2IX1 U3275 ( .D0(n17), .D1(n33), .S(n3853), .Y(n1) );
  MUX2IX1 U3276 ( .D0(n25), .D1(n41), .S(n3852), .Y(n9) );
  MUX2IX1 U3277 ( .D0(n8), .D1(n16), .S(SH[3]), .Y(B[7]) );
  MUX2IX1 U3278 ( .D0(n24), .D1(n40), .S(n3852), .Y(n8) );
  INVX1 U3279 ( .A(A[173]), .Y(n3813) );
  ENOX1 U3280 ( .A(n3986), .B(n3797), .C(n3958), .D(A[946]), .Y(n826) );
  INVX1 U3281 ( .A(A[434]), .Y(n3797) );
  AND2XL U3282 ( .A(n3976), .B(n3808), .Y(n637) );
  INVX1 U3283 ( .A(A[226]), .Y(n3808) );
  MUX2IX1 U3284 ( .D0(A[485]), .D1(A[997]), .S(n3932), .Y(n626) );
  MUX2IXL U3285 ( .D0(A[483]), .D1(A[995]), .S(n3932), .Y(n634) );
  NOR21XL U3286 ( .B(n3942), .A(A[539]), .Y(n1487) );
  NOR21XL U3287 ( .B(n3963), .A(A[656]), .Y(n997) );
  NOR21XL U3288 ( .B(n3935), .A(A[664]), .Y(n965) );
  MUX2IXL U3289 ( .D0(A[406]), .D1(A[918]), .S(n3926), .Y(n974) );
  NOR21XL U3290 ( .B(n3935), .A(A[662]), .Y(n973) );
  NOR21XL U3291 ( .B(n3935), .A(A[615]), .Y(n1177) );
  NOR21XL U3292 ( .B(n3935), .A(A[663]), .Y(n969) );
  NOR21XL U3293 ( .B(n3986), .A(A[657]), .Y(n993) );
  NOR21XL U3294 ( .B(n3942), .A(A[608]), .Y(n1205) );
  NOR21XL U3295 ( .B(n3993), .A(A[607]), .Y(n1209) );
  NOR21XL U3296 ( .B(n3943), .A(A[606]), .Y(n1213) );
  MUX2IXL U3297 ( .D0(A[486]), .D1(A[998]), .S(n3932), .Y(n622) );
  NOR21XL U3298 ( .B(n3940), .A(A[569]), .Y(n1335) );
  MUX2IXL U3299 ( .D0(A[313]), .D1(A[825]), .S(n3928), .Y(n1336) );
  NOR21XL U3300 ( .B(n3928), .A(A[974]), .Y(n710) );
  NOR21XL U3301 ( .B(n3990), .A(A[718]), .Y(n709) );
  NOR21XL U3302 ( .B(n3686), .A(A[968]), .Y(n734) );
  NOR21XL U3303 ( .B(n3990), .A(A[712]), .Y(n733) );
  MUX2IXL U3304 ( .D0(A[187]), .D1(A[699]), .S(n3928), .Y(n777) );
  NOR21XL U3305 ( .B(n3940), .A(A[568]), .Y(n1339) );
  MUX2IXL U3306 ( .D0(A[312]), .D1(A[824]), .S(n3928), .Y(n1340) );
  NOR21XL U3307 ( .B(n3993), .A(A[531]), .Y(n1519) );
  NOR21XL U3308 ( .B(n3938), .A(A[585]), .Y(n1281) );
  NOR21XL U3309 ( .B(n3941), .A(A[832]), .Y(n1308) );
  NOR21XL U3310 ( .B(n3937), .A(A[833]), .Y(n1305) );
  NOR21XL U3311 ( .B(n3937), .A(A[835]), .Y(n1299) );
  NOR21XL U3312 ( .B(n3938), .A(A[838]), .Y(n1290) );
  NOR21XL U3313 ( .B(n3938), .A(A[839]), .Y(n1287) );
  MUX2IXL U3314 ( .D0(A[272]), .D1(A[784]), .S(n3648), .Y(n1532) );
  MUX2IXL U3315 ( .D0(A[270]), .D1(A[782]), .S(n3648), .Y(n1540) );
  MUX2IXL U3316 ( .D0(A[273]), .D1(A[785]), .S(n3648), .Y(n1528) );
  MUX2IXL U3317 ( .D0(A[280]), .D1(A[792]), .S(n3963), .Y(n1500) );
  MUX2IX1 U3318 ( .D0(n3841), .D1(n3846), .S(n3874), .Y(n163) );
  NOR21XL U3319 ( .B(n3941), .A(A[563]), .Y(n1359) );
  MUX2IX1 U3320 ( .D0(n989), .D1(n3685), .S(n3886), .Y(n1721) );
  NOR21XL U3321 ( .B(n3992), .A(A[658]), .Y(n989) );
  MUX2IX1 U3322 ( .D0(n3829), .D1(n3661), .S(n3869), .Y(n211) );
  MUX2X1 U3323 ( .D0(n1198), .D1(n1197), .S(n3911), .Y(n3829) );
  NOR21XL U3324 ( .B(n3940), .A(A[566]), .Y(n1347) );
  NOR21XL U3325 ( .B(n3941), .A(A[560]), .Y(n1371) );
  NOR21XL U3326 ( .B(n3941), .A(A[561]), .Y(n1367) );
  MUX2IXL U3327 ( .D0(A[267]), .D1(A[779]), .S(n3930), .Y(n1552) );
  NOR21XL U3328 ( .B(n3940), .A(A[567]), .Y(n1343) );
  NOR21XL U3329 ( .B(n3942), .A(A[535]), .Y(n1503) );
  NOR21XL U3330 ( .B(n3992), .A(A[624]), .Y(n1141) );
  NOR21XL U3331 ( .B(n3835), .A(A[627]), .Y(n1129) );
  NOR21XL U3332 ( .B(n3990), .A(A[625]), .Y(n1137) );
  NOR21XL U3333 ( .B(n3686), .A(A[619]), .Y(n1161) );
  NOR21XL U3334 ( .B(n3992), .A(A[623]), .Y(n1145) );
  NOR21XL U3335 ( .B(n3943), .A(A[536]), .Y(n1499) );
  NOR21XL U3336 ( .B(n3943), .A(A[526]), .Y(n1539) );
  NOR21XL U3337 ( .B(n3936), .A(A[630]), .Y(n1117) );
  NOR21XL U3338 ( .B(n3936), .A(A[631]), .Y(n1113) );
  NOR21XL U3339 ( .B(n3943), .A(A[529]), .Y(n1527) );
  NOR21XL U3340 ( .B(n3943), .A(A[609]), .Y(n1201) );
  NOR21XL U3341 ( .B(n3936), .A(A[521]), .Y(n1559) );
  NOR21XL U3342 ( .B(n3943), .A(A[611]), .Y(n1193) );
  NOR21XL U3343 ( .B(n3992), .A(A[659]), .Y(n985) );
  NOR21XL U3344 ( .B(n3940), .A(A[571]), .Y(n1327) );
  NOR21XL U3345 ( .B(n3937), .A(A[520]), .Y(n1563) );
  NOR21XL U3346 ( .B(n3990), .A(A[528]), .Y(n1531) );
  NOR21XL U3347 ( .B(n3935), .A(A[665]), .Y(n961) );
  NOR21XL U3348 ( .B(n3925), .A(A[534]), .Y(n1507) );
  NOR21XL U3349 ( .B(n3993), .A(A[614]), .Y(n1181) );
  NOR21XL U3350 ( .B(n3925), .A(A[533]), .Y(n1511) );
  NOR21XL U3351 ( .B(n3993), .A(A[613]), .Y(n1185) );
  NOR21XL U3352 ( .B(n3993), .A(A[523]), .Y(n1551) );
  NOR21XL U3353 ( .B(n3934), .A(A[713]), .Y(n729) );
  NOR21XL U3354 ( .B(n3934), .A(A[667]), .Y(n953) );
  MUX2IX1 U3355 ( .D0(A[277]), .D1(A[789]), .S(n3932), .Y(n1512) );
  MUX2IXL U3356 ( .D0(A[307]), .D1(A[819]), .S(n3929), .Y(n1360) );
  MUX2IXL U3357 ( .D0(A[315]), .D1(A[827]), .S(n3927), .Y(n1328) );
  MUX2IXL U3358 ( .D0(A[279]), .D1(A[791]), .S(n3932), .Y(n1504) );
  MUX2IXL U3359 ( .D0(A[487]), .D1(A[999]), .S(n3932), .Y(n618) );
  MUX2IXL U3360 ( .D0(A[304]), .D1(A[816]), .S(n3929), .Y(n1372) );
  MUX2IXL U3361 ( .D0(A[278]), .D1(A[790]), .S(n3932), .Y(n1508) );
  MUX2IXL U3362 ( .D0(A[305]), .D1(A[817]), .S(n3929), .Y(n1368) );
  NOR21XL U3363 ( .B(n3943), .A(A[522]), .Y(n1555) );
  MUX2IXL U3364 ( .D0(A[185]), .D1(A[697]), .S(n3928), .Y(n785) );
  MUX2IXL U3365 ( .D0(A[311]), .D1(A[823]), .S(n3928), .Y(n1344) );
  MUX2IXL U3366 ( .D0(A[310]), .D1(A[822]), .S(n3928), .Y(n1348) );
  MUX2IXL U3367 ( .D0(A[121]), .D1(A[633]), .S(n3925), .Y(n1105) );
  MUX2IX1 U3368 ( .D0(n3831), .D1(n3839), .S(n3880), .Y(n235) );
  EORX1 U3369 ( .A(n521), .B(n3798), .C(n3824), .D(n3912), .Y(n3831) );
  MUX2IXL U3370 ( .D0(A[403]), .D1(A[915]), .S(n3926), .Y(n986) );
  MUX2IXL U3371 ( .D0(A[411]), .D1(A[923]), .S(n3926), .Y(n954) );
  MUX2IXL U3372 ( .D0(A[409]), .D1(A[921]), .S(n3926), .Y(n962) );
  MUX2IXL U3373 ( .D0(A[698]), .D1(A[186]), .S(n3851), .Y(n781) );
  MUX2IX1 U3374 ( .D0(n769), .D1(n770), .S(n3889), .Y(n1764) );
  MUX2IX1 U3375 ( .D0(A[189]), .D1(A[701]), .S(n3928), .Y(n769) );
  MUX2IXL U3376 ( .D0(A[474]), .D1(A[986]), .S(n3930), .Y(n670) );
  NOR21XL U3377 ( .B(n3938), .A(A[584]), .Y(n1284) );
  NAND2X1 U3378 ( .A(n758), .B(n3762), .Y(n1767) );
  MUX2IXL U3379 ( .D0(A[634]), .D1(A[122]), .S(n3964), .Y(n1101) );
  NOR21XL U3380 ( .B(n3835), .A(A[626]), .Y(n1133) );
  MUX2IX1 U3381 ( .D0(n3753), .D1(n3754), .S(n3880), .Y(n230) );
  AOI22X1 U3382 ( .A(n552), .B(n3687), .C(n551), .D(n3911), .Y(n3753) );
  MUX2X1 U3383 ( .D0(n1121), .D1(n1122), .S(n3883), .Y(n3754) );
  NOR21XL U3384 ( .B(n3934), .A(A[970]), .Y(n726) );
  NOR21XL U3385 ( .B(n3934), .A(A[714]), .Y(n725) );
  MUX2IXL U3386 ( .D0(A[794]), .D1(A[282]), .S(n3965), .Y(n3755) );
  NOR21XL U3387 ( .B(n3934), .A(A[666]), .Y(n957) );
  MUX2IXL U3388 ( .D0(n3827), .D1(n3828), .S(n3648), .Y(n3815) );
  INVX1 U3389 ( .A(A[922]), .Y(n3828) );
  AOI22BX1 U3390 ( .B(n3758), .A(n3687), .D(n3759), .C(n3915), .Y(n3757) );
  AOI22XL U3391 ( .A(n3973), .B(A[430]), .C(n3957), .D(A[942]), .Y(n3758) );
  AOI22XL U3392 ( .A(n3973), .B(A[174]), .C(n3957), .D(A[686]), .Y(n3759) );
  AOI22XL U3393 ( .A(n3982), .B(A[435]), .C(n3991), .D(A[947]), .Y(n3761) );
  AOI22XL U3394 ( .A(n3975), .B(A[164]), .C(n3955), .D(A[676]), .Y(n3763) );
  AO22X1 U3395 ( .A(n808), .B(n3899), .C(n807), .D(n3916), .Y(n1756) );
  AOI22XL U3396 ( .A(n3977), .B(A[302]), .C(n3961), .D(A[814]), .Y(n3765) );
  AOI22XL U3397 ( .A(n3980), .B(A[511]), .C(n3956), .D(A[1023]), .Y(n3768) );
  AOI22XL U3398 ( .A(n3980), .B(A[255]), .C(n3952), .D(A[767]), .Y(n3769) );
  AOI22XL U3399 ( .A(n3976), .B(A[399]), .C(n3963), .D(A[911]), .Y(n3771) );
  AOI22XL U3400 ( .A(n3971), .B(A[143]), .C(n3963), .D(A[655]), .Y(n3772) );
  NAND21X1 U3401 ( .B(n3896), .A(n1256), .Y(n1657) );
  MUX2X1 U3402 ( .D0(A[125]), .D1(A[637]), .S(n3925), .Y(n3799) );
  NOR21XL U3403 ( .B(n3938), .A(A[586]), .Y(n1278) );
  AOI22XL U3404 ( .A(n3966), .B(A[510]), .C(n3992), .D(A[1022]), .Y(n3774) );
  INVX1 U3405 ( .A(n1650), .Y(n308) );
  NOR21XL U3406 ( .B(n3938), .A(A[587]), .Y(n1275) );
  INVX1 U3407 ( .A(n1655), .Y(n313) );
  NOR21XL U3408 ( .B(n3938), .A(A[592]), .Y(n1262) );
  INVX1 U3409 ( .A(n1662), .Y(n320) );
  NOR21XL U3410 ( .B(n3939), .A(A[599]), .Y(n1241) );
  INVX1 U3411 ( .A(n1658), .Y(n316) );
  NOR21XL U3412 ( .B(n3939), .A(A[595]), .Y(n1253) );
  INVX1 U3413 ( .A(n1661), .Y(n319) );
  NOR21XL U3414 ( .B(n3939), .A(A[598]), .Y(n1244) );
  NOR21XL U3415 ( .B(n3938), .A(A[593]), .Y(n1259) );
  MUX2IXL U3416 ( .D0(n3778), .D1(n3779), .S(n3892), .Y(n3777) );
  OR2XL U3417 ( .A(n3945), .B(A[232]), .Y(n3778) );
  MUX2XL U3418 ( .D0(A[488]), .D1(A[1000]), .S(n3648), .Y(n3779) );
  MUX2IXL U3419 ( .D0(A[494]), .D1(A[1006]), .S(n3930), .Y(n590) );
  MUX2IXL U3420 ( .D0(A[287]), .D1(A[799]), .S(n3989), .Y(n1472) );
  NOR21XL U3421 ( .B(n3942), .A(A[543]), .Y(n1471) );
  MUX2IXL U3422 ( .D0(A[472]), .D1(A[984]), .S(n3929), .Y(n678) );
  NOR21XL U3423 ( .B(n3963), .A(A[975]), .Y(n706) );
  NOR21XL U3424 ( .B(n3986), .A(A[719]), .Y(n705) );
  OR2XL U3425 ( .A(n3947), .B(A[360]), .Y(n3781) );
  MUX2XL U3426 ( .D0(n1237), .D1(n1238), .S(n3888), .Y(n3782) );
  NOR21XL U3427 ( .B(n3939), .A(A[601]), .Y(n1233) );
  NOR21XL U3428 ( .B(n3941), .A(A[603]), .Y(n1225) );
  MUX2IXL U3429 ( .D0(A[319]), .D1(A[831]), .S(n3927), .Y(n1312) );
  NOR21XL U3430 ( .B(n3939), .A(A[575]), .Y(n1311) );
  MUX2IXL U3431 ( .D0(A[318]), .D1(A[830]), .S(n3927), .Y(n1316) );
  NOR21XL U3432 ( .B(n3939), .A(A[574]), .Y(n1315) );
  MUX2X1 U3433 ( .D0(n1153), .D1(n1154), .S(n3882), .Y(n3783) );
  NOR21XL U3434 ( .B(n3937), .A(A[617]), .Y(n1169) );
  NOR21XL U3435 ( .B(n3941), .A(A[542]), .Y(n1475) );
  MUX2IXL U3436 ( .D0(A[286]), .D1(A[798]), .S(n3937), .Y(n1476) );
  NOR21XL U3437 ( .B(n3934), .A(A[669]), .Y(n945) );
  MUX2IXL U3438 ( .D0(A[415]), .D1(A[927]), .S(n3927), .Y(n938) );
  NOR21XL U3439 ( .B(n3990), .A(A[671]), .Y(n937) );
  MUX2IXL U3440 ( .D0(A[414]), .D1(A[926]), .S(n3927), .Y(n942) );
  NOR21XL U3441 ( .B(n3686), .A(A[670]), .Y(n941) );
  MUX2IXL U3442 ( .D0(A[271]), .D1(A[783]), .S(n3648), .Y(n1536) );
  NOR21XL U3443 ( .B(n3942), .A(A[527]), .Y(n1535) );
  MUX2IXL U3444 ( .D0(A[127]), .D1(A[639]), .S(n3925), .Y(n1081) );
  MUX2IXL U3445 ( .D0(A[479]), .D1(A[991]), .S(n3933), .Y(n650) );
  MUX2IXL U3446 ( .D0(A[478]), .D1(A[990]), .S(n3686), .Y(n654) );
  MUX2IXL U3447 ( .D0(A[473]), .D1(A[985]), .S(n3929), .Y(n674) );
  MUX2IXL U3448 ( .D0(A[475]), .D1(A[987]), .S(n3686), .Y(n666) );
  NOR21XL U3449 ( .B(n3934), .A(A[971]), .Y(n722) );
  NOR21XL U3450 ( .B(n3934), .A(A[715]), .Y(n721) );
  MUX2IXL U3451 ( .D0(A[489]), .D1(A[1001]), .S(n3648), .Y(n610) );
  MUX2IXL U3452 ( .D0(A[126]), .D1(A[638]), .S(n3925), .Y(n1085) );
  NOR2XL U3453 ( .A(n3965), .B(A[602]), .Y(n3788) );
  NOR2XL U3454 ( .A(n3965), .B(A[618]), .Y(n3789) );
  INVX1 U3455 ( .A(A[418]), .Y(n3821) );
  INVX1 U3456 ( .A(A[410]), .Y(n3827) );
  INVX1 U3457 ( .A(A[700]), .Y(n3804) );
  INVX1 U3458 ( .A(A[170]), .Y(n3807) );
  NOR21XL U3459 ( .B(n3940), .A(A[572]), .Y(n1323) );
  NOR21XL U3460 ( .B(n3940), .A(A[573]), .Y(n1319) );
  AOI22X1 U3461 ( .A(n558), .B(n3901), .C(n557), .D(n3915), .Y(n3791) );
  INVX1 U3462 ( .A(n1659), .Y(n317) );
  INVX1 U3463 ( .A(SH[8]), .Y(n3923) );
  INVXL U3464 ( .A(n3991), .Y(n3972) );
  AOI22XL U3465 ( .A(n3980), .B(A[509]), .C(n3956), .D(A[1021]), .Y(n3795) );
  OA22X1 U3466 ( .A(n3796), .B(n3901), .C(n3823), .D(n3915), .Y(n3830) );
  AOI22X1 U3467 ( .A(n3972), .B(A[242]), .C(n3954), .D(A[754]), .Y(n3796) );
  INVXL U3468 ( .A(n3918), .Y(n3914) );
  MUX2IX1 U3469 ( .D0(n3810), .D1(n3799), .S(n3798), .Y(n3809) );
  INVX1 U3470 ( .A(n3923), .Y(n3919) );
  INVXL U3471 ( .A(n3923), .Y(n3920) );
  INVXL U3472 ( .A(n3922), .Y(n3921) );
  INVXL U3473 ( .A(n3919), .Y(n3911) );
  INVXL U3474 ( .A(n3919), .Y(n3910) );
  INVX1 U3475 ( .A(n3812), .Y(n3903) );
  INVX1 U3476 ( .A(n3812), .Y(n3904) );
  INVXL U3477 ( .A(SH[9]), .Y(n3997) );
  INVXL U3478 ( .A(n3920), .Y(n3909) );
  MUX2IX1 U3479 ( .D0(n79), .D1(n111), .S(n3855), .Y(n47) );
  MUX2IX1 U3480 ( .D0(n3703), .D1(n3676), .S(n3878), .Y(n127) );
  MUX2IX1 U3481 ( .D0(A[636]), .D1(A[124]), .S(n3976), .Y(n1093) );
  MUX2X1 U3482 ( .D0(A[284]), .D1(A[796]), .S(n3990), .Y(n3832) );
  INVX2 U3483 ( .A(n3993), .Y(n3966) );
  MUX2IX1 U3484 ( .D0(A[916]), .D1(A[404]), .S(n3976), .Y(n982) );
  AOI22X1 U3485 ( .A(n904), .B(n3898), .C(n903), .D(n3909), .Y(n3806) );
  OAI22AXL U3486 ( .D(A[682]), .C(n3971), .A(n3988), .B(n3807), .Y(n873) );
  INVXL U3487 ( .A(n3991), .Y(n3971) );
  AOI22X1 U3488 ( .A(n3978), .B(A[301]), .C(n3961), .D(A[813]), .Y(n3847) );
  INVX1 U3489 ( .A(n3992), .Y(n3974) );
  INVX1 U3490 ( .A(n3966), .Y(n3942) );
  EORX1 U3491 ( .A(n1407), .B(n3917), .C(n3811), .D(n3915), .Y(n3834) );
  AOI22X1 U3492 ( .A(n3969), .B(A[298]), .C(n3956), .D(A[810]), .Y(n3811) );
  INVX1 U3493 ( .A(n3998), .Y(n3987) );
  OAI22AXL U3494 ( .D(A[685]), .C(n3971), .A(n3960), .B(n3813), .Y(n855) );
  MUX2X1 U3495 ( .D0(A[826]), .D1(A[314]), .S(n3965), .Y(n3820) );
  AOI22X1 U3496 ( .A(n3974), .B(A[426]), .C(n3957), .D(A[938]), .Y(n3814) );
  NOR2XL U3497 ( .A(n3965), .B(A[538]), .Y(n1491) );
  MUX2IX1 U3498 ( .D0(A[788]), .D1(A[276]), .S(n3976), .Y(n1516) );
  MUX2AX2 U3499 ( .D0(n3815), .D1(n957), .S(n3916), .Y(n3837) );
  MUX2X1 U3500 ( .D0(A[818]), .D1(A[306]), .S(n3965), .Y(n3826) );
  NAND2X1 U3501 ( .A(n3802), .B(n3879), .Y(n115) );
  OA22X1 U3502 ( .A(n3818), .B(n3817), .C(n3819), .D(n3897), .Y(n3816) );
  AOI22XL U3503 ( .A(n3970), .B(A[290]), .C(n3835), .D(A[802]), .Y(n3818) );
  AOI22XL U3504 ( .A(n3851), .B(A[34]), .C(n3835), .D(A[546]), .Y(n3819) );
  MUX2AX2 U3505 ( .D0(n3820), .D1(n1331), .S(n3917), .Y(n3836) );
  EORX1 U3506 ( .A(n1034), .B(n3898), .C(n3822), .D(n3901), .Y(n3845) );
  AOI22X1 U3507 ( .A(n3977), .B(A[138]), .C(n3962), .D(A[650]), .Y(n3822) );
  AOI22X1 U3508 ( .A(n3972), .B(A[498]), .C(n3954), .D(A[1010]), .Y(n3823) );
  AOI22AX1 U3509 ( .A(n825), .B(n3915), .D(n3912), .C(n826), .Y(n3846) );
  AOI22X1 U3510 ( .A(n3971), .B(A[506]), .C(n3988), .D(A[1018]), .Y(n3824) );
  MUX2AX2 U3511 ( .D0(n3826), .D1(n1363), .S(n3912), .Y(n3841) );
  INVXL U3512 ( .A(n3919), .Y(n3915) );
  INVXL U3513 ( .A(n3996), .Y(n3992) );
  INVXL U3514 ( .A(n3998), .Y(n3835) );
  MUX2IXL U3515 ( .D0(n3746), .D1(n3677), .S(n3878), .Y(n124) );
  MUX2IX1 U3516 ( .D0(n174), .D1(n238), .S(n3859), .Y(n110) );
  AOI22X1 U3517 ( .A(n1022), .B(n3897), .C(n1021), .D(n3912), .Y(n3833) );
  AO22AX1 U3518 ( .A(n3960), .B(A[556]), .C(A[44]), .D(n3960), .Y(n1395) );
  INVX1 U3519 ( .A(n3998), .Y(n3995) );
  INVXL U3520 ( .A(n3986), .Y(n3983) );
  AO22X1 U3521 ( .A(n3981), .B(A[180]), .C(n3835), .D(A[692]), .Y(n813) );
  BUFX1 U3522 ( .A(n3996), .Y(n3851) );
  MUX2IXL U3523 ( .D0(A[994]), .D1(A[482]), .S(n3964), .Y(n638) );
  INVXL U3524 ( .A(SH[8]), .Y(n3924) );
  MUX2IXL U3525 ( .D0(A[786]), .D1(A[274]), .S(n3964), .Y(n1524) );
  MUX2X2 U3526 ( .D0(n1166), .D1(n3789), .S(n3917), .Y(n3842) );
  INVX1 U3527 ( .A(n3997), .Y(n3989) );
  MUX2X2 U3528 ( .D0(n1555), .D1(n1556), .S(n3891), .Y(n3843) );
  OA22X1 U3529 ( .A(n3849), .B(n3912), .C(n3850), .D(n3919), .Y(n3848) );
  INVXL U3530 ( .A(n3996), .Y(n3991) );
  MUX2IX1 U3531 ( .D0(n6), .D1(n14), .S(SH[3]), .Y(B[5]) );
  MUX2IX1 U3532 ( .D0(n3809), .D1(n3794), .S(n3867), .Y(n238) );
endmodule


module regbank_a0_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module regbank_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regbank_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_49 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10776;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_49 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10776), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10776), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10776), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10776), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10776), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10776), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10776), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10776), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10776), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_50 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10794;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_50 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10794), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10794), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10794), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10794), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10794), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10794), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10794), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10794), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10794), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_51 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10812;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_51 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10812), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10812), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10812), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10812), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10812), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10812), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10812), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10812), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10812), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_52 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10830;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_52 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10830), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10830), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10830), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10830), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10830), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10830), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10830), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10830), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10830), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_53 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10848;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_53 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10848), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10848), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10848), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10848), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10848), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10848), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10848), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10848), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10848), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_0000001f ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10866;

  SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10866), .TE(test_se) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10866), .XS(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10866), .XS(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10866), .XS(arstz), .Q(rdat[1]) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10866), .XS(arstz), .Q(rdat[0]) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10866), .XS(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10866), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10866), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10866), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000004 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10884;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10884), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10884), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10884), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10884), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10884), .XR(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10884), .XS(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10884), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10884), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10884), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_4_00000004 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10902;

  SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10902), .TE(test_se) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10902), .XS(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10902), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10902), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10902), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_54 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10920;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_54 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10920), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10920), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10920), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10920), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10920), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10920), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10920), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10920), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10920), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_55 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10938;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_55 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10938), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10938), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10938), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10938), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10938), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10938), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10938), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10938), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10938), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_55 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_2 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_2 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[2]), .Y(n11) );
  INVX1 U4 ( .A(set2[4]), .Y(n1) );
  INVX1 U5 ( .A(set2[5]), .Y(n2) );
  INVX1 U6 ( .A(set2[7]), .Y(n12) );
  INVX1 U7 ( .A(set2[0]), .Y(n13) );
  INVX1 U8 ( .A(set2[1]), .Y(n14) );
  INVX1 U9 ( .A(set2[3]), .Y(n15) );
  NAND3X1 U10 ( .A(n16), .B(n12), .C(n2), .Y(n21) );
  AOI211X1 U11 ( .C(n1), .D(n10), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U12 ( .A(rdat[4]), .Y(n10) );
  AOI211X1 U13 ( .C(n11), .D(n9), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U14 ( .A(rdat[2]), .Y(n9) );
  AOI211X1 U15 ( .C(n2), .D(n8), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U16 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U17 ( .C(n13), .D(n7), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U18 ( .A(rdat[0]), .Y(n7) );
  AOI211X1 U19 ( .C(n14), .D(n6), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U20 ( .A(rdat[1]), .Y(n6) );
  AOI211X1 U21 ( .C(n16), .D(n4), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U22 ( .A(rdat[6]), .Y(n4) );
  AOI211X1 U23 ( .C(n12), .D(n3), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U24 ( .A(rdat[7]), .Y(n3) );
  AOI211X1 U25 ( .C(n15), .D(n5), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U26 ( .A(rdat[3]), .Y(n5) );
  NAND4X1 U27 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U28 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U29 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U30 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR2X1 U31 ( .A(rdat[3]), .B(n15), .Y(irq[3]) );
  NOR2X1 U32 ( .A(rdat[2]), .B(n11), .Y(irq[2]) );
  NOR2X1 U33 ( .A(rdat[5]), .B(n2), .Y(irq[5]) );
  NOR2X1 U34 ( .A(rdat[4]), .B(n1), .Y(irq[4]) );
  NOR2X1 U35 ( .A(rdat[0]), .B(n13), .Y(irq[0]) );
  NOR2X1 U36 ( .A(rdat[7]), .B(n12), .Y(irq[7]) );
  NOR2X1 U37 ( .A(rdat[1]), .B(n14), .Y(irq[1]) );
  NOR2X1 U38 ( .A(rdat[6]), .B(n16), .Y(irq[6]) );
  INVX1 U39 ( .A(set2[6]), .Y(n16) );
endmodule


module glreg_WIDTH8_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10956;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10956), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10956), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10956), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10956), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10956), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10956), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10956), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10956), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10956), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_8 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR3XL U7 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_9 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR3XL U7 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_10 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR3XL U7 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n2), .Y(n8) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_11 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_12 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_13 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n4, n5, n6, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n5), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n6), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n4), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n4) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n6) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n5) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_1_, db_cnt_0_, N13, N14, N15, N16, net10974, n7, n5,
         n6, n1, n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_0 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net10974), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N16), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net10974), .XR(rstz), .Q(test_so) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N15), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net10974), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N14), .SIN(o_dbc), .SMC(test_se), .C(net10974), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n7), .SIN(d_org_0_), .SMC(test_se), .C(net10974), 
        .XR(rstz), .Q(o_dbc) );
  OAI22X1 U3 ( .A(n1), .B(n3), .C(n6), .D(n2), .Y(N16) );
  INVX1 U4 ( .A(N14), .Y(n3) );
  NAND4X1 U5 ( .A(n5), .B(n4), .C(n2), .D(n1), .Y(N13) );
  XNOR2XL U6 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  NOR4XL U7 ( .A(n1), .B(n4), .C(n5), .D(db_cnt_1_), .Y(o_chg) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n4) );
  AO22AXL U9 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  INVX1 U10 ( .A(test_so), .Y(n1) );
  NAND31X1 U11 ( .C(n5), .A(n1), .B(db_cnt_0_), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt_0_), .Y(N14) );
  OAI22X1 U13 ( .A(n2), .B(n3), .C(db_cnt_1_), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt_1_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_1_, db_cnt_0_, N13, N14, N15, N16, net10992, n7, n5,
         n6, n1, n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_1 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net10992), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N16), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net10992), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N15), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net10992), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N14), .SIN(o_dbc), .SMC(test_se), .C(net10992), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n7), .SIN(d_org_0_), .SMC(test_se), .C(net10992), 
        .XR(rstz), .Q(o_dbc) );
  OAI22X1 U3 ( .A(n1), .B(n4), .C(n6), .D(n2), .Y(N16) );
  INVX1 U4 ( .A(N14), .Y(n4) );
  NAND4X1 U5 ( .A(n5), .B(n3), .C(n2), .D(n1), .Y(N13) );
  XNOR2XL U6 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  NOR4XL U7 ( .A(n1), .B(n3), .C(n5), .D(db_cnt_1_), .Y(o_chg) );
  INVX1 U8 ( .A(test_so), .Y(n1) );
  INVX1 U9 ( .A(db_cnt_0_), .Y(n3) );
  AO22AXL U10 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  NAND31X1 U11 ( .C(n5), .A(n1), .B(db_cnt_0_), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt_0_), .Y(N14) );
  OAI22X1 U13 ( .A(n2), .B(n4), .C(db_cnt_1_), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt_1_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_1_, db_cnt_0_, N13, N14, N15, N16, net11010, n7, n5,
         n6, n1, n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_2 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net11010), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N16), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11010), .XR(rstz), .Q(test_so) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N15), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11010), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N14), .SIN(o_dbc), .SMC(test_se), .C(net11010), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n7), .SIN(d_org_0_), .SMC(test_se), .C(net11010), 
        .XR(rstz), .Q(o_dbc) );
  NOR4XL U3 ( .A(n1), .B(n3), .C(n5), .D(db_cnt_1_), .Y(o_chg) );
  OAI22X1 U4 ( .A(n1), .B(n4), .C(n6), .D(n2), .Y(N16) );
  INVX1 U5 ( .A(N14), .Y(n4) );
  NAND4X1 U6 ( .A(n5), .B(n3), .C(n2), .D(n1), .Y(N13) );
  XNOR2XL U7 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n3) );
  AO22AXL U9 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  INVX1 U10 ( .A(test_so), .Y(n1) );
  NAND31X1 U11 ( .C(n5), .A(n1), .B(db_cnt_0_), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt_0_), .Y(N14) );
  OAI22X1 U13 ( .A(n2), .B(n4), .C(db_cnt_1_), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt_1_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_1_, db_cnt_0_, N13, N14, N15, N16, net11028, n7, n5,
         n6, n1, n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_3 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net11028), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N16), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11028), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N15), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11028), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N14), .SIN(o_dbc), .SMC(test_se), .C(net11028), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n7), .SIN(d_org_0_), .SMC(test_se), .C(net11028), 
        .XR(rstz), .Q(o_dbc) );
  NOR4XL U3 ( .A(n1), .B(n4), .C(n5), .D(db_cnt_1_), .Y(o_chg) );
  OAI22X1 U4 ( .A(n1), .B(n3), .C(n6), .D(n2), .Y(N16) );
  INVX1 U5 ( .A(N14), .Y(n3) );
  NAND4X1 U6 ( .A(n5), .B(n4), .C(n2), .D(n1), .Y(N13) );
  XNOR2XL U7 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  INVX1 U8 ( .A(test_so), .Y(n1) );
  INVX1 U9 ( .A(db_cnt_0_), .Y(n4) );
  AO22AXL U10 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  NAND31X1 U11 ( .C(n5), .A(n1), .B(db_cnt_0_), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt_0_), .Y(N14) );
  OAI22X1 U13 ( .A(n2), .B(n3), .C(db_cnt_1_), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt_1_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_4 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_1_, db_cnt_0_, N13, N14, N15, N16, net11046, n7, n5,
         n6, n1, n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_4 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net11046), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N16), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11046), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N15), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11046), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N14), .SIN(o_dbc), .SMC(test_se), .C(net11046), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n7), .SIN(d_org_0_), .SMC(test_se), .C(net11046), 
        .XR(rstz), .Q(o_dbc) );
  OAI22X1 U3 ( .A(n1), .B(n3), .C(n6), .D(n2), .Y(N16) );
  INVX1 U4 ( .A(N14), .Y(n3) );
  NAND4X1 U5 ( .A(n5), .B(n4), .C(n2), .D(n1), .Y(N13) );
  XNOR2XL U6 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  NOR4XL U7 ( .A(n1), .B(n4), .C(n5), .D(db_cnt_1_), .Y(o_chg) );
  INVX1 U8 ( .A(test_so), .Y(n1) );
  INVX1 U9 ( .A(db_cnt_0_), .Y(n4) );
  AO22AXL U10 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  NAND31X1 U11 ( .C(n5), .A(n1), .B(db_cnt_0_), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt_0_), .Y(N14) );
  OAI22X1 U13 ( .A(n2), .B(n3), .C(db_cnt_1_), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt_1_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N16, N17, N18, N19, N20,
         net11064, n12, n3, n4, n5, n6, n7, n8, n9, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_2 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net11064), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N20), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11064), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N18), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11064), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N17), .SIN(o_dbc), .SMC(test_se), .C(net11064), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N19), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11064), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n12), .SIN(d_org_0_), .SMC(test_se), .C(net11064), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n6), .Y(n1) );
  NOR2X1 U4 ( .A(n3), .B(n4), .Y(o_chg) );
  NOR21XL U5 ( .B(n3), .A(n4), .Y(n6) );
  XNOR2XL U6 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  NAND4X1 U7 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(db_cnt_0_), .Y(n3) );
  OAI22X1 U8 ( .A(db_cnt_2_), .B(n5), .C(n7), .D(n2), .Y(N19) );
  AOI21BBXL U9 ( .B(n1), .C(db_cnt_1_), .A(N17), .Y(n7) );
  AO22AXL U10 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR2X1 U11 ( .A(n1), .B(db_cnt_0_), .Y(N17) );
  NAND3X1 U12 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(n6), .Y(n5) );
  ENOX1 U13 ( .A(n2), .B(n5), .C(test_so), .D(n6), .Y(N20) );
  NOR2X1 U14 ( .A(n8), .B(n1), .Y(N18) );
  XNOR2XL U15 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n8) );
  NAND31X1 U16 ( .C(db_cnt_0_), .A(n4), .B(n9), .Y(N16) );
  NOR3XL U17 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n9) );
  INVX1 U18 ( .A(db_cnt_2_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N19,
         net11082, n13, n6, n7, n8, n9, n10, n11, n12, n14, n1, n2, n3, n4, n5
;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11082), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11082), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11082), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11082), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(n1), .SIN(db_cnt_1_), .SMC(test_se), .C(net11082), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11082), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n2) );
  NOR2X1 U4 ( .A(n2), .B(n11), .Y(n9) );
  NOR21XL U5 ( .B(n6), .A(n7), .Y(n8) );
  NOR2X1 U6 ( .A(n3), .B(n4), .Y(n11) );
  AOI211X1 U7 ( .C(n3), .D(n4), .A(n2), .B(n11), .Y(N17) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  GEN2XL U9 ( .D(n8), .E(n5), .C(n9), .B(test_so), .A(n10), .Y(N19) );
  NOR42XL U10 ( .C(n11), .D(db_cnt_2_), .A(n2), .B(test_so), .Y(n10) );
  INVX1 U11 ( .A(n12), .Y(n1) );
  AOI32X1 U12 ( .A(n11), .B(n5), .C(n8), .D(db_cnt_2_), .E(n9), .Y(n12) );
  AO22AXL U13 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U14 ( .A(n6), .B(n7), .Y(o_chg) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  NAND4X1 U16 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(n3), .Y(n6) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n5) );
  INVX1 U18 ( .A(db_cnt_1_), .Y(n4) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n2), .Y(N16) );
  NAND3X1 U20 ( .A(n7), .B(n3), .C(n14), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N19,
         net11100, n13, n6, n7, n8, n9, n10, n11, n12, n14, n1, n2, n3, n4, n5
;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11100), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11100), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11100), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11100), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(n1), .SIN(db_cnt_1_), .SMC(test_se), .C(net11100), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11100), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n2) );
  NOR2X1 U4 ( .A(n2), .B(n11), .Y(n9) );
  NOR21XL U5 ( .B(n6), .A(n7), .Y(n8) );
  NOR2X1 U6 ( .A(n3), .B(n4), .Y(n11) );
  AOI211X1 U7 ( .C(n3), .D(n4), .A(n2), .B(n11), .Y(N17) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  GEN2XL U9 ( .D(n8), .E(n5), .C(n9), .B(test_so), .A(n10), .Y(N19) );
  NOR42XL U10 ( .C(n11), .D(db_cnt_2_), .A(n2), .B(test_so), .Y(n10) );
  INVX1 U11 ( .A(n12), .Y(n1) );
  AOI32X1 U12 ( .A(n11), .B(n5), .C(n8), .D(db_cnt_2_), .E(n9), .Y(n12) );
  AO22AXL U13 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U14 ( .A(n6), .B(n7), .Y(o_chg) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  NAND4X1 U16 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(n3), .Y(n6) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n5) );
  INVX1 U18 ( .A(db_cnt_1_), .Y(n4) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n2), .Y(N16) );
  NAND3X1 U20 ( .A(n7), .B(n3), .C(n14), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N19,
         net11118, n13, n6, n7, n8, n9, n10, n11, n12, n14, n1, n2, n3, n4, n5
;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11118), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11118), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11118), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11118), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(n1), .SIN(db_cnt_1_), .SMC(test_se), .C(net11118), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11118), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n2) );
  NOR2X1 U4 ( .A(n2), .B(n11), .Y(n9) );
  NOR21XL U5 ( .B(n6), .A(n7), .Y(n8) );
  NOR2X1 U6 ( .A(n3), .B(n4), .Y(n11) );
  AOI211X1 U7 ( .C(n3), .D(n4), .A(n2), .B(n11), .Y(N17) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  GEN2XL U9 ( .D(n8), .E(n5), .C(n9), .B(test_so), .A(n10), .Y(N19) );
  NOR42XL U10 ( .C(n11), .D(db_cnt_2_), .A(n2), .B(test_so), .Y(n10) );
  INVX1 U11 ( .A(n12), .Y(n1) );
  AOI32X1 U12 ( .A(n11), .B(n5), .C(n8), .D(db_cnt_2_), .E(n9), .Y(n12) );
  AO22AXL U13 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U14 ( .A(n6), .B(n7), .Y(o_chg) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  NAND4X1 U16 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(n3), .Y(n6) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n5) );
  INVX1 U18 ( .A(db_cnt_1_), .Y(n4) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n2), .Y(N16) );
  NAND3X1 U20 ( .A(n7), .B(n3), .C(n14), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000028 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11136;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11136), .TE(test_se) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11136), .XS(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11136), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11136), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11136), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11136), .XR(arstz), .Q(rdat[1]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11136), .XS(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11136), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11136), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_56 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11154;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_56 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11154), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11154), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11154), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11154), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11154), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11154), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11154), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11154), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11154), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_56 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_57 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11172;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_57 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11172), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11172), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11172), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11172), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11172), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11172), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11172), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11172), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11172), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_57 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_58 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11190;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_58 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11190), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11190), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11190), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11190), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11190), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11190), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11190), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11190), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11190), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_58 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_59 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11208;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_59 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11208), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11208), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11208), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11208), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11208), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11208), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11208), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11208), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11208), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_59 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_60 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11226;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_60 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11226), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11226), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11226), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11226), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11226), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11226), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11226), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11226), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11226), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_60 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_61 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11244;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_61 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11244), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11244), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11244), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11244), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11244), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11244), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11244), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11244), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11244), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_61 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_62 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11262;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_62 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11262), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11262), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11262), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11262), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11262), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11262), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11262), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11262), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11262), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_62 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_63 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11280;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_63 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11280), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11280), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11280), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11280), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11280), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11280), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11280), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11280), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11280), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_63 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11298;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11298), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11298), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11298), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11298), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11298), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_64 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11316;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_64 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11316), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11316), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11316), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11316), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11316), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11316), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11316), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11316), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11316), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_64 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_3 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_3 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[0]), .Y(n13) );
  INVX1 U4 ( .A(set2[1]), .Y(n12) );
  INVX1 U5 ( .A(set2[2]), .Y(n15) );
  INVX1 U6 ( .A(set2[3]), .Y(n11) );
  INVX1 U7 ( .A(set2[4]), .Y(n16) );
  NAND3X1 U8 ( .A(n14), .B(n9), .C(n10), .Y(n21) );
  AOI211X1 U9 ( .C(n16), .D(n8), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U10 ( .A(rdat[4]), .Y(n8) );
  AOI211X1 U11 ( .C(n13), .D(n7), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U12 ( .A(rdat[0]), .Y(n7) );
  AOI211X1 U13 ( .C(n12), .D(n6), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U14 ( .A(rdat[1]), .Y(n6) );
  AOI211X1 U15 ( .C(n15), .D(n5), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U16 ( .A(rdat[2]), .Y(n5) );
  AOI211X1 U17 ( .C(n10), .D(n3), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U18 ( .A(rdat[5]), .Y(n3) );
  AOI211X1 U19 ( .C(n14), .D(n2), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U20 ( .A(rdat[6]), .Y(n2) );
  AOI211X1 U21 ( .C(n9), .D(n1), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U22 ( .A(rdat[7]), .Y(n1) );
  AOI211X1 U23 ( .C(n11), .D(n4), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U24 ( .A(rdat[3]), .Y(n4) );
  NAND4X1 U25 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U26 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U27 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U28 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR2X1 U29 ( .A(rdat[0]), .B(n13), .Y(irq[0]) );
  NOR2X1 U30 ( .A(rdat[1]), .B(n12), .Y(irq[1]) );
  NOR2X1 U31 ( .A(rdat[2]), .B(n15), .Y(irq[2]) );
  NOR2X1 U32 ( .A(rdat[3]), .B(n11), .Y(irq[3]) );
  INVX1 U33 ( .A(set2[6]), .Y(n14) );
  INVX1 U34 ( .A(set2[7]), .Y(n9) );
  INVX1 U35 ( .A(set2[5]), .Y(n10) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n16), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n14), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[5]), .B(n10), .Y(irq[5]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n9), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11334;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11334), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11334), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11334), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11334), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11334), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11334), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11334), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11334), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11334), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_65 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11352;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_65 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11352), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11352), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11352), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11352), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11352), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11352), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11352), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11352), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11352), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_65 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_66 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11370;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_66 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11370), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11370), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11370), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11370), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11370), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11370), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11370), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11370), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11370), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_66 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000032 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11388;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11388), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11388), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11388), .XR(arstz), .Q(rdat[7]) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11388), .XS(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11388), .XR(arstz), .Q(rdat[2]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11388), .XS(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11388), .XR(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11388), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11388), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000098 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11406;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11406), .TE(test_se) );
  SDFFSQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11406), .XS(arstz), .Q(rdat[7]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11406), .XS(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11406), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11406), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11406), .XR(arstz), .Q(rdat[1]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11406), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11406), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11406), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_000000f0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11424;

  SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11424), .TE(test_se) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11424), .XS(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11424), .XS(arstz), .Q(rdat[7]) );
  SDFFSQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11424), .XS(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11424), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11424), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11424), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11424), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11424), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH1_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH1_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH2_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2, n3, n1;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(n3), .SIN(rdat[0]), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[1]) );
  INVX1 U2 ( .A(we), .Y(n1) );
  AO22XL U3 ( .A(we), .B(wdat[1]), .C(rdat[1]), .D(n1), .Y(n3) );
  AO22XL U4 ( .A(wdat[0]), .B(we), .C(rdat[0]), .D(n1), .Y(n2) );
endmodule


module glreg_WIDTH3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [2:0] wdat;
  output [2:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11442;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11442), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11442), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11442), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11442), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000011 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11460;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11460), .TE(test_se) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11460), .XS(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11460), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11460), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11460), .XR(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11460), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11460), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11460), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11460), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000001 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11478;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11478), .TE(test_se) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11478), .XS(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11478), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11478), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11478), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11478), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11478), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11478), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11478), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_67 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11496;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_67 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11496), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11496), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11496), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11496), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11496), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11496), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11496), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11496), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11496), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_67 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_4 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_4 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[0]), .Y(n13) );
  INVX1 U4 ( .A(set2[7]), .Y(n12) );
  NAND3X1 U5 ( .A(n11), .B(n12), .C(n10), .Y(n21) );
  INVX1 U6 ( .A(set2[3]), .Y(n14) );
  INVX1 U7 ( .A(set2[1]), .Y(n16) );
  INVX1 U8 ( .A(set2[5]), .Y(n10) );
  INVX1 U9 ( .A(set2[4]), .Y(n9) );
  INVX1 U10 ( .A(set2[6]), .Y(n11) );
  INVX1 U11 ( .A(set2[2]), .Y(n15) );
  NAND4X1 U12 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U13 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U14 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U15 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U16 ( .C(n10), .D(n1), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U17 ( .A(rdat[5]), .Y(n1) );
  AOI211X1 U18 ( .C(n12), .D(n8), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U19 ( .A(rdat[7]), .Y(n8) );
  AOI211X1 U20 ( .C(n9), .D(n7), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U21 ( .A(rdat[4]), .Y(n7) );
  AOI211X1 U22 ( .C(n11), .D(n6), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U23 ( .A(rdat[6]), .Y(n6) );
  AOI211X1 U24 ( .C(n13), .D(n5), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U25 ( .A(rdat[0]), .Y(n5) );
  AOI211X1 U26 ( .C(n15), .D(n4), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U27 ( .A(rdat[2]), .Y(n4) );
  AOI211X1 U28 ( .C(n16), .D(n3), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U29 ( .A(rdat[1]), .Y(n3) );
  AOI211X1 U30 ( .C(n14), .D(n2), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U31 ( .A(rdat[3]), .Y(n2) );
  NOR2X1 U32 ( .A(rdat[7]), .B(n12), .Y(irq[7]) );
  NOR2X1 U33 ( .A(rdat[6]), .B(n11), .Y(irq[6]) );
  NOR2X1 U34 ( .A(rdat[3]), .B(n14), .Y(irq[3]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n15), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n13), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[4]), .B(n9), .Y(irq[4]) );
  NOR2X1 U38 ( .A(rdat[1]), .B(n16), .Y(irq[1]) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n10), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11514;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11514), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11514), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11514), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11514), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11514), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11514), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11514), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11514), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11514), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_68 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11532;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_68 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11532), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11532), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11532), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11532), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11532), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11532), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11532), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11532), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11532), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_68 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_7_70 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11550;

  SNPS_CLOCK_GATE_HIGH_glreg_7_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11550), .TE(test_se) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11550), .XS(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11550), .XS(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11550), .XS(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11550), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11550), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11550), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11550), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_7_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_1_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n1;

  SDFFSQX1 mem_reg_0_ ( .D(n1), .SIN(test_si), .SMC(test_se), .C(clk), .XS(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n1) );
endmodule


module glreg_WIDTH1_6 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_6_00000018 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11568;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11568), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11568), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11568), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11568), .XR(arstz), .Q(rdat[2]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11568), .XS(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11568), .XR(arstz), .Q(rdat[1]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11568), .XS(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_69 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11586;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_69 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11586), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11586), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11586), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11586), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11586), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11586), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11586), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11586), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11586), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_69 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_70 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11604;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11604), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11604), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11604), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11604), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11604), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11604), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11604), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11604), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11604), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_71 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11622;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_71 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11622), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11622), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11622), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11622), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11622), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11622), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11622), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11622), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11622), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_71 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_72 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11640;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_72 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11640), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11640), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11640), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11640), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11640), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11640), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11640), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11640), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11640), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_72 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_73 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11658;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_73 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11658), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11658), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11658), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11658), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11658), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11658), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11658), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11658), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11658), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_73 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11676;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11676), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11676), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11676), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11676), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11676), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11676), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_74 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11694;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_74 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11694), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11694), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11694), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11694), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11694), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11694), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11694), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11694), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11694), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_74 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_75 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11712;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_75 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11712), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11712), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11712), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11712), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11712), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11712), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11712), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11712), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11712), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_75 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_76 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11730;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_76 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11730), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11730), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11730), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11730), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11730), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11730), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11730), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11730), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11730), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_76 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_77 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11748;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_77 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11748), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11748), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11748), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11748), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11748), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11748), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11748), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11748), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11748), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_77 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_5 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_5 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[1]), .Y(n14) );
  INVX1 U3 ( .A(set2[4]), .Y(n2) );
  NOR3XL U4 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NAND3X1 U5 ( .A(n16), .B(n1), .C(n3), .Y(n21) );
  NAND4X1 U6 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U7 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U8 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  NOR4XL U9 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  INVX1 U10 ( .A(set2[3]), .Y(n4) );
  INVX1 U11 ( .A(set2[0]), .Y(n15) );
  INVX1 U12 ( .A(set2[2]), .Y(n5) );
  INVX1 U13 ( .A(set2[5]), .Y(n3) );
  NOR2X1 U14 ( .A(rdat[4]), .B(n2), .Y(irq[4]) );
  NOR2X1 U15 ( .A(rdat[5]), .B(n3), .Y(irq[5]) );
  AOI211X1 U16 ( .C(n2), .D(n12), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U17 ( .A(rdat[4]), .Y(n12) );
  AOI211X1 U18 ( .C(n3), .D(n8), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U19 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U20 ( .C(n14), .D(n13), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U21 ( .A(rdat[1]), .Y(n13) );
  AOI211X1 U22 ( .C(n4), .D(n11), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U23 ( .A(rdat[3]), .Y(n11) );
  AOI211X1 U24 ( .C(n15), .D(n10), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U25 ( .A(rdat[0]), .Y(n10) );
  AOI211X1 U26 ( .C(n5), .D(n9), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U27 ( .A(rdat[2]), .Y(n9) );
  AOI211X1 U28 ( .C(n16), .D(n7), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U29 ( .A(rdat[6]), .Y(n7) );
  AOI211X1 U30 ( .C(n1), .D(n6), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U31 ( .A(rdat[7]), .Y(n6) );
  NOR2X1 U32 ( .A(rdat[2]), .B(n5), .Y(irq[2]) );
  NOR2X1 U33 ( .A(rdat[3]), .B(n4), .Y(irq[3]) );
  INVX1 U34 ( .A(set2[6]), .Y(n16) );
  NOR2X1 U35 ( .A(rdat[6]), .B(n16), .Y(irq[6]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n15), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[1]), .B(n14), .Y(irq[1]) );
  INVX1 U38 ( .A(set2[7]), .Y(n1) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n1), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11766;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11766), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11766), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11766), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11766), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11766), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11766), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11766), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11766), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11766), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_6 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_6 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[3]), .Y(n4) );
  INVX1 U3 ( .A(set2[7]), .Y(n2) );
  INVX1 U4 ( .A(set2[6]), .Y(n5) );
  NOR4XL U5 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NAND4X1 U6 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR3XL U7 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U8 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U9 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U10 ( .A(set2[1]), .Y(n1) );
  INVX1 U11 ( .A(set2[2]), .Y(n3) );
  NAND3X1 U12 ( .A(n5), .B(n2), .C(n16), .Y(n21) );
  INVX1 U13 ( .A(set2[4]), .Y(n6) );
  INVX1 U14 ( .A(set2[0]), .Y(n15) );
  AOI211X1 U15 ( .C(n15), .D(n14), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U16 ( .A(rdat[0]), .Y(n14) );
  AOI211X1 U17 ( .C(n1), .D(n13), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U18 ( .A(rdat[1]), .Y(n13) );
  AOI211X1 U19 ( .C(n3), .D(n12), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U20 ( .A(rdat[2]), .Y(n12) );
  AOI211X1 U21 ( .C(n6), .D(n10), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U22 ( .A(rdat[4]), .Y(n10) );
  AOI211X1 U23 ( .C(n16), .D(n9), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U24 ( .A(rdat[5]), .Y(n9) );
  AOI211X1 U25 ( .C(n5), .D(n8), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U26 ( .A(rdat[6]), .Y(n8) );
  AOI211X1 U27 ( .C(n2), .D(n7), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U28 ( .A(rdat[7]), .Y(n7) );
  AOI211X1 U29 ( .C(n4), .D(n11), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U30 ( .A(rdat[3]), .Y(n11) );
  NOR2X1 U31 ( .A(rdat[0]), .B(n15), .Y(irq[0]) );
  NOR2X1 U32 ( .A(rdat[1]), .B(n1), .Y(irq[1]) );
  NOR2X1 U33 ( .A(rdat[6]), .B(n5), .Y(irq[6]) );
  NOR2X1 U34 ( .A(rdat[7]), .B(n2), .Y(irq[7]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n3), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[3]), .B(n4), .Y(irq[3]) );
  NOR2X1 U37 ( .A(rdat[4]), .B(n6), .Y(irq[4]) );
  INVX1 U38 ( .A(set2[5]), .Y(n16) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_6 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11784;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11784), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11784), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11784), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11784), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11784), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11784), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11784), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11784), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11784), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_78 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11802;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_78 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11802), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11802), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11802), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11802), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11802), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11802), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11802), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11802), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11802), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_78 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_79 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11820;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_79 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11820), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11820), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11820), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11820), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11820), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11820), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11820), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11820), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11820), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_79 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ictlr_a0 ( bkpt_ena, bkpt_pc, memaddr_c, memaddr, mcu_psr_c, mcu_psw, 
        hit_ps_c, hit_ps, mempsack, memdatao, o_set_hold, o_bkp_hold, 
        o_ofs_inc, o_inst, d_inst, sfr_psrack, sfr_psofs, sfr_psr, sfr_psw, 
        dw_rst, dw_ena, sfr_wdat, pmem_pgm, pmem_re, pmem_csb, pmem_clk, 
        pmem_a, pmem_q0, pmem_q1, pmem_twlb, wd_twlb, we_twlb, pwrdn_rst, 
        r_pwdn_en, r_multi, r_hold_mcu, clk, srst, test_si3, test_si2, 
        test_si1, test_so2, test_so1, test_se );
  input [14:0] bkpt_pc;
  input [14:0] memaddr_c;
  input [14:0] memaddr;
  input [7:0] memdatao;
  output [7:0] o_inst;
  output [7:0] d_inst;
  input [14:0] sfr_psofs;
  input [7:0] sfr_wdat;
  output [1:0] pmem_clk;
  output [15:0] pmem_a;
  input [7:0] pmem_q0;
  input [7:0] pmem_q1;
  output [1:0] pmem_twlb;
  input [1:0] wd_twlb;
  input bkpt_ena, mcu_psr_c, mcu_psw, hit_ps_c, hit_ps, sfr_psr, sfr_psw,
         dw_rst, dw_ena, we_twlb, pwrdn_rst, r_pwdn_en, r_multi, r_hold_mcu,
         clk, srst, test_si3, test_si2, test_si1, test_se;
  output mempsack, o_set_hold, o_bkp_hold, o_ofs_inc, sfr_psrack, pmem_pgm,
         pmem_re, pmem_csb, test_so2, test_so1;
  wire   N152, N153, N154, c_buf_22__7_, c_buf_22__6_, c_buf_22__5_,
         c_buf_22__4_, c_buf_22__3_, c_buf_22__2_, c_buf_22__1_, c_buf_22__0_,
         c_buf_21__7_, c_buf_21__6_, c_buf_21__5_, c_buf_21__4_, c_buf_21__3_,
         c_buf_21__2_, c_buf_21__1_, c_buf_21__0_, c_buf_20__7_, c_buf_20__6_,
         c_buf_20__5_, c_buf_20__4_, c_buf_20__3_, c_buf_20__2_, c_buf_20__1_,
         c_buf_20__0_, c_buf_19__7_, c_buf_19__6_, c_buf_19__5_, c_buf_19__4_,
         c_buf_19__3_, c_buf_19__2_, c_buf_19__1_, c_buf_19__0_, c_buf_18__7_,
         c_buf_18__6_, c_buf_18__5_, c_buf_18__4_, c_buf_18__3_, c_buf_18__2_,
         c_buf_18__1_, c_buf_18__0_, c_buf_17__7_, c_buf_17__6_, c_buf_17__5_,
         c_buf_17__4_, c_buf_17__3_, c_buf_17__2_, c_buf_17__1_, c_buf_17__0_,
         c_buf_16__7_, c_buf_16__6_, c_buf_16__5_, c_buf_16__4_, c_buf_16__3_,
         c_buf_16__2_, c_buf_16__1_, c_buf_16__0_, wspp_cnt_5_, wspp_cnt_4_,
         wspp_cnt_3_, wspp_cnt_2_, wspp_cnt_1_, wspp_cnt_0_, d_psrd, r_rdy,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617,
         N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628,
         N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639,
         N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650,
         N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661,
         N662, N757, N759, N786, N787, N788, N789, N790, N791, N792, N793,
         N795, N796, N797, N798, N799, N800, N801, N820, N821, N822, N823,
         N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834,
         N835, N836, N837, N838, N839, N840, N842, N843, N844, N845, N846,
         N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863,
         N864, N865, N866, N867, N868, N874, N875, N876, N877, N878, N879,
         N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890,
         N891, N892, N893, N894, N895, N896, N897, N898, N899, un_hold,
         net11846, net11852, net11857, net11862, net11867, net11872, net11877,
         net11882, net11887, net11892, net11897, net11902, net11907, net11912,
         net11917, net11922, net11927, net11932, net11937, net11942, net11947,
         net11952, net11957, net11962, net11967, net11972, net11977, net11982,
         net11987, net11992, n93, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n801, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n400, n401,
         n412, n442, n446, n448, n453, n520, n531, n532, n533, n534, n535,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n569, n570,
         n675, n717, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n397, n398, n399, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n443, n444, n445, n447, n449, n450,
         n451, n452, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n536, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852;
  wire   [3:0] d_hold;
  wire   [1:0] dummy;
  wire   [3:0] cs_ft;
  wire   [4:0] c_ptr;
  wire   [14:0] c_adr;
  wire   [14:13] adr_p;
  wire   [7:0] rd_buf;
  wire   [7:0] dbg_01;
  wire   [7:0] dbg_02;
  wire   [7:0] dbg_03;
  wire   [7:0] dbg_04;
  wire   [7:0] dbg_05;
  wire   [7:0] dbg_06;
  wire   [7:0] dbg_07;
  wire   [7:0] dbg_08;
  wire   [7:0] dbg_09;
  wire   [7:0] dbg_0a;
  wire   [7:0] dbg_0b;
  wire   [7:0] dbg_0c;
  wire   [7:0] dbg_0d;
  wire   [7:0] dbg_0e;
  wire   [7:0] dbg_0f;
  wire   [7:0] wr_buf;
  wire   [14:0] pre_1_adr;
  wire   [4:1] popptr;
  wire   [4:1] sub_313_carry;

  FAD1X1 sub_313_U2_1 ( .A(memaddr[1]), .B(n686), .CI(sub_313_carry[1]), .CO(
        sub_313_carry[2]), .SO(popptr[1]) );
  FAD1X1 sub_313_U2_2 ( .A(memaddr[2]), .B(n684), .CI(sub_313_carry[2]), .CO(
        sub_313_carry[3]), .SO(popptr[2]) );
  FAD1X1 sub_313_U2_3 ( .A(memaddr[3]), .B(n683), .CI(sub_313_carry[3]), .CO(
        sub_313_carry[4]), .SO(popptr[3]) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 clk_gate_wspp_cnt_reg ( .CLK(clk), .EN(N899), 
        .ENCLK(net11846), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 clk_gate_a_bit_reg ( .CLK(clk), .EN(N898), 
        .ENCLK(net11852), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 clk_gate_adr_p_reg ( .CLK(clk), .EN(N853), 
        .ENCLK(net11857), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 clk_gate_c_buf_reg_23_ ( .CLK(clk), .EN(
        N897), .ENCLK(net11862), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 clk_gate_c_buf_reg_22_ ( .CLK(clk), .EN(
        N896), .ENCLK(net11867), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 clk_gate_c_buf_reg_21_ ( .CLK(clk), .EN(
        N895), .ENCLK(net11872), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 clk_gate_c_buf_reg_20_ ( .CLK(clk), .EN(
        N894), .ENCLK(net11877), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 clk_gate_c_buf_reg_19_ ( .CLK(clk), .EN(
        N893), .ENCLK(net11882), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 clk_gate_c_buf_reg_18_ ( .CLK(clk), .EN(
        N892), .ENCLK(net11887), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 clk_gate_c_buf_reg_17_ ( .CLK(clk), .EN(
        N891), .ENCLK(net11892), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 clk_gate_c_buf_reg_16_ ( .CLK(clk), .EN(
        N890), .ENCLK(net11897), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 clk_gate_c_buf_reg_15_ ( .CLK(clk), .EN(
        N889), .ENCLK(net11902), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 clk_gate_c_buf_reg_14_ ( .CLK(clk), .EN(
        N888), .ENCLK(net11907), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 clk_gate_c_buf_reg_13_ ( .CLK(clk), .EN(
        N887), .ENCLK(net11912), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 clk_gate_c_buf_reg_12_ ( .CLK(clk), .EN(
        N886), .ENCLK(net11917), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 clk_gate_c_buf_reg_11_ ( .CLK(clk), .EN(
        N885), .ENCLK(net11922), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 clk_gate_c_buf_reg_10_ ( .CLK(clk), .EN(
        N884), .ENCLK(net11927), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 clk_gate_c_buf_reg_9_ ( .CLK(clk), .EN(N883), .ENCLK(net11932), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 clk_gate_c_buf_reg_8_ ( .CLK(clk), .EN(N882), .ENCLK(net11937), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 clk_gate_c_buf_reg_7_ ( .CLK(clk), .EN(N881), .ENCLK(net11942), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 clk_gate_c_buf_reg_6_ ( .CLK(clk), .EN(N880), .ENCLK(net11947), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 clk_gate_c_buf_reg_5_ ( .CLK(clk), .EN(N879), 
        .ENCLK(net11952), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 clk_gate_c_buf_reg_4_ ( .CLK(clk), .EN(N878), 
        .ENCLK(net11957), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 clk_gate_c_buf_reg_3_ ( .CLK(clk), .EN(N877), 
        .ENCLK(net11962), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 clk_gate_c_buf_reg_2_ ( .CLK(clk), .EN(N876), 
        .ENCLK(net11967), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 clk_gate_c_buf_reg_1_ ( .CLK(clk), .EN(N875), 
        .ENCLK(net11972), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 clk_gate_c_buf_reg_0_ ( .CLK(clk), .EN(N874), 
        .ENCLK(net11977), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 clk_gate_c_ptr_reg ( .CLK(clk), .EN(n93), 
        .ENCLK(net11982), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 clk_gate_c_adr_reg ( .CLK(clk), .EN(N825), 
        .ENCLK(net11987), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 clk_gate_cs_ft_reg ( .CLK(clk), .EN(N820), 
        .ENCLK(net11992), .TE(test_se) );
  ictlr_a0_DW01_inc_1 add_242 ( .A(c_adr), .SUM({N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431}) );
  ictlr_a0_DW01_inc_2 r492 ( .A({adr_p, pmem_a[15:9], pmem_a[5:0]}), .SUM(
        pre_1_adr) );
  SDFFQX2 a_bit_reg_2_ ( .D(N759), .SIN(pmem_a[7]), .SMC(test_se), .C(net11852), .Q(pmem_a[8]) );
  SDFFQX2 a_bit_reg_0_ ( .D(N757), .SIN(test_si2), .SMC(test_se), .C(net11852), 
        .Q(pmem_a[6]) );
  SDFFQX1 wspp_cnt_reg_2_ ( .D(N797), .SIN(wspp_cnt_1_), .SMC(test_se), .C(
        net11846), .Q(wspp_cnt_2_) );
  SDFFQX1 wspp_cnt_reg_0_ ( .D(N795), .SIN(un_hold), .SMC(test_se), .C(
        net11846), .Q(wspp_cnt_0_) );
  SDFFQX1 wspp_cnt_reg_1_ ( .D(N796), .SIN(wspp_cnt_0_), .SMC(test_se), .C(
        net11846), .Q(wspp_cnt_1_) );
  SDFFQX1 d_hold_reg_3_ ( .D(N154), .SIN(d_hold[2]), .SMC(test_se), .C(clk), 
        .Q(d_hold[3]) );
  SDFFQX1 d_hold_reg_2_ ( .D(N153), .SIN(d_hold[1]), .SMC(test_se), .C(clk), 
        .Q(d_hold[2]) );
  SDFFQX1 d_hold_reg_1_ ( .D(N152), .SIN(d_hold[0]), .SMC(test_se), .C(clk), 
        .Q(d_hold[1]) );
  SDFFQX1 dummy_reg_0_ ( .D(n651), .SIN(n19), .SMC(test_se), .C(clk), .Q(
        dummy[0]) );
  SDFFQX1 d_hold_reg_0_ ( .D(n801), .SIN(cs_ft[3]), .SMC(test_se), .C(clk), 
        .Q(d_hold[0]) );
  SDFFQX1 dummy_reg_1_ ( .D(n650), .SIN(dummy[0]), .SMC(test_se), .C(clk), .Q(
        dummy[1]) );
  SDFFQX2 adr_p_reg_3_ ( .D(N857), .SIN(pmem_a[2]), .SMC(test_se), .C(net11857), .Q(pmem_a[3]) );
  SDFFQX2 adr_p_reg_4_ ( .D(N858), .SIN(pmem_a[3]), .SMC(test_se), .C(net11857), .Q(pmem_a[4]) );
  SDFFQX2 adr_p_reg_5_ ( .D(N859), .SIN(pmem_a[4]), .SMC(test_se), .C(net11857), .Q(pmem_a[5]) );
  SDFFQX1 d_psrd_reg ( .D(n649), .SIN(d_hold[3]), .SMC(test_se), .C(net11992), 
        .Q(d_psrd) );
  SDFFQX2 adr_p_reg_1_ ( .D(N855), .SIN(pmem_a[0]), .SMC(test_se), .C(net11857), .Q(pmem_a[1]) );
  SDFFQX2 adr_p_reg_2_ ( .D(N856), .SIN(pmem_a[1]), .SMC(test_se), .C(net11857), .Q(pmem_a[2]) );
  SDFFQX1 c_adr_reg_14_ ( .D(N840), .SIN(c_adr[13]), .SMC(test_se), .C(
        net11987), .Q(c_adr[14]) );
  SDFFQX1 c_adr_reg_13_ ( .D(N839), .SIN(c_adr[12]), .SMC(test_se), .C(
        net11987), .Q(c_adr[13]) );
  SDFFQX1 c_adr_reg_12_ ( .D(N838), .SIN(c_adr[11]), .SMC(test_se), .C(
        net11987), .Q(c_adr[12]) );
  SDFFQX1 c_adr_reg_11_ ( .D(N837), .SIN(c_adr[10]), .SMC(test_se), .C(
        net11987), .Q(c_adr[11]) );
  SDFFQX1 c_adr_reg_10_ ( .D(N836), .SIN(c_adr[9]), .SMC(test_se), .C(net11987), .Q(c_adr[10]) );
  SDFFQX1 c_adr_reg_8_ ( .D(N834), .SIN(c_adr[7]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[8]) );
  SDFFQX1 c_adr_reg_9_ ( .D(N835), .SIN(c_adr[8]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[9]) );
  SDFFQX1 c_adr_reg_7_ ( .D(N833), .SIN(c_adr[6]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[7]) );
  SDFFQX1 c_adr_reg_6_ ( .D(N832), .SIN(c_adr[5]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[6]) );
  SDFFQX1 c_adr_reg_5_ ( .D(N831), .SIN(c_adr[4]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[5]) );
  SDFFQX1 c_ptr_reg_4_ ( .D(N846), .SIN(c_ptr[3]), .SMC(test_se), .C(net11982), 
        .Q(c_ptr[4]) );
  SDFFQX1 c_ptr_reg_3_ ( .D(N845), .SIN(c_ptr[2]), .SMC(test_se), .C(net11982), 
        .Q(c_ptr[3]) );
  SDFFQX1 pgm_p_reg ( .D(n644), .SIN(dummy[1]), .SMC(test_se), .C(net11992), 
        .Q(pmem_pgm) );
  SDFFQX1 c_ptr_reg_2_ ( .D(N844), .SIN(c_ptr[1]), .SMC(test_se), .C(net11982), 
        .Q(c_ptr[2]) );
  SDFFQX1 c_ptr_reg_1_ ( .D(N843), .SIN(c_ptr[0]), .SMC(test_se), .C(net11982), 
        .Q(c_ptr[1]) );
  SDFFQX1 c_ptr_reg_0_ ( .D(N842), .SIN(wr_buf[7]), .SMC(test_se), .C(net11982), .Q(c_ptr[0]) );
  SDFFQX1 un_hold_reg ( .D(n717), .SIN(pmem_re), .SMC(test_se), .C(clk), .Q(
        un_hold) );
  SDFFQX1 c_buf_reg_15__6_ ( .D(N605), .SIN(dbg_0f[5]), .SMC(test_se), .C(
        net11902), .Q(dbg_0f[6]) );
  SDFFQX1 c_buf_reg_15__4_ ( .D(N603), .SIN(dbg_0f[3]), .SMC(test_se), .C(
        net11902), .Q(dbg_0f[4]) );
  SDFFQX1 c_buf_reg_15__3_ ( .D(N602), .SIN(dbg_0f[2]), .SMC(test_se), .C(
        net11902), .Q(dbg_0f[3]) );
  SDFFQX1 c_buf_reg_15__2_ ( .D(N601), .SIN(dbg_0f[1]), .SMC(test_se), .C(
        net11902), .Q(dbg_0f[2]) );
  SDFFQX1 c_buf_reg_15__1_ ( .D(N600), .SIN(dbg_0f[0]), .SMC(test_se), .C(
        net11902), .Q(dbg_0f[1]) );
  SDFFQX1 c_buf_reg_15__0_ ( .D(N599), .SIN(dbg_0e[7]), .SMC(test_se), .C(
        net11902), .Q(dbg_0f[0]) );
  SDFFQX1 c_buf_reg_12__6_ ( .D(N581), .SIN(dbg_0c[5]), .SMC(test_se), .C(
        net11917), .Q(dbg_0c[6]) );
  SDFFQX1 c_buf_reg_12__4_ ( .D(N579), .SIN(dbg_0c[3]), .SMC(test_se), .C(
        net11917), .Q(dbg_0c[4]) );
  SDFFQX1 c_buf_reg_12__3_ ( .D(N578), .SIN(dbg_0c[2]), .SMC(test_se), .C(
        net11917), .Q(dbg_0c[3]) );
  SDFFQX1 c_buf_reg_12__2_ ( .D(N577), .SIN(dbg_0c[1]), .SMC(test_se), .C(
        net11917), .Q(dbg_0c[2]) );
  SDFFQX1 c_buf_reg_12__1_ ( .D(N576), .SIN(dbg_0c[0]), .SMC(test_se), .C(
        net11917), .Q(dbg_0c[1]) );
  SDFFQX1 c_buf_reg_12__0_ ( .D(N575), .SIN(dbg_0b[7]), .SMC(test_se), .C(
        net11917), .Q(dbg_0c[0]) );
  SDFFQX1 c_buf_reg_16__6_ ( .D(N613), .SIN(c_buf_16__5_), .SMC(test_se), .C(
        net11897), .Q(c_buf_16__6_) );
  SDFFQX1 c_buf_reg_16__4_ ( .D(N611), .SIN(c_buf_16__3_), .SMC(test_se), .C(
        net11897), .Q(c_buf_16__4_) );
  SDFFQX1 c_buf_reg_16__3_ ( .D(N610), .SIN(c_buf_16__2_), .SMC(test_se), .C(
        net11897), .Q(c_buf_16__3_) );
  SDFFQX1 c_buf_reg_16__2_ ( .D(N609), .SIN(c_buf_16__1_), .SMC(test_se), .C(
        net11897), .Q(c_buf_16__2_) );
  SDFFQX1 c_buf_reg_16__1_ ( .D(N608), .SIN(c_buf_16__0_), .SMC(test_se), .C(
        net11897), .Q(c_buf_16__1_) );
  SDFFQX1 c_buf_reg_16__0_ ( .D(N607), .SIN(dbg_0f[7]), .SMC(test_se), .C(
        net11897), .Q(c_buf_16__0_) );
  SDFFQX1 c_buf_reg_13__6_ ( .D(N589), .SIN(dbg_0d[5]), .SMC(test_se), .C(
        net11912), .Q(dbg_0d[6]) );
  SDFFQX1 c_buf_reg_13__4_ ( .D(N587), .SIN(dbg_0d[3]), .SMC(test_se), .C(
        net11912), .Q(dbg_0d[4]) );
  SDFFQX1 c_buf_reg_13__3_ ( .D(N586), .SIN(dbg_0d[2]), .SMC(test_se), .C(
        net11912), .Q(dbg_0d[3]) );
  SDFFQX1 c_buf_reg_13__2_ ( .D(N585), .SIN(dbg_0d[1]), .SMC(test_se), .C(
        net11912), .Q(dbg_0d[2]) );
  SDFFQX1 c_buf_reg_13__1_ ( .D(N584), .SIN(dbg_0d[0]), .SMC(test_se), .C(
        net11912), .Q(dbg_0d[1]) );
  SDFFQX1 c_buf_reg_13__0_ ( .D(N583), .SIN(dbg_0c[7]), .SMC(test_se), .C(
        net11912), .Q(dbg_0d[0]) );
  SDFFQX1 c_buf_reg_17__6_ ( .D(N621), .SIN(c_buf_17__5_), .SMC(test_se), .C(
        net11892), .Q(c_buf_17__6_) );
  SDFFQX1 c_buf_reg_17__5_ ( .D(N620), .SIN(c_buf_17__4_), .SMC(test_se), .C(
        net11892), .Q(c_buf_17__5_) );
  SDFFQX1 c_buf_reg_17__4_ ( .D(N619), .SIN(c_buf_17__3_), .SMC(test_se), .C(
        net11892), .Q(c_buf_17__4_) );
  SDFFQX1 c_buf_reg_17__3_ ( .D(N618), .SIN(c_buf_17__2_), .SMC(test_se), .C(
        net11892), .Q(c_buf_17__3_) );
  SDFFQX1 c_buf_reg_17__2_ ( .D(N617), .SIN(c_buf_17__1_), .SMC(test_se), .C(
        net11892), .Q(c_buf_17__2_) );
  SDFFQX1 c_buf_reg_17__1_ ( .D(N616), .SIN(c_buf_17__0_), .SMC(test_se), .C(
        net11892), .Q(c_buf_17__1_) );
  SDFFQX1 c_buf_reg_17__0_ ( .D(N615), .SIN(c_buf_16__7_), .SMC(test_se), .C(
        net11892), .Q(c_buf_17__0_) );
  SDFFQX1 c_buf_reg_14__6_ ( .D(N597), .SIN(dbg_0e[5]), .SMC(test_se), .C(
        net11907), .Q(dbg_0e[6]) );
  SDFFQX1 c_buf_reg_14__5_ ( .D(N596), .SIN(dbg_0e[4]), .SMC(test_se), .C(
        net11907), .Q(dbg_0e[5]) );
  SDFFQX1 c_buf_reg_14__4_ ( .D(N595), .SIN(dbg_0e[3]), .SMC(test_se), .C(
        net11907), .Q(dbg_0e[4]) );
  SDFFQX1 c_buf_reg_14__3_ ( .D(N594), .SIN(dbg_0e[2]), .SMC(test_se), .C(
        net11907), .Q(dbg_0e[3]) );
  SDFFQX1 c_buf_reg_14__2_ ( .D(N593), .SIN(dbg_0e[1]), .SMC(test_se), .C(
        net11907), .Q(dbg_0e[2]) );
  SDFFQX1 c_buf_reg_14__1_ ( .D(N592), .SIN(dbg_0e[0]), .SMC(test_se), .C(
        net11907), .Q(dbg_0e[1]) );
  SDFFQX1 c_buf_reg_14__0_ ( .D(N591), .SIN(dbg_0d[7]), .SMC(test_se), .C(
        net11907), .Q(dbg_0e[0]) );
  SDFFQX1 re_p_reg ( .D(n647), .SIN(pmem_twlb[1]), .SMC(test_se), .C(clk), .Q(
        pmem_re) );
  SDFFQX1 adr_p_reg_14_ ( .D(N868), .SIN(adr_p[13]), .SMC(test_se), .C(
        net11857), .Q(adr_p[14]) );
  SDFFQX1 c_buf_reg_22__0_ ( .D(N655), .SIN(c_buf_21__7_), .SMC(test_se), .C(
        net11867), .Q(c_buf_22__0_) );
  SDFFQX1 c_buf_reg_21__0_ ( .D(N647), .SIN(c_buf_20__7_), .SMC(test_se), .C(
        net11872), .Q(c_buf_21__0_) );
  SDFFQX1 c_buf_reg_23__1_ ( .D(N787), .SIN(wr_buf[0]), .SMC(test_se), .C(
        net11862), .Q(wr_buf[1]) );
  SDFFQX1 c_buf_reg_23__0_ ( .D(N786), .SIN(c_buf_22__7_), .SMC(test_se), .C(
        net11862), .Q(wr_buf[0]) );
  SDFFQX1 c_buf_reg_23__4_ ( .D(N790), .SIN(wr_buf[3]), .SMC(test_se), .C(
        net11862), .Q(wr_buf[4]) );
  SDFFQX1 c_buf_reg_23__6_ ( .D(N792), .SIN(wr_buf[5]), .SMC(test_se), .C(
        net11862), .Q(wr_buf[6]) );
  SDFFQX1 c_buf_reg_23__2_ ( .D(N788), .SIN(wr_buf[1]), .SMC(test_se), .C(
        net11862), .Q(wr_buf[2]) );
  SDFFQX1 c_buf_reg_23__3_ ( .D(N789), .SIN(wr_buf[2]), .SMC(test_se), .C(
        net11862), .Q(wr_buf[3]) );
  SDFFQX2 adr_p_reg_6_ ( .D(N860), .SIN(pmem_a[5]), .SMC(test_se), .C(net11857), .Q(pmem_a[9]) );
  SDFFQX1 c_buf_reg_15__5_ ( .D(N604), .SIN(dbg_0f[4]), .SMC(test_se), .C(
        net11902), .Q(dbg_0f[5]) );
  SDFFQX1 c_buf_reg_12__5_ ( .D(N580), .SIN(dbg_0c[4]), .SMC(test_se), .C(
        net11917), .Q(dbg_0c[5]) );
  SDFFQX1 c_buf_reg_13__5_ ( .D(N588), .SIN(dbg_0d[4]), .SMC(test_se), .C(
        net11912), .Q(dbg_0d[5]) );
  SDFFQX1 c_buf_reg_16__5_ ( .D(N612), .SIN(c_buf_16__4_), .SMC(test_se), .C(
        net11897), .Q(c_buf_16__5_) );
  SDFFQX1 c_buf_reg_0__6_ ( .D(N485), .SIN(rd_buf[5]), .SMC(test_se), .C(
        net11977), .Q(rd_buf[6]) );
  SDFFQX1 c_buf_reg_0__3_ ( .D(N482), .SIN(rd_buf[2]), .SMC(test_se), .C(
        net11977), .Q(rd_buf[3]) );
  SDFFQX1 c_buf_reg_0__2_ ( .D(N481), .SIN(rd_buf[1]), .SMC(test_se), .C(
        net11977), .Q(rd_buf[2]) );
  SDFFQX1 c_buf_reg_0__1_ ( .D(N480), .SIN(rd_buf[0]), .SMC(test_se), .C(
        net11977), .Q(rd_buf[1]) );
  SDFFQX1 c_buf_reg_0__4_ ( .D(N483), .SIN(rd_buf[3]), .SMC(test_se), .C(
        net11977), .Q(rd_buf[4]) );
  SDFFQX1 c_buf_reg_0__0_ ( .D(N479), .SIN(c_adr[14]), .SMC(test_se), .C(
        net11977), .Q(rd_buf[0]) );
  SDFFQX1 adr_p_reg_13_ ( .D(N867), .SIN(pmem_a[14]), .SMC(test_se), .C(
        net11857), .Q(adr_p[13]) );
  SDFFQX1 c_buf_reg_5__6_ ( .D(N525), .SIN(dbg_05[5]), .SMC(test_se), .C(
        net11952), .Q(dbg_05[6]) );
  SDFFQX1 c_buf_reg_2__6_ ( .D(N501), .SIN(dbg_02[5]), .SMC(test_se), .C(
        net11967), .Q(dbg_02[6]) );
  SDFFQX1 c_buf_reg_5__4_ ( .D(N523), .SIN(dbg_05[3]), .SMC(test_se), .C(
        net11952), .Q(dbg_05[4]) );
  SDFFQX1 c_buf_reg_2__4_ ( .D(N499), .SIN(dbg_02[3]), .SMC(test_se), .C(
        net11967), .Q(dbg_02[4]) );
  SDFFQX1 c_buf_reg_5__3_ ( .D(N522), .SIN(dbg_05[2]), .SMC(test_se), .C(
        net11952), .Q(dbg_05[3]) );
  SDFFQX1 c_buf_reg_2__3_ ( .D(N498), .SIN(dbg_02[2]), .SMC(test_se), .C(
        net11967), .Q(dbg_02[3]) );
  SDFFQX1 c_buf_reg_5__2_ ( .D(N521), .SIN(dbg_05[1]), .SMC(test_se), .C(
        net11952), .Q(dbg_05[2]) );
  SDFFQX1 c_buf_reg_2__2_ ( .D(N497), .SIN(dbg_02[1]), .SMC(test_se), .C(
        net11967), .Q(dbg_02[2]) );
  SDFFQX1 c_buf_reg_5__1_ ( .D(N520), .SIN(dbg_05[0]), .SMC(test_se), .C(
        net11952), .Q(dbg_05[1]) );
  SDFFQX1 c_buf_reg_2__1_ ( .D(N496), .SIN(dbg_02[0]), .SMC(test_se), .C(
        net11967), .Q(dbg_02[1]) );
  SDFFQX1 c_buf_reg_5__0_ ( .D(N519), .SIN(dbg_04[7]), .SMC(test_se), .C(
        net11952), .Q(dbg_05[0]) );
  SDFFQX1 c_buf_reg_2__0_ ( .D(N495), .SIN(dbg_01[7]), .SMC(test_se), .C(
        net11967), .Q(dbg_02[0]) );
  SDFFQX1 c_buf_reg_3__6_ ( .D(N509), .SIN(dbg_03[5]), .SMC(test_se), .C(
        net11962), .Q(dbg_03[6]) );
  SDFFQX1 c_buf_reg_3__4_ ( .D(N507), .SIN(dbg_03[3]), .SMC(test_se), .C(
        net11962), .Q(dbg_03[4]) );
  SDFFQX1 c_buf_reg_3__3_ ( .D(N506), .SIN(dbg_03[2]), .SMC(test_se), .C(
        net11962), .Q(dbg_03[3]) );
  SDFFQX1 c_buf_reg_3__2_ ( .D(N505), .SIN(dbg_03[1]), .SMC(test_se), .C(
        net11962), .Q(dbg_03[2]) );
  SDFFQX1 c_buf_reg_3__1_ ( .D(N504), .SIN(dbg_03[0]), .SMC(test_se), .C(
        net11962), .Q(dbg_03[1]) );
  SDFFQX1 c_buf_reg_3__0_ ( .D(N503), .SIN(dbg_02[7]), .SMC(test_se), .C(
        net11962), .Q(dbg_03[0]) );
  SDFFQX1 c_buf_reg_4__6_ ( .D(N517), .SIN(dbg_04[5]), .SMC(test_se), .C(
        net11957), .Q(dbg_04[6]) );
  SDFFQX1 c_buf_reg_1__6_ ( .D(N493), .SIN(dbg_01[5]), .SMC(test_se), .C(
        net11972), .Q(dbg_01[6]) );
  SDFFQX1 c_buf_reg_4__4_ ( .D(N515), .SIN(dbg_04[3]), .SMC(test_se), .C(
        net11957), .Q(dbg_04[4]) );
  SDFFQX1 c_buf_reg_1__4_ ( .D(N491), .SIN(dbg_01[3]), .SMC(test_se), .C(
        net11972), .Q(dbg_01[4]) );
  SDFFQX1 c_buf_reg_4__3_ ( .D(N514), .SIN(dbg_04[2]), .SMC(test_se), .C(
        net11957), .Q(dbg_04[3]) );
  SDFFQX1 c_buf_reg_1__3_ ( .D(N490), .SIN(dbg_01[2]), .SMC(test_se), .C(
        net11972), .Q(dbg_01[3]) );
  SDFFQX1 c_buf_reg_4__2_ ( .D(N513), .SIN(dbg_04[1]), .SMC(test_se), .C(
        net11957), .Q(dbg_04[2]) );
  SDFFQX1 c_buf_reg_1__2_ ( .D(N489), .SIN(dbg_01[1]), .SMC(test_se), .C(
        net11972), .Q(dbg_01[2]) );
  SDFFQX1 c_buf_reg_4__1_ ( .D(N512), .SIN(dbg_04[0]), .SMC(test_se), .C(
        net11957), .Q(dbg_04[1]) );
  SDFFQX1 c_buf_reg_1__1_ ( .D(N488), .SIN(dbg_01[0]), .SMC(test_se), .C(
        net11972), .Q(dbg_01[1]) );
  SDFFQX1 c_buf_reg_4__0_ ( .D(N511), .SIN(dbg_03[7]), .SMC(test_se), .C(
        net11957), .Q(dbg_04[0]) );
  SDFFQX1 c_buf_reg_1__0_ ( .D(N487), .SIN(rd_buf[7]), .SMC(test_se), .C(
        net11972), .Q(dbg_01[0]) );
  SDFFQX1 c_buf_reg_6__6_ ( .D(N533), .SIN(dbg_06[5]), .SMC(test_se), .C(
        net11947), .Q(dbg_06[6]) );
  SDFFQX1 c_buf_reg_6__4_ ( .D(N531), .SIN(dbg_06[3]), .SMC(test_se), .C(
        net11947), .Q(dbg_06[4]) );
  SDFFQX1 c_buf_reg_6__3_ ( .D(N530), .SIN(dbg_06[2]), .SMC(test_se), .C(
        net11947), .Q(dbg_06[3]) );
  SDFFQX1 c_buf_reg_6__2_ ( .D(N529), .SIN(dbg_06[1]), .SMC(test_se), .C(
        net11947), .Q(dbg_06[2]) );
  SDFFQX1 c_buf_reg_6__1_ ( .D(N528), .SIN(dbg_06[0]), .SMC(test_se), .C(
        net11947), .Q(dbg_06[1]) );
  SDFFQX1 c_buf_reg_6__0_ ( .D(N527), .SIN(dbg_05[7]), .SMC(test_se), .C(
        net11947), .Q(dbg_06[0]) );
  SDFFQX1 c_buf_reg_11__4_ ( .D(N571), .SIN(dbg_0b[3]), .SMC(test_se), .C(
        net11922), .Q(dbg_0b[4]) );
  SDFFQX1 c_buf_reg_11__3_ ( .D(N570), .SIN(dbg_0b[2]), .SMC(test_se), .C(
        net11922), .Q(dbg_0b[3]) );
  SDFFQX1 c_buf_reg_11__2_ ( .D(N569), .SIN(dbg_0b[1]), .SMC(test_se), .C(
        net11922), .Q(dbg_0b[2]) );
  SDFFQX1 c_buf_reg_11__1_ ( .D(N568), .SIN(dbg_0b[0]), .SMC(test_se), .C(
        net11922), .Q(dbg_0b[1]) );
  SDFFQX1 c_buf_reg_11__0_ ( .D(N567), .SIN(dbg_0a[7]), .SMC(test_se), .C(
        net11922), .Q(dbg_0b[0]) );
  SDFFQX1 c_buf_reg_10__6_ ( .D(N565), .SIN(dbg_0a[5]), .SMC(test_se), .C(
        net11927), .Q(dbg_0a[6]) );
  SDFFQX1 c_buf_reg_10__4_ ( .D(N563), .SIN(dbg_0a[3]), .SMC(test_se), .C(
        net11927), .Q(dbg_0a[4]) );
  SDFFQX1 c_buf_reg_10__3_ ( .D(N562), .SIN(dbg_0a[2]), .SMC(test_se), .C(
        net11927), .Q(dbg_0a[3]) );
  SDFFQX1 c_buf_reg_10__2_ ( .D(N561), .SIN(dbg_0a[1]), .SMC(test_se), .C(
        net11927), .Q(dbg_0a[2]) );
  SDFFQX1 c_buf_reg_10__1_ ( .D(N560), .SIN(dbg_0a[0]), .SMC(test_se), .C(
        net11927), .Q(dbg_0a[1]) );
  SDFFQX1 c_buf_reg_10__0_ ( .D(N559), .SIN(dbg_09[7]), .SMC(test_se), .C(
        net11927), .Q(dbg_0a[0]) );
  SDFFQX1 c_buf_reg_7__4_ ( .D(N539), .SIN(dbg_07[3]), .SMC(test_se), .C(
        net11942), .Q(dbg_07[4]) );
  SDFFQX1 c_buf_reg_22__6_ ( .D(N661), .SIN(c_buf_22__5_), .SMC(test_se), .C(
        net11867), .Q(c_buf_22__6_) );
  SDFFQX1 c_buf_reg_22__4_ ( .D(N659), .SIN(c_buf_22__3_), .SMC(test_se), .C(
        net11867), .Q(c_buf_22__4_) );
  SDFFQX1 c_buf_reg_22__3_ ( .D(N658), .SIN(c_buf_22__2_), .SMC(test_se), .C(
        net11867), .Q(c_buf_22__3_) );
  SDFFQX1 c_buf_reg_22__2_ ( .D(N657), .SIN(c_buf_22__1_), .SMC(test_se), .C(
        net11867), .Q(c_buf_22__2_) );
  SDFFQX1 c_buf_reg_22__1_ ( .D(N656), .SIN(c_buf_22__0_), .SMC(test_se), .C(
        net11867), .Q(c_buf_22__1_) );
  SDFFQX1 c_buf_reg_21__6_ ( .D(N653), .SIN(c_buf_21__5_), .SMC(test_se), .C(
        net11872), .Q(c_buf_21__6_) );
  SDFFQX1 c_buf_reg_21__4_ ( .D(N651), .SIN(c_buf_21__3_), .SMC(test_se), .C(
        net11872), .Q(c_buf_21__4_) );
  SDFFQX1 c_buf_reg_21__3_ ( .D(N650), .SIN(c_buf_21__2_), .SMC(test_se), .C(
        net11872), .Q(c_buf_21__3_) );
  SDFFQX1 c_buf_reg_21__2_ ( .D(N649), .SIN(c_buf_21__1_), .SMC(test_se), .C(
        net11872), .Q(c_buf_21__2_) );
  SDFFQX1 c_buf_reg_21__1_ ( .D(N648), .SIN(c_buf_21__0_), .SMC(test_se), .C(
        net11872), .Q(c_buf_21__1_) );
  SDFFQX1 c_buf_reg_20__6_ ( .D(N645), .SIN(c_buf_20__5_), .SMC(test_se), .C(
        net11877), .Q(c_buf_20__6_) );
  SDFFQX1 c_buf_reg_20__5_ ( .D(N644), .SIN(c_buf_20__4_), .SMC(test_se), .C(
        net11877), .Q(c_buf_20__5_) );
  SDFFQX1 c_buf_reg_20__4_ ( .D(N643), .SIN(c_buf_20__3_), .SMC(test_se), .C(
        net11877), .Q(c_buf_20__4_) );
  SDFFQX1 c_buf_reg_20__3_ ( .D(N642), .SIN(c_buf_20__2_), .SMC(test_se), .C(
        net11877), .Q(c_buf_20__3_) );
  SDFFQX1 c_buf_reg_20__2_ ( .D(N641), .SIN(c_buf_20__1_), .SMC(test_se), .C(
        net11877), .Q(c_buf_20__2_) );
  SDFFQX1 c_buf_reg_20__1_ ( .D(N640), .SIN(c_buf_20__0_), .SMC(test_se), .C(
        net11877), .Q(c_buf_20__1_) );
  SDFFQX1 c_buf_reg_20__0_ ( .D(N639), .SIN(c_buf_19__7_), .SMC(test_se), .C(
        net11877), .Q(c_buf_20__0_) );
  SDFFQX1 c_buf_reg_19__6_ ( .D(N637), .SIN(c_buf_19__5_), .SMC(test_se), .C(
        net11882), .Q(c_buf_19__6_) );
  SDFFQX1 c_buf_reg_19__4_ ( .D(N635), .SIN(c_buf_19__3_), .SMC(test_se), .C(
        net11882), .Q(c_buf_19__4_) );
  SDFFQX1 c_buf_reg_19__3_ ( .D(N634), .SIN(c_buf_19__2_), .SMC(test_se), .C(
        net11882), .Q(c_buf_19__3_) );
  SDFFQX1 c_buf_reg_19__2_ ( .D(N633), .SIN(c_buf_19__1_), .SMC(test_se), .C(
        net11882), .Q(c_buf_19__2_) );
  SDFFQX1 c_buf_reg_19__1_ ( .D(N632), .SIN(c_buf_19__0_), .SMC(test_se), .C(
        net11882), .Q(c_buf_19__1_) );
  SDFFQX1 c_buf_reg_19__0_ ( .D(N631), .SIN(c_buf_18__7_), .SMC(test_se), .C(
        net11882), .Q(c_buf_19__0_) );
  SDFFQX1 c_buf_reg_18__6_ ( .D(N629), .SIN(c_buf_18__5_), .SMC(test_se), .C(
        net11887), .Q(c_buf_18__6_) );
  SDFFQX1 c_buf_reg_18__4_ ( .D(N627), .SIN(c_buf_18__3_), .SMC(test_se), .C(
        net11887), .Q(c_buf_18__4_) );
  SDFFQX1 c_buf_reg_18__3_ ( .D(N626), .SIN(c_buf_18__2_), .SMC(test_se), .C(
        net11887), .Q(c_buf_18__3_) );
  SDFFQX1 c_buf_reg_18__2_ ( .D(N625), .SIN(c_buf_18__1_), .SMC(test_se), .C(
        net11887), .Q(c_buf_18__2_) );
  SDFFQX1 c_buf_reg_18__1_ ( .D(N624), .SIN(c_buf_18__0_), .SMC(test_se), .C(
        net11887), .Q(c_buf_18__1_) );
  SDFFQX1 c_buf_reg_18__0_ ( .D(N623), .SIN(c_buf_17__7_), .SMC(test_se), .C(
        net11887), .Q(c_buf_18__0_) );
  SDFFQX1 c_buf_reg_11__6_ ( .D(N573), .SIN(dbg_0b[5]), .SMC(test_se), .C(
        net11922), .Q(dbg_0b[6]) );
  SDFFQX1 c_buf_reg_11__5_ ( .D(N572), .SIN(dbg_0b[4]), .SMC(test_se), .C(
        net11922), .Q(dbg_0b[5]) );
  SDFFQX1 c_buf_reg_10__5_ ( .D(N564), .SIN(dbg_0a[4]), .SMC(test_se), .C(
        net11927), .Q(dbg_0a[5]) );
  SDFFQX1 c_buf_reg_9__6_ ( .D(N557), .SIN(dbg_09[5]), .SMC(test_se), .C(
        net11932), .Q(dbg_09[6]) );
  SDFFQX1 c_buf_reg_9__5_ ( .D(N556), .SIN(dbg_09[4]), .SMC(test_se), .C(
        net11932), .Q(dbg_09[5]) );
  SDFFQX1 c_buf_reg_9__4_ ( .D(N555), .SIN(dbg_09[3]), .SMC(test_se), .C(
        net11932), .Q(dbg_09[4]) );
  SDFFQX1 c_buf_reg_9__3_ ( .D(N554), .SIN(dbg_09[2]), .SMC(test_se), .C(
        net11932), .Q(dbg_09[3]) );
  SDFFQX1 c_buf_reg_9__2_ ( .D(N553), .SIN(dbg_09[1]), .SMC(test_se), .C(
        net11932), .Q(dbg_09[2]) );
  SDFFQX1 c_buf_reg_9__1_ ( .D(N552), .SIN(dbg_09[0]), .SMC(test_se), .C(
        net11932), .Q(dbg_09[1]) );
  SDFFQX1 c_buf_reg_9__0_ ( .D(N551), .SIN(dbg_08[7]), .SMC(test_se), .C(
        net11932), .Q(dbg_09[0]) );
  SDFFQX1 c_buf_reg_8__6_ ( .D(N549), .SIN(dbg_08[5]), .SMC(test_se), .C(
        net11937), .Q(dbg_08[6]) );
  SDFFQX1 c_buf_reg_8__4_ ( .D(N547), .SIN(dbg_08[3]), .SMC(test_se), .C(
        net11937), .Q(dbg_08[4]) );
  SDFFQX1 c_buf_reg_8__3_ ( .D(N546), .SIN(dbg_08[2]), .SMC(test_se), .C(
        net11937), .Q(dbg_08[3]) );
  SDFFQX1 c_buf_reg_8__2_ ( .D(N545), .SIN(dbg_08[1]), .SMC(test_se), .C(
        net11937), .Q(dbg_08[2]) );
  SDFFQX1 c_buf_reg_8__1_ ( .D(N544), .SIN(dbg_08[0]), .SMC(test_se), .C(
        net11937), .Q(dbg_08[1]) );
  SDFFQX1 c_buf_reg_8__0_ ( .D(N543), .SIN(dbg_07[7]), .SMC(test_se), .C(
        net11937), .Q(dbg_08[0]) );
  SDFFQX1 c_buf_reg_7__6_ ( .D(N541), .SIN(dbg_07[5]), .SMC(test_se), .C(
        net11942), .Q(dbg_07[6]) );
  SDFFQX1 c_buf_reg_7__5_ ( .D(N540), .SIN(dbg_07[4]), .SMC(test_se), .C(
        net11942), .Q(dbg_07[5]) );
  SDFFQX1 c_buf_reg_7__3_ ( .D(N538), .SIN(dbg_07[2]), .SMC(test_se), .C(
        net11942), .Q(dbg_07[3]) );
  SDFFQX1 c_buf_reg_7__2_ ( .D(N537), .SIN(dbg_07[1]), .SMC(test_se), .C(
        net11942), .Q(dbg_07[2]) );
  SDFFQX1 c_buf_reg_7__1_ ( .D(N536), .SIN(dbg_07[0]), .SMC(test_se), .C(
        net11942), .Q(dbg_07[1]) );
  SDFFQX1 c_buf_reg_7__0_ ( .D(N535), .SIN(dbg_06[7]), .SMC(test_se), .C(
        net11942), .Q(dbg_07[0]) );
  SDFFQX1 c_buf_reg_22__5_ ( .D(N660), .SIN(c_buf_22__4_), .SMC(test_se), .C(
        net11867), .Q(c_buf_22__5_) );
  SDFFQX1 c_buf_reg_21__5_ ( .D(N652), .SIN(c_buf_21__4_), .SMC(test_se), .C(
        net11872), .Q(c_buf_21__5_) );
  SDFFQX1 c_buf_reg_19__5_ ( .D(N636), .SIN(c_buf_19__4_), .SMC(test_se), .C(
        net11882), .Q(c_buf_19__5_) );
  SDFFQX1 c_buf_reg_18__5_ ( .D(N628), .SIN(c_buf_18__4_), .SMC(test_se), .C(
        net11887), .Q(c_buf_18__5_) );
  SDFFQX1 c_buf_reg_23__5_ ( .D(N791), .SIN(wr_buf[4]), .SMC(test_se), .C(
        net11862), .Q(wr_buf[5]) );
  SDFFQX1 wspp_cnt_reg_6_ ( .D(N801), .SIN(wspp_cnt_5_), .SMC(test_se), .C(
        net11846), .Q(test_so2) );
  SDFFQX2 adr_p_reg_12_ ( .D(N866), .SIN(test_si3), .SMC(test_se), .C(net11857), .Q(pmem_a[15]) );
  SDFFQX2 adr_p_reg_11_ ( .D(N865), .SIN(pmem_a[13]), .SMC(test_se), .C(
        net11857), .Q(pmem_a[14]) );
  SDFFQX2 adr_p_reg_10_ ( .D(N864), .SIN(pmem_a[12]), .SMC(test_se), .C(
        net11857), .Q(pmem_a[13]) );
  SDFFQX2 adr_p_reg_8_ ( .D(N862), .SIN(pmem_a[10]), .SMC(test_se), .C(
        net11857), .Q(pmem_a[11]) );
  SDFFQX2 adr_p_reg_9_ ( .D(N863), .SIN(pmem_a[11]), .SMC(test_se), .C(
        net11857), .Q(pmem_a[12]) );
  SDFFQX2 adr_p_reg_7_ ( .D(N861), .SIN(pmem_a[9]), .SMC(test_se), .C(net11857), .Q(pmem_a[10]) );
  SDFFQX1 c_buf_reg_15__7_ ( .D(N606), .SIN(dbg_0f[6]), .SMC(test_se), .C(
        net11902), .Q(dbg_0f[7]) );
  SDFFQX1 c_buf_reg_12__7_ ( .D(N582), .SIN(dbg_0c[6]), .SMC(test_se), .C(
        net11917), .Q(dbg_0c[7]) );
  SDFFQX1 c_buf_reg_16__7_ ( .D(N614), .SIN(c_buf_16__6_), .SMC(test_se), .C(
        net11897), .Q(c_buf_16__7_) );
  SDFFQX1 c_buf_reg_13__7_ ( .D(N590), .SIN(dbg_0d[6]), .SMC(test_se), .C(
        net11912), .Q(dbg_0d[7]) );
  SDFFQX1 c_buf_reg_14__7_ ( .D(N598), .SIN(dbg_0e[6]), .SMC(test_se), .C(
        net11907), .Q(dbg_0e[7]) );
  SDFFQX1 c_buf_reg_17__7_ ( .D(N622), .SIN(c_buf_17__6_), .SMC(test_se), .C(
        net11892), .Q(c_buf_17__7_) );
  SDFFQX1 r_twlb_reg_0_ ( .D(n646), .SIN(r_rdy), .SMC(test_se), .C(clk), .Q(
        pmem_twlb[0]) );
  SDFFQX1 r_twlb_reg_1_ ( .D(n645), .SIN(pmem_twlb[0]), .SMC(test_se), .C(clk), 
        .Q(pmem_twlb[1]) );
  SDFFQX1 wspp_cnt_reg_5_ ( .D(N800), .SIN(wspp_cnt_4_), .SMC(test_se), .C(
        net11846), .Q(wspp_cnt_5_) );
  SDFFQX1 wspp_cnt_reg_3_ ( .D(N798), .SIN(wspp_cnt_2_), .SMC(test_se), .C(
        net11846), .Q(wspp_cnt_3_) );
  SDFFQX1 c_buf_reg_0__5_ ( .D(N484), .SIN(rd_buf[4]), .SMC(test_se), .C(
        net11977), .Q(rd_buf[5]) );
  SDFFQX1 c_buf_reg_3__5_ ( .D(N508), .SIN(dbg_03[4]), .SMC(test_se), .C(
        net11962), .Q(dbg_03[5]) );
  SDFFQX1 c_buf_reg_6__5_ ( .D(N532), .SIN(dbg_06[4]), .SMC(test_se), .C(
        net11947), .Q(dbg_06[5]) );
  SDFFQX1 c_buf_reg_5__5_ ( .D(N524), .SIN(dbg_05[4]), .SMC(test_se), .C(
        net11952), .Q(dbg_05[5]) );
  SDFFQX1 c_buf_reg_2__5_ ( .D(N500), .SIN(dbg_02[4]), .SMC(test_se), .C(
        net11967), .Q(dbg_02[5]) );
  SDFFQX1 c_buf_reg_4__5_ ( .D(N516), .SIN(dbg_04[4]), .SMC(test_se), .C(
        net11957), .Q(dbg_04[5]) );
  SDFFQX1 c_buf_reg_1__5_ ( .D(N492), .SIN(dbg_01[4]), .SMC(test_se), .C(
        net11972), .Q(dbg_01[5]) );
  SDFFQX1 c_buf_reg_8__5_ ( .D(N548), .SIN(dbg_08[4]), .SMC(test_se), .C(
        net11937), .Q(dbg_08[5]) );
  SDFFQX1 c_buf_reg_10__7_ ( .D(N566), .SIN(dbg_0a[6]), .SMC(test_se), .C(
        net11927), .Q(dbg_0a[7]) );
  SDFFQX1 c_buf_reg_7__7_ ( .D(N542), .SIN(dbg_07[6]), .SMC(test_se), .C(
        net11942), .Q(dbg_07[7]) );
  SDFFQX1 c_buf_reg_22__7_ ( .D(N662), .SIN(c_buf_22__6_), .SMC(test_se), .C(
        net11867), .Q(c_buf_22__7_) );
  SDFFQX1 c_buf_reg_21__7_ ( .D(N654), .SIN(c_buf_21__6_), .SMC(test_se), .C(
        net11872), .Q(c_buf_21__7_) );
  SDFFQX1 c_buf_reg_19__7_ ( .D(N638), .SIN(c_buf_19__6_), .SMC(test_se), .C(
        net11882), .Q(c_buf_19__7_) );
  SDFFQX1 c_buf_reg_18__7_ ( .D(N630), .SIN(c_buf_18__6_), .SMC(test_se), .C(
        net11887), .Q(c_buf_18__7_) );
  SDFFQX1 c_buf_reg_23__7_ ( .D(N793), .SIN(wr_buf[6]), .SMC(test_se), .C(
        net11862), .Q(wr_buf[7]) );
  SDFFQX1 wspp_cnt_reg_4_ ( .D(N799), .SIN(wspp_cnt_3_), .SMC(test_se), .C(
        net11846), .Q(wspp_cnt_4_) );
  SDFFQX1 c_buf_reg_0__7_ ( .D(N486), .SIN(rd_buf[6]), .SMC(test_se), .C(
        net11977), .Q(rd_buf[7]) );
  SDFFQX1 c_buf_reg_5__7_ ( .D(N526), .SIN(dbg_05[6]), .SMC(test_se), .C(
        net11952), .Q(dbg_05[7]) );
  SDFFQX1 c_buf_reg_2__7_ ( .D(N502), .SIN(dbg_02[6]), .SMC(test_se), .C(
        net11967), .Q(dbg_02[7]) );
  SDFFQX1 c_buf_reg_3__7_ ( .D(N510), .SIN(dbg_03[6]), .SMC(test_se), .C(
        net11962), .Q(dbg_03[7]) );
  SDFFQX1 c_buf_reg_4__7_ ( .D(N518), .SIN(dbg_04[6]), .SMC(test_se), .C(
        net11957), .Q(dbg_04[7]) );
  SDFFQX1 c_buf_reg_1__7_ ( .D(N494), .SIN(dbg_01[6]), .SMC(test_se), .C(
        net11972), .Q(dbg_01[7]) );
  SDFFQX1 c_buf_reg_6__7_ ( .D(N534), .SIN(dbg_06[6]), .SMC(test_se), .C(
        net11947), .Q(dbg_06[7]) );
  SDFFQX1 c_buf_reg_11__7_ ( .D(N574), .SIN(dbg_0b[6]), .SMC(test_se), .C(
        net11922), .Q(dbg_0b[7]) );
  SDFFQX1 c_buf_reg_8__7_ ( .D(N550), .SIN(dbg_08[6]), .SMC(test_se), .C(
        net11937), .Q(dbg_08[7]) );
  SDFFQX1 c_buf_reg_20__7_ ( .D(N646), .SIN(c_buf_20__6_), .SMC(test_se), .C(
        net11877), .Q(c_buf_20__7_) );
  SDFFQX1 c_buf_reg_9__7_ ( .D(N558), .SIN(dbg_09[6]), .SMC(test_se), .C(
        net11932), .Q(dbg_09[7]) );
  SDFFQX1 r_rdy_reg ( .D(n648), .SIN(pmem_pgm), .SMC(test_se), .C(clk), .Q(
        r_rdy) );
  SDFFQX1 cs_ft_reg_2_ ( .D(N823), .SIN(cs_ft[1]), .SMC(test_se), .C(net11992), 
        .Q(cs_ft[2]) );
  SDFFQX1 cs_ft_reg_3_ ( .D(N824), .SIN(cs_ft[2]), .SMC(test_se), .C(net11992), 
        .Q(cs_ft[3]) );
  SDFFQX1 c_adr_reg_4_ ( .D(N830), .SIN(c_adr[3]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[4]) );
  SDFFQX1 c_adr_reg_2_ ( .D(N828), .SIN(c_adr[1]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[2]) );
  SDFFQX1 c_adr_reg_3_ ( .D(N829), .SIN(c_adr[2]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[3]) );
  SDFFQX1 cs_ft_reg_1_ ( .D(N822), .SIN(cs_ft[0]), .SMC(test_se), .C(net11992), 
        .Q(cs_ft[1]) );
  SDFFQX1 cs_ft_reg_0_ ( .D(N821), .SIN(c_ptr[4]), .SMC(test_se), .C(net11992), 
        .Q(cs_ft[0]) );
  SDFFQX1 c_adr_reg_1_ ( .D(N827), .SIN(c_adr[0]), .SMC(test_se), .C(net11987), 
        .Q(c_adr[1]) );
  SDFFQX1 c_adr_reg_0_ ( .D(N826), .SIN(adr_p[14]), .SMC(test_se), .C(net11987), .Q(c_adr[0]) );
  SDFFNQXL ck_n_reg_1_ ( .D(n642), .SIN(pmem_clk[0]), .SMC(test_se), .XC(clk), 
        .Q(pmem_clk[1]) );
  SDFFNQXL ck_n_reg_0_ ( .D(n641), .SIN(test_si1), .SMC(test_se), .XC(clk), 
        .Q(pmem_clk[0]) );
  SDFFNQX1 cs_n_reg ( .D(n643), .SIN(pmem_clk[1]), .SMC(test_se), .XC(clk), 
        .Q(test_so1) );
  SDFFQX2 adr_p_reg_0_ ( .D(N854), .SIN(pmem_a[8]), .SMC(test_se), .C(net11857), .Q(pmem_a[0]) );
  SDFFQX2 a_bit_reg_1_ ( .D(n705), .SIN(pmem_a[6]), .SMC(test_se), .C(net11852), .Q(pmem_a[7]) );
  AO21X1 U3 ( .B(n134), .C(c_adr[8]), .A(c_adr[9]), .Y(n132) );
  NAND21X1 U4 ( .B(pwrdn_rst), .A(n84), .Y(n61) );
  NOR21XL U5 ( .B(n618), .A(n28), .Y(n642) );
  AO21X1 U6 ( .B(n661), .C(n622), .A(n621), .Y(n647) );
  INVXL U7 ( .A(n665), .Y(n1) );
  INVXL U8 ( .A(n1), .Y(n2) );
  INVX1 U9 ( .A(n604), .Y(n3) );
  INVX1 U10 ( .A(n604), .Y(n4) );
  INVX1 U11 ( .A(n596), .Y(n5) );
  INVX1 U12 ( .A(n601), .Y(n6) );
  INVX1 U13 ( .A(n601), .Y(n7) );
  INVX1 U14 ( .A(n611), .Y(n8) );
  INVX1 U15 ( .A(n600), .Y(n9) );
  INVX1 U16 ( .A(n600), .Y(n10) );
  INVX1 U17 ( .A(n599), .Y(n11) );
  INVX1 U18 ( .A(n599), .Y(n12) );
  INVX1 U19 ( .A(n673), .Y(n13) );
  BUFX3 U20 ( .A(n657), .Y(n14) );
  INVX1 U21 ( .A(n607), .Y(n15) );
  INVX1 U22 ( .A(n598), .Y(n16) );
  INVX1 U23 ( .A(n598), .Y(n17) );
  INVX1 U24 ( .A(n656), .Y(n18) );
  NAND21X1 U25 ( .B(pwrdn_rst), .A(n84), .Y(n656) );
  INVX1 U26 ( .A(n679), .Y(n19) );
  INVX1 U27 ( .A(n572), .Y(n20) );
  INVX1 U28 ( .A(n572), .Y(n21) );
  INVX1 U29 ( .A(n431), .Y(n22) );
  NAND2X1 U30 ( .A(n541), .B(n602), .Y(n45) );
  INVX1 U31 ( .A(n45), .Y(n23) );
  INVX1 U32 ( .A(n45), .Y(n24) );
  INVX1 U33 ( .A(n45), .Y(n25) );
  INVX1 U34 ( .A(n571), .Y(n26) );
  INVX1 U35 ( .A(n571), .Y(n27) );
  AOI211XL U36 ( .C(memaddr_c[0]), .D(n411), .A(n410), .B(n409), .Y(n424) );
  OA22XL U37 ( .A(memaddr_c[0]), .B(n411), .C(memaddr_c[1]), .D(n140), .Y(n145) );
  AOI21XL U38 ( .B(memaddr_c[5]), .C(n657), .A(n60), .Y(n34) );
  OA22XL U39 ( .A(memaddr_c[1]), .B(n686), .C(memaddr_c[0]), .D(n685), .Y(n96)
         );
  NAND2XL U40 ( .A(n153), .B(memaddr_c[5]), .Y(n416) );
  AND2X1 U41 ( .A(n618), .B(n500), .Y(n641) );
  AOI21X1 U42 ( .B(n499), .C(n490), .A(n489), .Y(n28) );
  NAND21XL U43 ( .B(c_adr[3]), .A(memaddr_c[3]), .Y(n91) );
  INVX1 U44 ( .A(n460), .Y(n62) );
  INVX1 U45 ( .A(n460), .Y(n63) );
  INVX1 U46 ( .A(n460), .Y(n578) );
  INVX1 U47 ( .A(n401), .Y(n690) );
  NAND21X1 U48 ( .B(n577), .A(n64), .Y(n460) );
  AOI21X1 U49 ( .B(n592), .C(we_twlb), .A(N853), .Y(n29) );
  INVX1 U50 ( .A(n82), .Y(n76) );
  INVX1 U51 ( .A(n82), .Y(n74) );
  INVX1 U52 ( .A(n82), .Y(n75) );
  INVX1 U53 ( .A(n82), .Y(n73) );
  INVX1 U54 ( .A(n515), .Y(n71) );
  INVX1 U55 ( .A(n515), .Y(n70) );
  INVX1 U56 ( .A(n82), .Y(n69) );
  INVX1 U57 ( .A(n82), .Y(n68) );
  INVX1 U58 ( .A(n515), .Y(n67) );
  INVX1 U59 ( .A(n82), .Y(n72) );
  INVX1 U60 ( .A(n82), .Y(n65) );
  INVX1 U61 ( .A(n515), .Y(n66) );
  INVX1 U62 ( .A(n515), .Y(n77) );
  INVX1 U63 ( .A(n82), .Y(n80) );
  INVX1 U64 ( .A(n515), .Y(n78) );
  INVX1 U65 ( .A(n515), .Y(n79) );
  INVX1 U66 ( .A(n515), .Y(n81) );
  INVX1 U67 ( .A(n510), .Y(n438) );
  NAND21X1 U68 ( .B(n573), .A(n592), .Y(n436) );
  INVX1 U69 ( .A(n522), .Y(n584) );
  INVX1 U70 ( .A(n622), .Y(n662) );
  NAND21X1 U71 ( .B(n612), .A(n661), .Y(n557) );
  AND2X1 U72 ( .A(n367), .B(n372), .Y(n281) );
  INVX1 U73 ( .A(n577), .Y(n525) );
  AND2X1 U74 ( .A(n374), .B(n367), .Y(n291) );
  INVX1 U75 ( .A(n574), .Y(n661) );
  INVX1 U76 ( .A(n575), .Y(n615) );
  NAND21X1 U77 ( .B(n574), .A(n573), .Y(n575) );
  NOR2X1 U78 ( .A(dw_rst), .B(n83), .Y(n401) );
  INVX1 U79 ( .A(n84), .Y(n83) );
  NAND21X1 U80 ( .B(n62), .A(n634), .Y(n665) );
  NAND6XL U81 ( .A(n427), .B(n426), .C(n425), .D(n424), .E(n423), .F(n422), 
        .Y(n437) );
  INVX1 U82 ( .A(n407), .Y(n425) );
  AND4X1 U83 ( .A(n421), .B(n420), .C(n419), .D(n418), .Y(n422) );
  AND4X1 U84 ( .A(n417), .B(n416), .C(n415), .D(n414), .Y(n423) );
  INVX1 U85 ( .A(n656), .Y(n618) );
  INVX1 U86 ( .A(n82), .Y(n64) );
  INVX1 U87 ( .A(n629), .Y(n82) );
  INVX1 U88 ( .A(n431), .Y(n659) );
  NAND21X1 U89 ( .B(n412), .A(n64), .Y(n431) );
  NAND32X1 U90 ( .B(n659), .C(n464), .A(n510), .Y(N853) );
  AO21X1 U91 ( .B(n445), .C(n457), .A(n63), .Y(N878) );
  AO21X1 U92 ( .B(n445), .C(n639), .A(n63), .Y(N881) );
  AO21X1 U93 ( .B(n449), .C(n457), .A(n63), .Y(N882) );
  AO21X1 U94 ( .B(n449), .C(n639), .A(n63), .Y(N885) );
  AO21X1 U95 ( .B(n46), .C(n457), .A(n63), .Y(N886) );
  AO21X1 U96 ( .B(n46), .C(n639), .A(n62), .Y(N889) );
  AO21X1 U97 ( .B(n458), .C(n457), .A(n62), .Y(N894) );
  INVX1 U98 ( .A(n462), .Y(n458) );
  NAND21X1 U99 ( .B(n566), .A(n504), .Y(n510) );
  OAI211X1 U100 ( .C(n617), .D(n491), .A(n503), .B(n506), .Y(n536) );
  AO21X1 U101 ( .B(n438), .C(n437), .A(n464), .Y(n93) );
  INVX1 U102 ( .A(n634), .Y(n655) );
  INVX1 U103 ( .A(n414), .Y(n172) );
  INVX1 U104 ( .A(n427), .Y(n161) );
  INVX1 U105 ( .A(n420), .Y(n171) );
  INVX1 U106 ( .A(n617), .Y(n619) );
  NAND32X1 U107 ( .B(n574), .C(n459), .A(n589), .Y(n522) );
  INVX1 U108 ( .A(n459), .Y(n612) );
  INVX1 U109 ( .A(n631), .Y(n592) );
  INVX1 U110 ( .A(n413), .Y(n417) );
  AO21X1 U111 ( .B(n676), .C(n459), .A(n630), .Y(n622) );
  NAND2X1 U112 ( .A(n363), .B(n365), .Y(n270) );
  NAND2X1 U113 ( .A(n368), .B(n366), .Y(n273) );
  NAND2X1 U114 ( .A(n363), .B(n366), .Y(n269) );
  NAND2X1 U115 ( .A(n368), .B(n364), .Y(n272) );
  NAND2X1 U116 ( .A(n368), .B(n367), .Y(n275) );
  NAND2X1 U117 ( .A(n363), .B(n364), .Y(n271) );
  NAND2X1 U118 ( .A(n363), .B(n367), .Y(n274) );
  NAND2X1 U119 ( .A(n368), .B(n365), .Y(n277) );
  AND2X1 U120 ( .A(n373), .B(n366), .Y(n289) );
  AND2X1 U121 ( .A(n364), .B(n373), .Y(n290) );
  NOR2X1 U122 ( .A(n692), .B(n695), .Y(n372) );
  NAND2X1 U123 ( .A(n366), .B(n372), .Y(n284) );
  NAND2X1 U124 ( .A(n369), .B(n364), .Y(n276) );
  NAND2X1 U125 ( .A(n369), .B(n367), .Y(n279) );
  NAND2X1 U126 ( .A(n373), .B(n367), .Y(n287) );
  NAND2X1 U127 ( .A(n373), .B(n365), .Y(n286) );
  NAND2X1 U128 ( .A(n369), .B(n366), .Y(n280) );
  NAND2X1 U129 ( .A(n364), .B(n372), .Y(n288) );
  NAND2X1 U130 ( .A(n365), .B(n372), .Y(n285) );
  AND2X1 U131 ( .A(n374), .B(n364), .Y(n294) );
  AND2X1 U132 ( .A(n374), .B(n365), .Y(n292) );
  AND2X1 U133 ( .A(n374), .B(n366), .Y(n293) );
  NOR2X1 U134 ( .A(n697), .B(n696), .Y(n367) );
  NAND2X1 U135 ( .A(n369), .B(n365), .Y(n278) );
  NOR2X1 U136 ( .A(n693), .B(n695), .Y(n374) );
  NAND21X1 U137 ( .B(n60), .A(n676), .Y(n574) );
  INVX1 U138 ( .A(n583), .Y(n597) );
  INVX1 U139 ( .A(n596), .Y(n667) );
  INVX1 U140 ( .A(n589), .Y(n573) );
  INVX1 U141 ( .A(n250), .Y(o_ofs_inc) );
  INVX1 U142 ( .A(srst), .Y(n84) );
  INVX1 U143 ( .A(n150), .Y(n151) );
  INVX1 U144 ( .A(n130), .Y(n169) );
  INVX1 U145 ( .A(n210), .Y(n243) );
  INVX1 U146 ( .A(n242), .Y(n245) );
  INVX1 U147 ( .A(n412), .Y(n673) );
  INVX1 U148 ( .A(n475), .Y(n482) );
  NAND21X1 U149 ( .B(n490), .A(n484), .Y(n475) );
  INVX1 U150 ( .A(n453), .Y(n674) );
  INVX1 U151 ( .A(n491), .Y(n620) );
  INVX1 U152 ( .A(n529), .Y(n508) );
  NOR2X1 U153 ( .A(n668), .B(n674), .Y(n554) );
  INVX1 U154 ( .A(n506), .Y(n507) );
  INVX1 U155 ( .A(n637), .Y(n652) );
  GEN2XL U156 ( .D(memaddr_c[1]), .E(n686), .C(n96), .B(n95), .A(n100), .Y(n97) );
  INVX1 U157 ( .A(n90), .Y(n100) );
  NAND21X1 U158 ( .B(n566), .A(n564), .Y(n617) );
  OA222X1 U159 ( .A(n145), .B(n413), .C(memaddr_c[3]), .D(n144), .E(
        memaddr_c[2]), .F(n143), .Y(n152) );
  INVX1 U160 ( .A(n142), .Y(n143) );
  INVX1 U161 ( .A(n148), .Y(n144) );
  NAND32X1 U162 ( .B(n433), .C(n617), .A(n432), .Y(n579) );
  INVX1 U163 ( .A(n437), .Y(n433) );
  OAI22X1 U164 ( .A(n150), .B(n149), .C(n148), .D(n147), .Y(n407) );
  INVX1 U165 ( .A(memaddr_c[3]), .Y(n147) );
  INVXL U166 ( .A(memaddr_c[4]), .Y(n149) );
  AO22AXL U167 ( .A(n140), .B(memaddr_c[1]), .C(memaddr_c[2]), .D(n142), .Y(
        n413) );
  OAI2B11X1 U168 ( .D(n432), .C(n561), .A(n518), .B(n564), .Y(n519) );
  OA222X1 U169 ( .A(memaddr_c[8]), .B(n159), .C(n158), .D(n157), .E(
        memaddr_c[7]), .F(n156), .Y(n160) );
  INVX1 U170 ( .A(n419), .Y(n158) );
  AOI32X1 U171 ( .A(n415), .B(n416), .C(n155), .D(n51), .E(n154), .Y(n157) );
  AO21X1 U172 ( .B(n408), .C(n606), .A(n409), .Y(n179) );
  NAND2X1 U173 ( .A(n30), .B(n91), .Y(n95) );
  OAI22XL U174 ( .A(memaddr_c[2]), .B(n684), .C(memaddr_c[3]), .D(n683), .Y(
        n30) );
  INVX1 U175 ( .A(n515), .Y(n629) );
  XOR2X1 U176 ( .A(memaddr_c[14]), .B(n408), .Y(n410) );
  OA21X1 U177 ( .B(memaddr_c[10]), .C(n167), .A(n166), .Y(n173) );
  AOI32X1 U178 ( .A(n418), .B(n421), .C(n165), .D(n57), .E(n164), .Y(n166) );
  INVX1 U179 ( .A(memaddr_c[11]), .Y(n164) );
  OAI22X1 U180 ( .A(memaddr_c[9]), .B(n162), .C(n161), .D(n160), .Y(n165) );
  INVX1 U181 ( .A(n429), .Y(n561) );
  NAND32X1 U182 ( .B(n487), .C(n437), .A(n428), .Y(n429) );
  INVX1 U183 ( .A(n513), .Y(n566) );
  INVX1 U184 ( .A(n177), .Y(n409) );
  OAI211X1 U185 ( .C(n408), .D(n606), .A(n426), .B(n176), .Y(n177) );
  AO21X1 U186 ( .B(n59), .C(n175), .A(n174), .Y(n176) );
  OAI32X1 U187 ( .A(n173), .B(n172), .C(n171), .D(memaddr_c[12]), .E(n170), 
        .Y(n174) );
  INVX1 U188 ( .A(n664), .Y(n607) );
  OR2X1 U189 ( .A(n577), .B(n576), .Y(n634) );
  OAI211X1 U190 ( .C(n412), .D(n576), .A(n436), .B(n435), .Y(n464) );
  INVX1 U191 ( .A(n91), .Y(n94) );
  AND2XL U192 ( .A(memaddr_c[4]), .B(n99), .Y(n92) );
  NAND2X1 U193 ( .A(n156), .B(memaddr_c[7]), .Y(n419) );
  NAND21X1 U194 ( .B(n511), .A(n456), .Y(n462) );
  NAND41X1 U195 ( .D(n22), .A(n31), .B(n501), .C(n18), .Y(N825) );
  NAND3X1 U196 ( .A(n438), .B(n679), .C(n437), .Y(n31) );
  INVX1 U197 ( .A(n571), .Y(n595) );
  NAND21X1 U198 ( .B(n603), .A(n539), .Y(n571) );
  INVX1 U199 ( .A(n572), .Y(n623) );
  NAND21X1 U200 ( .B(n603), .A(n543), .Y(n572) );
  INVX1 U201 ( .A(n599), .Y(n625) );
  NAND21X1 U202 ( .B(n603), .A(n551), .Y(n599) );
  INVX1 U203 ( .A(n600), .Y(n626) );
  NAND21X1 U204 ( .B(n603), .A(n549), .Y(n600) );
  INVX1 U205 ( .A(n601), .Y(n627) );
  NAND21X1 U206 ( .B(n603), .A(n547), .Y(n601) );
  INVX1 U207 ( .A(n598), .Y(n624) );
  NAND21X1 U208 ( .B(n603), .A(n553), .Y(n598) );
  INVX1 U209 ( .A(n604), .Y(n628) );
  NAND21X1 U210 ( .B(n603), .A(n545), .Y(n604) );
  OAI21BBX1 U211 ( .A(N432), .B(n659), .C(n32), .Y(N827) );
  AOI21X1 U212 ( .B(memaddr_c[1]), .C(n657), .A(n60), .Y(n32) );
  OAI21BBX1 U213 ( .A(N434), .B(n659), .C(n33), .Y(N829) );
  AOI21X1 U214 ( .B(memaddr_c[3]), .C(n657), .A(n60), .Y(n33) );
  OAI21BBX1 U215 ( .A(N436), .B(n659), .C(n34), .Y(N831) );
  OAI21BBX1 U216 ( .A(N438), .B(n22), .C(n35), .Y(N833) );
  AOI21XL U217 ( .B(memaddr_c[7]), .C(n14), .A(n61), .Y(n35) );
  OAI21BBX1 U218 ( .A(N440), .B(n659), .C(n36), .Y(N835) );
  AOI21X1 U219 ( .B(memaddr_c[9]), .C(n657), .A(n60), .Y(n36) );
  OAI21BBX1 U220 ( .A(N442), .B(n659), .C(n37), .Y(N837) );
  AOI21X1 U221 ( .B(memaddr_c[11]), .C(n657), .A(n60), .Y(n37) );
  OAI21BBX1 U222 ( .A(N444), .B(n22), .C(n38), .Y(N839) );
  AOI21XL U223 ( .B(memaddr_c[13]), .C(n14), .A(n61), .Y(n38) );
  OAI21BBX1 U224 ( .A(N443), .B(n659), .C(n39), .Y(N838) );
  AOI21X1 U225 ( .B(memaddr_c[12]), .C(n657), .A(n60), .Y(n39) );
  OAI21BBX1 U226 ( .A(N433), .B(n659), .C(n40), .Y(N828) );
  AOI21XL U227 ( .B(memaddr_c[2]), .C(n657), .A(n60), .Y(n40) );
  OAI21BBX1 U228 ( .A(N435), .B(n22), .C(n41), .Y(N830) );
  AOI21XL U229 ( .B(memaddr_c[4]), .C(n14), .A(n61), .Y(n41) );
  OAI21BBX1 U230 ( .A(N437), .B(n22), .C(n42), .Y(N832) );
  AOI21XL U231 ( .B(memaddr_c[6]), .C(n14), .A(n60), .Y(n42) );
  OAI21BBX1 U232 ( .A(N441), .B(n22), .C(n43), .Y(N836) );
  AOI21XL U233 ( .B(memaddr_c[10]), .C(n14), .A(n61), .Y(n43) );
  OAI21BBX1 U234 ( .A(N439), .B(n22), .C(n44), .Y(N834) );
  AOI21XL U235 ( .B(memaddr_c[8]), .C(n14), .A(n61), .Y(n44) );
  AO21X1 U236 ( .B(n445), .C(n636), .A(n63), .Y(N879) );
  AO21X1 U237 ( .B(n445), .C(n635), .A(n63), .Y(N880) );
  AO21X1 U238 ( .B(n449), .C(n636), .A(n63), .Y(N883) );
  AO21X1 U239 ( .B(n449), .C(n635), .A(n63), .Y(N884) );
  AO21X1 U240 ( .B(n46), .C(n636), .A(n63), .Y(N887) );
  AO21X1 U241 ( .B(n46), .C(n635), .A(n62), .Y(N888) );
  AO21X1 U242 ( .B(n455), .C(n457), .A(n62), .Y(N890) );
  AO21X1 U243 ( .B(n455), .C(n636), .A(n62), .Y(N891) );
  AO21X1 U244 ( .B(n455), .C(n635), .A(n62), .Y(N892) );
  AO21X1 U245 ( .B(n455), .C(n639), .A(n62), .Y(N893) );
  AO21X1 U246 ( .B(n636), .C(n458), .A(n62), .Y(N895) );
  AO21X1 U247 ( .B(n635), .C(n458), .A(n62), .Y(N896) );
  AO21X1 U248 ( .B(n443), .C(n457), .A(n578), .Y(N874) );
  AO21X1 U249 ( .B(n443), .C(n639), .A(n578), .Y(N877) );
  AO21X1 U250 ( .B(n443), .C(n636), .A(n578), .Y(N875) );
  AO21X1 U251 ( .B(n443), .C(n635), .A(n578), .Y(N876) );
  INVX1 U252 ( .A(n602), .Y(n603) );
  OAI211X1 U253 ( .C(n463), .D(n462), .A(n471), .B(n461), .Y(N897) );
  AND2X1 U254 ( .A(n522), .B(n460), .Y(n461) );
  NAND21X1 U255 ( .B(n57), .A(memaddr_c[11]), .Y(n414) );
  NAND2X1 U256 ( .A(n159), .B(memaddr_c[8]), .Y(n427) );
  NAND21X1 U257 ( .B(n504), .A(n501), .Y(n657) );
  NAND2X1 U258 ( .A(n170), .B(memaddr_c[12]), .Y(n420) );
  OA21X1 U259 ( .B(n636), .C(n635), .A(n655), .Y(N843) );
  INVX1 U260 ( .A(memaddr_c[9]), .Y(n89) );
  INVX1 U261 ( .A(n444), .Y(n445) );
  NAND32X1 U262 ( .B(n511), .C(n450), .A(n451), .Y(n444) );
  INVX1 U263 ( .A(n447), .Y(n449) );
  NAND32X1 U264 ( .B(n451), .C(n450), .A(n511), .Y(n447) );
  NOR3XL U265 ( .A(n511), .B(n451), .C(n450), .Y(n46) );
  INVX1 U266 ( .A(n111), .Y(n108) );
  AND2X1 U267 ( .A(n655), .B(n680), .Y(N842) );
  NAND2X1 U268 ( .A(n162), .B(memaddr_c[9]), .Y(n418) );
  NAND21X1 U269 ( .B(n59), .A(memaddr_c[13]), .Y(n426) );
  NAND2X1 U270 ( .A(n167), .B(memaddr_c[10]), .Y(n421) );
  INVX1 U271 ( .A(memaddr_c[13]), .Y(n175) );
  NAND6XL U272 ( .A(n13), .B(n581), .C(n197), .D(n560), .E(n436), .F(n196), 
        .Y(N820) );
  AOI33X1 U273 ( .A(n620), .B(n660), .C(n521), .D(n55), .E(n672), .F(n670), 
        .Y(n196) );
  AND3X1 U274 ( .A(n187), .B(n662), .C(n674), .Y(n197) );
  INVX1 U275 ( .A(n536), .Y(n187) );
  INVX1 U276 ( .A(memaddr_c[14]), .Y(n606) );
  INVX1 U277 ( .A(n219), .Y(n124) );
  AO21X1 U278 ( .B(sfr_psr), .C(n194), .A(n564), .Y(n459) );
  NAND21X1 U279 ( .B(n192), .A(n612), .Y(n631) );
  XNOR3X1 U280 ( .A(n230), .B(n229), .C(memaddr_c[3]), .Y(n234) );
  XOR3X1 U281 ( .A(n226), .B(n225), .C(memaddr_c[1]), .Y(n236) );
  XOR2X1 U282 ( .A(memaddr_c[8]), .B(n246), .Y(n247) );
  AO21X1 U283 ( .B(n584), .C(n687), .A(n597), .Y(n586) );
  XNOR2XL U284 ( .A(n224), .B(n47), .Y(n237) );
  NAND2X1 U285 ( .A(n223), .B(n222), .Y(n47) );
  NOR3XL U286 ( .A(popptr[3]), .B(popptr[4]), .C(popptr[2]), .Y(n363) );
  NOR3XL U287 ( .A(popptr[3]), .B(popptr[4]), .C(n695), .Y(n368) );
  NOR4XL U288 ( .A(n265), .B(n266), .C(n267), .D(n268), .Y(n264) );
  OAI222XL U289 ( .A(n278), .B(n842), .C(n279), .D(n841), .E(n280), .F(n850), 
        .Y(n265) );
  OAI222XL U290 ( .A(n275), .B(n844), .C(n276), .D(n843), .E(n277), .F(n835), 
        .Y(n266) );
  OAI222XL U291 ( .A(n272), .B(n832), .C(n273), .D(n829), .E(n274), .F(n831), 
        .Y(n267) );
  INVX1 U292 ( .A(popptr[2]), .Y(n695) );
  INVX1 U293 ( .A(popptr[3]), .Y(n693) );
  NOR2X1 U294 ( .A(n693), .B(popptr[2]), .Y(n369) );
  INVX1 U295 ( .A(popptr[4]), .Y(n692) );
  NOR2X1 U296 ( .A(n692), .B(popptr[2]), .Y(n373) );
  INVX1 U297 ( .A(n564), .Y(n660) );
  OAI211X1 U298 ( .C(n472), .D(n471), .A(n522), .B(n557), .Y(N898) );
  AND2X1 U299 ( .A(n528), .B(n529), .Y(n472) );
  NAND32X1 U300 ( .B(n87), .C(n183), .A(n428), .Y(n250) );
  INVX1 U301 ( .A(popptr[1]), .Y(n697) );
  NOR2X1 U302 ( .A(n697), .B(n375), .Y(n365) );
  NOR2X1 U303 ( .A(n375), .B(popptr[1]), .Y(n364) );
  NOR2X1 U304 ( .A(n696), .B(popptr[1]), .Y(n366) );
  NOR4XL U305 ( .A(n349), .B(n350), .C(n351), .D(n352), .Y(n348) );
  OAI222XL U306 ( .A(n278), .B(n767), .C(n279), .D(n761), .E(n280), .F(n814), 
        .Y(n349) );
  OAI222XL U307 ( .A(n275), .B(n827), .C(n276), .D(n821), .E(n277), .F(n754), 
        .Y(n350) );
  OAI222XL U308 ( .A(n272), .B(n740), .C(n273), .D(n721), .E(n274), .F(n730), 
        .Y(n351) );
  NOR4XL U309 ( .A(n319), .B(n320), .C(n321), .D(n322), .Y(n318) );
  OAI222XL U310 ( .A(n278), .B(n764), .C(n279), .D(n758), .E(n280), .F(n811), 
        .Y(n319) );
  OAI222XL U311 ( .A(n275), .B(n769), .C(n276), .D(n818), .E(n277), .F(n751), 
        .Y(n320) );
  OAI222XL U312 ( .A(n272), .B(n734), .C(n273), .D(n714), .E(n274), .F(n727), 
        .Y(n321) );
  NOR4XL U313 ( .A(n309), .B(n310), .C(n311), .D(n312), .Y(n308) );
  OAI222XL U314 ( .A(n278), .B(n808), .C(n279), .D(n807), .E(n280), .F(n810), 
        .Y(n309) );
  OAI222XL U315 ( .A(n275), .B(n824), .C(n276), .D(n817), .E(n277), .F(n750), 
        .Y(n310) );
  OAI222XL U316 ( .A(n272), .B(n772), .C(n273), .D(n770), .E(n274), .F(n726), 
        .Y(n311) );
  NOR4XL U317 ( .A(n329), .B(n330), .C(n331), .D(n332), .Y(n328) );
  OAI222XL U318 ( .A(n278), .B(n765), .C(n279), .D(n759), .E(n280), .F(n812), 
        .Y(n329) );
  OAI222XL U319 ( .A(n275), .B(n825), .C(n276), .D(n819), .E(n277), .F(n752), 
        .Y(n330) );
  OAI222XL U320 ( .A(n272), .B(n736), .C(n273), .D(n716), .E(n274), .F(n728), 
        .Y(n331) );
  NOR4XL U321 ( .A(n359), .B(n360), .C(n361), .D(n362), .Y(n358) );
  OAI222XL U322 ( .A(n278), .B(n768), .C(n279), .D(n762), .E(n280), .F(n815), 
        .Y(n359) );
  OAI222XL U323 ( .A(n275), .B(n828), .C(n276), .D(n822), .E(n277), .F(n755), 
        .Y(n360) );
  OAI222XL U324 ( .A(n272), .B(n742), .C(n273), .D(n723), .E(n274), .F(n731), 
        .Y(n361) );
  NOR4XL U325 ( .A(n339), .B(n340), .C(n341), .D(n342), .Y(n338) );
  OAI222XL U326 ( .A(n278), .B(n766), .C(n279), .D(n760), .E(n280), .F(n813), 
        .Y(n339) );
  OAI222XL U327 ( .A(n275), .B(n826), .C(n276), .D(n820), .E(n277), .F(n753), 
        .Y(n340) );
  OAI222XL U328 ( .A(n272), .B(n738), .C(n273), .D(n719), .E(n274), .F(n729), 
        .Y(n341) );
  NOR4XL U329 ( .A(n299), .B(n300), .C(n301), .D(n302), .Y(n298) );
  OAI222XL U330 ( .A(n278), .B(n763), .C(n279), .D(n806), .E(n280), .F(n809), 
        .Y(n299) );
  OAI222XL U331 ( .A(n275), .B(n823), .C(n276), .D(n816), .E(n277), .F(n749), 
        .Y(n300) );
  OAI222XL U332 ( .A(n272), .B(n732), .C(n273), .D(n712), .E(n274), .F(n725), 
        .Y(n301) );
  INVX1 U333 ( .A(n375), .Y(n696) );
  NAND21X1 U334 ( .B(n687), .A(n661), .Y(n596) );
  NAND21XL U335 ( .B(pwrdn_rst), .A(n84), .Y(n60) );
  INVX1 U336 ( .A(n609), .Y(n587) );
  INVX1 U337 ( .A(n580), .Y(n567) );
  AO21X1 U338 ( .B(n661), .C(n687), .A(n597), .Y(n666) );
  NAND21X1 U339 ( .B(n184), .A(n86), .Y(n529) );
  NAND32X1 U340 ( .B(n428), .C(n184), .A(n183), .Y(n506) );
  AO21XL U341 ( .B(n852), .C(n674), .A(n61), .Y(n523) );
  NAND2X1 U342 ( .A(n560), .B(n852), .Y(n495) );
  NAND2X1 U343 ( .A(n487), .B(n529), .Y(n496) );
  INVX1 U344 ( .A(n483), .Y(n490) );
  ENOX1 U345 ( .A(n250), .B(n679), .C(n679), .D(sfr_psr), .Y(sfr_psrack) );
  NAND2X1 U346 ( .A(n48), .B(n193), .Y(n589) );
  NAND4X1 U347 ( .A(sfr_psw), .B(n678), .C(n194), .D(n677), .Y(n48) );
  NAND32X1 U348 ( .B(n183), .C(n184), .A(n428), .Y(n491) );
  NAND21X1 U349 ( .B(n428), .A(n185), .Y(n503) );
  AOI21BBXL U350 ( .B(n49), .C(n50), .A(n60), .Y(N899) );
  AOI21X1 U351 ( .B(n687), .C(n473), .A(n674), .Y(n49) );
  AOI21X1 U352 ( .B(n55), .C(n670), .A(n852), .Y(n50) );
  INVX1 U353 ( .A(n400), .Y(n689) );
  AO21X1 U354 ( .B(n135), .C(n207), .A(n134), .Y(n156) );
  AO21X1 U355 ( .B(n141), .C(n203), .A(n202), .Y(n146) );
  AO21X1 U356 ( .B(n675), .C(n199), .A(n198), .Y(n139) );
  NOR2X1 U357 ( .A(n685), .B(n680), .Y(n675) );
  AO21X1 U358 ( .B(n201), .C(n139), .A(n200), .Y(n141) );
  AOI21AX1 U359 ( .B(n136), .C(n206), .A(n135), .Y(n51) );
  INVX1 U360 ( .A(n133), .Y(n134) );
  AOI21X1 U361 ( .B(n146), .C(n205), .A(n204), .Y(n52) );
  NAND32X1 U362 ( .B(n246), .C(n208), .A(n134), .Y(n131) );
  AO21X1 U363 ( .B(n131), .C(n209), .A(n168), .Y(n167) );
  OR2X1 U364 ( .A(n163), .B(n211), .Y(n130) );
  XNOR2XL U365 ( .A(n228), .B(n139), .Y(n142) );
  XNOR2XL U366 ( .A(n232), .B(n146), .Y(n150) );
  XNOR2XL U367 ( .A(n230), .B(n141), .Y(n148) );
  XOR2X1 U368 ( .A(n138), .B(n226), .Y(n140) );
  INVX1 U369 ( .A(n163), .Y(n168) );
  INVX1 U370 ( .A(n137), .Y(n226) );
  NAND21X1 U371 ( .B(n198), .A(n199), .Y(n137) );
  NAND2X1 U372 ( .A(n138), .B(n225), .Y(n411) );
  AO21X1 U373 ( .B(n231), .C(n205), .A(n204), .Y(n216) );
  OR2X1 U374 ( .A(n209), .B(n224), .Y(n210) );
  NAND32X1 U375 ( .B(n246), .C(n207), .A(n245), .Y(n241) );
  NAND21X1 U376 ( .B(n211), .A(n243), .Y(n217) );
  AO21X1 U377 ( .B(n227), .C(n201), .A(n200), .Y(n229) );
  AO21X1 U378 ( .B(n225), .C(n199), .A(n198), .Y(n227) );
  AO21X1 U379 ( .B(n229), .C(n203), .A(n202), .Y(n231) );
  OR2X1 U380 ( .A(n208), .B(n241), .Y(n224) );
  OR2X1 U381 ( .A(n206), .B(n212), .Y(n242) );
  AND3X1 U382 ( .A(o_inst[2]), .B(o_inst[4]), .C(o_inst[3]), .Y(n258) );
  AO21X1 U383 ( .B(n184), .C(n87), .A(n188), .Y(n412) );
  NAND21X1 U384 ( .B(n687), .A(hit_ps), .Y(n193) );
  INVX1 U385 ( .A(n430), .Y(n457) );
  INVX1 U386 ( .A(n434), .Y(n518) );
  NAND21X1 U387 ( .B(n679), .A(n504), .Y(n582) );
  NAND21X1 U388 ( .B(n194), .A(n193), .Y(n521) );
  INVX1 U389 ( .A(n581), .Y(n504) );
  INVX1 U390 ( .A(n498), .Y(n484) );
  NOR21XL U391 ( .B(r_hold_mcu), .A(n83), .Y(n801) );
  INVX1 U392 ( .A(n192), .Y(n676) );
  NAND21X1 U393 ( .B(n508), .A(n493), .Y(n453) );
  NAND21X1 U394 ( .B(n620), .A(n560), .Y(n568) );
  INVX1 U395 ( .A(n691), .Y(n669) );
  INVX1 U396 ( .A(n528), .Y(n668) );
  NAND21X1 U397 ( .B(n511), .A(n639), .Y(n637) );
  INVX1 U398 ( .A(n463), .Y(n639) );
  NAND2X1 U399 ( .A(n676), .B(n687), .Y(n537) );
  INVX1 U400 ( .A(n709), .Y(n671) );
  INVX1 U401 ( .A(n534), .Y(n708) );
  INVX1 U402 ( .A(n533), .Y(n707) );
  INVX1 U403 ( .A(n852), .Y(n672) );
  NAND31X1 U404 ( .C(o_ofs_inc), .A(test_so1), .B(n491), .Y(n492) );
  GEN2XL U405 ( .D(c_adr[8]), .E(n113), .C(n112), .B(n111), .A(n110), .Y(n114)
         );
  INVX1 U406 ( .A(memaddr_c[8]), .Y(n113) );
  AND2X1 U407 ( .A(c_adr[9]), .B(n89), .Y(n112) );
  AOI211X1 U408 ( .C(memaddr_c[8]), .D(n246), .A(n109), .B(n108), .Y(n110) );
  AO2222XL U409 ( .A(memaddr[13]), .B(n667), .C(sfr_psofs[13]), .D(n666), .E(
        pre_1_adr[13]), .F(n665), .G(memaddr_c[13]), .H(n664), .Y(N867) );
  AO2222XL U410 ( .A(memaddr[12]), .B(n667), .C(sfr_psofs[12]), .D(n666), .E(
        pre_1_adr[12]), .F(n2), .G(memaddr_c[12]), .H(n664), .Y(N866) );
  AO2222XL U411 ( .A(memaddr[11]), .B(n667), .C(sfr_psofs[11]), .D(n666), .E(
        pre_1_adr[11]), .F(n665), .G(memaddr_c[11]), .H(n664), .Y(N865) );
  AO2222XL U412 ( .A(memaddr[10]), .B(n667), .C(sfr_psofs[10]), .D(n666), .E(
        pre_1_adr[10]), .F(n2), .G(memaddr_c[10]), .H(n664), .Y(N864) );
  AO2222XL U413 ( .A(memaddr[9]), .B(n667), .C(sfr_psofs[9]), .D(n666), .E(
        pre_1_adr[9]), .F(n665), .G(memaddr_c[9]), .H(n664), .Y(N863) );
  AO2222XL U414 ( .A(memaddr[8]), .B(n667), .C(sfr_psofs[8]), .D(n666), .E(
        pre_1_adr[8]), .F(n2), .G(memaddr_c[8]), .H(n664), .Y(N862) );
  AO2222XL U415 ( .A(memaddr[7]), .B(n667), .C(sfr_psofs[7]), .D(n666), .E(
        pre_1_adr[7]), .F(n665), .G(memaddr_c[7]), .H(n664), .Y(N861) );
  AO2222XL U416 ( .A(memaddr[5]), .B(n667), .C(sfr_psofs[5]), .D(n666), .E(
        pre_1_adr[5]), .F(n2), .G(memaddr_c[5]), .H(n664), .Y(N859) );
  AO2222XL U417 ( .A(memaddr[3]), .B(n667), .C(sfr_psofs[3]), .D(n666), .E(
        pre_1_adr[3]), .F(n665), .G(memaddr_c[3]), .H(n15), .Y(N857) );
  AO2222XL U418 ( .A(memaddr[1]), .B(n667), .C(sfr_psofs[1]), .D(n8), .E(
        pre_1_adr[1]), .F(n2), .G(memaddr_c[1]), .H(n15), .Y(N855) );
  AO2222XL U419 ( .A(memaddr[0]), .B(n5), .C(sfr_psofs[0]), .D(n8), .E(
        pre_1_adr[0]), .F(n2), .G(memaddr_c[0]), .H(n15), .Y(N854) );
  OR2X1 U420 ( .A(d_psrd), .B(n519), .Y(n515) );
  OAI211X1 U421 ( .C(n181), .D(n180), .A(n179), .B(n178), .Y(n513) );
  NAND43X1 U422 ( .B(c_ptr[2]), .C(c_ptr[3]), .D(c_ptr[4]), .A(n457), .Y(n178)
         );
  INVX1 U423 ( .A(n218), .Y(n181) );
  AOI211X1 U424 ( .C(c_adr[13]), .D(n175), .A(n124), .B(n123), .Y(n180) );
  OAI221X1 U425 ( .A(n118), .B(n222), .C(memaddr_c[11]), .D(n117), .E(n116), 
        .Y(n119) );
  INVX1 U426 ( .A(c_adr[11]), .Y(n117) );
  NAND32X1 U427 ( .B(n115), .C(n118), .A(n114), .Y(n116) );
  INVX1 U428 ( .A(n223), .Y(n115) );
  NAND2X1 U429 ( .A(n2), .B(pre_1_adr[14]), .Y(n605) );
  AO21X1 U430 ( .B(n594), .C(n615), .A(n593), .Y(n645) );
  AND3X1 U431 ( .A(wd_twlb[1]), .B(we_twlb), .C(n612), .Y(n594) );
  MUX2X1 U432 ( .D0(n613), .D1(pmem_twlb[1]), .S(n29), .Y(n593) );
  AO21X1 U433 ( .B(n616), .C(n615), .A(n614), .Y(n646) );
  AND3X1 U434 ( .A(wd_twlb[0]), .B(we_twlb), .C(n612), .Y(n616) );
  MUX2X1 U435 ( .D0(n613), .D1(pmem_twlb[0]), .S(n29), .Y(n614) );
  OA21X1 U436 ( .B(c_adr[13]), .C(n175), .A(n122), .Y(n123) );
  OAI22X1 U437 ( .A(memaddr_c[12]), .B(n121), .C(n120), .D(n129), .Y(n122) );
  AND2X1 U438 ( .A(n120), .B(n129), .Y(n121) );
  INVX1 U439 ( .A(n119), .Y(n120) );
  OAI211X1 U440 ( .C(pre_1_adr[13]), .D(n605), .A(n591), .B(n590), .Y(n613) );
  AOI33X1 U441 ( .A(n589), .B(n588), .C(n587), .D(sfr_psofs[14]), .E(n586), 
        .F(n585), .Y(n590) );
  NAND32XL U442 ( .B(memaddr_c[13]), .C(n606), .A(n664), .Y(n591) );
  INVX1 U443 ( .A(sfr_psofs[13]), .Y(n585) );
  AOI21X1 U444 ( .B(c_adr[7]), .C(n107), .A(n106), .Y(n109) );
  INVX1 U445 ( .A(memaddr_c[7]), .Y(n107) );
  GEN2XL U446 ( .D(c_adr[5]), .E(n105), .C(n104), .B(n103), .A(n102), .Y(n106)
         );
  INVXL U447 ( .A(memaddr_c[5]), .Y(n105) );
  OAI31XL U448 ( .A(n496), .B(n495), .C(n488), .D(n506), .Y(n489) );
  INVX1 U449 ( .A(pmem_clk[1]), .Y(n488) );
  AO21X1 U450 ( .B(n499), .C(n498), .A(n497), .Y(n500) );
  OAI31XL U451 ( .A(n496), .B(n495), .C(n494), .D(n506), .Y(n497) );
  INVX1 U452 ( .A(pmem_clk[0]), .Y(n494) );
  OAI211X1 U453 ( .C(n611), .D(n610), .A(n609), .B(n608), .Y(N868) );
  INVX1 U454 ( .A(sfr_psofs[14]), .Y(n610) );
  INVX1 U455 ( .A(n666), .Y(n611) );
  OA21X1 U456 ( .B(n607), .C(n606), .A(n605), .Y(n608) );
  NAND32X1 U457 ( .B(d_psrd), .C(n579), .A(n673), .Y(n501) );
  NAND21XL U458 ( .B(c_adr[5]), .A(memaddr_c[5]), .Y(n90) );
  NAND31X1 U459 ( .C(d_psrd), .A(n579), .B(n434), .Y(n576) );
  NAND21X1 U460 ( .B(d_psrd), .A(n576), .Y(n602) );
  NAND21X1 U461 ( .B(c_adr[7]), .A(memaddr_c[7]), .Y(n101) );
  AO21X1 U462 ( .B(n64), .C(dbg_0a[7]), .A(n595), .Y(N558) );
  AO21X1 U463 ( .B(dbg_0d[7]), .C(n629), .A(n26), .Y(N582) );
  AO21X1 U464 ( .B(dbg_0e[7]), .C(n629), .A(n27), .Y(N590) );
  AO21X1 U465 ( .B(c_buf_16__7_), .C(n629), .A(n595), .Y(N606) );
  AO21X1 U466 ( .B(c_buf_17__7_), .C(n629), .A(n26), .Y(N614) );
  AO21X1 U467 ( .B(n77), .C(c_buf_18__7_), .A(n27), .Y(N622) );
  AO21X1 U468 ( .B(n77), .C(c_buf_19__7_), .A(n595), .Y(N630) );
  AO21X1 U469 ( .B(n74), .C(c_buf_20__7_), .A(n26), .Y(N638) );
  AO21X1 U470 ( .B(n76), .C(c_buf_21__7_), .A(n27), .Y(N646) );
  AO21X1 U471 ( .B(n75), .C(c_buf_22__7_), .A(n595), .Y(N654) );
  AO21X1 U472 ( .B(wr_buf[7]), .C(n629), .A(n26), .Y(N662) );
  AO21X1 U473 ( .B(n76), .C(dbg_08[7]), .A(n27), .Y(N542) );
  AO21X1 U474 ( .B(n76), .C(dbg_09[7]), .A(n595), .Y(N550) );
  AO21X1 U475 ( .B(n74), .C(dbg_0b[7]), .A(n26), .Y(N566) );
  AO21X1 U476 ( .B(dbg_0c[7]), .C(n81), .A(n27), .Y(N574) );
  AO21X1 U477 ( .B(dbg_0f[7]), .C(n81), .A(n595), .Y(N598) );
  AO21X1 U478 ( .B(c_buf_17__5_), .C(n81), .A(n623), .Y(N612) );
  AO21X1 U479 ( .B(n74), .C(c_buf_19__5_), .A(n20), .Y(N628) );
  AO21X1 U480 ( .B(n76), .C(c_buf_20__5_), .A(n21), .Y(N636) );
  AO21X1 U481 ( .B(n74), .C(c_buf_22__5_), .A(n623), .Y(N652) );
  AO21X1 U482 ( .B(n73), .C(wr_buf[5]), .A(n20), .Y(N660) );
  AO21X1 U483 ( .B(n76), .C(dbg_07[7]), .A(n26), .Y(N534) );
  AO21X1 U484 ( .B(n74), .C(dbg_01[7]), .A(n27), .Y(N486) );
  AO21X1 U485 ( .B(n76), .C(dbg_02[7]), .A(n595), .Y(N494) );
  AO21X1 U486 ( .B(n76), .C(dbg_05[7]), .A(n26), .Y(N518) );
  AO21X1 U487 ( .B(n73), .C(dbg_04[7]), .A(n27), .Y(N510) );
  AO21X1 U488 ( .B(n76), .C(dbg_03[7]), .A(n595), .Y(N502) );
  AO21X1 U489 ( .B(n76), .C(dbg_06[7]), .A(n26), .Y(N526) );
  AO21X1 U490 ( .B(n74), .C(dbg_08[0]), .A(n624), .Y(N535) );
  AO21X1 U491 ( .B(n76), .C(dbg_08[1]), .A(n625), .Y(N536) );
  AO21X1 U492 ( .B(n75), .C(dbg_08[2]), .A(n626), .Y(N537) );
  AO21X1 U493 ( .B(n74), .C(dbg_08[3]), .A(n627), .Y(N538) );
  AO21X1 U494 ( .B(n75), .C(dbg_08[5]), .A(n21), .Y(N540) );
  AO21X1 U495 ( .B(n73), .C(dbg_08[6]), .A(n24), .Y(N541) );
  AO21X1 U496 ( .B(n74), .C(dbg_09[0]), .A(n16), .Y(N543) );
  AO21X1 U497 ( .B(n75), .C(dbg_09[1]), .A(n11), .Y(N544) );
  AO21X1 U498 ( .B(n75), .C(dbg_09[2]), .A(n9), .Y(N545) );
  AO21X1 U499 ( .B(n74), .C(dbg_09[3]), .A(n6), .Y(N546) );
  AO21X1 U500 ( .B(n75), .C(dbg_09[4]), .A(n628), .Y(N547) );
  AO21X1 U501 ( .B(n74), .C(dbg_09[5]), .A(n623), .Y(N548) );
  AO21X1 U502 ( .B(n73), .C(dbg_09[6]), .A(n25), .Y(N549) );
  AO21X1 U503 ( .B(n73), .C(dbg_0a[0]), .A(n17), .Y(N551) );
  AO21X1 U504 ( .B(n75), .C(dbg_0a[1]), .A(n12), .Y(N552) );
  AO21X1 U505 ( .B(n73), .C(dbg_0a[2]), .A(n10), .Y(N553) );
  AO21X1 U506 ( .B(n73), .C(dbg_0a[3]), .A(n7), .Y(N554) );
  AO21X1 U507 ( .B(n75), .C(dbg_0a[4]), .A(n3), .Y(N555) );
  AO21X1 U508 ( .B(n75), .C(dbg_0a[5]), .A(n20), .Y(N556) );
  AO21X1 U509 ( .B(n73), .C(dbg_0a[6]), .A(n24), .Y(N557) );
  AO21X1 U510 ( .B(n75), .C(dbg_0b[5]), .A(n21), .Y(N564) );
  AO21X1 U511 ( .B(dbg_0c[5]), .C(n79), .A(n623), .Y(N572) );
  AO21X1 U512 ( .B(dbg_0c[6]), .C(n81), .A(n25), .Y(N573) );
  AO21X1 U513 ( .B(dbg_0d[0]), .C(n79), .A(n624), .Y(N575) );
  AO21X1 U514 ( .B(dbg_0d[1]), .C(n81), .A(n625), .Y(N576) );
  AO21X1 U515 ( .B(dbg_0d[2]), .C(n81), .A(n626), .Y(N577) );
  AO21X1 U516 ( .B(dbg_0d[3]), .C(n79), .A(n627), .Y(N578) );
  AO21X1 U517 ( .B(dbg_0d[4]), .C(n78), .A(n4), .Y(N579) );
  AO21X1 U518 ( .B(dbg_0d[5]), .C(n81), .A(n20), .Y(N580) );
  AO21X1 U519 ( .B(dbg_0d[6]), .C(n78), .A(n23), .Y(N581) );
  AO21X1 U520 ( .B(dbg_0e[0]), .C(n78), .A(n16), .Y(N583) );
  AO21X1 U521 ( .B(dbg_0e[1]), .C(n78), .A(n11), .Y(N584) );
  AO21X1 U522 ( .B(dbg_0e[2]), .C(n80), .A(n9), .Y(N585) );
  AO21X1 U523 ( .B(dbg_0e[3]), .C(n78), .A(n6), .Y(N586) );
  AO21X1 U524 ( .B(dbg_0e[4]), .C(n78), .A(n628), .Y(N587) );
  AO21X1 U525 ( .B(dbg_0e[5]), .C(n80), .A(n21), .Y(N588) );
  AO21X1 U526 ( .B(dbg_0e[6]), .C(n78), .A(n23), .Y(N589) );
  AO21X1 U527 ( .B(dbg_0f[0]), .C(n78), .A(n17), .Y(N591) );
  AO21X1 U528 ( .B(dbg_0f[1]), .C(n80), .A(n12), .Y(N592) );
  AO21X1 U529 ( .B(dbg_0f[2]), .C(n80), .A(n10), .Y(N593) );
  AO21X1 U530 ( .B(dbg_0f[3]), .C(n77), .A(n7), .Y(N594) );
  AO21X1 U531 ( .B(dbg_0f[4]), .C(n80), .A(n3), .Y(N595) );
  AO21X1 U532 ( .B(dbg_0f[5]), .C(n77), .A(n623), .Y(N596) );
  AO21X1 U533 ( .B(dbg_0f[6]), .C(n80), .A(n23), .Y(N597) );
  AO21X1 U534 ( .B(c_buf_16__0_), .C(n80), .A(n624), .Y(N599) );
  AO21X1 U535 ( .B(c_buf_16__1_), .C(n77), .A(n625), .Y(N600) );
  AO21X1 U536 ( .B(c_buf_16__2_), .C(n77), .A(n626), .Y(N601) );
  AO21X1 U537 ( .B(c_buf_16__3_), .C(n79), .A(n627), .Y(N602) );
  AO21X1 U538 ( .B(c_buf_16__4_), .C(n77), .A(n4), .Y(N603) );
  AO21X1 U539 ( .B(c_buf_16__5_), .C(n80), .A(n20), .Y(N604) );
  AO21X1 U540 ( .B(c_buf_16__6_), .C(n79), .A(n23), .Y(N605) );
  AO21X1 U541 ( .B(c_buf_17__0_), .C(n81), .A(n16), .Y(N607) );
  AO21X1 U542 ( .B(c_buf_17__1_), .C(n77), .A(n11), .Y(N608) );
  AO21X1 U543 ( .B(c_buf_17__2_), .C(n79), .A(n9), .Y(N609) );
  AO21X1 U544 ( .B(c_buf_17__3_), .C(n77), .A(n6), .Y(N610) );
  AO21X1 U545 ( .B(c_buf_17__4_), .C(n77), .A(n628), .Y(N611) );
  AO21X1 U546 ( .B(c_buf_17__6_), .C(n79), .A(n23), .Y(N613) );
  AO21X1 U547 ( .B(n73), .C(c_buf_18__0_), .A(n17), .Y(N615) );
  AO21X1 U548 ( .B(n73), .C(c_buf_18__1_), .A(n12), .Y(N616) );
  AO21X1 U549 ( .B(n72), .C(c_buf_18__2_), .A(n10), .Y(N617) );
  AO21X1 U550 ( .B(n72), .C(c_buf_18__3_), .A(n7), .Y(N618) );
  AO21X1 U551 ( .B(n72), .C(c_buf_18__4_), .A(n3), .Y(N619) );
  AO21X1 U552 ( .B(n72), .C(c_buf_18__5_), .A(n21), .Y(N620) );
  AO21X1 U553 ( .B(n72), .C(c_buf_18__6_), .A(n25), .Y(N621) );
  AO21X1 U554 ( .B(n72), .C(c_buf_19__0_), .A(n624), .Y(N623) );
  AO21X1 U555 ( .B(n72), .C(c_buf_19__1_), .A(n625), .Y(N624) );
  AO21X1 U556 ( .B(n72), .C(c_buf_19__2_), .A(n626), .Y(N625) );
  AO21X1 U557 ( .B(n72), .C(c_buf_19__3_), .A(n627), .Y(N626) );
  AO21X1 U558 ( .B(n71), .C(c_buf_19__4_), .A(n4), .Y(N627) );
  AO21X1 U559 ( .B(n71), .C(c_buf_19__6_), .A(n24), .Y(N629) );
  AO21X1 U560 ( .B(n71), .C(c_buf_20__0_), .A(n16), .Y(N631) );
  AO21X1 U561 ( .B(n71), .C(c_buf_20__1_), .A(n11), .Y(N632) );
  AO21X1 U562 ( .B(n71), .C(c_buf_20__2_), .A(n9), .Y(N633) );
  AO21X1 U563 ( .B(n71), .C(c_buf_20__3_), .A(n6), .Y(N634) );
  AO21X1 U564 ( .B(n71), .C(c_buf_20__4_), .A(n628), .Y(N635) );
  AO21X1 U565 ( .B(n71), .C(c_buf_20__6_), .A(n25), .Y(N637) );
  AO21X1 U566 ( .B(n71), .C(c_buf_21__0_), .A(n17), .Y(N639) );
  AO21X1 U567 ( .B(n71), .C(c_buf_21__1_), .A(n12), .Y(N640) );
  AO21X1 U568 ( .B(n70), .C(c_buf_21__2_), .A(n10), .Y(N641) );
  AO21X1 U569 ( .B(n70), .C(c_buf_21__3_), .A(n7), .Y(N642) );
  AO21X1 U570 ( .B(n70), .C(c_buf_21__4_), .A(n3), .Y(N643) );
  AO21X1 U571 ( .B(n70), .C(c_buf_21__5_), .A(n623), .Y(N644) );
  AO21X1 U572 ( .B(n70), .C(c_buf_21__6_), .A(n24), .Y(N645) );
  AO21X1 U573 ( .B(n70), .C(c_buf_22__0_), .A(n624), .Y(N647) );
  AO21X1 U574 ( .B(n70), .C(c_buf_22__1_), .A(n625), .Y(N648) );
  AO21X1 U575 ( .B(n70), .C(c_buf_22__2_), .A(n626), .Y(N649) );
  AO21X1 U576 ( .B(n70), .C(c_buf_22__3_), .A(n627), .Y(N650) );
  AO21X1 U577 ( .B(n70), .C(c_buf_22__4_), .A(n4), .Y(N651) );
  AO21X1 U578 ( .B(n69), .C(c_buf_22__6_), .A(n25), .Y(N653) );
  AO21X1 U579 ( .B(wr_buf[0]), .C(n80), .A(n16), .Y(N655) );
  AO21X1 U580 ( .B(n69), .C(wr_buf[1]), .A(n11), .Y(N656) );
  AO21X1 U581 ( .B(wr_buf[2]), .C(n81), .A(n9), .Y(N657) );
  AO21X1 U582 ( .B(wr_buf[3]), .C(n80), .A(n6), .Y(N658) );
  AO21X1 U583 ( .B(wr_buf[4]), .C(n78), .A(n628), .Y(N659) );
  AO21X1 U584 ( .B(wr_buf[6]), .C(n78), .A(n23), .Y(N661) );
  AO21X1 U585 ( .B(n69), .C(dbg_02[5]), .A(n20), .Y(N492) );
  AO21X1 U586 ( .B(n69), .C(dbg_05[5]), .A(n21), .Y(N516) );
  AO21X1 U587 ( .B(n69), .C(dbg_03[5]), .A(n623), .Y(N500) );
  AO21X1 U588 ( .B(n69), .C(dbg_06[5]), .A(n20), .Y(N524) );
  AO21X1 U589 ( .B(n69), .C(dbg_08[4]), .A(n3), .Y(N539) );
  AO21X1 U590 ( .B(n69), .C(dbg_0b[0]), .A(n17), .Y(N559) );
  AO21X1 U591 ( .B(n69), .C(dbg_0b[1]), .A(n12), .Y(N560) );
  AO21X1 U592 ( .B(n69), .C(dbg_0b[2]), .A(n10), .Y(N561) );
  AO21X1 U593 ( .B(n68), .C(dbg_0b[3]), .A(n7), .Y(N562) );
  AO21X1 U594 ( .B(n68), .C(dbg_0b[4]), .A(n4), .Y(N563) );
  AO21X1 U595 ( .B(n68), .C(dbg_0b[6]), .A(n24), .Y(N565) );
  AO21X1 U596 ( .B(dbg_0c[0]), .C(n79), .A(n624), .Y(N567) );
  AO21X1 U597 ( .B(dbg_0c[1]), .C(n629), .A(n625), .Y(N568) );
  AO21X1 U598 ( .B(dbg_0c[2]), .C(n79), .A(n626), .Y(N569) );
  AO21X1 U599 ( .B(dbg_0c[3]), .C(n79), .A(n627), .Y(N570) );
  AO21X1 U600 ( .B(dbg_0c[4]), .C(n81), .A(n628), .Y(N571) );
  AO21X1 U601 ( .B(n68), .C(dbg_01[0]), .A(n16), .Y(N479) );
  AO21X1 U602 ( .B(n68), .C(dbg_01[4]), .A(n3), .Y(N483) );
  AO21X1 U603 ( .B(n68), .C(dbg_07[0]), .A(n17), .Y(N527) );
  AO21X1 U604 ( .B(n68), .C(dbg_07[1]), .A(n11), .Y(N528) );
  AO21X1 U605 ( .B(n68), .C(dbg_07[2]), .A(n9), .Y(N529) );
  AO21X1 U606 ( .B(n68), .C(dbg_07[3]), .A(n6), .Y(N530) );
  AO21X1 U607 ( .B(n68), .C(dbg_07[4]), .A(n4), .Y(N531) );
  AO21X1 U608 ( .B(n67), .C(dbg_07[5]), .A(n21), .Y(N532) );
  AO21X1 U609 ( .B(n67), .C(dbg_07[6]), .A(n25), .Y(N533) );
  AO21X1 U610 ( .B(n67), .C(dbg_01[1]), .A(n12), .Y(N480) );
  AO21X1 U611 ( .B(n67), .C(dbg_01[2]), .A(n10), .Y(N481) );
  AO21X1 U612 ( .B(n67), .C(dbg_01[3]), .A(n7), .Y(N482) );
  AO21X1 U613 ( .B(n67), .C(dbg_01[5]), .A(n623), .Y(N484) );
  AO21X1 U614 ( .B(n67), .C(dbg_01[6]), .A(n23), .Y(N485) );
  AO21X1 U615 ( .B(n67), .C(dbg_02[0]), .A(n624), .Y(N487) );
  AO21X1 U616 ( .B(n67), .C(dbg_05[0]), .A(n16), .Y(N511) );
  AO21X1 U617 ( .B(n67), .C(dbg_02[1]), .A(n625), .Y(N488) );
  AO21X1 U618 ( .B(n66), .C(dbg_05[1]), .A(n11), .Y(N512) );
  AO21X1 U619 ( .B(n66), .C(dbg_02[2]), .A(n626), .Y(N489) );
  AO21X1 U620 ( .B(n66), .C(dbg_05[2]), .A(n9), .Y(N513) );
  AO21X1 U621 ( .B(n66), .C(dbg_02[3]), .A(n627), .Y(N490) );
  AO21X1 U622 ( .B(n72), .C(dbg_05[3]), .A(n6), .Y(N514) );
  AO21X1 U623 ( .B(n66), .C(dbg_02[4]), .A(n628), .Y(N491) );
  AO21X1 U624 ( .B(n66), .C(dbg_05[4]), .A(n3), .Y(N515) );
  AO21X1 U625 ( .B(n66), .C(dbg_02[6]), .A(n24), .Y(N493) );
  AO21X1 U626 ( .B(n66), .C(dbg_05[6]), .A(n25), .Y(N517) );
  AO21X1 U627 ( .B(n66), .C(dbg_04[0]), .A(n17), .Y(N503) );
  AO21X1 U628 ( .B(n65), .C(dbg_04[1]), .A(n12), .Y(N504) );
  AO21X1 U629 ( .B(n65), .C(dbg_04[2]), .A(n10), .Y(N505) );
  AO21X1 U630 ( .B(n65), .C(dbg_04[3]), .A(n7), .Y(N506) );
  AO21X1 U631 ( .B(n65), .C(dbg_04[4]), .A(n4), .Y(N507) );
  AO21X1 U632 ( .B(n65), .C(dbg_04[5]), .A(n20), .Y(N508) );
  AO21X1 U633 ( .B(n65), .C(dbg_04[6]), .A(n24), .Y(N509) );
  AO21X1 U634 ( .B(n65), .C(dbg_03[0]), .A(n624), .Y(N495) );
  AO21X1 U635 ( .B(n65), .C(dbg_06[0]), .A(n16), .Y(N519) );
  AO21X1 U636 ( .B(n65), .C(dbg_03[1]), .A(n625), .Y(N496) );
  AO21X1 U637 ( .B(n65), .C(dbg_06[1]), .A(n11), .Y(N520) );
  AO21X1 U638 ( .B(n64), .C(dbg_03[2]), .A(n626), .Y(N497) );
  AO21X1 U639 ( .B(n64), .C(dbg_06[2]), .A(n9), .Y(N521) );
  AO21X1 U640 ( .B(n64), .C(dbg_03[3]), .A(n627), .Y(N498) );
  AO21X1 U641 ( .B(n64), .C(dbg_06[3]), .A(n6), .Y(N522) );
  AO21X1 U642 ( .B(n64), .C(dbg_03[4]), .A(n628), .Y(N499) );
  AO21X1 U643 ( .B(n64), .C(dbg_06[4]), .A(n3), .Y(N523) );
  AO21X1 U644 ( .B(n64), .C(dbg_03[6]), .A(n25), .Y(N501) );
  AO21X1 U645 ( .B(n66), .C(dbg_06[6]), .A(n24), .Y(N525) );
  AO21X1 U646 ( .B(N431), .C(n659), .A(n502), .Y(N826) );
  AO21X1 U647 ( .B(N445), .C(n659), .A(n658), .Y(N840) );
  OA21X1 U648 ( .B(c_adr[6]), .C(n154), .A(n101), .Y(n103) );
  INVX1 U649 ( .A(n452), .Y(n456) );
  NAND43X1 U650 ( .B(c_ptr[3]), .C(n603), .D(n512), .A(n525), .Y(n452) );
  AND3X1 U651 ( .A(c_adr[6]), .B(n154), .C(n101), .Y(n102) );
  OAI21X1 U652 ( .B(n517), .C(n61), .A(n516), .Y(N822) );
  AND4X1 U653 ( .A(n510), .B(n582), .C(n560), .D(n509), .Y(n517) );
  GEN2XL U654 ( .D(n603), .E(n515), .C(n514), .B(n617), .A(n577), .Y(n516) );
  AOI221XL U655 ( .A(n508), .B(mcu_psw), .C(n668), .D(n669), .E(n507), .Y(n509) );
  INVX1 U656 ( .A(n454), .Y(n455) );
  NAND21X1 U657 ( .B(c_ptr[2]), .A(n456), .Y(n454) );
  AND2X1 U658 ( .A(n561), .B(n567), .Y(n565) );
  INVX1 U659 ( .A(n568), .Y(n562) );
  NAND32X1 U660 ( .B(c_ptr[4]), .C(n577), .A(n602), .Y(n450) );
  NAND21X1 U661 ( .B(c_adr[9]), .A(memaddr_c[9]), .Y(n111) );
  INVX1 U662 ( .A(n557), .Y(n558) );
  NAND32X1 U663 ( .B(n672), .C(n536), .A(n530), .Y(n559) );
  AOI32X1 U664 ( .A(n529), .B(mcu_psw), .C(n453), .D(n528), .E(n669), .Y(n530)
         );
  GEN2XL U665 ( .D(n527), .E(n526), .C(n19), .B(n525), .A(n524), .Y(N824) );
  NAND21X1 U666 ( .B(n584), .A(n523), .Y(n524) );
  AND3X1 U667 ( .A(n518), .B(cs_ft[0]), .C(n617), .Y(n527) );
  OA21X1 U668 ( .B(r_pwdn_en), .C(n521), .A(n519), .Y(n526) );
  INVX1 U669 ( .A(n439), .Y(n443) );
  NAND32X1 U670 ( .B(c_ptr[3]), .C(n450), .A(n511), .Y(n439) );
  INVX1 U671 ( .A(n88), .Y(n118) );
  NAND21X1 U672 ( .B(c_adr[11]), .A(memaddr_c[11]), .Y(n88) );
  AND2X1 U673 ( .A(n655), .B(n654), .Y(N846) );
  XOR2X1 U674 ( .A(c_ptr[4]), .B(n653), .Y(n654) );
  AND2X1 U675 ( .A(n652), .B(c_ptr[3]), .Y(n653) );
  AND2X1 U676 ( .A(n638), .B(n655), .Y(N845) );
  XOR2X1 U677 ( .A(c_ptr[3]), .B(n652), .Y(n638) );
  AND2X1 U678 ( .A(n640), .B(n655), .Y(N844) );
  XOR2X1 U679 ( .A(c_ptr[2]), .B(n639), .Y(n640) );
  INVX1 U680 ( .A(test_so1), .Y(pmem_csb) );
  NAND21X1 U681 ( .B(c_adr[10]), .A(memaddr_c[10]), .Y(n223) );
  NAND21X1 U682 ( .B(memaddr_c[10]), .A(c_adr[10]), .Y(n222) );
  MUX2IX1 U683 ( .D0(n53), .D1(n54), .S(n620), .Y(n621) );
  NAND2X1 U684 ( .A(pmem_re), .B(n662), .Y(n53) );
  NAND2XL U685 ( .A(n619), .B(n618), .Y(n54) );
  NOR5X1 U686 ( .A(c_ptr[3]), .B(n513), .C(n637), .D(n19), .E(n512), .Y(n514)
         );
  NAND42X1 U687 ( .C(n406), .D(n405), .A(n404), .B(n403), .Y(n432) );
  NOR32XL U688 ( .B(n402), .C(n399), .A(n398), .Y(n403) );
  XNOR3X1 U689 ( .A(c_adr[11]), .B(n210), .C(memaddr_c[11]), .Y(n406) );
  NOR8XL U690 ( .A(n240), .B(n239), .C(n238), .D(n237), .E(n236), .F(n235), 
        .G(n234), .H(n233), .Y(n404) );
  NAND31X1 U691 ( .C(n215), .A(n214), .B(n213), .Y(n405) );
  NOR32XL U692 ( .B(c_adr[13]), .C(c_adr[14]), .A(n217), .Y(n215) );
  XOR3X1 U693 ( .A(c_adr[13]), .B(n217), .C(memaddr_c[13]), .Y(n213) );
  NAND21X1 U694 ( .B(c_adr[14]), .A(memaddr_c[14]), .Y(n218) );
  NAND21X1 U695 ( .B(memaddr_c[14]), .A(c_adr[14]), .Y(n219) );
  AND2X1 U696 ( .A(hit_ps_c), .B(mcu_psr_c), .Y(n564) );
  NAND21X1 U697 ( .B(n397), .A(n249), .Y(n398) );
  XOR2X1 U698 ( .A(n248), .B(n247), .Y(n249) );
  XOR3X1 U699 ( .A(n244), .B(memaddr_c[12]), .C(c_adr[12]), .Y(n397) );
  AND2X1 U700 ( .A(n245), .B(c_adr[7]), .Y(n248) );
  XOR2X1 U701 ( .A(n221), .B(n220), .Y(n238) );
  NAND21X1 U702 ( .B(n217), .A(c_adr[13]), .Y(n221) );
  AND2X1 U703 ( .A(n219), .B(n218), .Y(n220) );
  XOR3X1 U704 ( .A(c_adr[9]), .B(n241), .C(memaddr_c[9]), .Y(n402) );
  XOR3X1 U705 ( .A(c_adr[7]), .B(n242), .C(memaddr_c[7]), .Y(n399) );
  XNOR3XL U706 ( .A(c_ptr[0]), .B(memaddr_c[0]), .C(c_adr[0]), .Y(n240) );
  XOR3XL U707 ( .A(memaddr_c[5]), .B(c_adr[5]), .C(n216), .Y(n239) );
  XNOR3X1 U708 ( .A(memaddr[4]), .B(c_adr[4]), .C(sub_313_carry[4]), .Y(
        popptr[4]) );
  INVX1 U709 ( .A(memaddr[0]), .Y(n698) );
  OAI222XL U710 ( .A(n269), .B(n833), .C(n270), .D(n830), .E(n271), .F(n834), 
        .Y(n268) );
  INVX1 U711 ( .A(dbg_01[7]), .Y(n833) );
  INVX1 U712 ( .A(dbg_02[7]), .Y(n830) );
  NAND4X1 U713 ( .A(n261), .B(n262), .C(n263), .D(n264), .Y(o_inst[7]) );
  AOI222XL U714 ( .A(dbg_0e[7]), .B(n292), .C(dbg_0d[7]), .D(n293), .E(
        dbg_0c[7]), .F(n294), .Y(n261) );
  AOI222XL U715 ( .A(c_buf_17__7_), .B(n289), .C(c_buf_16__7_), .D(n290), .E(
        dbg_0f[7]), .F(n291), .Y(n262) );
  AOI211X1 U716 ( .C(wr_buf[7]), .D(n281), .A(n282), .B(n283), .Y(n263) );
  NAND2X1 U717 ( .A(c_adr[0]), .B(n698), .Y(sub_313_carry[1]) );
  MUX2X1 U718 ( .D0(n663), .D1(n19), .S(n662), .Y(n649) );
  AND2X1 U719 ( .A(n661), .B(n660), .Y(n663) );
  OAI22X1 U720 ( .A(mcu_psw), .B(n851), .C(n250), .D(n687), .Y(mempsack) );
  OAI222XL U721 ( .A(n286), .B(n849), .C(n287), .D(n848), .E(n288), .F(n847), 
        .Y(n282) );
  INVX1 U722 ( .A(c_buf_18__7_), .Y(n849) );
  INVX1 U723 ( .A(c_buf_19__7_), .Y(n848) );
  INVX1 U724 ( .A(c_buf_20__7_), .Y(n847) );
  MUX2X1 U725 ( .D0(n661), .D1(pmem_pgm), .S(n633), .Y(n644) );
  AND2X1 U726 ( .A(n632), .B(n631), .Y(n633) );
  INVX1 U727 ( .A(n630), .Y(n632) );
  OAI22X1 U728 ( .A(n284), .B(n846), .C(n285), .D(n845), .Y(n283) );
  INVX1 U729 ( .A(c_buf_21__7_), .Y(n846) );
  INVX1 U730 ( .A(c_buf_22__7_), .Y(n845) );
  INVX1 U731 ( .A(c_adr[1]), .Y(n686) );
  NAND21X1 U732 ( .B(cs_ft[0]), .A(cs_ft[1]), .Y(n87) );
  NAND21X1 U733 ( .B(d_psrd), .A(n525), .Y(n580) );
  OAI222XL U734 ( .A(n269), .B(n741), .C(n270), .D(n722), .E(n271), .F(n748), 
        .Y(n352) );
  INVX1 U735 ( .A(dbg_01[1]), .Y(n741) );
  INVX1 U736 ( .A(dbg_02[1]), .Y(n722) );
  OAI222XL U737 ( .A(n269), .B(n735), .C(n270), .D(n715), .E(n271), .F(n756), 
        .Y(n322) );
  INVX1 U738 ( .A(dbg_01[4]), .Y(n735) );
  INVX1 U739 ( .A(dbg_02[4]), .Y(n715) );
  OAI222XL U740 ( .A(n269), .B(n773), .C(n270), .D(n771), .E(n271), .F(n745), 
        .Y(n312) );
  INVX1 U741 ( .A(dbg_01[5]), .Y(n773) );
  INVX1 U742 ( .A(dbg_02[5]), .Y(n771) );
  OAI222XL U743 ( .A(n269), .B(n737), .C(n270), .D(n718), .E(n271), .F(n746), 
        .Y(n332) );
  INVX1 U744 ( .A(dbg_01[3]), .Y(n737) );
  INVX1 U745 ( .A(dbg_02[3]), .Y(n718) );
  OAI222XL U746 ( .A(n269), .B(n743), .C(n270), .D(n724), .E(n271), .F(n757), 
        .Y(n362) );
  INVX1 U747 ( .A(dbg_01[0]), .Y(n743) );
  INVX1 U748 ( .A(dbg_02[0]), .Y(n724) );
  OAI222XL U749 ( .A(n269), .B(n739), .C(n270), .D(n720), .E(n271), .F(n747), 
        .Y(n342) );
  INVX1 U750 ( .A(dbg_01[2]), .Y(n739) );
  INVX1 U751 ( .A(dbg_02[2]), .Y(n720) );
  OAI222XL U752 ( .A(n269), .B(n733), .C(n270), .D(n713), .E(n271), .F(n744), 
        .Y(n302) );
  INVX1 U753 ( .A(dbg_01[6]), .Y(n733) );
  INVX1 U754 ( .A(dbg_02[6]), .Y(n713) );
  OAI222XL U755 ( .A(n286), .B(n804), .C(n287), .D(n797), .E(n288), .F(n791), 
        .Y(n353) );
  INVX1 U756 ( .A(c_buf_18__1_), .Y(n804) );
  INVX1 U757 ( .A(c_buf_19__1_), .Y(n797) );
  INVX1 U758 ( .A(c_buf_20__1_), .Y(n791) );
  OAI222XL U759 ( .A(n286), .B(n800), .C(n287), .D(n794), .E(n288), .F(n788), 
        .Y(n323) );
  INVX1 U760 ( .A(c_buf_18__4_), .Y(n800) );
  INVX1 U761 ( .A(c_buf_19__4_), .Y(n794) );
  INVX1 U762 ( .A(c_buf_20__4_), .Y(n788) );
  OAI222XL U763 ( .A(n286), .B(n840), .C(n287), .D(n839), .E(n288), .F(n787), 
        .Y(n313) );
  INVX1 U764 ( .A(c_buf_18__5_), .Y(n840) );
  INVX1 U765 ( .A(c_buf_19__5_), .Y(n839) );
  INVX1 U766 ( .A(c_buf_20__5_), .Y(n787) );
  OAI222XL U767 ( .A(n286), .B(n802), .C(n287), .D(n795), .E(n288), .F(n789), 
        .Y(n333) );
  INVX1 U768 ( .A(c_buf_18__3_), .Y(n802) );
  INVX1 U769 ( .A(c_buf_19__3_), .Y(n795) );
  INVX1 U770 ( .A(c_buf_20__3_), .Y(n789) );
  OAI222XL U771 ( .A(n286), .B(n805), .C(n287), .D(n798), .E(n288), .F(n792), 
        .Y(n370) );
  INVX1 U772 ( .A(c_buf_18__0_), .Y(n805) );
  INVX1 U773 ( .A(c_buf_19__0_), .Y(n798) );
  INVX1 U774 ( .A(c_buf_20__0_), .Y(n792) );
  OAI222XL U775 ( .A(n286), .B(n803), .C(n287), .D(n796), .E(n288), .F(n790), 
        .Y(n343) );
  INVX1 U776 ( .A(c_buf_18__2_), .Y(n803) );
  INVX1 U777 ( .A(c_buf_19__2_), .Y(n796) );
  INVX1 U778 ( .A(c_buf_20__2_), .Y(n790) );
  OAI222XL U779 ( .A(n286), .B(n799), .C(n287), .D(n793), .E(n288), .F(n786), 
        .Y(n303) );
  INVX1 U780 ( .A(c_buf_18__6_), .Y(n799) );
  INVX1 U781 ( .A(c_buf_19__6_), .Y(n793) );
  INVX1 U782 ( .A(c_buf_20__6_), .Y(n786) );
  OAI22X1 U783 ( .A(n284), .B(n784), .C(n285), .D(n778), .Y(n354) );
  INVX1 U784 ( .A(c_buf_21__1_), .Y(n784) );
  INVX1 U785 ( .A(c_buf_22__1_), .Y(n778) );
  OAI22X1 U786 ( .A(n284), .B(n781), .C(n285), .D(n775), .Y(n324) );
  INVX1 U787 ( .A(c_buf_21__4_), .Y(n781) );
  INVX1 U788 ( .A(c_buf_22__4_), .Y(n775) );
  OAI22X1 U789 ( .A(n284), .B(n838), .C(n285), .D(n837), .Y(n314) );
  INVX1 U790 ( .A(c_buf_21__5_), .Y(n838) );
  INVX1 U791 ( .A(c_buf_22__5_), .Y(n837) );
  OAI22X1 U792 ( .A(n284), .B(n782), .C(n285), .D(n776), .Y(n334) );
  INVX1 U793 ( .A(c_buf_21__3_), .Y(n782) );
  INVX1 U794 ( .A(c_buf_22__3_), .Y(n776) );
  OAI22X1 U795 ( .A(n284), .B(n783), .C(n285), .D(n777), .Y(n344) );
  INVX1 U796 ( .A(c_buf_21__2_), .Y(n783) );
  INVX1 U797 ( .A(c_buf_22__2_), .Y(n777) );
  OAI22X1 U798 ( .A(n284), .B(n780), .C(n285), .D(n774), .Y(n304) );
  INVX1 U799 ( .A(c_buf_21__6_), .Y(n780) );
  INVX1 U800 ( .A(c_buf_22__6_), .Y(n774) );
  INVX1 U801 ( .A(c_adr[2]), .Y(n684) );
  INVX1 U802 ( .A(c_adr[3]), .Y(n683) );
  NAND4X1 U803 ( .A(n295), .B(n296), .C(n297), .D(n298), .Y(o_inst[6]) );
  AOI222XL U804 ( .A(dbg_0e[6]), .B(n292), .C(dbg_0d[6]), .D(n293), .E(
        dbg_0c[6]), .F(n294), .Y(n295) );
  AOI222XL U805 ( .A(c_buf_17__6_), .B(n289), .C(c_buf_16__6_), .D(n290), .E(
        dbg_0f[6]), .F(n291), .Y(n296) );
  AOI211X1 U806 ( .C(wr_buf[6]), .D(n281), .A(n303), .B(n304), .Y(n297) );
  NAND4X1 U807 ( .A(n355), .B(n356), .C(n357), .D(n358), .Y(o_inst[0]) );
  AOI222XL U808 ( .A(dbg_0e[0]), .B(n292), .C(dbg_0d[0]), .D(n293), .E(
        dbg_0c[0]), .F(n294), .Y(n355) );
  AOI222XL U809 ( .A(c_buf_17__0_), .B(n289), .C(c_buf_16__0_), .D(n290), .E(
        dbg_0f[0]), .F(n291), .Y(n356) );
  AOI211X1 U810 ( .C(wr_buf[0]), .D(n281), .A(n370), .B(n371), .Y(n357) );
  NAND4X1 U811 ( .A(n335), .B(n336), .C(n337), .D(n338), .Y(o_inst[2]) );
  AOI222XL U812 ( .A(dbg_0e[2]), .B(n292), .C(dbg_0d[2]), .D(n293), .E(
        dbg_0c[2]), .F(n294), .Y(n335) );
  AOI222XL U813 ( .A(c_buf_17__2_), .B(n289), .C(c_buf_16__2_), .D(n290), .E(
        dbg_0f[2]), .F(n291), .Y(n336) );
  AOI211X1 U814 ( .C(wr_buf[2]), .D(n281), .A(n343), .B(n344), .Y(n337) );
  NAND4X1 U815 ( .A(n305), .B(n306), .C(n307), .D(n308), .Y(o_inst[5]) );
  AOI222XL U816 ( .A(dbg_0e[5]), .B(n292), .C(dbg_0d[5]), .D(n293), .E(
        dbg_0c[5]), .F(n294), .Y(n305) );
  AOI222XL U817 ( .A(c_buf_17__5_), .B(n289), .C(c_buf_16__5_), .D(n290), .E(
        dbg_0f[5]), .F(n291), .Y(n306) );
  AOI211X1 U818 ( .C(wr_buf[5]), .D(n281), .A(n313), .B(n314), .Y(n307) );
  NAND4X1 U819 ( .A(n345), .B(n346), .C(n347), .D(n348), .Y(o_inst[1]) );
  AOI222XL U820 ( .A(dbg_0e[1]), .B(n292), .C(dbg_0d[1]), .D(n293), .E(
        dbg_0c[1]), .F(n294), .Y(n345) );
  AOI222XL U821 ( .A(c_buf_17__1_), .B(n289), .C(c_buf_16__1_), .D(n290), .E(
        dbg_0f[1]), .F(n291), .Y(n346) );
  AOI211X1 U822 ( .C(wr_buf[1]), .D(n281), .A(n353), .B(n354), .Y(n347) );
  NAND4X1 U823 ( .A(n315), .B(n316), .C(n317), .D(n318), .Y(o_inst[4]) );
  AOI222XL U824 ( .A(dbg_0e[4]), .B(n292), .C(dbg_0d[4]), .D(n293), .E(
        dbg_0c[4]), .F(n294), .Y(n315) );
  AOI222XL U825 ( .A(c_buf_17__4_), .B(n289), .C(c_buf_16__4_), .D(n290), .E(
        dbg_0f[4]), .F(n291), .Y(n316) );
  AOI211X1 U826 ( .C(wr_buf[4]), .D(n281), .A(n323), .B(n324), .Y(n317) );
  NAND4X1 U827 ( .A(n325), .B(n326), .C(n327), .D(n328), .Y(o_inst[3]) );
  AOI222XL U828 ( .A(dbg_0e[3]), .B(n292), .C(dbg_0d[3]), .D(n293), .E(
        dbg_0c[3]), .F(n294), .Y(n325) );
  AOI222XL U829 ( .A(c_buf_17__3_), .B(n289), .C(c_buf_16__3_), .D(n290), .E(
        dbg_0f[3]), .F(n291), .Y(n326) );
  AOI211X1 U830 ( .C(wr_buf[3]), .D(n281), .A(n333), .B(n334), .Y(n327) );
  OAI21X1 U831 ( .B(c_adr[0]), .C(n698), .A(sub_313_carry[1]), .Y(n375) );
  INVX1 U832 ( .A(cs_ft[2]), .Y(n428) );
  INVX1 U833 ( .A(mcu_psw), .Y(n687) );
  INVX1 U834 ( .A(cs_ft[3]), .Y(n183) );
  OAI22X1 U835 ( .A(n284), .B(n785), .C(n285), .D(n779), .Y(n371) );
  INVX1 U836 ( .A(c_buf_21__0_), .Y(n785) );
  INVX1 U837 ( .A(c_buf_22__0_), .Y(n779) );
  INVX1 U838 ( .A(r_rdy), .Y(n851) );
  NAND21X1 U839 ( .B(n596), .A(memaddr[14]), .Y(n609) );
  INVX1 U840 ( .A(rd_buf[7]), .Y(n834) );
  INVX1 U841 ( .A(dbg_04[7]), .Y(n832) );
  INVX1 U842 ( .A(dbg_05[7]), .Y(n829) );
  INVX1 U843 ( .A(dbg_08[7]), .Y(n843) );
  INVX1 U844 ( .A(dbg_0b[7]), .Y(n841) );
  INVX1 U845 ( .A(dbg_03[7]), .Y(n831) );
  INVX1 U846 ( .A(dbg_06[7]), .Y(n835) );
  INVX1 U847 ( .A(dbg_09[7]), .Y(n850) );
  NOR4XL U848 ( .A(wspp_cnt_5_), .B(wspp_cnt_3_), .C(wspp_cnt_4_), .D(test_so2), .Y(n55) );
  NAND32X1 U849 ( .B(n504), .C(n520), .A(n503), .Y(n505) );
  OAI31XL U850 ( .A(n691), .B(wr_buf[0]), .C(n668), .D(n852), .Y(n520) );
  INVX1 U851 ( .A(n486), .Y(n499) );
  OAI31XL U852 ( .A(pmem_re), .B(n442), .C(n485), .D(n495), .Y(n486) );
  AOI221XL U853 ( .A(n836), .B(wspp_cnt_5_), .C(n446), .D(test_so2), .E(n55), 
        .Y(n485) );
  OAI21X1 U854 ( .B(n448), .C(wspp_cnt_4_), .A(r_multi), .Y(n442) );
  AOI21BBXL U855 ( .B(wspp_cnt_3_), .C(n55), .A(test_so2), .Y(n448) );
  INVX1 U856 ( .A(rd_buf[5]), .Y(n745) );
  INVX1 U857 ( .A(dbg_04[5]), .Y(n772) );
  INVX1 U858 ( .A(dbg_07[7]), .Y(n844) );
  INVX1 U859 ( .A(dbg_0a[7]), .Y(n842) );
  INVX1 U860 ( .A(dbg_05[5]), .Y(n770) );
  INVX1 U861 ( .A(dbg_08[5]), .Y(n817) );
  INVX1 U862 ( .A(dbg_03[5]), .Y(n726) );
  INVX1 U863 ( .A(dbg_06[5]), .Y(n750) );
  NAND32X1 U864 ( .B(cs_ft[1]), .C(cs_ft[0]), .A(n86), .Y(n852) );
  NAND2X1 U865 ( .A(d_psrd), .B(n834), .Y(d_inst[7]) );
  NAND32X1 U866 ( .B(n191), .C(n190), .A(n189), .Y(n560) );
  INVX1 U867 ( .A(cs_ft[1]), .Y(n191) );
  INVX1 U868 ( .A(n188), .Y(n189) );
  NAND21X1 U869 ( .B(cs_ft[2]), .A(n183), .Y(n188) );
  NAND21X1 U870 ( .B(cs_ft[1]), .A(cs_ft[0]), .Y(n184) );
  XNOR2XL U871 ( .A(wspp_cnt_5_), .B(wspp_cnt_3_), .Y(n446) );
  NOR4XL U872 ( .A(pmem_a[11]), .B(pmem_a[10]), .C(adr_p[13]), .D(n570), .Y(
        n569) );
  OR4X1 U873 ( .A(pmem_a[15]), .B(pmem_a[14]), .C(pmem_a[13]), .D(pmem_a[12]), 
        .Y(n570) );
  MUX2IX1 U874 ( .D0(adr_p[13]), .D1(n474), .S(adr_p[14]), .Y(n483) );
  AND2X1 U875 ( .A(pmem_a[9]), .B(n569), .Y(n474) );
  INVX1 U876 ( .A(n85), .Y(n86) );
  NAND21X1 U877 ( .B(n428), .A(cs_ft[3]), .Y(n85) );
  OR2X1 U878 ( .A(cs_ft[3]), .B(n87), .Y(n487) );
  INVX1 U879 ( .A(cs_ft[0]), .Y(n190) );
  INVX1 U880 ( .A(rd_buf[1]), .Y(n748) );
  INVX1 U881 ( .A(rd_buf[3]), .Y(n746) );
  INVX1 U882 ( .A(rd_buf[2]), .Y(n747) );
  INVX1 U883 ( .A(rd_buf[6]), .Y(n744) );
  INVX1 U884 ( .A(rd_buf[4]), .Y(n756) );
  INVX1 U885 ( .A(rd_buf[0]), .Y(n757) );
  INVX1 U886 ( .A(wspp_cnt_4_), .Y(n836) );
  INVX1 U887 ( .A(dbg_04[1]), .Y(n740) );
  INVX1 U888 ( .A(dbg_07[1]), .Y(n827) );
  INVX1 U889 ( .A(dbg_0a[1]), .Y(n767) );
  INVX1 U890 ( .A(dbg_04[4]), .Y(n734) );
  INVX1 U891 ( .A(dbg_07[4]), .Y(n769) );
  INVX1 U892 ( .A(dbg_0a[4]), .Y(n764) );
  INVX1 U893 ( .A(dbg_07[5]), .Y(n824) );
  INVX1 U894 ( .A(dbg_0a[5]), .Y(n808) );
  INVX1 U895 ( .A(dbg_04[3]), .Y(n736) );
  INVX1 U896 ( .A(dbg_07[3]), .Y(n825) );
  INVX1 U897 ( .A(dbg_0a[3]), .Y(n765) );
  INVX1 U898 ( .A(dbg_04[0]), .Y(n742) );
  INVX1 U899 ( .A(dbg_07[0]), .Y(n828) );
  INVX1 U900 ( .A(dbg_0a[0]), .Y(n768) );
  INVX1 U901 ( .A(dbg_04[2]), .Y(n738) );
  INVX1 U902 ( .A(dbg_07[2]), .Y(n826) );
  INVX1 U903 ( .A(dbg_0a[2]), .Y(n766) );
  INVX1 U904 ( .A(dbg_04[6]), .Y(n732) );
  INVX1 U905 ( .A(dbg_07[6]), .Y(n823) );
  INVX1 U906 ( .A(dbg_0a[6]), .Y(n763) );
  INVX1 U907 ( .A(dbg_05[1]), .Y(n721) );
  INVX1 U908 ( .A(dbg_08[1]), .Y(n821) );
  INVX1 U909 ( .A(dbg_0b[1]), .Y(n761) );
  INVX1 U910 ( .A(dbg_05[4]), .Y(n714) );
  INVX1 U911 ( .A(dbg_08[4]), .Y(n818) );
  INVX1 U912 ( .A(dbg_0b[4]), .Y(n758) );
  INVX1 U913 ( .A(dbg_0b[5]), .Y(n807) );
  INVX1 U914 ( .A(dbg_05[3]), .Y(n716) );
  INVX1 U915 ( .A(dbg_08[3]), .Y(n819) );
  INVX1 U916 ( .A(dbg_0b[3]), .Y(n759) );
  INVX1 U917 ( .A(dbg_05[0]), .Y(n723) );
  INVX1 U918 ( .A(dbg_08[0]), .Y(n822) );
  INVX1 U919 ( .A(dbg_0b[0]), .Y(n762) );
  INVX1 U920 ( .A(dbg_05[2]), .Y(n719) );
  INVX1 U921 ( .A(dbg_08[2]), .Y(n820) );
  INVX1 U922 ( .A(dbg_0b[2]), .Y(n760) );
  INVX1 U923 ( .A(dbg_05[6]), .Y(n712) );
  INVX1 U924 ( .A(dbg_08[6]), .Y(n816) );
  INVX1 U925 ( .A(dbg_0b[6]), .Y(n806) );
  INVX1 U926 ( .A(dbg_03[1]), .Y(n730) );
  INVX1 U927 ( .A(dbg_06[1]), .Y(n754) );
  INVX1 U928 ( .A(dbg_09[1]), .Y(n814) );
  INVX1 U929 ( .A(dbg_03[4]), .Y(n727) );
  INVX1 U930 ( .A(dbg_06[4]), .Y(n751) );
  INVX1 U931 ( .A(dbg_09[4]), .Y(n811) );
  INVX1 U932 ( .A(dbg_09[5]), .Y(n810) );
  INVX1 U933 ( .A(dbg_03[3]), .Y(n728) );
  INVX1 U934 ( .A(dbg_06[3]), .Y(n752) );
  INVX1 U935 ( .A(dbg_09[3]), .Y(n812) );
  INVX1 U936 ( .A(dbg_03[0]), .Y(n731) );
  INVX1 U937 ( .A(dbg_06[0]), .Y(n755) );
  INVX1 U938 ( .A(dbg_09[0]), .Y(n815) );
  INVX1 U939 ( .A(dbg_03[2]), .Y(n729) );
  INVX1 U940 ( .A(dbg_06[2]), .Y(n753) );
  INVX1 U941 ( .A(dbg_09[2]), .Y(n813) );
  INVX1 U942 ( .A(dbg_03[6]), .Y(n725) );
  INVX1 U943 ( .A(dbg_06[6]), .Y(n749) );
  INVX1 U944 ( .A(dbg_09[6]), .Y(n809) );
  OAI22AX1 U945 ( .D(n569), .C(pmem_a[9]), .A(adr_p[14]), .B(adr_p[13]), .Y(
        n498) );
  INVX1 U946 ( .A(n254), .Y(o_bkp_hold) );
  INVX1 U947 ( .A(memaddr[12]), .Y(n694) );
  XNOR2XL U948 ( .A(memaddr[10]), .B(bkpt_pc[10]), .Y(n393) );
  XNOR2XL U949 ( .A(memaddr[7]), .B(bkpt_pc[7]), .Y(n385) );
  XOR2X1 U950 ( .A(bkpt_pc[9]), .B(memaddr[9]), .Y(n381) );
  XOR2X1 U951 ( .A(bkpt_pc[8]), .B(memaddr[8]), .Y(n380) );
  XOR2X1 U952 ( .A(bkpt_pc[13]), .B(memaddr[13]), .Y(n388) );
  XNOR2XL U953 ( .A(bkpt_pc[12]), .B(n694), .Y(n389) );
  INVX1 U954 ( .A(n182), .Y(n185) );
  NAND32X1 U955 ( .B(cs_ft[3]), .C(cs_ft[1]), .A(n190), .Y(n182) );
  NAND2X1 U956 ( .A(n376), .B(n377), .Y(n254) );
  NOR4XL U957 ( .A(n378), .B(n379), .C(n380), .D(n381), .Y(n377) );
  NOR4XL U958 ( .A(n386), .B(n387), .C(n388), .D(n389), .Y(n376) );
  NAND3X1 U959 ( .A(n711), .B(r_rdy), .C(bkpt_ena), .Y(n379) );
  NAND4X1 U960 ( .A(n393), .B(n394), .C(n395), .D(n396), .Y(n386) );
  XNOR2XL U961 ( .A(memaddr[4]), .B(bkpt_pc[4]), .Y(n396) );
  XNOR2XL U962 ( .A(memaddr[5]), .B(bkpt_pc[5]), .Y(n395) );
  XNOR2XL U963 ( .A(memaddr[0]), .B(bkpt_pc[0]), .Y(n394) );
  NAND4X1 U964 ( .A(n382), .B(n383), .C(n384), .D(n385), .Y(n378) );
  XNOR2XL U965 ( .A(memaddr[3]), .B(bkpt_pc[3]), .Y(n382) );
  XNOR2XL U966 ( .A(memaddr[1]), .B(bkpt_pc[1]), .Y(n383) );
  XNOR2XL U967 ( .A(memaddr[6]), .B(bkpt_pc[6]), .Y(n384) );
  NAND3X1 U968 ( .A(n390), .B(n391), .C(n392), .Y(n387) );
  XNOR2XL U969 ( .A(memaddr[14]), .B(bkpt_pc[14]), .Y(n390) );
  XNOR2XL U970 ( .A(memaddr[2]), .B(bkpt_pc[2]), .Y(n391) );
  XNOR2XL U971 ( .A(memaddr[11]), .B(bkpt_pc[11]), .Y(n392) );
  NAND2X1 U972 ( .A(d_psrd), .B(n747), .Y(d_inst[2]) );
  NOR2X1 U973 ( .A(n679), .B(n756), .Y(d_inst[4]) );
  NAND2X1 U974 ( .A(d_psrd), .B(n745), .Y(d_inst[5]) );
  NAND2X1 U975 ( .A(n19), .B(n744), .Y(d_inst[6]) );
  NAND2X1 U976 ( .A(n19), .B(n746), .Y(d_inst[3]) );
  NAND2X1 U977 ( .A(n19), .B(n748), .Y(d_inst[1]) );
  NOR2X1 U978 ( .A(n679), .B(n757), .Y(d_inst[0]) );
  NAND43X1 U979 ( .B(cs_ft[2]), .C(cs_ft[0]), .D(cs_ft[1]), .A(cs_ft[3]), .Y(
        n493) );
  INVX1 U980 ( .A(un_hold), .Y(n711) );
  NAND3X1 U981 ( .A(n401), .B(sfr_psw), .C(dw_ena), .Y(n400) );
  OAI33XL U982 ( .A(n400), .B(dummy[1]), .C(dummy[0]), .D(n678), .E(n689), .F(
        n690), .Y(n651) );
  OAI33XL U983 ( .A(n400), .B(dummy[1]), .C(n678), .D(n677), .E(n689), .F(n690), .Y(n650) );
  NAND21X1 U984 ( .B(n136), .A(c_adr[6]), .Y(n135) );
  NAND21X1 U985 ( .B(n52), .A(c_adr[5]), .Y(n136) );
  NAND21X1 U986 ( .B(n135), .A(c_adr[7]), .Y(n133) );
  OR2X1 U987 ( .A(c_adr[1]), .B(c_ptr[1]), .Y(n199) );
  INVX1 U988 ( .A(c_ptr[0]), .Y(n680) );
  INVX1 U989 ( .A(c_adr[0]), .Y(n685) );
  INVX1 U990 ( .A(n125), .Y(n198) );
  NAND21X1 U991 ( .B(n686), .A(c_ptr[1]), .Y(n125) );
  NAND21X1 U992 ( .B(n131), .A(c_adr[10]), .Y(n163) );
  OAI21BX1 U993 ( .C(n52), .B(c_adr[5]), .A(n136), .Y(n153) );
  XOR2X1 U994 ( .A(n133), .B(c_adr[8]), .Y(n159) );
  NAND2X1 U995 ( .A(n131), .B(n132), .Y(n162) );
  OR2X1 U996 ( .A(n169), .B(n56), .Y(n170) );
  AOI21X1 U997 ( .B(n168), .C(c_adr[11]), .A(c_adr[12]), .Y(n56) );
  NAND21X1 U998 ( .B(c_adr[2]), .A(n511), .Y(n201) );
  INVX1 U999 ( .A(c_ptr[2]), .Y(n511) );
  OAI222XL U1000 ( .A(n699), .B(n412), .C(sfr_wdat[7]), .D(n537), .E(
        memdatao[7]), .F(n538), .Y(N793) );
  INVX1 U1001 ( .A(n539), .Y(n699) );
  OAI221X1 U1002 ( .A(sfr_wdat[1]), .B(n537), .C(n704), .D(n412), .E(n550), 
        .Y(N787) );
  EORX1 U1003 ( .A(wr_buf[2]), .B(n453), .C(memdatao[1]), .D(n538), .Y(n550)
         );
  INVX1 U1004 ( .A(n551), .Y(n704) );
  OAI221X1 U1005 ( .A(sfr_wdat[5]), .B(n537), .C(n701), .D(n412), .E(n542), 
        .Y(N791) );
  EORX1 U1006 ( .A(wr_buf[6]), .B(n453), .C(memdatao[5]), .D(n538), .Y(n542)
         );
  INVX1 U1007 ( .A(n543), .Y(n701) );
  OAI221X1 U1008 ( .A(sfr_wdat[3]), .B(n537), .C(n702), .D(n412), .E(n546), 
        .Y(N789) );
  EORX1 U1009 ( .A(wr_buf[4]), .B(n453), .C(memdatao[3]), .D(n538), .Y(n546)
         );
  INVX1 U1010 ( .A(n547), .Y(n702) );
  OAI221X1 U1011 ( .A(sfr_wdat[2]), .B(n537), .C(n703), .D(n412), .E(n548), 
        .Y(N788) );
  EORX1 U1012 ( .A(wr_buf[3]), .B(n453), .C(memdatao[2]), .D(n538), .Y(n548)
         );
  INVX1 U1013 ( .A(n549), .Y(n703) );
  OAI221X1 U1014 ( .A(sfr_wdat[6]), .B(n537), .C(n700), .D(n13), .E(n540), .Y(
        N792) );
  EORX1 U1015 ( .A(wr_buf[7]), .B(n453), .C(memdatao[6]), .D(n538), .Y(n540)
         );
  INVX1 U1016 ( .A(n541), .Y(n700) );
  OAI221X1 U1017 ( .A(memdatao[0]), .B(n538), .C(n674), .D(n682), .E(n552), 
        .Y(N786) );
  EORX1 U1018 ( .A(n673), .B(n553), .C(sfr_wdat[0]), .D(n537), .Y(n552) );
  OAI221X1 U1019 ( .A(memdatao[4]), .B(n538), .C(n674), .D(n681), .E(n544), 
        .Y(N790) );
  EORX1 U1020 ( .A(n673), .B(n545), .C(sfr_wdat[4]), .D(n537), .Y(n544) );
  XNOR2XL U1021 ( .A(n163), .B(c_adr[11]), .Y(n57) );
  INVX1 U1022 ( .A(n126), .Y(n200) );
  NAND21X1 U1023 ( .B(n684), .A(c_ptr[2]), .Y(n126) );
  NAND21X1 U1024 ( .B(n680), .A(c_adr[0]), .Y(n138) );
  XOR2X1 U1025 ( .A(n451), .B(c_adr[3]), .Y(n230) );
  XNOR2XL U1026 ( .A(c_adr[14]), .B(n58), .Y(n408) );
  NAND2X1 U1027 ( .A(c_adr[13]), .B(n169), .Y(n58) );
  XOR2X1 U1028 ( .A(n511), .B(c_adr[2]), .Y(n228) );
  XOR2X1 U1029 ( .A(n512), .B(c_adr[4]), .Y(n232) );
  NAND21X1 U1030 ( .B(c_adr[3]), .A(n451), .Y(n203) );
  INVX1 U1031 ( .A(c_ptr[3]), .Y(n451) );
  INVX1 U1032 ( .A(c_ptr[4]), .Y(n512) );
  XNOR2XL U1033 ( .A(n130), .B(c_adr[13]), .Y(n59) );
  INVX1 U1034 ( .A(n127), .Y(n202) );
  NAND21X1 U1035 ( .B(n683), .A(c_ptr[3]), .Y(n127) );
  NAND21X1 U1036 ( .B(c_adr[0]), .A(n680), .Y(n225) );
  NAND21X1 U1037 ( .B(c_adr[4]), .A(n512), .Y(n205) );
  INVX1 U1038 ( .A(n128), .Y(n204) );
  NAND21X1 U1039 ( .B(n512), .A(c_adr[4]), .Y(n128) );
  INVX1 U1040 ( .A(c_adr[4]), .Y(n99) );
  INVX1 U1041 ( .A(c_adr[6]), .Y(n206) );
  NAND2X1 U1042 ( .A(n216), .B(c_adr[5]), .Y(n212) );
  AND2X1 U1043 ( .A(n243), .B(c_adr[11]), .Y(n244) );
  INVX1 U1044 ( .A(c_adr[8]), .Y(n246) );
  INVX1 U1045 ( .A(c_adr[7]), .Y(n207) );
  INVX1 U1046 ( .A(c_adr[9]), .Y(n208) );
  INVX1 U1047 ( .A(c_adr[10]), .Y(n209) );
  NAND21X1 U1048 ( .B(n129), .A(c_adr[11]), .Y(n211) );
  NOR43XL U1049 ( .B(o_inst[6]), .C(o_inst[5]), .D(o_inst[7]), .A(n260), .Y(
        n259) );
  NAND32X1 U1050 ( .B(memaddr[10]), .C(memaddr[11]), .A(n698), .Y(n260) );
  AND3X1 U1051 ( .A(o_inst[0]), .B(o_inst[1]), .C(r_rdy), .Y(n257) );
  OAI31XL U1052 ( .A(n251), .B(n252), .C(n253), .D(n254), .Y(o_set_hold) );
  NAND42X1 U1053 ( .C(memaddr[14]), .D(memaddr[13]), .A(n694), .B(n255), .Y(
        n253) );
  NAND43X1 U1054 ( .B(memaddr[5]), .C(memaddr[6]), .D(memaddr[4]), .A(n256), 
        .Y(n252) );
  NAND3X1 U1055 ( .A(n257), .B(n258), .C(n259), .Y(n251) );
  INVX1 U1056 ( .A(c_adr[12]), .Y(n129) );
  INVX1 U1057 ( .A(n186), .Y(n194) );
  NAND5XL U1058 ( .A(d_hold[1]), .B(d_hold[3]), .C(d_hold[2]), .D(d_hold[0]), 
        .E(r_hold_mcu), .Y(n186) );
  NAND43X1 U1059 ( .B(c_ptr[2]), .C(n430), .D(n451), .A(c_ptr[4]), .Y(n434) );
  NAND21X1 U1060 ( .B(n487), .A(cs_ft[2]), .Y(n581) );
  NAND21X1 U1061 ( .B(c_ptr[1]), .A(n680), .Y(n430) );
  INVX1 U1062 ( .A(d_psrd), .Y(n679) );
  NAND21X1 U1063 ( .B(n482), .A(n477), .Y(n541) );
  MUX2X1 U1064 ( .D0(pmem_q0[6]), .D1(pmem_q1[6]), .S(n484), .Y(n477) );
  NAND21X1 U1065 ( .B(n482), .A(n476), .Y(n539) );
  MUX2X1 U1066 ( .D0(pmem_q0[7]), .D1(pmem_q1[7]), .S(n484), .Y(n476) );
  NAND21X1 U1067 ( .B(n482), .A(n481), .Y(n551) );
  MUX2X1 U1068 ( .D0(pmem_q0[1]), .D1(pmem_q1[1]), .S(n484), .Y(n481) );
  NAND21X1 U1069 ( .B(n482), .A(n478), .Y(n543) );
  MUX2X1 U1070 ( .D0(pmem_q0[5]), .D1(pmem_q1[5]), .S(n484), .Y(n478) );
  NAND21X1 U1071 ( .B(n482), .A(n479), .Y(n547) );
  MUX2X1 U1072 ( .D0(pmem_q0[3]), .D1(pmem_q1[3]), .S(n484), .Y(n479) );
  NAND21X1 U1073 ( .B(n482), .A(n480), .Y(n549) );
  MUX2X1 U1074 ( .D0(pmem_q0[2]), .D1(pmem_q1[2]), .S(n484), .Y(n480) );
  NAND21X1 U1075 ( .B(cs_ft[2]), .A(n185), .Y(n192) );
  OAI31XL U1076 ( .A(n711), .B(n83), .C(r_rdy), .D(n688), .Y(n717) );
  INVX1 U1077 ( .A(n801), .Y(n688) );
  INVX1 U1078 ( .A(dummy[0]), .Y(n678) );
  INVX1 U1079 ( .A(dummy[1]), .Y(n677) );
  NAND21X1 U1080 ( .B(mcu_psw), .A(n453), .Y(n691) );
  NOR21XL U1081 ( .B(n554), .A(pmem_a[6]), .Y(N757) );
  INVX1 U1082 ( .A(memaddr[13]), .Y(n588) );
  NAND5XL U1083 ( .A(n681), .B(n682), .C(n470), .D(n469), .E(n468), .Y(n528)
         );
  INVX1 U1084 ( .A(wr_buf[4]), .Y(n470) );
  INVX1 U1085 ( .A(wr_buf[6]), .Y(n469) );
  AND4X1 U1086 ( .A(n467), .B(n466), .C(n473), .D(n465), .Y(n468) );
  INVX1 U1087 ( .A(n556), .Y(n705) );
  AOI32X1 U1088 ( .A(pmem_a[6]), .B(n706), .C(n554), .D(pmem_a[7]), .E(N757), 
        .Y(n556) );
  OAI22X1 U1089 ( .A(pmem_q0[0]), .B(n484), .C(pmem_q1[0]), .D(n483), .Y(n553)
         );
  OAI22X1 U1090 ( .A(pmem_q0[4]), .B(n484), .C(pmem_q1[4]), .D(n483), .Y(n545)
         );
  NOR3XL U1091 ( .A(memaddr[7]), .B(memaddr[9]), .C(memaddr[8]), .Y(n256) );
  NOR3XL U1092 ( .A(memaddr[1]), .B(memaddr[3]), .C(memaddr[2]), .Y(n255) );
  INVX1 U1093 ( .A(wr_buf[7]), .Y(n465) );
  NAND21X1 U1094 ( .B(n680), .A(c_ptr[1]), .Y(n463) );
  OR2X1 U1095 ( .A(wspp_cnt_0_), .B(wspp_cnt_1_), .Y(n709) );
  GEN2XL U1096 ( .D(n554), .E(n706), .C(N757), .B(pmem_a[8]), .A(n555), .Y(
        N759) );
  NOR42XL U1097 ( .C(pmem_a[6]), .D(n554), .A(n706), .B(pmem_a[8]), .Y(n555)
         );
  GEN2XL U1098 ( .D(wspp_cnt_1_), .E(wspp_cnt_0_), .C(n671), .B(n672), .A(n669), .Y(N796) );
  GEN2XL U1099 ( .D(wspp_cnt_2_), .E(n709), .C(n670), .B(n672), .A(n669), .Y(
        N797) );
  GEN2XL U1100 ( .D(wspp_cnt_4_), .E(n708), .C(n533), .B(n672), .A(n669), .Y(
        N799) );
  GEN2XL U1101 ( .D(wspp_cnt_5_), .E(n707), .C(n532), .B(n672), .A(n669), .Y(
        N800) );
  NOR2X1 U1102 ( .A(n195), .B(wspp_cnt_3_), .Y(n534) );
  NOR2X1 U1103 ( .A(n708), .B(wspp_cnt_4_), .Y(n533) );
  INVX1 U1104 ( .A(n195), .Y(n670) );
  NAND21X1 U1105 ( .B(wspp_cnt_2_), .A(n671), .Y(n195) );
  NAND2X1 U1106 ( .A(n676), .B(mcu_psw), .Y(n538) );
  OAI21X1 U1107 ( .B(wspp_cnt_0_), .C(n852), .A(n691), .Y(N795) );
  OAI21X1 U1108 ( .B(n531), .C(n852), .A(n691), .Y(N801) );
  XNOR2XL U1109 ( .A(test_so2), .B(n532), .Y(n531) );
  NOR2X1 U1110 ( .A(n707), .B(wspp_cnt_5_), .Y(n532) );
  INVX1 U1111 ( .A(wr_buf[0]), .Y(n473) );
  INVX1 U1112 ( .A(wr_buf[5]), .Y(n681) );
  INVX1 U1113 ( .A(wr_buf[1]), .Y(n682) );
  INVX1 U1114 ( .A(wr_buf[2]), .Y(n467) );
  INVX1 U1115 ( .A(wr_buf[3]), .Y(n466) );
  NOR21XL U1116 ( .B(d_hold[1]), .A(n83), .Y(N153) );
  NOR21XL U1117 ( .B(d_hold[2]), .A(n83), .Y(N154) );
  INVX1 U1118 ( .A(pmem_a[7]), .Y(n706) );
  INVX1 U1119 ( .A(n441), .Y(n635) );
  NAND21X1 U1120 ( .B(c_ptr[0]), .A(c_ptr[1]), .Y(n441) );
  INVX1 U1121 ( .A(n440), .Y(n636) );
  NAND21X1 U1122 ( .B(c_ptr[1]), .A(c_ptr[0]), .Y(n440) );
  NOR2X1 U1123 ( .A(n83), .B(n710), .Y(N152) );
  INVX1 U1124 ( .A(d_hold[0]), .Y(n710) );
  NOR2X1 U1125 ( .A(n535), .B(n852), .Y(N798) );
  AOI21X1 U1126 ( .B(wspp_cnt_3_), .C(n195), .A(n534), .Y(n535) );
  AO2222XL U1127 ( .A(memaddr[6]), .B(n5), .C(sfr_psofs[6]), .D(n8), .E(
        pre_1_adr[6]), .F(n665), .G(memaddr_c[6]), .H(n15), .Y(N860) );
  XOR3XL U1128 ( .A(memaddr_c[6]), .B(c_adr[6]), .C(n212), .Y(n214) );
  NAND21XL U1129 ( .B(n51), .A(memaddr_c[6]), .Y(n415) );
  INVXL U1130 ( .A(memaddr_c[6]), .Y(n154) );
  AO2222XL U1131 ( .A(memaddr[2]), .B(n5), .C(sfr_psofs[2]), .D(n8), .E(
        pre_1_adr[2]), .F(n2), .G(memaddr_c[2]), .H(n15), .Y(N856) );
  XNOR3XL U1132 ( .A(n228), .B(n227), .C(memaddr_c[2]), .Y(n235) );
  GEN2XL U1133 ( .D(memaddr_c[2]), .E(n684), .C(n94), .B(n95), .A(n92), .Y(n98) );
  AOI31XL U1134 ( .A(n493), .B(n503), .C(n492), .D(n61), .Y(n643) );
  AO21XL U1135 ( .B(memaddr_c[0]), .C(n657), .A(n61), .Y(n502) );
  AO21XL U1136 ( .B(memaddr_c[14]), .C(n657), .A(n61), .Y(n658) );
  NAND21XL U1137 ( .B(n691), .A(n18), .Y(n471) );
  AO21XL U1138 ( .B(n18), .C(n559), .A(n558), .Y(N823) );
  AO21XL U1139 ( .B(n618), .C(n505), .A(n567), .Y(N821) );
  AND4XL U1140 ( .A(n618), .B(r_rdy), .C(n412), .D(n562), .Y(n563) );
  GEN3XL U1141 ( .F(n618), .G(n568), .E(n567), .D(n566), .C(n565), .B(n564), 
        .A(n563), .Y(n648) );
  NAND21XL U1142 ( .B(o_ofs_inc), .A(n618), .Y(n630) );
  NAND21XL U1143 ( .B(n582), .A(n618), .Y(n583) );
  AND3XL U1144 ( .A(n618), .B(n582), .C(n501), .Y(n435) );
  NAND21XL U1145 ( .B(n412), .A(n618), .Y(n577) );
  OAI32XL U1146 ( .A(n581), .B(d_psrd), .C(n656), .D(n580), .E(n579), .Y(n664)
         );
  AO2222XL U1147 ( .A(memaddr[4]), .B(n5), .C(sfr_psofs[4]), .D(n8), .E(
        pre_1_adr[4]), .F(n665), .G(memaddr_c[4]), .H(n15), .Y(N858) );
  XNOR3XL U1148 ( .A(n232), .B(n231), .C(memaddr_c[4]), .Y(n233) );
  OAI32XL U1149 ( .A(n100), .B(memaddr_c[4]), .C(n99), .D(n98), .E(n97), .Y(
        n104) );
  OAI222XL U1150 ( .A(memaddr_c[5]), .B(n153), .C(n152), .D(n407), .E(
        memaddr_c[4]), .F(n151), .Y(n155) );
endmodule


module ictlr_a0_DW01_inc_2 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module ictlr_a0_DW01_inc_1 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mcu51_a0 ( bclki2c, pc_ini, slp2wakeup, r_hold_mcu, wdt_slow, wdtov, 
        mdubsy, cs_run, t0_intr, clki2c, clkmdu, clkur0, clktm0, clktm1, 
        clkwdt, i2c_autoack, i2c_con_ens1, clkcpu, clkper, reset, ro, port0i, 
        exint_9, exint, clkcpuen, clkperen, port0o, port0ff, rxd0o, txd0, 
        rxd0i, rxd0oe, scli, sdai, sclo, sdao, waitstaten, mempsack, memack, 
        memdatai, memdatao, memaddr, mempswr, mempsrd, memwr, memrd, 
        memdatao_comb, memaddr_comb, mempswr_comb, mempsrd_comb, memwr_comb, 
        memrd_comb, ramdatai, ramdatao, ramaddr, ramwe, ramoe, dbgpo, sfrack, 
        sfrdatai, sfrdatao, sfraddr, sfrwe, sfroe, esfrm_wrdata, esfrm_addr, 
        esfrm_we, esfrm_oe, esfrm_rddata, test_si2, test_si1, test_so1, 
        test_se );
  input [15:0] pc_ini;
  output [1:0] wdtov;
  input [7:0] port0i;
  input [7:0] exint;
  output [7:0] port0o;
  output [7:0] port0ff;
  input [7:0] memdatai;
  output [7:0] memdatao;
  output [15:0] memaddr;
  output [7:0] memdatao_comb;
  output [15:0] memaddr_comb;
  input [7:0] ramdatai;
  output [7:0] ramdatao;
  output [7:0] ramaddr;
  output [31:0] dbgpo;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  output [6:0] sfraddr;
  input [7:0] esfrm_wrdata;
  input [6:0] esfrm_addr;
  output [7:0] esfrm_rddata;
  input bclki2c, slp2wakeup, r_hold_mcu, wdt_slow, clki2c, clkmdu, clkur0,
         clktm0, clktm1, clkwdt, i2c_autoack, clkcpu, clkper, reset, exint_9,
         rxd0i, scli, sdai, mempsack, memack, sfrack, esfrm_we, esfrm_oe,
         test_si2, test_si1, test_se;
  output mdubsy, cs_run, t0_intr, i2c_con_ens1, ro, clkcpuen, clkperen, rxd0o,
         txd0, rxd0oe, sclo, sdao, waitstaten, mempswr, mempsrd, memwr, memrd,
         mempswr_comb, mempsrd_comb, memwr_comb, memrd_comb, ramwe, ramoe,
         sfrwe, sfroe, test_so1;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         t0_tf1, t1_tf1, t0_tr1, t1_tr1, stop_flag, idle_flag, isfrwait,
         sfroe_s, sfroe_mcu51_per, sfrwe_s, sfrwe_mcu51_per, newinstr,
         intcall_int, cpu_resume, rmwinstr, pmw, p2sel, gf0, c, ac, ov, f0, f1,
         p, rsttowdt, rsttosrst, rst, int0ff, int1ff, rxd0ff, sdaiff,
         rsttowdtff, rsttosrstff, resetff, smod, ip0wdts, wdt_tm, bd, ie0, it0,
         ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9, isr_tm,
         i2c_int, i2ccon_o_7, tf1_gate, riti0_gate, iex7_gate, iex2_gate,
         srstflag, int_vect_8b, int_vect_93, int_vect_9b, int_vect_a3, wdts,
         srst, pmuintreq_rev, pmuintreq, t1ov, t0ack, t1ack, isr_irq, int0ack,
         int1ack, iex7ack, iex2ack, iex3ack, iex4ack, iex5ack, iex6ack,
         iex8ack, iex9ack, n11, n110, n75, n76, n98, n104, n105, n107, n3, n7,
         n8, n9, n10, n12, n1, n2, n4, n5, n6, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n45, n46, n47, n49, n50, n52, n53, n55, n57, n58, n59, n60, n61,
         n63, n65, n67, n69, n71, n73, n77, n79, n80, n81, n82, n84, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5;
  wire   [13:0] timer_1ms;
  wire   [5:0] ien2;
  wire   [6:0] ramsfraddr;
  wire   [4:0] intvect_int;
  wire   [7:0] ckcon;
  wire   [7:0] dph;
  wire   [7:0] dpl;
  wire   [3:0] dps;
  wire   [7:0] p2;
  wire   [5:0] dpc;
  wire   [7:0] sp;
  wire   [7:0] acc_s;
  wire   [7:0] b;
  wire   [1:0] rs;
  wire   [7:0] arcon;
  wire   [7:0] md0;
  wire   [7:0] md1;
  wire   [7:0] md2;
  wire   [7:0] md3;
  wire   [7:0] md4;
  wire   [7:0] md5;
  wire   [3:0] t0_tmod;
  wire   [7:0] tl0;
  wire   [7:0] th0;
  wire   [3:0] t1_tmod;
  wire   [7:0] tl1;
  wire   [7:0] th1;
  wire   [7:0] wdtrel;
  wire   [6:5] t2con;
  wire   [7:0] s0con;
  wire   [7:0] s0buf;
  wire   [7:0] s0rell;
  wire   [7:0] s0relh;
  wire   [7:0] ien0;
  wire   [5:0] ien1;
  wire   [5:0] ip0;
  wire   [5:0] ip1;
  wire   [7:0] i2cdat_o;
  wire   [7:0] i2cadr_o;
  wire   [5:0] i2ccon_o;
  wire   [7:0] i2csta_o;
  wire   [3:0] isreg;

  INVX1 U40 ( .A(n76), .Y(n75) );
  INVX1 U41 ( .A(reset), .Y(n76) );
  INVX8 U52 ( .A(n76), .Y(n3) );
  mcu51_cpu_a0 u_cpu ( .clkcpu(clkcpu), .rst(n84), .mempsack(mempsack), 
        .memack(memack), .memdatai(memdatai), .memaddr(memaddr), .mempsrd(
        mempsrd), .mempswr(mempswr), .memrd(memrd), .memwr(memwr), 
        .memaddr_comb(memaddr_comb), .mempsrd_comb(mempsrd_comb), 
        .mempswr_comb(mempswr_comb), .memrd_comb(memrd_comb), .memwr_comb(
        memwr_comb), .cpu_hold(r_hold_mcu), .cpu_resume(cpu_resume), .irq(
        dbgpo[20]), .intvect(intvect_int), .intcall(intcall_int), .retiinstr(
        dbgpo[21]), .newinstr(newinstr), .rmwinstr(rmwinstr), .waitstaten(
        waitstaten), .ramdatai(ramdatai), .sfrdatai(esfrm_rddata), 
        .ramsfraddr({SYNOPSYS_UNCONNECTED_1, ramsfraddr}), .ramdatao(memdatao), 
        .ramoe(), .ramwe(), .sfroe(sfroe_s), .sfrwe(sfrwe_s), .sfroe_r(), 
        .sfrwe_r(), .sfroe_comb_s(), .sfrwe_comb_s(), .pc_o(dbgpo[15:0]), 
        .pc_ini(pc_ini), .cs_run(cs_run), .instr(dbgpo[31:24]), .codefetch_s(), 
        .sfrack(sfrack), .ramsfraddr_comb(ramaddr), .ramdatao_comb(ramdatao), 
        .ramoe_comb(ramoe), .ramwe_comb(ramwe), .ckcon(ckcon), .pmw(pmw), 
        .p2sel(p2sel), .gf0(gf0), .stop(stop_flag), .idle(idle_flag), .acc(
        acc_s), .b(b), .rs(rs), .c(c), .ac(ac), .ov(ov), .p(p), .f0(f0), .f1(
        f1), .dph(dph), .dpl(dpl), .dps(dps), .dpc(dpc), .p2(p2), .sp(sp), 
        .test_si(timer_1ms[13]), .test_so(n107), .test_se(test_se) );
  syncneg_a0 u_syncneg ( .clk(clkper), .reset(n75), .rsttowdt(rsttowdt), 
        .rsttosrst(rsttosrst), .rst(rst), .int0(exint[0]), .int1(exint[1]), 
        .port0i(port0i), .rxd0i(rxd0i), .sdai(sdai), .int0ff(int0ff), .int1ff(
        int1ff), .port0ff(port0ff), .t0ff(), .t1ff(), .rxd0ff(rxd0ff), 
        .sdaiff(sdaiff), .rsttowdtff(rsttowdtff), .rsttosrstff(rsttosrstff), 
        .rstff(n98), .resetff(resetff), .test_si(srstflag), .test_se(test_se)
         );
  sfrmux_a0 u_sfrmux ( .isfrwait(isfrwait), .sfraddr({n59, sfraddr[5], n55, 
        n53, n50, n47, n45}), .c(c), .ac(ac), .f0(f0), .rs(rs), .ov(ov), .f1(
        f1), .p(p), .acc(acc_s), .b(b), .dpl(dpl), .dph(dph), .dps(dps), .dpc(
        dpc), .p2(p2), .sp(sp), .smod(smod), .pmw(pmw), .p2sel(p2sel), .gf0(
        gf0), .stop(stop_flag), .idle(idle_flag), .ckcon(ckcon), .port0(port0o), .port0ff(port0ff), .rmwinstr(rmwinstr), .arcon(arcon), .md0(md0), .md1(md1), 
        .md2(md2), .md3(md3), .md4(md4), .md5(md5), .t0_tmod(t0_tmod), 
        .t0_tf0(dbgpo[17]), .t0_tf1(t0_tf1), .t0_tr0(dbgpo[16]), .t0_tr1(
        t0_tr1), .tl0(tl0), .th0(th0), .t1_tmod(t1_tmod), .t1_tf1(t1_tf1), 
        .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1), .wdtrel(wdtrel), .ip0wdts(
        ip0wdts), .wdt_tm(wdt_tm), .t2con({1'b0, t2con, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .s0con(s0con), .s0buf(s0buf), .s0rell(s0rell), .s0relh(s0relh), 
        .bd(bd), .ie0(ie0), .it0(it0), .ie1(ie1), .it1(it1), .iex2(iex2), 
        .iex3(iex3), .iex4(iex4), .iex5(iex5), .iex6(iex6), .iex7(iex7), 
        .iex8(iex8), .iex9(iex9), .iex10(1'b0), .iex11(1'b0), .iex12(1'b0), 
        .ien0({ien0[7], 1'b0, ien0[5:0]}), .ien1(ien1), .ien2(ien2), .ip0(ip0), 
        .ip1(ip1), .isr_tm(isr_tm), .i2c_int(i2c_int), .i2cdat_o(i2cdat_o), 
        .i2cadr_o(i2cadr_o), .i2ccon_o({i2ccon_o_7, i2c_con_ens1, i2ccon_o}), 
        .i2csta_o({i2csta_o[7:3], 1'b0, 1'b0, 1'b0}), .sfrdatai(sfrdatai), 
        .tf1_gate(tf1_gate), .riti0_gate(riti0_gate), .iex7_gate(iex7_gate), 
        .iex2_gate(iex2_gate), .srstflag(srstflag), .int_vect_8b(int_vect_8b), 
        .int_vect_93(int_vect_93), .int_vect_9b(int_vect_9b), .int_vect_a3(
        int_vect_a3), .ext_sfr_sel(), .sfrdatao(esfrm_rddata) );
  pmurstctrl_a0 u_pmurstctrl ( .resetff(resetff), .wdts(wdts), .srst(srst), 
        .pmuintreq(pmuintreq_rev), .stop(stop_flag), .idle(idle_flag), 
        .clkcpu_en(clkcpuen), .clkper_en(clkperen), .cpu_resume(cpu_resume), 
        .rsttowdt(rsttowdt), .rsttosrst(rsttosrst), .rst(rst) );
  wakeupctrl_a0 u_wakeupctrl ( .irq(dbgpo[20]), .int0ff(exint[0]), .int1ff(
        exint[1]), .it0(it0), .it1(it1), .isreg(isreg), .intprior0({ip0[2], 
        ip0[0]}), .intprior1({ip1[2], ip1[0]}), .eal(ien0[7]), .eint0(ien0[0]), 
        .eint1(ien0[2]), .pmuintreq(pmuintreq) );
  mdu_a0 u_mdu ( .clkper(clkmdu), .rst(ro), .mdubsy(mdubsy), .sfrdatai(
        sfrdatao), .sfraddr({n61, n58, n55, n53, n6, n46, sfraddr[0]}), 
        .sfrwe(n40), .sfroe(sfroe_mcu51_per), .arcon(arcon), .md0(md0), .md1(
        md1), .md2(md2), .md3(md3), .md4(md4), .md5(md5), .test_si(isr_tm), 
        .test_so(n104), .test_se(test_se) );
  ports_a0 u_ports ( .clkper(clkper), .rst(n84), .port0(port0o), .sfrdatai({
        sfrdatao[7], n18, n21, n17, sfrdatao[3:0]}), .sfraddr({n61, n58, 
        sfraddr[4:3], n50, n110, n14}), .sfrwe(n40), .test_si(n104), .test_se(
        test_se) );
  serial0_a0 u_serial0 ( .t_shift_clk(), .r_shift_clk(), .clkper(clkur0), 
        .rst(n84), .newinstr(newinstr), .rxd0ff(rxd0ff), .t1ov(t1ov), .rxd0o(
        rxd0o), .rxd0oe(rxd0oe), .txd0(txd0), .sfrdatai({n79, sfrdatao[6:4], 
        n15, n20, n19, n16}), .sfraddr({n61, n57, n4, n52, n5, n46, n36}), 
        .sfrwe(n41), .s0con(s0con), .s0buf(s0buf), .s0rell(s0rell), .s0relh(
        s0relh), .smod(smod), .bd(bd), .test_si(port0o[7]), .test_se(test_se)
         );
  timer0_a0 u_timer0 ( .clkper(clktm0), .rst(n82), .newinstr(newinstr), .t0ff(
        1'b0), .t0ack(t0ack), .t1ack(t1ack), .int0ff(int0ff), .t0_tf0(
        dbgpo[17]), .t0_tf1(t0_tf1), .sfrdatai(sfrdatao), .sfraddr({n60, n57, 
        n4, sfraddr[3], n5, n47, n45}), .sfrwe(n40), .t0_tmod(t0_tmod), 
        .t0_tr0(dbgpo[16]), .t0_tr1(t0_tr1), .tl0(tl0), .th0(th0), .test_si(
        sdaiff), .test_se(test_se) );
  timer1_a0 u_timer1 ( .clkper(clktm1), .rst(n80), .newinstr(newinstr), .t1ff(
        1'b0), .t1ack(t1ack), .int1ff(int1ff), .t1_tf1(t1_tf1), .t1ov(t1ov), 
        .sfrdatai({n79, sfrdatao[6:4], n15, sfrdatao[2:1], n16}), .sfraddr({
        n60, n57, n4, n52, n6, n110, n14}), .sfrwe(n41), .t1_tmod(t1_tmod), 
        .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1), .test_si(tl0[7]), .test_se(
        test_se) );
  watchdog_a0 u_watchdog ( .wdt_slow(wdt_slow), .clkwdt(clkwdt), .clkper(
        clkper), .resetff(rsttowdtff), .newinstr(newinstr), .wdts_s(wdtov), 
        .wdts(wdts), .ip0wdts(ip0wdts), .wdt_tm(wdt_tm), .sfrdatai({
        sfrdatao[7:6], n21, n17, sfrdatao[3:0]}), .sfraddr({n61, n57, n4, n52, 
        n6, sfraddr[1:0]}), .sfrwe(n41), .wdtrel(wdtrel), .test_si(tl1[7]), 
        .test_se(test_se) );
  isr_a0 u_isr ( .clkper(clkper), .rst(n81), .intcall(intcall_int), 
        .retiinstr(dbgpo[21]), .int_vect_03(ie0), .int_vect_0b(dbgpo[17]), 
        .t0ff(1'b0), .int_vect_13(ie1), .int_vect_1b(tf1_gate), .t1ff(1'b0), 
        .int_vect_23(riti0_gate), .i2c_int(i2c_int), .rxd0ff(rxd0ff), 
        .int_vect_43(iex7_gate), .sdaiff(sdaiff), .int_vect_4b(iex2_gate), 
        .int_vect_53(iex3), .int_vect_5b(iex4), .int_vect_63(iex5), 
        .int_vect_6b(iex6), .int_vect_8b(int_vect_8b), .int_vect_93(
        int_vect_93), .int_vect_9b(int_vect_9b), .int_vect_a3(int_vect_a3), 
        .int_vect_ab(1'b0), .irq(isr_irq), .intvect(intvect_int), .int_ack_03(
        int0ack), .int_ack_0b(t0ack), .int_ack_13(int1ack), .int_ack_1b(t1ack), 
        .int_ack_43(iex7ack), .int_ack_4b(iex2ack), .int_ack_53(iex3ack), 
        .int_ack_5b(iex4ack), .int_ack_63(iex5ack), .int_ack_6b(iex6ack), 
        .int_ack_8b(iex8ack), .int_ack_93(iex9ack), .int_ack_9b(), 
        .int_ack_a3(), .int_ack_ab(), .is_reg(isreg), .ip0(ip0), .ip1(ip1), 
        .ien0({ien0[7], SYNOPSYS_UNCONNECTED_2, ien0[5:0]}), .ien1(ien1), 
        .ien2(ien2), .isr_tm(isr_tm), .sfraddr({n60, n58, n55, n53, 
        sfraddr[2:1], n36}), .sfrdatai({sfrdatao[7], n18, n21, sfrdatao[4:0]}), 
        .sfrwe(n41), .test_si(n105), .test_se(test_se) );
  extint_a0 u_extint ( .clkper(clkper), .rst(n82), .newinstr(newinstr), 
        .int0ff(int0ff), .int0ack(int0ack), .int1ff(int1ff), .int1ack(int1ack), 
        .int2ff(exint[2]), .iex2ack(iex2ack), .int3ff(exint[3]), .iex3ack(
        iex3ack), .int4ff(exint[4]), .iex4ack(iex4ack), .int5ff(exint[5]), 
        .iex5ack(iex5ack), .int6ff(exint[6]), .iex6ack(iex6ack), .int7ff(
        exint[7]), .iex7ack(iex7ack), .int8ff(n11), .iex8ack(iex8ack), 
        .int9ff(exint_9), .iex9ack(iex9ack), .ie0(ie0), .it0(it0), .ie1(ie1), 
        .it1(it1), .i2fr(t2con[5]), .iex2(iex2), .i3fr(t2con[6]), .iex3(iex3), 
        .iex4(iex4), .iex5(iex5), .iex6(iex6), .iex7(iex7), .iex8(iex8), 
        .iex9(iex9), .iex10(), .iex11(), .iex12(), .sfraddr({n60, n58, 
        sfraddr[4:3], n50, sfraddr[1], n36}), .sfrdatai({n79, n18, sfrdatao[5], 
        n17, n15, n20, n19, n16}), .sfrwe(n40), .test_si(n107), .test_se(
        test_se) );
  i2c_a0 u_i2c ( .clk(clki2c), .rst(n84), .bclksel(bclki2c), .scli(scli), 
        .sdai(sdai), .sclo(sclo), .sdao(sdao), .intack(i2c_autoack), .si(
        i2c_int), .sfrwe(n40), .sfraddr({n60, n58, n4, n52, sfraddr[2], n46, 
        n14}), .sfrdatai({sfrdatao[7], n18, n21, sfrdatao[4:3], n20, 
        sfrdatao[1:0]}), .i2cdat_o(i2cdat_o), .i2cadr_o(i2cadr_o), .i2ccon_o({
        i2ccon_o_7, i2c_con_ens1, i2ccon_o}), .i2csta_o({i2csta_o[7:3], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5}), .test_si2(test_si2), .test_si1(it1), .test_so2(n105), .test_so1(test_so1), 
        .test_se(test_se) );
  softrstctrl_a0 u_softrstctrl ( .clkcpu(clkcpu), .resetff(rsttosrstff), 
        .newinstr(newinstr), .srstreq(srst), .srstflag(srstflag), .sfrdatai({
        n79, n18, n21, n17, sfrdatao[3:0]}), .sfraddr({n61, n58, sfraddr[4], 
        n52, n6, sfraddr[1], n14}), .sfrwe(n41), .test_si(txd0), .test_se(
        test_se) );
  mcu51_a0_DW01_inc_0 add_268 ( .A(timer_1ms), .SUM({N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7}) );
  SDFFQX1 timer_1ms_reg_9_ ( .D(N30), .SIN(timer_1ms[8]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[9]) );
  SDFFQX1 timer_1ms_reg_13_ ( .D(N34), .SIN(timer_1ms[12]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[13]) );
  SDFFQX1 timer_1ms_reg_12_ ( .D(N33), .SIN(timer_1ms[11]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[12]) );
  SDFFQX1 timer_1ms_reg_8_ ( .D(N29), .SIN(timer_1ms[7]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[8]) );
  SDFFQX1 timer_1ms_reg_10_ ( .D(N31), .SIN(timer_1ms[9]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[10]) );
  SDFFQX1 timer_1ms_reg_6_ ( .D(N27), .SIN(timer_1ms[5]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[6]) );
  SDFFQX1 timer_1ms_reg_11_ ( .D(N32), .SIN(timer_1ms[10]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[11]) );
  SDFFQX1 timer_1ms_reg_7_ ( .D(N28), .SIN(timer_1ms[6]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[7]) );
  SDFFQX1 timer_1ms_reg_5_ ( .D(N26), .SIN(timer_1ms[4]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[5]) );
  SDFFQX1 timer_1ms_reg_4_ ( .D(N25), .SIN(timer_1ms[3]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[4]) );
  SDFFQX1 timer_1ms_reg_3_ ( .D(N24), .SIN(timer_1ms[2]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[3]) );
  SDFFQX1 timer_1ms_reg_2_ ( .D(N23), .SIN(timer_1ms[1]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[2]) );
  SDFFQX1 timer_1ms_reg_1_ ( .D(N22), .SIN(timer_1ms[0]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[1]) );
  SDFFQX1 timer_1ms_reg_0_ ( .D(N21), .SIN(test_si1), .SMC(test_se), .C(clkper), .Q(timer_1ms[0]) );
  INVXL U3 ( .A(n39), .Y(sfraddr[4]) );
  MUX2IX2 U4 ( .D0(esfrm_addr[0]), .D1(ramsfraddr[0]), .S(n92), .Y(n88) );
  MUX2IX2 U5 ( .D0(esfrm_addr[6]), .D1(ramsfraddr[6]), .S(n92), .Y(n91) );
  MUX2IX1 U6 ( .D0(esfrm_addr[1]), .D1(ramsfraddr[1]), .S(n92), .Y(n89) );
  INVX1 U7 ( .A(n91), .Y(n59) );
  INVX3 U8 ( .A(n1), .Y(n53) );
  INVXL U9 ( .A(n91), .Y(n61) );
  INVXL U10 ( .A(n91), .Y(n60) );
  INVX3 U11 ( .A(n91), .Y(sfraddr[6]) );
  INVX1 U12 ( .A(esfrm_we), .Y(n94) );
  INVX1 U13 ( .A(n93), .Y(n96) );
  INVX1 U14 ( .A(n90), .Y(sfraddr[5]) );
  AO21X1 U15 ( .B(n96), .C(n95), .A(esfrm_we), .Y(sfrwe) );
  NAND21X1 U16 ( .B(esfrm_oe), .A(n94), .Y(isfrwait) );
  MUX2IX1 U17 ( .D0(ramsfraddr[2]), .D1(esfrm_addr[2]), .S(n34), .Y(n33) );
  INVX3 U18 ( .A(isfrwait), .Y(n92) );
  INVX1 U19 ( .A(n33), .Y(n50) );
  INVX1 U20 ( .A(n35), .Y(n45) );
  MUX2IX1 U21 ( .D0(esfrm_addr[3]), .D1(ramsfraddr[3]), .S(n92), .Y(n1) );
  INVXL U22 ( .A(n1), .Y(sfraddr[3]) );
  MUX2IX1 U23 ( .D0(esfrm_wrdata[7]), .D1(memdatao[7]), .S(n13), .Y(n2) );
  INVX1 U24 ( .A(n89), .Y(n47) );
  INVX1 U25 ( .A(n35), .Y(sfraddr[0]) );
  INVXL U26 ( .A(n39), .Y(n4) );
  BUFX3 U27 ( .A(n32), .Y(n49) );
  INVX1 U28 ( .A(n49), .Y(n5) );
  INVX1 U29 ( .A(n49), .Y(n6) );
  INVX1 U30 ( .A(n34), .Y(n13) );
  INVXL U31 ( .A(n35), .Y(n14) );
  INVXL U32 ( .A(n33), .Y(sfraddr[2]) );
  NAND21XL U33 ( .B(isfrwait), .A(sfrwe_s), .Y(n93) );
  MUX2XL U34 ( .D0(esfrm_wrdata[3]), .D1(memdatao[3]), .S(n92), .Y(n15) );
  MUX2XL U35 ( .D0(esfrm_wrdata[0]), .D1(memdatao[0]), .S(n92), .Y(n16) );
  MUX2XL U36 ( .D0(esfrm_wrdata[4]), .D1(memdatao[4]), .S(n13), .Y(n17) );
  MUX2XL U37 ( .D0(esfrm_wrdata[6]), .D1(memdatao[6]), .S(n13), .Y(n18) );
  MUX2XL U38 ( .D0(esfrm_wrdata[1]), .D1(memdatao[1]), .S(n13), .Y(n19) );
  MUX2XL U39 ( .D0(esfrm_wrdata[2]), .D1(memdatao[2]), .S(n13), .Y(n20) );
  MUX2XL U42 ( .D0(esfrm_wrdata[5]), .D1(memdatao[5]), .S(n13), .Y(n21) );
  BUFX3 U43 ( .A(sfrwe_mcu51_per), .Y(n40) );
  BUFX3 U44 ( .A(sfrwe_mcu51_per), .Y(n41) );
  INVX1 U45 ( .A(n89), .Y(n46) );
  BUFX3 U46 ( .A(ramdatao[0]), .Y(memdatao_comb[0]) );
  BUFX3 U47 ( .A(ramdatao[1]), .Y(memdatao_comb[1]) );
  BUFX3 U48 ( .A(ramdatao[3]), .Y(memdatao_comb[3]) );
  BUFX3 U49 ( .A(ramdatao[2]), .Y(memdatao_comb[2]) );
  BUFX3 U50 ( .A(ramdatao[4]), .Y(memdatao_comb[4]) );
  BUFX3 U51 ( .A(ramdatao[5]), .Y(memdatao_comb[5]) );
  BUFX3 U53 ( .A(ramdatao[6]), .Y(memdatao_comb[6]) );
  BUFX3 U54 ( .A(ramdatao[7]), .Y(memdatao_comb[7]) );
  INVX1 U55 ( .A(n89), .Y(n110) );
  INVX1 U56 ( .A(n39), .Y(n55) );
  INVX1 U57 ( .A(n69), .Y(sfrdatao[3]) );
  INVX1 U58 ( .A(n86), .Y(ro) );
  INVX1 U59 ( .A(n63), .Y(sfrdatao[0]) );
  INVX1 U60 ( .A(n71), .Y(sfrdatao[4]) );
  INVX1 U61 ( .A(n77), .Y(sfrdatao[6]) );
  INVX1 U62 ( .A(n73), .Y(sfrdatao[5]) );
  INVX1 U63 ( .A(n2), .Y(sfrdatao[7]) );
  INVX1 U64 ( .A(n65), .Y(sfrdatao[1]) );
  INVX1 U65 ( .A(n67), .Y(sfrdatao[2]) );
  NAND21XL U66 ( .B(esfrm_oe), .A(n97), .Y(sfroe_mcu51_per) );
  INVXL U67 ( .A(n1), .Y(n52) );
  INVX1 U68 ( .A(n86), .Y(dbgpo[22]) );
  NOR21XL U69 ( .B(N19), .A(n42), .Y(N33) );
  INVX1 U70 ( .A(n86), .Y(n84) );
  NOR21XL U71 ( .B(N18), .A(n43), .Y(N32) );
  NOR21XL U72 ( .B(N17), .A(n42), .Y(N31) );
  NOR21XL U73 ( .B(N16), .A(n43), .Y(N30) );
  INVX1 U74 ( .A(n87), .Y(n80) );
  INVX1 U75 ( .A(n87), .Y(n81) );
  INVX1 U76 ( .A(n87), .Y(n82) );
  NOR21XL U77 ( .B(N8), .A(n43), .Y(N22) );
  NOR21XL U78 ( .B(N9), .A(n42), .Y(N23) );
  NOR21XL U79 ( .B(N10), .A(n43), .Y(N24) );
  NOR21XL U80 ( .B(N11), .A(n42), .Y(N25) );
  NOR21XL U81 ( .B(N14), .A(n43), .Y(N28) );
  NOR21XL U82 ( .B(N13), .A(n42), .Y(N27) );
  NOR21XL U83 ( .B(N12), .A(n43), .Y(N26) );
  NOR21XL U84 ( .B(N15), .A(n42), .Y(N29) );
  BUFX3 U85 ( .A(n7), .Y(n42) );
  BUFX3 U86 ( .A(n7), .Y(n43) );
  BUFX3 U87 ( .A(rxd0i), .Y(dbgpo[23]) );
  INVX1 U88 ( .A(n2), .Y(n79) );
  MUX2IXL U89 ( .D0(esfrm_addr[4]), .D1(ramsfraddr[4]), .S(n92), .Y(n39) );
  INVX1 U90 ( .A(n15), .Y(n69) );
  INVX1 U91 ( .A(n98), .Y(n86) );
  INVX1 U92 ( .A(n16), .Y(n63) );
  AO21XL U93 ( .B(sfroe_s), .C(n95), .A(esfrm_oe), .Y(sfroe) );
  INVX1 U94 ( .A(sfroe_s), .Y(n97) );
  INVX1 U95 ( .A(n17), .Y(n71) );
  INVX1 U96 ( .A(n19), .Y(n65) );
  INVX1 U97 ( .A(n18), .Y(n77) );
  INVX1 U98 ( .A(n21), .Y(n73) );
  INVX1 U99 ( .A(n20), .Y(n67) );
  NOR21XL U100 ( .B(isr_irq), .A(r_hold_mcu), .Y(dbgpo[20]) );
  OR2X1 U101 ( .A(pmuintreq), .B(slp2wakeup), .Y(pmuintreq_rev) );
  OR2X1 U102 ( .A(t0_tf1), .B(t1_tf1), .Y(dbgpo[19]) );
  OR2X1 U103 ( .A(t0_tr1), .B(t1_tr1), .Y(dbgpo[18]) );
  NOR21XL U104 ( .B(N20), .A(n43), .Y(N34) );
  INVX1 U105 ( .A(n98), .Y(n87) );
  NAND32X1 U106 ( .B(n11), .C(n3), .A(ien2[1]), .Y(n7) );
  NOR21XL U107 ( .B(N7), .A(n42), .Y(N21) );
  NAND43X1 U108 ( .B(timer_1ms[8]), .C(timer_1ms[5]), .D(timer_1ms[12]), .A(
        timer_1ms[0]), .Y(n10) );
  NOR4XL U109 ( .A(n8), .B(n9), .C(n10), .D(n12), .Y(n11) );
  NAND4X1 U110 ( .A(timer_1ms[4]), .B(timer_1ms[3]), .C(timer_1ms[2]), .D(
        timer_1ms[1]), .Y(n8) );
  NAND3X1 U111 ( .A(timer_1ms[7]), .B(timer_1ms[6]), .C(timer_1ms[9]), .Y(n9)
         );
  NAND3X1 U112 ( .A(timer_1ms[11]), .B(timer_1ms[10]), .C(timer_1ms[13]), .Y(
        n12) );
  AND2X1 U113 ( .A(ien0[0]), .B(dbgpo[17]), .Y(t0_intr) );
  INVXL U114 ( .A(n89), .Y(sfraddr[1]) );
  INVXL U115 ( .A(n50), .Y(n32) );
  INVXL U116 ( .A(n92), .Y(n34) );
  BUFX3 U117 ( .A(n88), .Y(n35) );
  INVXL U118 ( .A(n35), .Y(n36) );
  INVXL U119 ( .A(sfraddr[5]), .Y(n37) );
  BUFXL U120 ( .A(n37), .Y(n38) );
  INVXL U130 ( .A(n38), .Y(n57) );
  INVXL U131 ( .A(n38), .Y(n58) );
  MUX2IXL U132 ( .D0(esfrm_addr[5]), .D1(ramsfraddr[5]), .S(n92), .Y(n90) );
  NAND21XL U133 ( .B(n96), .A(n94), .Y(sfrwe_mcu51_per) );
  INVX8 U134 ( .A(n3), .Y(n95) );
endmodule


module mcu51_a0_DW01_inc_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;

  wire   [13:2] carry;

  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module softrstctrl_a0 ( clkcpu, resetff, newinstr, srstreq, srstflag, sfrdatai, 
        sfraddr, sfrwe, test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkcpu, resetff, newinstr, sfrwe, test_si, test_se;
  output srstreq, srstflag;
  wire   srst_ff0, srst_ff1, N37, N38, N41, net12009, n24, n25, n26, n27, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n28, n29,
         n30, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [3:0] srst_count;

  SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 clk_gate_srst_count_reg ( .CLK(clkcpu), 
        .EN(N37), .ENCLK(net12009), .TE(test_se) );
  SDFFQX1 srst_ff1_reg ( .D(n24), .SIN(srst_ff0), .SMC(test_se), .C(clkcpu), 
        .Q(srst_ff1) );
  SDFFQX1 srst_count_reg_1_ ( .D(n6), .SIN(srst_count[0]), .SMC(test_se), .C(
        net12009), .Q(srst_count[1]) );
  SDFFQX1 srst_count_reg_3_ ( .D(N41), .SIN(srst_count[2]), .SMC(test_se), .C(
        net12009), .Q(srst_count[3]) );
  SDFFQX1 srst_ff0_reg ( .D(n26), .SIN(srst_count[3]), .SMC(test_se), .C(
        clkcpu), .Q(srst_ff0) );
  SDFFQX1 srst_count_reg_0_ ( .D(N38), .SIN(test_si), .SMC(test_se), .C(
        net12009), .Q(srst_count[0]) );
  SDFFQX1 srst_count_reg_2_ ( .D(n4), .SIN(srst_count[1]), .SMC(test_se), .C(
        net12009), .Q(srst_count[2]) );
  SDFFQX1 srst_r_reg ( .D(n27), .SIN(srst_ff1), .SMC(test_se), .C(clkcpu), .Q(
        srstreq) );
  SDFFQX1 srstflag_reg ( .D(n25), .SIN(srstreq), .SMC(test_se), .C(clkcpu), 
        .Q(srstflag) );
  INVX1 U3 ( .A(n15), .Y(n2) );
  NAND42X1 U4 ( .C(sfraddr[3]), .D(n20), .A(sfraddr[0]), .B(n21), .Y(n15) );
  NAND2X1 U5 ( .A(sfraddr[2]), .B(sfraddr[1]), .Y(n20) );
  AND4X1 U6 ( .A(sfrwe), .B(sfraddr[6]), .C(sfraddr[5]), .D(sfraddr[4]), .Y(
        n21) );
  NAND2X1 U7 ( .A(sfrdatai[0]), .B(n2), .Y(n12) );
  INVX1 U8 ( .A(newinstr), .Y(n3) );
  NOR2X1 U9 ( .A(n16), .B(n5), .Y(n22) );
  INVX1 U10 ( .A(n28), .Y(n5) );
  INVX1 U11 ( .A(n16), .Y(n9) );
  NAND2X1 U12 ( .A(n10), .B(n16), .Y(N37) );
  NOR2X1 U13 ( .A(resetff), .B(n18), .Y(n24) );
  AOI22AXL U14 ( .A(srst_ff0), .B(n2), .D(n19), .C(n8), .Y(n18) );
  AOI32X1 U15 ( .A(srst_ff1), .B(n3), .C(n15), .D(srst_ff0), .E(newinstr), .Y(
        n19) );
  NOR2X1 U16 ( .A(resetff), .B(n11), .Y(n27) );
  AOI32X1 U17 ( .A(n12), .B(n13), .C(srstreq), .D(srst_ff1), .E(n1), .Y(n11)
         );
  NAND3X1 U18 ( .A(srst_count[2]), .B(n5), .C(srst_count[3]), .Y(n13) );
  INVX1 U19 ( .A(n12), .Y(n1) );
  AOI21X1 U20 ( .B(n12), .C(n14), .A(resetff), .Y(n26) );
  NAND4X1 U21 ( .A(srst_ff0), .B(n15), .C(n3), .D(n8), .Y(n14) );
  NAND2X1 U22 ( .A(n16), .B(n17), .Y(n25) );
  OAI211X1 U23 ( .C(sfrdatai[0]), .D(n15), .A(n10), .B(srstflag), .Y(n17) );
  GEN2XL U24 ( .D(n9), .E(n7), .C(n22), .B(srst_count[3]), .A(n23), .Y(N41) );
  NOR4XL U25 ( .A(srst_count[3]), .B(n28), .C(n7), .D(n16), .Y(n23) );
  NAND2X1 U26 ( .A(srstreq), .B(n10), .Y(n16) );
  NAND2X1 U27 ( .A(srst_count[1]), .B(srst_count[0]), .Y(n28) );
  INVX1 U28 ( .A(resetff), .Y(n10) );
  INVX1 U29 ( .A(srst_count[2]), .Y(n7) );
  INVX1 U30 ( .A(srstreq), .Y(n8) );
  INVX1 U31 ( .A(n30), .Y(n6) );
  OAI211X1 U32 ( .C(srst_count[0]), .D(srst_count[1]), .A(n9), .B(n28), .Y(n30) );
  INVX1 U33 ( .A(n29), .Y(n4) );
  AOI32X1 U34 ( .A(n9), .B(n7), .C(n5), .D(srst_count[2]), .E(n22), .Y(n29) );
  NOR2X1 U35 ( .A(srst_count[0]), .B(n16), .Y(N38) );
endmodule


module SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2c_a0 ( clk, rst, bclksel, scli, sdai, sclo, sdao, intack, si, sfrwe, 
        sfraddr, sfrdatai, i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o, test_si2, 
        test_si1, test_so2, test_so1, test_se );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  output [7:0] i2cdat_o;
  output [7:0] i2cadr_o;
  output [7:0] i2ccon_o;
  output [7:0] i2csta_o;
  input clk, rst, bclksel, scli, sdai, intack, sfrwe, test_si2, test_si1,
         test_se;
  output sclo, sdao, si, test_so2, test_so1;
  wire   scli_ff, N180, sdai_ff, N181, sclo_int, wait_for_setup_r, adrcomp,
         adrcompen, nedetect, ack_bit, bsd7, pedetect, N224, N225, N226, N227,
         N232, N233, N234, sclint, ack, sdaint, bsd7_tmp, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N332, N333, N335, N336, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N406, N407, N408,
         N409, N410, N412, N413, N414, sdai_ff_reg0_1_, sdai_ff_reg0_0_, N431,
         N432, N433, N468, N469, N470, N471, N491, N492, N493, N494, N495,
         busfree, N510, N511, rst_delay, clk_count1_ov, N653, N654, N655, N656,
         N657, clk_count2_ov, N685, N686, N687, N688, N689, N690, clkint,
         clkint_ff, N700, N746, N747, N748, N749, N1022, N1023, N1024, N1025,
         N1026, N1027, N1063, N1064, N1065, sclscl, starto_en, N1124, N1125,
         N1126, net12048, net12054, net12059, net12064, net12069, net12074,
         net12079, net12084, net12089, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n282,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454;
  wire   [2:0] fsmmod;
  wire   [4:0] fsmsta;
  wire   [3:0] framesync;
  wire   [2:0] fsmdet;
  wire   [2:0] setup_counter_r;
  wire   [2:0] scli_ff_reg0;
  wire   [2:0] indelay;
  wire   [2:0] fsmsync;
  wire   [1:0] bclkcnt;
  wire   [3:0] clk_count1;
  wire   [3:0] clk_count2;

  SNPS_CLOCK_GATE_HIGH_i2c_a0_0 clk_gate_i2ccon_reg ( .CLK(clk), .EN(N224), 
        .ENCLK(net12048), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_8 clk_gate_i2cdat_reg ( .CLK(clk), .EN(N296), 
        .ENCLK(net12054), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_7 clk_gate_setup_counter_r_reg ( .CLK(clk), .EN(
        N332), .ENCLK(net12059), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_6 clk_gate_i2cadr_reg ( .CLK(clk), .EN(N342), 
        .ENCLK(net12064), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_5 clk_gate_indelay_reg ( .CLK(clk), .EN(N468), 
        .ENCLK(net12069), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_4 clk_gate_framesync_reg ( .CLK(clk), .EN(N491), 
        .ENCLK(net12074), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_3 clk_gate_clk_count1_reg ( .CLK(clk), .EN(N653), 
        .ENCLK(net12079), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_2 clk_gate_clk_count2_reg ( .CLK(clk), .EN(N689), 
        .ENCLK(net12084), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_1 clk_gate_fsmsta_reg ( .CLK(clk), .EN(N1022), 
        .ENCLK(net12089), .TE(test_se) );
  SDFFQX1 scli_ff_reg ( .D(N180), .SIN(rst_delay), .SMC(test_se), .C(clk), .Q(
        scli_ff) );
  SDFFQX1 sdai_ff_reg ( .D(N181), .SIN(sclscl), .SMC(test_se), .C(clk), .Q(
        sdai_ff) );
  SDFFQX1 clk_count2_ov_reg ( .D(N690), .SIN(clk_count1[3]), .SMC(test_se), 
        .C(clk), .Q(clk_count2_ov) );
  SDFFQX1 sdai_ff_reg_reg_2_ ( .D(N433), .SIN(sdai_ff_reg0_1_), .SMC(test_se), 
        .C(clk), .Q(test_so1) );
  SDFFQX1 sdai_ff_reg_reg_1_ ( .D(N432), .SIN(sdai_ff_reg0_0_), .SMC(test_se), 
        .C(clk), .Q(sdai_ff_reg0_1_) );
  SDFFQX1 clk_count1_ov_reg ( .D(n505), .SIN(busfree), .SMC(test_se), .C(clk), 
        .Q(clk_count1_ov) );
  SDFFQX1 rst_delay_reg ( .D(n26), .SIN(pedetect), .SMC(test_se), .C(clk), .Q(
        rst_delay) );
  SDFFQX1 ack_bit_reg ( .D(n494), .SIN(test_si1), .SMC(test_se), .C(net12048), 
        .Q(ack_bit) );
  SDFFQX1 bsd7_reg ( .D(n491), .SIN(bclkcnt[1]), .SMC(test_se), .C(clk), .Q(
        bsd7) );
  SDFFQX1 clk_count2_reg_3_ ( .D(N688), .SIN(clk_count2[2]), .SMC(test_se), 
        .C(net12084), .Q(clk_count2[3]) );
  SDFFQX1 sdai_ff_reg_reg_0_ ( .D(N431), .SIN(sdai_ff), .SMC(test_se), .C(clk), 
        .Q(sdai_ff_reg0_0_) );
  SDFFQX1 sclscl_reg ( .D(n50), .SIN(sclo_int), .SMC(test_se), .C(clk), .Q(
        sclscl) );
  SDFFQX1 setup_counter_r_reg_2_ ( .D(N335), .SIN(setup_counter_r[1]), .SMC(
        test_se), .C(net12059), .Q(setup_counter_r[2]) );
  SDFFQX1 clk_count2_reg_1_ ( .D(N686), .SIN(clk_count2[0]), .SMC(test_se), 
        .C(net12084), .Q(clk_count2[1]) );
  SDFFQX1 clk_count2_reg_2_ ( .D(N687), .SIN(clk_count2[1]), .SMC(test_se), 
        .C(net12084), .Q(clk_count2[2]) );
  SDFFQX1 bclkcnt_reg_1_ ( .D(N511), .SIN(bclkcnt[0]), .SMC(test_se), .C(clk), 
        .Q(bclkcnt[1]) );
  SDFFQX1 indelay_reg_2_ ( .D(N471), .SIN(indelay[1]), .SMC(test_se), .C(
        net12069), .Q(indelay[2]) );
  SDFFQX1 bclkcnt_reg_0_ ( .D(N510), .SIN(adrcompen), .SMC(test_se), .C(clk), 
        .Q(bclkcnt[0]) );
  SDFFQX1 clkint_ff_reg ( .D(N700), .SIN(clk_count2[3]), .SMC(test_se), .C(clk), .Q(clkint_ff) );
  SDFFQX1 setup_counter_r_reg_0_ ( .D(N333), .SIN(sdao), .SMC(test_se), .C(
        net12059), .Q(setup_counter_r[0]) );
  SDFFQX1 write_data_r_reg ( .D(n500), .SIN(wait_for_setup_r), .SMC(test_se), 
        .C(clk), .Q(test_so2) );
  SDFFQX1 clk_count2_reg_0_ ( .D(N685), .SIN(clk_count2_ov), .SMC(test_se), 
        .C(net12084), .Q(clk_count2[0]) );
  SDFFQX1 bsd7_tmp_reg ( .D(n492), .SIN(bsd7), .SMC(test_se), .C(clk), .Q(
        bsd7_tmp) );
  SDFFQX1 busfree_reg ( .D(n506), .SIN(bsd7_tmp), .SMC(test_se), .C(clk), .Q(
        busfree) );
  SDFFQX1 indelay_reg_1_ ( .D(N470), .SIN(indelay[0]), .SMC(test_se), .C(
        net12069), .Q(indelay[1]) );
  SDFFQX1 clkint_reg ( .D(n504), .SIN(clkint_ff), .SMC(test_se), .C(clk), .Q(
        clkint) );
  SDFFQX1 indelay_reg_0_ ( .D(N469), .SIN(i2csta_o[7]), .SMC(test_se), .C(
        net12069), .Q(indelay[0]) );
  SDFFQX1 starto_en_reg ( .D(n490), .SIN(setup_counter_r[2]), .SMC(test_se), 
        .C(clk), .Q(starto_en) );
  SDFFQX1 scli_ff_reg_reg_1_ ( .D(N413), .SIN(scli_ff_reg0[0]), .SMC(test_se), 
        .C(clk), .Q(scli_ff_reg0[1]) );
  SDFFQX1 scli_ff_reg_reg_0_ ( .D(N412), .SIN(scli_ff), .SMC(test_se), .C(clk), 
        .Q(scli_ff_reg0[0]) );
  SDFFQX1 setup_counter_r_reg_1_ ( .D(n42), .SIN(setup_counter_r[0]), .SMC(
        test_se), .C(net12059), .Q(setup_counter_r[1]) );
  SDFFQX1 scli_ff_reg_reg_2_ ( .D(N414), .SIN(scli_ff_reg0[1]), .SMC(test_se), 
        .C(clk), .Q(scli_ff_reg0[2]) );
  SDFFQX1 fsmsync_reg_1_ ( .D(N747), .SIN(fsmsync[0]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[1]) );
  SDFFQX1 fsmsync_reg_0_ ( .D(N746), .SIN(fsmsta[4]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[0]) );
  SDFFQX1 fsmsync_reg_2_ ( .D(N748), .SIN(fsmsync[1]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[2]) );
  SDFFQX1 pedetect_reg ( .D(n497), .SIN(nedetect), .SMC(test_se), .C(clk), .Q(
        pedetect) );
  SDFFQX1 nedetect_reg ( .D(n498), .SIN(indelay[2]), .SMC(test_se), .C(clk), 
        .Q(nedetect) );
  SDFFQX1 sclint_reg ( .D(n499), .SIN(scli_ff_reg0[2]), .SMC(test_se), .C(clk), 
        .Q(sclint) );
  SDFFQX1 clk_count1_reg_2_ ( .D(N656), .SIN(clk_count1[1]), .SMC(test_se), 
        .C(net12079), .Q(clk_count1[2]) );
  SDFFQX1 clk_count1_reg_3_ ( .D(N657), .SIN(clk_count1[2]), .SMC(test_se), 
        .C(net12079), .Q(clk_count1[3]) );
  SDFFQX1 adrcompen_reg ( .D(n496), .SIN(adrcomp), .SMC(test_se), .C(clk), .Q(
        adrcompen) );
  SDFFQX1 adrcomp_reg ( .D(n501), .SIN(ack), .SMC(test_se), .C(clk), .Q(
        adrcomp) );
  SDFFQX1 clk_count1_reg_1_ ( .D(N655), .SIN(clk_count1[0]), .SMC(test_se), 
        .C(net12079), .Q(clk_count1[1]) );
  SDFFQX1 clk_count1_reg_0_ ( .D(N654), .SIN(clk_count1_ov), .SMC(test_se), 
        .C(net12079), .Q(clk_count1[0]) );
  SDFFQX1 ack_reg ( .D(n493), .SIN(ack_bit), .SMC(test_se), .C(clk), .Q(ack)
         );
  SDFFQX1 sdaint_reg ( .D(n507), .SIN(test_si2), .SMC(test_se), .C(clk), .Q(
        sdaint) );
  SDFFQX1 fsmdet_reg_0_ ( .D(N1063), .SIN(framesync[3]), .SMC(test_se), .C(clk), .Q(fsmdet[0]) );
  SDFFQX1 fsmdet_reg_1_ ( .D(N1064), .SIN(fsmdet[0]), .SMC(test_se), .C(clk), 
        .Q(fsmdet[1]) );
  SDFFQX1 framesync_reg_3_ ( .D(N495), .SIN(framesync[2]), .SMC(test_se), .C(
        net12074), .Q(framesync[3]) );
  SDFFQX1 fsmmod_reg_0_ ( .D(N1124), .SIN(fsmdet[2]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[0]) );
  SDFFQX1 fsmmod_reg_1_ ( .D(N1125), .SIN(fsmmod[0]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[1]) );
  SDFFQX1 fsmdet_reg_2_ ( .D(N1065), .SIN(fsmdet[1]), .SMC(test_se), .C(clk), 
        .Q(fsmdet[2]) );
  SDFFQX1 fsmmod_reg_2_ ( .D(N1126), .SIN(fsmmod[1]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[2]) );
  SDFFQX1 framesync_reg_1_ ( .D(N493), .SIN(framesync[0]), .SMC(test_se), .C(
        net12074), .Q(framesync[1]) );
  SDFFQX1 framesync_reg_2_ ( .D(N494), .SIN(framesync[1]), .SMC(test_se), .C(
        net12074), .Q(framesync[2]) );
  SDFFQX1 framesync_reg_0_ ( .D(N492), .SIN(clkint), .SMC(test_se), .C(
        net12074), .Q(framesync[0]) );
  SDFFQX1 fsmsta_reg_4_ ( .D(N1027), .SIN(n9), .SMC(test_se), .C(net12089), 
        .Q(fsmsta[4]) );
  SDFFQX1 fsmsta_reg_0_ ( .D(N1023), .SIN(fsmmod[2]), .SMC(test_se), .C(
        net12089), .Q(fsmsta[0]) );
  SDFFQX1 fsmsta_reg_2_ ( .D(N1025), .SIN(fsmsta[1]), .SMC(test_se), .C(
        net12089), .Q(fsmsta[2]) );
  SDFFQX1 fsmsta_reg_1_ ( .D(N1024), .SIN(fsmsta[0]), .SMC(test_se), .C(
        net12089), .Q(fsmsta[1]) );
  SDFFQX1 fsmsta_reg_3_ ( .D(N1026), .SIN(fsmsta[2]), .SMC(test_se), .C(
        net12089), .Q(fsmsta[3]) );
  SDFFQX1 wait_for_setup_r_reg ( .D(N336), .SIN(starto_en), .SMC(test_se), .C(
        clk), .Q(wait_for_setup_r) );
  SDFFQX1 sclo_int_reg ( .D(N749), .SIN(sclint), .SMC(test_se), .C(clk), .Q(
        sclo_int) );
  SDFFQX1 sdao_int_reg ( .D(n502), .SIN(sdaint), .SMC(test_se), .C(clk), .Q(
        sdao) );
  SDFFQX1 i2csta_reg_4_ ( .D(N410), .SIN(i2csta_o[6]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[7]) );
  SDFFQX1 i2csta_reg_3_ ( .D(N409), .SIN(i2csta_o[5]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[6]) );
  SDFFQX1 i2cdat_reg_7_ ( .D(N304), .SIN(i2cdat_o[6]), .SMC(test_se), .C(
        net12054), .Q(i2cdat_o[7]) );
  SDFFQX1 i2cadr_reg_3_ ( .D(N346), .SIN(i2cadr_o[2]), .SMC(test_se), .C(
        net12064), .Q(i2cadr_o[3]) );
  SDFFQX1 i2ccon_reg_5_ ( .D(N232), .SIN(i2ccon_o[4]), .SMC(test_se), .C(
        net12048), .Q(i2ccon_o[5]) );
  SDFFQX1 i2cdat_reg_6_ ( .D(N303), .SIN(i2cdat_o[5]), .SMC(test_se), .C(
        net12054), .Q(i2cdat_o[6]) );
  SDFFQX1 i2cadr_reg_1_ ( .D(N344), .SIN(i2cadr_o[0]), .SMC(test_se), .C(
        net12064), .Q(i2cadr_o[1]) );
  SDFFQX1 i2cdat_reg_3_ ( .D(N300), .SIN(i2cdat_o[2]), .SMC(test_se), .C(
        net12054), .Q(i2cdat_o[3]) );
  SDFFQX1 i2ccon_reg_1_ ( .D(N226), .SIN(i2ccon_o[0]), .SMC(test_se), .C(
        net12048), .Q(i2ccon_o[1]) );
  SDFFQX1 i2ccon_reg_6_ ( .D(N233), .SIN(i2ccon_o[5]), .SMC(test_se), .C(
        net12048), .Q(i2ccon_o[6]) );
  SDFFQX1 i2cadr_reg_0_ ( .D(N343), .SIN(fsmsync[2]), .SMC(test_se), .C(
        net12064), .Q(i2cadr_o[0]) );
  SDFFQX1 i2cdat_reg_0_ ( .D(N297), .SIN(i2ccon_o[7]), .SMC(test_se), .C(
        net12054), .Q(i2cdat_o[0]) );
  SDFFQX1 i2ccon_reg_0_ ( .D(N225), .SIN(i2cadr_o[7]), .SMC(test_se), .C(
        net12048), .Q(i2ccon_o[0]) );
  SDFFQX1 i2ccon_reg_7_ ( .D(N234), .SIN(i2ccon_o[6]), .SMC(test_se), .C(
        net12048), .Q(i2ccon_o[7]) );
  SDFFQX1 i2cdat_reg_1_ ( .D(N298), .SIN(i2cdat_o[0]), .SMC(test_se), .C(
        net12054), .Q(i2cdat_o[1]) );
  SDFFQX1 i2ccon_reg_3_ ( .D(n495), .SIN(i2ccon_o[2]), .SMC(test_se), .C(clk), 
        .Q(i2ccon_o[3]) );
  SDFFQX1 i2csta_reg_2_ ( .D(N408), .SIN(i2csta_o[4]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[5]) );
  SDFFQX1 i2csta_reg_0_ ( .D(N406), .SIN(i2cdat_o[7]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[3]) );
  SDFFQX1 i2csta_reg_1_ ( .D(N407), .SIN(i2csta_o[3]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[4]) );
  SDFFQX1 i2cadr_reg_5_ ( .D(N348), .SIN(i2cadr_o[4]), .SMC(test_se), .C(
        net12064), .Q(i2cadr_o[5]) );
  SDFFQX1 i2cadr_reg_4_ ( .D(N347), .SIN(i2cadr_o[3]), .SMC(test_se), .C(
        net12064), .Q(i2cadr_o[4]) );
  SDFFQX1 i2cadr_reg_6_ ( .D(N349), .SIN(i2cadr_o[5]), .SMC(test_se), .C(
        net12064), .Q(i2cadr_o[6]) );
  SDFFQX1 i2cadr_reg_7_ ( .D(N350), .SIN(i2cadr_o[6]), .SMC(test_se), .C(
        net12064), .Q(i2cadr_o[7]) );
  SDFFQX1 i2cadr_reg_2_ ( .D(N345), .SIN(i2cadr_o[1]), .SMC(test_se), .C(
        net12064), .Q(i2cadr_o[2]) );
  SDFFQX1 i2cdat_reg_5_ ( .D(N302), .SIN(i2cdat_o[4]), .SMC(test_se), .C(
        net12054), .Q(i2cdat_o[5]) );
  SDFFQX1 i2cdat_reg_4_ ( .D(N301), .SIN(i2cdat_o[3]), .SMC(test_se), .C(
        net12054), .Q(i2cdat_o[4]) );
  SDFFQX1 i2ccon_reg_2_ ( .D(N227), .SIN(i2ccon_o[1]), .SMC(test_se), .C(
        net12048), .Q(i2ccon_o[2]) );
  SDFFQX1 i2cdat_reg_2_ ( .D(N299), .SIN(i2cdat_o[1]), .SMC(test_se), .C(
        net12054), .Q(i2cdat_o[2]) );
  SDFFQX1 i2ccon_reg_4_ ( .D(n503), .SIN(si), .SMC(test_se), .C(clk), .Q(
        i2ccon_o[4]) );
  INVX1 U3 ( .A(1'b1), .Y(i2csta_o[0]) );
  INVX1 U5 ( .A(1'b1), .Y(i2csta_o[1]) );
  INVX1 U7 ( .A(1'b1), .Y(i2csta_o[2]) );
  BUFX3 U9 ( .A(n443), .Y(n7) );
  INVX1 U10 ( .A(si), .Y(n8) );
  INVX1 U11 ( .A(n439), .Y(n9) );
  INVX1 U12 ( .A(n193), .Y(n10) );
  BUFX3 U13 ( .A(i2ccon_o[3]), .Y(si) );
  INVX1 U14 ( .A(n85), .Y(n12) );
  NAND2X1 U15 ( .A(framesync[3]), .B(n207), .Y(n13) );
  NOR4XL U16 ( .A(n110), .B(n443), .C(fsmsta[0]), .D(fsmsta[3]), .Y(n162) );
  INVX1 U17 ( .A(n29), .Y(n24) );
  INVX1 U18 ( .A(n28), .Y(n23) );
  INVX1 U19 ( .A(n29), .Y(n25) );
  INVX1 U20 ( .A(n224), .Y(n36) );
  INVX1 U21 ( .A(n135), .Y(n33) );
  NAND2X1 U22 ( .A(n24), .B(n135), .Y(N224) );
  OAI21X1 U23 ( .B(n309), .C(n15), .A(n31), .Y(N343) );
  OAI21X1 U24 ( .B(n18), .C(n309), .A(n25), .Y(N346) );
  OAI21X1 U25 ( .B(n22), .C(n309), .A(n25), .Y(N350) );
  NOR2X1 U26 ( .A(n309), .B(n16), .Y(N344) );
  NOR2X1 U27 ( .A(n309), .B(n20), .Y(N348) );
  NOR2X1 U28 ( .A(n309), .B(n17), .Y(N345) );
  NOR2X1 U29 ( .A(n309), .B(n21), .Y(N349) );
  NOR2X1 U30 ( .A(n19), .B(n309), .Y(N347) );
  NAND2X1 U31 ( .A(n24), .B(n309), .Y(N342) );
  NOR2X1 U32 ( .A(n27), .B(n15), .Y(N225) );
  NOR2X1 U33 ( .A(n27), .B(n21), .Y(N233) );
  NOR2X1 U34 ( .A(n27), .B(n17), .Y(N227) );
  NOR2X1 U35 ( .A(n27), .B(n16), .Y(N226) );
  NOR2X1 U36 ( .A(n27), .B(n22), .Y(N234) );
  NOR2X1 U37 ( .A(n27), .B(n20), .Y(N232) );
  INVX1 U38 ( .A(n30), .Y(n29) );
  INVX1 U39 ( .A(n30), .Y(n28) );
  INVX1 U40 ( .A(n431), .Y(n86) );
  INVX1 U41 ( .A(n31), .Y(n26) );
  INVX1 U42 ( .A(n31), .Y(n27) );
  NAND42X1 U43 ( .C(sfraddr[0]), .D(sfraddr[2]), .A(sfraddr[1]), .B(n311), .Y(
        n224) );
  NOR42XL U44 ( .C(sfraddr[4]), .D(sfraddr[3]), .A(sfraddr[5]), .B(n329), .Y(
        n311) );
  NAND2X1 U45 ( .A(sfrwe), .B(sfraddr[6]), .Y(n329) );
  AOI21X1 U46 ( .B(n224), .C(n228), .A(n318), .Y(n214) );
  NOR2X1 U47 ( .A(n35), .B(n322), .Y(n318) );
  NAND42X1 U48 ( .C(sfraddr[0]), .D(sfraddr[1]), .A(sfraddr[2]), .B(n311), .Y(
        n135) );
  NAND3X1 U49 ( .A(n33), .B(n25), .C(sfrdatai[3]), .Y(n198) );
  NAND4X1 U50 ( .A(sfraddr[0]), .B(sfraddr[1]), .C(n310), .D(n311), .Y(n309)
         );
  NOR2X1 U51 ( .A(sfraddr[2]), .B(n26), .Y(n310) );
  INVX1 U52 ( .A(sfrdatai[7]), .Y(n22) );
  INVX1 U53 ( .A(sfrdatai[4]), .Y(n19) );
  NAND21X1 U54 ( .B(sdai), .A(n23), .Y(N181) );
  INVX1 U55 ( .A(sfrdatai[5]), .Y(n20) );
  INVX1 U56 ( .A(sfrdatai[6]), .Y(n21) );
  INVX1 U57 ( .A(sfrdatai[1]), .Y(n16) );
  INVX1 U58 ( .A(sfrdatai[2]), .Y(n17) );
  INVX1 U59 ( .A(sfrdatai[0]), .Y(n15) );
  INVX1 U60 ( .A(sfrdatai[3]), .Y(n18) );
  INVX1 U61 ( .A(n324), .Y(n111) );
  NOR32XL U62 ( .B(n86), .C(n433), .A(n157), .Y(n357) );
  NAND2X1 U63 ( .A(n201), .B(n24), .Y(n431) );
  NAND2X1 U64 ( .A(n152), .B(n97), .Y(n376) );
  NOR2X1 U65 ( .A(n88), .B(n210), .Y(n322) );
  INVX1 U66 ( .A(rst), .Y(n30) );
  INVX1 U67 ( .A(n403), .Y(n82) );
  INVX1 U68 ( .A(n228), .Y(n89) );
  AND2X1 U69 ( .A(n385), .B(n386), .Y(n361) );
  NAND41X1 U70 ( .D(n161), .A(n363), .B(n325), .C(n364), .Y(n358) );
  OAI21X1 U71 ( .B(n365), .C(n362), .A(n97), .Y(n363) );
  NAND41X1 U72 ( .D(n357), .A(n77), .B(n403), .C(n430), .Y(N1022) );
  NOR2X1 U73 ( .A(n39), .B(n431), .Y(n430) );
  INVX1 U74 ( .A(rst), .Y(n31) );
  NAND2X1 U75 ( .A(n147), .B(n143), .Y(n145) );
  INVX1 U76 ( .A(n369), .Y(n77) );
  INVX1 U77 ( .A(n132), .Y(n68) );
  INVX1 U78 ( .A(n393), .Y(n98) );
  INVX1 U79 ( .A(n192), .Y(n101) );
  INVX1 U80 ( .A(n251), .Y(n103) );
  NAND2X1 U81 ( .A(n24), .B(n105), .Y(n238) );
  INVX1 U82 ( .A(n308), .Y(n437) );
  INVX1 U83 ( .A(n236), .Y(n435) );
  INVX1 U84 ( .A(n261), .Y(n52) );
  INVX1 U85 ( .A(n231), .Y(n71) );
  INVX1 U86 ( .A(n284), .Y(n37) );
  OAI21X1 U87 ( .B(n216), .C(n66), .A(n217), .Y(n492) );
  GEN2XL U88 ( .D(n22), .E(n35), .C(n181), .B(n31), .A(n34), .Y(n217) );
  INVX1 U89 ( .A(n216), .Y(n34) );
  OAI21BBX1 U90 ( .A(n36), .B(n215), .C(n218), .Y(n216) );
  OAI22AX1 U91 ( .D(n211), .C(n212), .A(n96), .B(n211), .Y(n493) );
  AND2X1 U92 ( .A(n213), .B(n94), .Y(n212) );
  OAI21X1 U93 ( .B(n214), .C(n80), .A(n213), .Y(n211) );
  NOR2X1 U94 ( .A(n26), .B(n215), .Y(n213) );
  INVX1 U95 ( .A(n226), .Y(n35) );
  OAI22AX1 U96 ( .D(n223), .C(n322), .A(n224), .B(n89), .Y(n320) );
  NOR2X1 U97 ( .A(n319), .B(n320), .Y(n317) );
  OAI32X1 U98 ( .A(n135), .B(n27), .C(n32), .D(n453), .E(n136), .Y(n503) );
  INVX1 U99 ( .A(n136), .Y(n32) );
  OAI221X1 U100 ( .A(n33), .B(n137), .C(n135), .D(n19), .E(n31), .Y(n136) );
  AOI21BBXL U101 ( .B(n123), .C(n122), .A(n119), .Y(n137) );
  AOI21X1 U102 ( .B(n319), .C(n36), .A(n320), .Y(n179) );
  OAI22X1 U103 ( .A(n317), .B(n16), .C(n214), .D(n451), .Y(N298) );
  OAI22X1 U104 ( .A(n317), .B(n18), .C(n214), .D(n447), .Y(N300) );
  OAI22X1 U105 ( .A(n317), .B(n17), .C(n214), .D(n454), .Y(N299) );
  OAI22X1 U106 ( .A(n317), .B(n15), .C(n214), .D(n96), .Y(N297) );
  AOI22X1 U107 ( .A(n88), .B(n223), .C(n215), .D(n224), .Y(n222) );
  NAND21X1 U108 ( .B(scli), .A(n23), .Y(N180) );
  NOR2X1 U109 ( .A(n442), .B(n443), .Y(n159) );
  OAI221X1 U110 ( .A(n374), .B(n377), .C(n393), .D(n302), .E(n407), .Y(n392)
         );
  AOI222XL U111 ( .A(n408), .B(n193), .C(n436), .D(n160), .E(n409), .F(n410), 
        .Y(n407) );
  INVX1 U112 ( .A(n303), .Y(n436) );
  OAI221X1 U113 ( .A(n13), .B(n384), .C(n10), .D(n296), .E(n383), .Y(n410) );
  INVX1 U114 ( .A(n193), .Y(n97) );
  NAND2X1 U115 ( .A(n398), .B(n159), .Y(n324) );
  NAND2X1 U116 ( .A(n328), .B(n443), .Y(n296) );
  NAND2X1 U117 ( .A(n111), .B(n439), .Y(n383) );
  NOR21XL U118 ( .B(n323), .A(n150), .Y(n228) );
  NAND42X1 U119 ( .C(n336), .D(n251), .A(n151), .B(n102), .Y(n164) );
  NAND42X1 U120 ( .C(n423), .D(n399), .A(n364), .B(n424), .Y(n406) );
  NAND4X1 U121 ( .A(n328), .B(n159), .C(n95), .D(n13), .Y(n424) );
  OAI22X1 U122 ( .A(n385), .B(n393), .C(n386), .D(n394), .Y(n423) );
  OAI211X1 U123 ( .C(n305), .D(n438), .A(n324), .B(n325), .Y(n150) );
  NOR2X1 U124 ( .A(n193), .B(n446), .Y(n393) );
  NOR4XL U125 ( .A(n431), .B(n80), .C(n157), .D(n433), .Y(n369) );
  NOR2X1 U126 ( .A(n104), .B(n107), .Y(n251) );
  AND2X1 U127 ( .A(n323), .B(n150), .Y(n210) );
  NOR2X1 U128 ( .A(n28), .B(n194), .Y(n121) );
  AOI21X1 U129 ( .B(n194), .C(n342), .A(n420), .Y(n201) );
  NAND4X1 U130 ( .A(n86), .B(n205), .C(n202), .D(n157), .Y(n403) );
  OAI21X1 U131 ( .B(n387), .C(n77), .A(n388), .Y(N1025) );
  OAI21BBX1 U132 ( .A(n166), .B(n96), .C(n357), .Y(n388) );
  NOR4XL U133 ( .A(n389), .B(n390), .C(n391), .D(n392), .Y(n387) );
  NOR2X1 U134 ( .A(n97), .B(n380), .Y(n391) );
  NOR2X1 U135 ( .A(n181), .B(n40), .Y(n215) );
  NAND3X1 U136 ( .A(n295), .B(n112), .C(n306), .Y(n384) );
  INVX1 U137 ( .A(n315), .Y(n43) );
  NAND2X1 U138 ( .A(n194), .B(n452), .Y(n180) );
  INVX1 U139 ( .A(n233), .Y(n452) );
  NAND3X1 U140 ( .A(n160), .B(n112), .C(n295), .Y(n325) );
  INVX1 U141 ( .A(n366), .Y(n39) );
  OAI211X1 U142 ( .C(n418), .D(n77), .A(n367), .B(n419), .Y(N1023) );
  NOR2X1 U143 ( .A(n420), .B(n39), .Y(n419) );
  NOR4XL U144 ( .A(n421), .B(n406), .C(n422), .D(n359), .Y(n418) );
  AOI21X1 U145 ( .B(n411), .C(n383), .A(n393), .Y(n422) );
  INVX1 U146 ( .A(n181), .Y(n88) );
  NAND2X1 U147 ( .A(n379), .B(n383), .Y(n408) );
  INVX1 U148 ( .A(n194), .Y(n87) );
  INVX1 U149 ( .A(n428), .Y(n108) );
  OAI211X1 U150 ( .C(n110), .D(n429), .A(n378), .B(n400), .Y(n428) );
  NAND2X1 U151 ( .A(n443), .B(n439), .Y(n429) );
  INVX1 U152 ( .A(n154), .Y(n102) );
  INVX1 U153 ( .A(n326), .Y(n113) );
  INVX1 U154 ( .A(n398), .Y(n110) );
  NOR21XL U155 ( .B(n151), .A(n152), .Y(n147) );
  NOR2X1 U156 ( .A(n276), .B(n26), .Y(n125) );
  INVX1 U157 ( .A(n206), .Y(n99) );
  NOR2X1 U158 ( .A(n74), .B(n69), .Y(n132) );
  OAI21X1 U159 ( .B(n149), .C(n97), .A(n150), .Y(n143) );
  NOR2X1 U160 ( .A(n453), .B(n164), .Y(n192) );
  AND3X1 U161 ( .A(n380), .B(n325), .C(n384), .Y(n411) );
  NAND2X1 U162 ( .A(n87), .B(n138), .Y(n157) );
  OAI31XL U163 ( .A(n376), .B(n96), .C(n109), .D(n435), .Y(n359) );
  OAI22X1 U164 ( .A(n393), .B(n386), .C(n374), .D(n378), .Y(n390) );
  NOR2X1 U165 ( .A(n79), .B(n81), .Y(n152) );
  AND2X1 U166 ( .A(n382), .B(n94), .Y(n399) );
  AOI21X1 U167 ( .B(n96), .C(n357), .A(n27), .Y(n367) );
  NOR3XL U168 ( .A(n80), .B(n162), .C(n376), .Y(n433) );
  AOI211X1 U169 ( .C(n109), .D(n164), .A(n165), .B(n79), .Y(n163) );
  OAI21X1 U170 ( .B(n166), .C(n96), .A(n167), .Y(n165) );
  OAI22X1 U171 ( .A(n166), .B(n450), .C(n168), .D(n169), .Y(n167) );
  NAND3X1 U172 ( .A(n170), .B(n171), .C(n172), .Y(n169) );
  OAI22AX1 U173 ( .D(n139), .C(n140), .A(n139), .B(n446), .Y(n502) );
  NOR32XL U174 ( .B(n452), .C(n141), .A(n142), .Y(n140) );
  NAND4X1 U175 ( .A(n452), .B(n141), .C(n148), .D(n147), .Y(n139) );
  AOI21X1 U176 ( .B(n81), .C(n153), .A(n154), .Y(n141) );
  NOR3XL U177 ( .A(n193), .B(n96), .C(n296), .Y(n382) );
  OAI31XL U178 ( .A(n80), .B(n186), .C(n182), .D(n187), .Y(n497) );
  NAND4X1 U179 ( .A(n24), .B(n85), .C(n183), .D(n188), .Y(n187) );
  NOR3XL U180 ( .A(n48), .B(n55), .C(n54), .Y(n188) );
  OAI31XL U181 ( .A(n44), .B(n313), .C(n43), .D(n312), .Y(N335) );
  AOI211X1 U182 ( .C(n52), .D(n57), .A(n260), .B(n263), .Y(N687) );
  AOI211X1 U183 ( .C(n56), .D(n53), .A(n260), .B(n261), .Y(N686) );
  AOI211X1 U184 ( .C(n74), .D(n69), .A(n267), .B(n132), .Y(N655) );
  NAND2X1 U185 ( .A(n306), .B(n159), .Y(n385) );
  NAND2X1 U186 ( .A(n425), .B(n443), .Y(n386) );
  NAND2X1 U187 ( .A(n97), .B(n446), .Y(n394) );
  NAND2X1 U188 ( .A(n377), .B(n378), .Y(n362) );
  NAND2X1 U189 ( .A(n54), .B(n23), .Y(N414) );
  NAND2X1 U190 ( .A(n55), .B(n24), .Y(N413) );
  NAND2X1 U191 ( .A(n379), .B(n380), .Y(n365) );
  NAND2X1 U192 ( .A(n43), .B(n312), .Y(N336) );
  NAND2X1 U193 ( .A(n24), .B(n118), .Y(n506) );
  OAI21X1 U194 ( .B(n119), .C(n120), .A(n121), .Y(n118) );
  OAI31XL U195 ( .A(n85), .B(n122), .C(n123), .D(n67), .Y(n120) );
  NAND2X1 U196 ( .A(n125), .B(n75), .Y(N700) );
  INVX1 U197 ( .A(n305), .Y(n434) );
  INVX1 U198 ( .A(n162), .Y(n109) );
  INVX1 U199 ( .A(n287), .Y(n100) );
  INVX1 U200 ( .A(n306), .Y(n438) );
  NOR2X1 U201 ( .A(n40), .B(n26), .Y(n300) );
  NAND21X1 U202 ( .B(n242), .A(n73), .Y(n240) );
  NOR2X1 U203 ( .A(n53), .B(n56), .Y(n261) );
  NOR2X1 U204 ( .A(n72), .B(n84), .Y(n231) );
  NOR2X1 U205 ( .A(n437), .B(n305), .Y(n236) );
  NOR2X1 U206 ( .A(n439), .B(n444), .Y(n308) );
  NOR2X1 U207 ( .A(n293), .B(n97), .Y(n284) );
  NOR2X1 U208 ( .A(n434), .B(n444), .Y(n161) );
  NOR2X1 U209 ( .A(n57), .B(n52), .Y(n263) );
  AOI21X1 U210 ( .B(n51), .C(n83), .A(n71), .Y(n257) );
  AOI21X1 U211 ( .B(n132), .C(n64), .A(n65), .Y(n126) );
  INVX1 U212 ( .A(n183), .Y(n47) );
  NAND2X1 U213 ( .A(n159), .B(n160), .Y(n364) );
  NOR2X1 U214 ( .A(n83), .B(n72), .Y(n244) );
  OAI21AX1 U215 ( .B(n85), .C(n47), .A(n182), .Y(n499) );
  INVX1 U216 ( .A(n409), .Y(n95) );
  INVX1 U217 ( .A(n297), .Y(n70) );
  NAND4X1 U218 ( .A(n300), .B(n301), .C(n302), .D(n440), .Y(N410) );
  NAND2X1 U219 ( .A(n161), .B(n7), .Y(n301) );
  NAND2X1 U220 ( .A(n122), .B(n63), .Y(n338) );
  INVX1 U221 ( .A(n253), .Y(n63) );
  INVX1 U222 ( .A(n243), .Y(n73) );
  INVX1 U223 ( .A(n160), .Y(n440) );
  NOR2X1 U224 ( .A(n299), .B(n70), .Y(N470) );
  XNOR2XL U225 ( .A(n58), .B(n59), .Y(n299) );
  INVX1 U226 ( .A(n245), .Y(n51) );
  NAND2X1 U227 ( .A(n297), .B(n51), .Y(N468) );
  INVX1 U228 ( .A(n153), .Y(n105) );
  INVX1 U229 ( .A(n122), .Y(n62) );
  INVX1 U230 ( .A(n339), .Y(n61) );
  INVX1 U231 ( .A(n258), .Y(n41) );
  INVX1 U232 ( .A(n295), .Y(n441) );
  NOR2X1 U233 ( .A(n93), .B(n92), .Y(n351) );
  NAND4X1 U234 ( .A(n291), .B(n121), .C(n293), .D(n99), .Y(N491) );
  INVX1 U235 ( .A(n133), .Y(n64) );
  AO22AXL U236 ( .A(n219), .B(n220), .C(bsd7), .D(n220), .Y(n491) );
  OAI211X1 U237 ( .C(n227), .D(n181), .A(n25), .B(n221), .Y(n219) );
  NAND3X1 U238 ( .A(n221), .B(n218), .C(n222), .Y(n220) );
  NOR2X1 U239 ( .A(n210), .B(n228), .Y(n221) );
  NOR2X1 U240 ( .A(i2ccon_o[3]), .B(n36), .Y(n226) );
  AND3X1 U241 ( .A(n180), .B(n225), .C(n25), .Y(n218) );
  NAND4X1 U242 ( .A(n226), .B(n88), .C(nedetect), .D(n80), .Y(n225) );
  AOI221XL U243 ( .A(i2cdat_o[7]), .B(n226), .C(sfrdatai[7]), .D(n223), .E(
        n229), .Y(n227) );
  AOI21X1 U244 ( .B(n85), .C(n66), .A(n40), .Y(n229) );
  NOR2X1 U245 ( .A(n224), .B(i2ccon_o[3]), .Y(n223) );
  OAI21X1 U246 ( .B(intack), .C(N224), .A(n198), .Y(n199) );
  OAI22AX1 U247 ( .D(i2cdat_o[3]), .C(n214), .A(n317), .B(n19), .Y(N301) );
  OAI22AX1 U248 ( .D(i2cdat_o[4]), .C(n214), .A(n317), .B(n20), .Y(N302) );
  OAI22AX1 U249 ( .D(i2cdat_o[5]), .C(n214), .A(n317), .B(n21), .Y(N303) );
  OAI22AX1 U250 ( .D(i2cdat_o[6]), .C(n214), .A(n317), .B(n22), .Y(N304) );
  OAI21X1 U251 ( .B(n177), .C(n178), .A(n179), .Y(n500) );
  NAND3X1 U252 ( .A(n452), .B(n33), .C(test_so2), .Y(n178) );
  NAND4X1 U253 ( .A(n180), .B(n89), .C(n35), .D(n181), .Y(n177) );
  ENOX1 U254 ( .A(n40), .B(n195), .C(n195), .D(n196), .Y(n495) );
  OAI21X1 U255 ( .B(n197), .C(N224), .A(n198), .Y(n196) );
  NAND2X1 U256 ( .A(n199), .B(n197), .Y(n195) );
  OAI21BBX1 U257 ( .A(n200), .B(n201), .C(i2ccon_o[6]), .Y(n197) );
  NAND3X1 U258 ( .A(n321), .B(n25), .C(n179), .Y(N296) );
  OAI21X1 U259 ( .B(n318), .C(n228), .A(pedetect), .Y(n321) );
  ENOX1 U260 ( .A(n208), .B(n209), .C(n208), .D(ack_bit), .Y(n494) );
  NOR2X1 U261 ( .A(n26), .B(sfrdatai[2]), .Y(n209) );
  AOI31X1 U262 ( .A(n210), .B(n33), .C(si), .D(n29), .Y(n208) );
  NOR2X1 U263 ( .A(wait_for_setup_r), .B(n445), .Y(sclo) );
  INVX1 U264 ( .A(sclo_int), .Y(n445) );
  NAND2X1 U265 ( .A(framesync[3]), .B(n207), .Y(n193) );
  NOR3XL U266 ( .A(fsmsta[3]), .B(fsmsta[4]), .C(fsmsta[2]), .Y(n328) );
  INVX1 U267 ( .A(fsmsta[1]), .Y(n443) );
  NOR2X1 U268 ( .A(n112), .B(fsmsta[4]), .Y(n398) );
  NOR3XL U269 ( .A(framesync[1]), .B(framesync[2]), .C(framesync[0]), .Y(n207)
         );
  INVX1 U270 ( .A(fsmsta[2]), .Y(n112) );
  OAI221X1 U271 ( .A(n401), .B(n77), .C(n81), .D(n366), .E(n402), .Y(N1024) );
  AOI31X1 U272 ( .A(n166), .B(n96), .C(n357), .D(n82), .Y(n402) );
  NOR4XL U273 ( .A(n404), .B(n405), .C(n392), .D(n406), .Y(n401) );
  ENOX1 U274 ( .A(n411), .B(n98), .C(n408), .D(sdao), .Y(n405) );
  INVX1 U275 ( .A(fsmsta[0]), .Y(n442) );
  OAI211X1 U276 ( .C(n258), .D(n432), .A(n157), .B(n86), .Y(n366) );
  NOR32XL U277 ( .B(n207), .C(n40), .A(framesync[3]), .Y(n432) );
  OAI31XL U278 ( .A(n327), .B(fsmsta[3]), .C(n159), .D(n282), .Y(n326) );
  INVX1 U279 ( .A(n328), .Y(n282) );
  OAI21X1 U280 ( .B(fsmsta[4]), .C(n443), .A(fsmsta[2]), .Y(n327) );
  AOI22AXL U281 ( .A(n44), .B(n313), .D(n316), .C(n184), .Y(n315) );
  NOR2X1 U282 ( .A(n26), .B(test_so2), .Y(n316) );
  NOR3XL U283 ( .A(n90), .B(fsmdet[2]), .C(n92), .Y(n194) );
  NOR2X1 U284 ( .A(n444), .B(fsmsta[3]), .Y(n160) );
  NOR2X1 U285 ( .A(n442), .B(fsmsta[1]), .Y(n295) );
  NOR2X1 U286 ( .A(n439), .B(fsmsta[4]), .Y(n306) );
  NOR3XL U287 ( .A(n106), .B(fsmmod[2]), .C(n104), .Y(n154) );
  NAND3X1 U288 ( .A(i2ccon_o[6]), .B(n326), .C(n121), .Y(n181) );
  INVX1 U289 ( .A(fsmsta[3]), .Y(n439) );
  AND3X1 U290 ( .A(n121), .B(i2ccon_o[6]), .C(n113), .Y(n323) );
  AOI21X1 U291 ( .B(n106), .C(fsmmod[2]), .A(n342), .Y(n151) );
  OAI221X1 U292 ( .A(n322), .B(n40), .C(n26), .D(i2ccon_o[6]), .E(n180), .Y(
        n319) );
  OAI21X1 U293 ( .B(framesync[3]), .C(n207), .A(n13), .Y(n205) );
  NAND2X1 U294 ( .A(n159), .B(fsmsta[2]), .Y(n303) );
  AOI221XL U295 ( .A(n365), .B(n193), .C(n374), .D(n362), .E(n375), .Y(n373)
         );
  OAI22X1 U296 ( .A(ack), .B(n376), .C(n439), .D(n434), .Y(n375) );
  NOR3XL U297 ( .A(n110), .B(fsmsta[0]), .C(n439), .Y(n425) );
  NAND2X1 U298 ( .A(i2ccon_o[6]), .B(n24), .Y(n233) );
  OAI21X1 U299 ( .B(n394), .C(n379), .A(n426), .Y(n421) );
  AOI33X1 U300 ( .A(sdaint), .B(n427), .C(n97), .D(n95), .E(n13), .F(n295), 
        .Y(n426) );
  OAI211X1 U301 ( .C(ack), .D(n296), .A(n377), .B(n108), .Y(n427) );
  NOR3XL U302 ( .A(fsmmod[0]), .B(fsmmod[2]), .C(n104), .Y(n336) );
  NAND2X1 U303 ( .A(sclint), .B(n24), .Y(n184) );
  NOR3XL U304 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(n106), .Y(n342) );
  INVX1 U305 ( .A(fsmsta[4]), .Y(n444) );
  NOR3XL U306 ( .A(n87), .B(fsmmod[0]), .C(n103), .Y(n420) );
  NAND3X1 U307 ( .A(n160), .B(n443), .C(fsmsta[2]), .Y(n378) );
  NAND2X1 U308 ( .A(n425), .B(fsmsta[1]), .Y(n379) );
  AOI32X1 U309 ( .A(pedetect), .B(n202), .C(n97), .D(n203), .E(n157), .Y(n200)
         );
  ENOX1 U310 ( .A(n204), .B(n81), .C(n202), .D(n205), .Y(n203) );
  NOR2X1 U311 ( .A(n206), .B(n207), .Y(n204) );
  INVX1 U312 ( .A(fsmmod[0]), .Y(n106) );
  OR2X1 U313 ( .A(n164), .B(adrcomp), .Y(n202) );
  INVX1 U314 ( .A(fsmmod[1]), .Y(n104) );
  OAI211X1 U315 ( .C(adrcomp), .D(n366), .A(n367), .B(n368), .Y(N1026) );
  AOI21X1 U316 ( .B(n369), .C(n370), .A(n82), .Y(n368) );
  NAND4X1 U317 ( .A(n371), .B(n435), .C(n372), .D(n373), .Y(n370) );
  OAI21BBX1 U318 ( .A(n384), .B(n361), .C(n98), .Y(n371) );
  NAND2X1 U319 ( .A(n328), .B(fsmsta[1]), .Y(n400) );
  INVX1 U320 ( .A(fsmmod[2]), .Y(n107) );
  INVX1 U321 ( .A(fsmdet[1]), .Y(n92) );
  NOR2X1 U322 ( .A(n43), .B(setup_counter_r[0]), .Y(N333) );
  INVX1 U323 ( .A(fsmdet[0]), .Y(n90) );
  INVX1 U324 ( .A(n314), .Y(n42) );
  AOI32X1 U325 ( .A(setup_counter_r[1]), .B(n315), .C(setup_counter_r[0]), .D(
        n46), .E(N333), .Y(n314) );
  INVX1 U326 ( .A(setup_counter_r[1]), .Y(n46) );
  NOR21XL U327 ( .B(framesync[3]), .A(n146), .Y(n206) );
  GEN2XL U328 ( .D(framesync[3]), .E(n283), .C(n149), .B(n284), .A(n285), .Y(
        N495) );
  AO2222XL U329 ( .A(n97), .B(n412), .C(n162), .D(n413), .E(n414), .F(n193), 
        .G(n415), .H(n305), .Y(n404) );
  AOI31X1 U330 ( .A(n440), .B(n438), .C(n437), .D(n443), .Y(n415) );
  OAI22X1 U331 ( .A(ack), .B(n296), .C(n417), .D(n378), .Y(n412) );
  OAI21X1 U332 ( .B(n108), .C(n95), .A(n400), .Y(n414) );
  NAND32X1 U333 ( .B(framesync[1]), .C(framesync[2]), .A(framesync[0]), .Y(
        n146) );
  INVX1 U334 ( .A(n273), .Y(n65) );
  OAI211X1 U335 ( .C(i2ccon_o[1]), .D(n274), .A(clk_count1[3]), .B(n275), .Y(
        n273) );
  AOI211X1 U336 ( .C(n74), .D(n69), .A(n133), .B(n449), .Y(n274) );
  AOI31X1 U337 ( .A(n133), .B(n449), .C(n68), .D(n272), .Y(n275) );
  OA21X1 U338 ( .B(n12), .C(n8), .A(n138), .Y(n291) );
  XNOR2XL U339 ( .A(i2cdat_o[2]), .B(i2cadr_o[3]), .Y(n176) );
  NOR2X1 U340 ( .A(n99), .B(i2ccon_o[3]), .Y(n258) );
  NOR2X1 U341 ( .A(fsmsta[2]), .B(fsmsta[0]), .Y(n305) );
  XNOR2XL U342 ( .A(i2cdat_o[1]), .B(i2cadr_o[2]), .Y(n170) );
  XNOR2XL U343 ( .A(i2cdat_o[0]), .B(i2cadr_o[1]), .Y(n171) );
  XNOR2XL U344 ( .A(i2cdat_o[4]), .B(i2cadr_o[5]), .Y(n172) );
  OAI32X1 U345 ( .A(n143), .B(ack_bit), .C(n78), .D(n144), .E(n145), .Y(n142)
         );
  INVX1 U346 ( .A(n147), .Y(n78) );
  AOI211X1 U347 ( .C(framesync[3]), .D(n146), .A(bsd7), .B(n113), .Y(n144) );
  INVX1 U348 ( .A(i2ccon_o[3]), .Y(n40) );
  NOR2X1 U349 ( .A(n446), .B(sdaint), .Y(n409) );
  NAND2X1 U350 ( .A(clk_count1[3]), .B(clk_count1[2]), .Y(n133) );
  NOR3XL U351 ( .A(n106), .B(fsmmod[1]), .C(n107), .Y(n115) );
  NAND2X1 U352 ( .A(framesync[1]), .B(framesync[0]), .Y(n287) );
  NOR3XL U353 ( .A(clk_count1[1]), .B(clk_count1[2]), .C(clk_count1[0]), .Y(
        n272) );
  AOI22X1 U354 ( .A(n381), .B(n95), .C(n382), .D(sdaint), .Y(n372) );
  OAI21X1 U355 ( .B(n193), .C(n383), .A(n384), .Y(n381) );
  NOR2X1 U356 ( .A(n343), .B(n333), .Y(N1124) );
  AOI221XL U357 ( .A(n115), .B(n334), .C(n342), .D(n60), .E(n345), .Y(n343) );
  OAI21X1 U358 ( .B(n346), .C(n339), .A(n347), .Y(n345) );
  OAI21BBX1 U359 ( .A(n338), .B(sclint), .C(n154), .Y(n347) );
  AOI21AX1 U360 ( .B(nedetect), .C(n149), .A(n145), .Y(n148) );
  NAND2X1 U361 ( .A(fsmdet[2]), .B(n352), .Y(n138) );
  NOR3XL U362 ( .A(i2ccon_o[2]), .B(sdaint), .C(n13), .Y(n374) );
  NAND3X1 U363 ( .A(n398), .B(n295), .C(fsmsta[3]), .Y(n380) );
  NOR2X1 U364 ( .A(n283), .B(framesync[3]), .Y(n149) );
  NAND4X1 U365 ( .A(n454), .B(n447), .C(n451), .D(n416), .Y(n166) );
  NOR4XL U366 ( .A(i2cdat_o[6]), .B(i2cdat_o[5]), .C(i2cdat_o[4]), .D(
        i2cdat_o[3]), .Y(n416) );
  AOI31X1 U367 ( .A(scli_ff_reg0[2]), .B(N414), .C(N413), .D(n47), .Y(n186) );
  OAI211X1 U368 ( .C(n385), .D(n394), .A(n395), .B(n396), .Y(n389) );
  AO21X1 U369 ( .B(n95), .C(n13), .A(n400), .Y(n395) );
  AOI211X1 U370 ( .C(n397), .D(n398), .A(n399), .B(n162), .Y(n396) );
  NOR2X1 U371 ( .A(fsmsta[3]), .B(fsmsta[1]), .Y(n397) );
  NAND2X1 U372 ( .A(clk_count1_ov), .B(n125), .Y(n260) );
  NAND2X1 U373 ( .A(n125), .B(n270), .Y(n267) );
  OAI211X1 U374 ( .C(i2ccon_o[7]), .D(n65), .A(n271), .B(n131), .Y(n270) );
  OAI21X1 U375 ( .B(n133), .C(n69), .A(n129), .Y(n271) );
  AOI33X1 U376 ( .A(n153), .B(n40), .C(starto_en), .D(n336), .E(n296), .F(n258), .Y(n346) );
  NAND3X1 U377 ( .A(n101), .B(n138), .C(i2ccon_o[6]), .Y(n119) );
  OAI22X1 U378 ( .A(n26), .B(n73), .C(n269), .D(n267), .Y(N656) );
  XNOR2XL U379 ( .A(n132), .B(clk_count1[2]), .Y(n269) );
  NOR2X1 U380 ( .A(n90), .B(fsmdet[1]), .Y(n352) );
  NAND3X1 U381 ( .A(nedetect), .B(n99), .C(n291), .Y(n293) );
  OAI211X1 U382 ( .C(n289), .D(n290), .A(n121), .B(n291), .Y(n285) );
  AOI211X1 U383 ( .C(i2ccon_o[5]), .D(n296), .A(i2ccon_o[4]), .B(i2ccon_o[3]), 
        .Y(n289) );
  EORX1 U384 ( .A(n206), .B(n292), .C(n293), .D(n13), .Y(n290) );
  OAI211X1 U385 ( .C(fsmsta[0]), .D(n112), .A(n441), .B(n294), .Y(n292) );
  NAND4X1 U386 ( .A(fsmsta[2]), .B(n160), .C(fsmsta[1]), .D(n442), .Y(n377) );
  INVX1 U387 ( .A(sdao), .Y(n446) );
  OAI31XL U388 ( .A(n450), .B(ack), .C(n166), .D(n76), .Y(n413) );
  INVX1 U389 ( .A(n376), .Y(n76) );
  OAI21X1 U390 ( .B(n183), .C(n184), .A(n185), .Y(n498) );
  NAND42X1 U391 ( .C(n186), .D(n47), .A(nedetect), .B(n23), .Y(n185) );
  GEN2XL U392 ( .D(n84), .E(n72), .C(n231), .B(n232), .A(n233), .Y(N749) );
  OAI211X1 U393 ( .C(n443), .D(n437), .A(si), .B(n234), .Y(n232) );
  AOI211X1 U394 ( .C(n235), .D(n444), .A(sclint), .B(n236), .Y(n234) );
  OAI21X1 U395 ( .B(fsmsta[2]), .C(n159), .A(fsmsta[3]), .Y(n235) );
  OAI21X1 U396 ( .B(rst_delay), .C(n277), .A(n31), .Y(N653) );
  NOR4XL U397 ( .A(n129), .B(n130), .C(n276), .D(n448), .Y(n277) );
  AOI211X1 U398 ( .C(n81), .D(n155), .A(n156), .B(n157), .Y(n501) );
  OAI211X1 U399 ( .C(n158), .D(n40), .A(n101), .B(n31), .Y(n156) );
  NAND4X1 U400 ( .A(nedetect), .B(n149), .C(i2ccon_o[2]), .D(n163), .Y(n155)
         );
  AOI211X1 U401 ( .C(n159), .D(n160), .A(n161), .B(n162), .Y(n158) );
  NAND3X1 U402 ( .A(n101), .B(n138), .C(n278), .Y(n276) );
  AOI21X1 U403 ( .B(n279), .C(n85), .A(n280), .Y(n278) );
  AOI21X1 U404 ( .B(n83), .C(n84), .A(fsmsync[1]), .Y(n280) );
  OAI22X1 U405 ( .A(n115), .B(n67), .C(n445), .D(n123), .Y(n279) );
  AOI21X1 U406 ( .B(fsmsta[3]), .C(fsmsta[1]), .A(n444), .Y(n294) );
  NAND3X1 U407 ( .A(n106), .B(n104), .C(fsmmod[2]), .Y(n123) );
  OAI2B11X1 U408 ( .D(test_so2), .C(sclint), .A(n43), .B(n25), .Y(N332) );
  INVX1 U409 ( .A(adrcomp), .Y(n81) );
  OAI211X1 U410 ( .C(n355), .D(n77), .A(n25), .B(n356), .Y(N1027) );
  NOR3XL U411 ( .A(n358), .B(n359), .C(n360), .Y(n355) );
  AOI22X1 U412 ( .A(n357), .B(ack), .C(n86), .D(n157), .Y(n356) );
  ENOX1 U413 ( .A(n361), .B(n98), .C(n95), .D(n362), .Y(n360) );
  NAND2X1 U414 ( .A(n111), .B(fsmsta[3]), .Y(n302) );
  INVX1 U415 ( .A(clk_count1[1]), .Y(n69) );
  OAI21AX1 U416 ( .B(framesync[0]), .C(n37), .A(n285), .Y(N492) );
  NAND2X1 U417 ( .A(framesync[2]), .B(n100), .Y(n283) );
  INVX1 U418 ( .A(clk_count1[0]), .Y(n74) );
  NAND4X1 U419 ( .A(n173), .B(n174), .C(n175), .D(n176), .Y(n168) );
  XNOR2XL U420 ( .A(i2cdat_o[6]), .B(i2cadr_o[7]), .Y(n173) );
  XNOR2XL U421 ( .A(i2cdat_o[5]), .B(i2cadr_o[6]), .Y(n174) );
  XNOR2XL U422 ( .A(i2cdat_o[3]), .B(i2cadr_o[4]), .Y(n175) );
  INVX1 U423 ( .A(i2ccon_o[0]), .Y(n449) );
  INVX1 U424 ( .A(adrcompen), .Y(n79) );
  NAND2X1 U425 ( .A(n134), .B(n125), .Y(n504) );
  XNOR2XL U426 ( .A(clkint), .B(clk_count2_ov), .Y(n134) );
  NOR2X1 U427 ( .A(clk_count1[0]), .B(n267), .Y(N654) );
  NOR2X1 U428 ( .A(n266), .B(n267), .Y(N657) );
  XNOR2XL U429 ( .A(clk_count1[3]), .B(n268), .Y(n266) );
  NOR21XL U430 ( .B(clk_count1[2]), .A(n68), .Y(n268) );
  NOR2X1 U431 ( .A(n264), .B(n260), .Y(N688) );
  XNOR2XL U432 ( .A(clk_count2[3]), .B(n263), .Y(n264) );
  NOR2X1 U433 ( .A(n259), .B(n260), .Y(N690) );
  AOI222XL U434 ( .A(n261), .B(n448), .C(i2ccon_o[7]), .D(n262), .E(
        clk_count2[3]), .F(n263), .Y(n259) );
  OAI21AX1 U435 ( .B(n449), .C(n56), .A(i2ccon_o[1]), .Y(n262) );
  AOI31X1 U436 ( .A(n55), .B(n48), .C(n54), .D(wait_for_setup_r), .Y(n183) );
  GEN2XL U437 ( .D(n297), .E(n58), .C(N469), .B(indelay[2]), .A(n298), .Y(N471) );
  NOR4XL U438 ( .A(indelay[2]), .B(n58), .C(n70), .D(n59), .Y(n298) );
  GEN2XL U439 ( .D(fsmsta[1]), .E(n442), .C(n295), .B(n437), .A(n38), .Y(N407)
         );
  INVX1 U440 ( .A(n300), .Y(n38) );
  AO33X1 U441 ( .A(clk_count1_ov), .B(n25), .C(rst_delay), .D(n124), .E(n45), 
        .F(n125), .Y(n505) );
  INVX1 U442 ( .A(rst_delay), .Y(n45) );
  OAI21X1 U443 ( .B(i2ccon_o[7]), .C(n126), .A(n127), .Y(n124) );
  AOI33X1 U444 ( .A(i2ccon_o[7]), .B(i2ccon_o[1]), .C(n128), .D(n129), .E(n64), 
        .F(clk_count1[1]), .Y(n127) );
  NAND21X1 U445 ( .B(clk_count1[3]), .A(n272), .Y(n131) );
  NOR21XL U446 ( .B(bclkcnt[1]), .A(n14), .Y(n130) );
  XNOR2XL U447 ( .A(bclksel), .B(bclkcnt[0]), .Y(n14) );
  NOR3XL U448 ( .A(fsmsync[2]), .B(n26), .C(n71), .Y(n297) );
  NOR3XL U449 ( .A(n84), .B(fsmsync[1]), .C(n83), .Y(n243) );
  NOR3XL U450 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(fsmmod[0]), .Y(n153) );
  NAND21X1 U451 ( .B(clk_count1_ov), .A(n125), .Y(N689) );
  NAND2X1 U452 ( .A(clkint_ff), .B(n75), .Y(n122) );
  OAI211X1 U453 ( .C(n109), .D(n344), .A(n138), .B(n452), .Y(n333) );
  NAND2X1 U454 ( .A(n97), .B(pedetect), .Y(n344) );
  NOR2X1 U455 ( .A(n75), .B(clkint_ff), .Y(n253) );
  AOI21X1 U456 ( .B(i2ccon_o[0]), .C(i2ccon_o[1]), .A(n448), .Y(n129) );
  NAND3X1 U457 ( .A(indelay[1]), .B(n59), .C(indelay[2]), .Y(n245) );
  NAND3X1 U458 ( .A(n62), .B(n453), .C(i2ccon_o[5]), .Y(n339) );
  AND3X1 U459 ( .A(n130), .B(n131), .C(i2ccon_o[0]), .Y(n128) );
  INVX1 U460 ( .A(sclint), .Y(n85) );
  INVX1 U461 ( .A(fsmsync[0]), .Y(n84) );
  INVX1 U462 ( .A(fsmsync[1]), .Y(n72) );
  INVX1 U463 ( .A(sdaint), .Y(n94) );
  NOR4XL U464 ( .A(n63), .B(n72), .C(fsmsync[0]), .D(fsmsync[2]), .Y(n242) );
  INVX1 U465 ( .A(pedetect), .Y(n80) );
  INVX1 U466 ( .A(ack), .Y(n96) );
  OAI221X1 U467 ( .A(fsmsta[1]), .B(n434), .C(fsmsta[0]), .D(n308), .E(n300), 
        .Y(N406) );
  INVX1 U468 ( .A(fsmsync[2]), .Y(n83) );
  OAI21X1 U469 ( .B(n37), .C(n288), .A(n121), .Y(N493) );
  OAI21X1 U470 ( .B(framesync[1]), .C(framesync[0]), .A(n287), .Y(n288) );
  OAI21X1 U471 ( .B(n286), .C(n37), .A(n121), .Y(N494) );
  XNOR2XL U472 ( .A(n100), .B(framesync[2]), .Y(n286) );
  OAI211X1 U473 ( .C(n9), .D(n303), .A(n300), .B(n304), .Y(N409) );
  AOI32X1 U474 ( .A(n9), .B(n7), .C(n305), .D(n306), .E(n303), .Y(n304) );
  AOI211X1 U475 ( .C(n49), .D(n122), .A(n230), .B(n115), .Y(n490) );
  INVX1 U476 ( .A(starto_en), .Y(n49) );
  OR2X1 U477 ( .A(n184), .B(n67), .Y(n230) );
  INVX1 U478 ( .A(clkint), .Y(n75) );
  AOI21X1 U479 ( .B(sclint), .C(n62), .A(n123), .Y(n335) );
  NOR3XL U480 ( .A(n105), .B(sdaint), .C(i2ccon_o[3]), .Y(n337) );
  INVX1 U481 ( .A(i2ccon_o[4]), .Y(n453) );
  AOI21X1 U482 ( .B(n254), .C(n255), .A(n238), .Y(N746) );
  AOI211X1 U483 ( .C(n244), .D(n94), .A(n256), .B(n257), .Y(n255) );
  AOI222XL U484 ( .A(n243), .B(si), .C(n240), .D(n453), .E(n242), .F(n41), .Y(
        n254) );
  NOR4XL U485 ( .A(sclint), .B(fsmsync[2]), .C(fsmsync[1]), .D(fsmsync[0]), 
        .Y(n256) );
  AOI21X1 U486 ( .B(n190), .C(n191), .A(n192), .Y(n496) );
  OAI211X1 U487 ( .C(n60), .D(n193), .A(n121), .B(adrcompen), .Y(n191) );
  NAND2X1 U488 ( .A(n194), .B(n23), .Y(n190) );
  AOI21X1 U489 ( .B(n353), .C(n354), .A(n184), .Y(N1063) );
  NAND2X1 U490 ( .A(n351), .B(n94), .Y(n354) );
  AOI32X1 U491 ( .A(n91), .B(n90), .C(sdaint), .D(n352), .E(n93), .Y(n353) );
  INVX1 U492 ( .A(n351), .Y(n91) );
  NAND3X1 U493 ( .A(n25), .B(n85), .C(test_so2), .Y(n312) );
  OAI21X1 U494 ( .B(n116), .C(n94), .A(n117), .Y(n507) );
  NOR3XL U495 ( .A(sdai_ff_reg0_0_), .B(test_so1), .C(sdai_ff_reg0_1_), .Y(
        n116) );
  AOI31X1 U496 ( .A(sdai_ff_reg0_1_), .B(sdai_ff_reg0_0_), .C(test_so1), .D(
        n29), .Y(n117) );
  AOI31X1 U497 ( .A(n246), .B(n247), .C(n248), .D(n238), .Y(N747) );
  OAI211X1 U498 ( .C(n40), .D(n63), .A(n84), .B(fsmsync[1]), .Y(n247) );
  AOI22X1 U499 ( .A(n243), .B(n40), .C(n231), .D(n245), .Y(n248) );
  AOI31X1 U500 ( .A(n72), .B(n83), .C(n249), .D(n244), .Y(n246) );
  AOI31X1 U501 ( .A(n330), .B(n331), .C(n332), .D(n333), .Y(N1126) );
  NAND3X1 U502 ( .A(n336), .B(i2ccon_o[4]), .C(n258), .Y(n331) );
  AOI221XL U503 ( .A(n251), .B(n60), .C(n115), .D(n334), .E(n335), .Y(n332) );
  AOI33X1 U504 ( .A(starto_en), .B(n61), .C(n337), .D(sclint), .E(n338), .F(
        n154), .Y(n330) );
  AOI31X1 U505 ( .A(n102), .B(n103), .C(n340), .D(n333), .Y(N1125) );
  AOI22X1 U506 ( .A(n336), .B(n341), .C(n342), .D(nedetect), .Y(n340) );
  NAND2X1 U507 ( .A(n258), .B(i2ccon_o[4]), .Y(n341) );
  INVX1 U508 ( .A(indelay[0]), .Y(n59) );
  INVX1 U509 ( .A(i2ccon_o[7]), .Y(n448) );
  INVX1 U510 ( .A(scli_ff_reg0[0]), .Y(n55) );
  INVX1 U511 ( .A(scli_ff_reg0[1]), .Y(n54) );
  INVX1 U512 ( .A(clk_count2[0]), .Y(n56) );
  INVX1 U513 ( .A(i2cdat_o[1]), .Y(n454) );
  OAI21BBX1 U514 ( .A(n56), .B(n125), .C(n265), .Y(N685) );
  NAND4X1 U515 ( .A(fsmsync[2]), .B(n84), .C(n72), .D(n23), .Y(n265) );
  NOR2X1 U516 ( .A(setup_counter_r[1]), .B(setup_counter_r[0]), .Y(n313) );
  NOR2X1 U517 ( .A(n70), .B(indelay[0]), .Y(N469) );
  INVX1 U518 ( .A(i2cdat_o[0]), .Y(n451) );
  NAND2X1 U519 ( .A(n24), .B(n189), .Y(n182) );
  NAND4X1 U520 ( .A(scli_ff_reg0[2]), .B(scli_ff_reg0[1]), .C(scli_ff_reg0[0]), 
        .D(n183), .Y(n189) );
  INVX1 U521 ( .A(i2cdat_o[2]), .Y(n447) );
  NAND2X1 U522 ( .A(n84), .B(n250), .Y(n249) );
  OAI211X1 U523 ( .C(n251), .D(n252), .A(sclint), .B(n253), .Y(n250) );
  AOI22X1 U524 ( .A(fsmmod[2]), .B(n106), .C(fsmmod[1]), .D(fsmmod[0]), .Y(
        n252) );
  INVX1 U525 ( .A(scli_ff_reg0[2]), .Y(n48) );
  NOR2X1 U526 ( .A(i2ccon_o[2]), .B(sdaint), .Y(n417) );
  NAND2X1 U527 ( .A(n300), .B(n307), .Y(N408) );
  OAI211X1 U528 ( .C(fsmsta[2]), .D(n159), .A(n437), .B(n303), .Y(n307) );
  NOR2X1 U529 ( .A(n348), .B(n184), .Y(N1065) );
  AOI221XL U530 ( .A(fsmdet[1]), .B(sdaint), .C(fsmdet[2]), .D(n92), .E(n194), 
        .Y(n348) );
  NOR2X1 U531 ( .A(n349), .B(n184), .Y(N1064) );
  AOI221XL U532 ( .A(fsmdet[2]), .B(fsmdet[0]), .C(n350), .D(n94), .E(n351), 
        .Y(n349) );
  OAI21AX1 U533 ( .B(fsmdet[2]), .C(fsmdet[0]), .A(n352), .Y(n350) );
  NOR2X1 U534 ( .A(n237), .B(n238), .Y(N748) );
  AOI221XL U535 ( .A(n239), .B(n85), .C(i2ccon_o[3]), .D(n240), .E(n241), .Y(
        n237) );
  OAI22X1 U539 ( .A(fsmsync[0]), .B(n83), .C(n245), .D(n71), .Y(n239) );
  GEN2XL U540 ( .D(n206), .E(n242), .C(n243), .B(i2ccon_o[4]), .A(n244), .Y(
        n241) );
  INVX1 U541 ( .A(busfree), .Y(n67) );
  INVX1 U542 ( .A(i2cadr_o[0]), .Y(n450) );
  INVX1 U543 ( .A(n114), .Y(n50) );
  OAI211X1 U544 ( .C(sclscl), .D(pedetect), .A(n115), .B(n31), .Y(n114) );
  INVX1 U545 ( .A(bsd7_tmp), .Y(n66) );
  NAND21X1 U546 ( .B(scli_ff), .A(n23), .Y(N412) );
  NAND21X1 U547 ( .B(sdai_ff), .A(n23), .Y(N431) );
  NAND21X1 U548 ( .B(sdai_ff_reg0_0_), .A(n23), .Y(N432) );
  NAND21X1 U549 ( .B(sdai_ff_reg0_1_), .A(n23), .Y(N433) );
  NOR3XL U550 ( .A(n281), .B(n27), .C(n130), .Y(N511) );
  XNOR2XL U551 ( .A(bclkcnt[1]), .B(bclkcnt[0]), .Y(n281) );
  INVX1 U552 ( .A(nedetect), .Y(n60) );
  NOR3XL U553 ( .A(n130), .B(n27), .C(bclkcnt[0]), .Y(N510) );
  INVX1 U554 ( .A(fsmdet[2]), .Y(n93) );
  NAND2X1 U555 ( .A(sclscl), .B(pedetect), .Y(n334) );
  INVX1 U556 ( .A(clk_count2[1]), .Y(n53) );
  INVX1 U557 ( .A(clk_count2[2]), .Y(n57) );
  INVX1 U558 ( .A(setup_counter_r[2]), .Y(n44) );
  INVX1 U559 ( .A(indelay[1]), .Y(n58) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module extint_a0 ( clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, 
        int2ff, iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, 
        int6ff, iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, 
        ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7, 
        iex8, iex9, iex10, iex11, iex12, sfraddr, sfrdatai, sfrwe, test_si, 
        test_se );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, int2ff,
         iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, int6ff,
         iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, sfrwe,
         test_si, test_se;
  output ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12;
  wire   int0_ff1, int0_fall, int0_clr, N23, int1_ff1, int1_fall, int1_clr,
         N51, int2_ff1, iex2_set, N71, int3_ff1, iex3_set, N90, iex4_set,
         int4_ff1, iex5_set, int5_ff1, iex6_set, int6_ff1, iex7_set, int7_ff1,
         iex8_set, int8_ff1, iex9_set, int9_ff1, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n77, n78, n79, n80,
         n81, n82, n83, n84;

  SDFFQX1 int4_ff1_reg ( .D(n19), .SIN(int3_ff1), .SMC(test_se), .C(clkper), 
        .Q(int4_ff1) );
  SDFFQX1 int5_ff1_reg ( .D(n13), .SIN(int4_ff1), .SMC(test_se), .C(clkper), 
        .Q(int5_ff1) );
  SDFFQX1 int6_ff1_reg ( .D(n11), .SIN(int5_ff1), .SMC(test_se), .C(clkper), 
        .Q(int6_ff1) );
  SDFFQX1 int7_ff1_reg ( .D(n12), .SIN(int6_ff1), .SMC(test_se), .C(clkper), 
        .Q(int7_ff1) );
  SDFFQX1 int8_ff1_reg ( .D(n84), .SIN(int7_ff1), .SMC(test_se), .C(clkper), 
        .Q(int8_ff1) );
  SDFFQX1 int9_ff1_reg ( .D(n10), .SIN(int8_ff1), .SMC(test_se), .C(clkper), 
        .Q(int9_ff1) );
  SDFFQX1 iex4_set_reg ( .D(n105), .SIN(iex4), .SMC(test_se), .C(clkper), .Q(
        iex4_set) );
  SDFFQX1 iex5_set_reg ( .D(n103), .SIN(iex5), .SMC(test_se), .C(clkper), .Q(
        iex5_set) );
  SDFFQX1 iex6_set_reg ( .D(n101), .SIN(iex6), .SMC(test_se), .C(clkper), .Q(
        iex6_set) );
  SDFFQX1 iex7_set_reg ( .D(n99), .SIN(iex7), .SMC(test_se), .C(clkper), .Q(
        iex7_set) );
  SDFFQX1 iex8_set_reg ( .D(n97), .SIN(iex8), .SMC(test_se), .C(clkper), .Q(
        iex8_set) );
  SDFFQX1 iex9_set_reg ( .D(n95), .SIN(iex9), .SMC(test_se), .C(clkper), .Q(
        iex9_set) );
  SDFFQX1 int0_ff1_reg ( .D(N23), .SIN(int0_fall), .SMC(test_se), .C(clkper), 
        .Q(int0_ff1) );
  SDFFQX1 iex2_set_reg ( .D(n110), .SIN(iex2), .SMC(test_se), .C(clkper), .Q(
        iex2_set) );
  SDFFQX1 iex3_set_reg ( .D(n107), .SIN(iex3), .SMC(test_se), .C(clkper), .Q(
        iex3_set) );
  SDFFQX1 int0_clr_reg ( .D(n118), .SIN(iex9_set), .SMC(test_se), .C(clkper), 
        .Q(int0_clr) );
  SDFFQX1 int1_clr_reg ( .D(n114), .SIN(int0_ff1), .SMC(test_se), .C(clkper), 
        .Q(int1_clr) );
  SDFFQX1 int2_ff1_reg ( .D(N71), .SIN(int1_ff1), .SMC(test_se), .C(clkper), 
        .Q(int2_ff1) );
  SDFFQX1 int3_ff1_reg ( .D(N90), .SIN(int2_ff1), .SMC(test_se), .C(clkper), 
        .Q(int3_ff1) );
  SDFFQX1 int1_ff1_reg ( .D(N51), .SIN(int1_fall), .SMC(test_se), .C(clkper), 
        .Q(int1_ff1) );
  SDFFQX1 int0_fall_reg ( .D(n116), .SIN(int0_clr), .SMC(test_se), .C(clkper), 
        .Q(int0_fall) );
  SDFFQX1 int1_fall_reg ( .D(n112), .SIN(int1_clr), .SMC(test_se), .C(clkper), 
        .Q(int1_fall) );
  SDFFQX1 iex9_s_reg ( .D(n94), .SIN(iex8_set), .SMC(test_se), .C(clkper), .Q(
        iex9) );
  SDFFQX1 iex8_s_reg ( .D(n96), .SIN(iex7_set), .SMC(test_se), .C(clkper), .Q(
        iex8) );
  SDFFQX1 i3fr_s_reg ( .D(n108), .SIN(i2fr), .SMC(test_se), .C(clkper), .Q(
        i3fr) );
  SDFFQX1 ie1_s_reg ( .D(n111), .SIN(ie0), .SMC(test_se), .C(clkper), .Q(ie1)
         );
  SDFFQX1 iex2_s_reg ( .D(n109), .SIN(ie1), .SMC(test_se), .C(clkper), .Q(iex2) );
  SDFFQX1 ie0_s_reg ( .D(n115), .SIN(i3fr), .SMC(test_se), .C(clkper), .Q(ie0)
         );
  SDFFQX1 it0_s_reg ( .D(n117), .SIN(int9_ff1), .SMC(test_se), .C(clkper), .Q(
        it0) );
  SDFFQX1 iex3_s_reg ( .D(n106), .SIN(iex2_set), .SMC(test_se), .C(clkper), 
        .Q(iex3) );
  SDFFQX1 iex4_s_reg ( .D(n104), .SIN(iex3_set), .SMC(test_se), .C(clkper), 
        .Q(iex4) );
  SDFFQX1 iex6_s_reg ( .D(n100), .SIN(iex5_set), .SMC(test_se), .C(clkper), 
        .Q(iex6) );
  SDFFQX1 i2fr_s_reg ( .D(n14), .SIN(test_si), .SMC(test_se), .C(clkper), .Q(
        i2fr) );
  SDFFQX1 iex7_s_reg ( .D(n98), .SIN(iex6_set), .SMC(test_se), .C(clkper), .Q(
        iex7) );
  SDFFQX1 iex5_s_reg ( .D(n102), .SIN(iex4_set), .SMC(test_se), .C(clkper), 
        .Q(iex5) );
  SDFFQX1 it1_s_reg ( .D(n113), .SIN(it0), .SMC(test_se), .C(clkper), .Q(it1)
         );
  INVX1 U3 ( .A(1'b1), .Y(iex12) );
  INVX1 U5 ( .A(1'b1), .Y(iex11) );
  INVX1 U7 ( .A(1'b1), .Y(iex10) );
  AND2X1 U9 ( .A(sfraddr[6]), .B(n63), .Y(n68) );
  INVX1 U10 ( .A(n34), .Y(n15) );
  INVX1 U11 ( .A(n52), .Y(n16) );
  NAND2X1 U12 ( .A(n75), .B(n9), .Y(n41) );
  NOR2X1 U13 ( .A(n75), .B(n7), .Y(n43) );
  INVX1 U14 ( .A(n46), .Y(n17) );
  INVX1 U15 ( .A(n8), .Y(n7) );
  AOI21X1 U16 ( .B(n68), .C(sfraddr[3]), .A(rst), .Y(n34) );
  NOR42XL U17 ( .C(sfrwe), .D(n76), .A(sfraddr[0]), .B(sfraddr[1]), .Y(n63) );
  NOR3XL U18 ( .A(sfraddr[2]), .B(sfraddr[5]), .C(sfraddr[4]), .Y(n76) );
  NOR32XL U19 ( .B(n63), .C(sfraddr[3]), .A(sfraddr[6]), .Y(n52) );
  NAND2X1 U20 ( .A(n49), .B(n50), .Y(n46) );
  AND4XL U21 ( .A(sfraddr[1]), .B(sfraddr[2]), .C(sfraddr[4]), .D(sfraddr[5]), 
        .Y(n49) );
  NOR43XL U22 ( .B(sfraddr[3]), .C(sfrwe), .D(sfraddr[0]), .A(sfraddr[6]), .Y(
        n50) );
  NAND21X1 U23 ( .B(sfraddr[3]), .A(n68), .Y(n75) );
  INVX1 U24 ( .A(n53), .Y(n18) );
  INVX1 U25 ( .A(n37), .Y(n12) );
  INVX1 U26 ( .A(rst), .Y(n8) );
  INVX1 U27 ( .A(rst), .Y(n9) );
  INVX1 U28 ( .A(n40), .Y(n84) );
  INVX1 U29 ( .A(n39), .Y(n13) );
  INVX1 U30 ( .A(n35), .Y(n10) );
  INVX1 U31 ( .A(n38), .Y(n19) );
  NOR2X1 U32 ( .A(n7), .B(newinstr), .Y(n53) );
  OAI22X1 U33 ( .A(n7), .B(n77), .C(n18), .D(n29), .Y(n114) );
  OAI22X1 U34 ( .A(rst), .B(n32), .C(n18), .D(n28), .Y(n118) );
  NAND2X1 U35 ( .A(int7ff), .B(n9), .Y(n37) );
  OR2X1 U36 ( .A(int2ff), .B(rst), .Y(N71) );
  INVX1 U37 ( .A(int0ack), .Y(n32) );
  INVX1 U38 ( .A(int1ack), .Y(n77) );
  INVX1 U39 ( .A(iex3ack), .Y(n79) );
  INVX1 U40 ( .A(iex2ack), .Y(n78) );
  OR2X1 U41 ( .A(int3ff), .B(rst), .Y(N90) );
  INVX1 U42 ( .A(n36), .Y(n11) );
  NAND2X1 U43 ( .A(int8ff), .B(n9), .Y(n40) );
  NOR2X1 U44 ( .A(n7), .B(n83), .Y(N23) );
  NOR2X1 U45 ( .A(n7), .B(n82), .Y(N51) );
  NAND2X1 U46 ( .A(int5ff), .B(n9), .Y(n39) );
  OAI32X1 U47 ( .A(n21), .B(iex5ack), .C(n18), .D(int5_ff1), .E(n39), .Y(n103)
         );
  INVX1 U48 ( .A(iex5_set), .Y(n21) );
  NAND2X1 U49 ( .A(int9ff), .B(n8), .Y(n35) );
  OAI32X1 U50 ( .A(n25), .B(iex9ack), .C(n18), .D(int9_ff1), .E(n35), .Y(n95)
         );
  INVX1 U51 ( .A(iex9_set), .Y(n25) );
  OAI21BBX1 U52 ( .A(n34), .B(i3fr), .C(n67), .Y(n108) );
  NAND3X1 U53 ( .A(n15), .B(n9), .C(sfrdatai[6]), .Y(n67) );
  INVX1 U54 ( .A(n33), .Y(n14) );
  AOI32X1 U55 ( .A(sfrdatai[5]), .B(n9), .C(n15), .D(n34), .E(i2fr), .Y(n33)
         );
  NAND2X1 U56 ( .A(int4ff), .B(n8), .Y(n38) );
  OAI32X1 U57 ( .A(n20), .B(iex4ack), .C(n18), .D(int4_ff1), .E(n38), .Y(n105)
         );
  INVX1 U58 ( .A(iex4_set), .Y(n20) );
  NOR2X1 U59 ( .A(n7), .B(n51), .Y(n117) );
  AOI22X1 U60 ( .A(n52), .B(sfrdatai[0]), .C(it0), .D(n16), .Y(n51) );
  NOR2X1 U61 ( .A(n7), .B(n58), .Y(n113) );
  AOI22X1 U62 ( .A(sfrdatai[2]), .B(n52), .C(it1), .D(n16), .Y(n58) );
  NOR2X1 U63 ( .A(n7), .B(n59), .Y(n111) );
  EORX1 U64 ( .A(sfrdatai[3]), .B(n52), .C(n60), .D(n52), .Y(n59) );
  AOI32X1 U65 ( .A(n29), .B(n77), .C(n61), .D(n82), .E(n30), .Y(n60) );
  ENOX1 U66 ( .A(n62), .B(n30), .C(n82), .D(int1_ff1), .Y(n61) );
  AND2X1 U67 ( .A(n54), .B(n9), .Y(n115) );
  ENOX1 U68 ( .A(n52), .B(n55), .C(sfrdatai[1]), .D(n52), .Y(n54) );
  AOI32X1 U69 ( .A(n28), .B(n32), .C(n56), .D(n83), .E(n31), .Y(n55) );
  ENOX1 U70 ( .A(n57), .B(n31), .C(n83), .D(int0_ff1), .Y(n56) );
  AOI21X1 U71 ( .B(n47), .C(n48), .A(rst), .Y(n94) );
  NAND2X1 U72 ( .A(sfrdatai[1]), .B(n17), .Y(n47) );
  OAI211X1 U73 ( .C(iex9), .D(iex9_set), .A(n46), .B(n80), .Y(n48) );
  INVX1 U74 ( .A(iex9ack), .Y(n80) );
  AOI21X1 U75 ( .B(n44), .C(n45), .A(rst), .Y(n96) );
  NAND2X1 U76 ( .A(n17), .B(sfrdatai[0]), .Y(n44) );
  OAI211X1 U77 ( .C(iex8), .D(iex8_set), .A(n46), .B(n81), .Y(n45) );
  INVX1 U78 ( .A(iex8ack), .Y(n81) );
  ENOX1 U79 ( .A(n41), .B(n42), .C(n43), .D(sfrdatai[0]), .Y(n98) );
  OAI21AX1 U80 ( .B(iex7), .C(iex7_set), .A(iex7ack), .Y(n42) );
  ENOX1 U81 ( .A(n41), .B(n72), .C(n43), .D(sfrdatai[3]), .Y(n104) );
  OAI21AX1 U82 ( .B(iex4), .C(iex4_set), .A(iex4ack), .Y(n72) );
  ENOX1 U83 ( .A(n41), .B(n74), .C(sfrdatai[5]), .D(n43), .Y(n100) );
  OAI21AX1 U84 ( .B(iex6), .C(iex6_set), .A(iex6ack), .Y(n74) );
  ENOX1 U85 ( .A(n41), .B(n73), .C(sfrdatai[4]), .D(n43), .Y(n102) );
  OAI21AX1 U86 ( .B(iex5), .C(iex5_set), .A(iex5ack), .Y(n73) );
  ENOX1 U87 ( .A(n41), .B(n71), .C(n43), .D(sfrdatai[2]), .Y(n106) );
  OAI21X1 U88 ( .B(iex3), .C(iex3_set), .A(n79), .Y(n71) );
  ENOX1 U89 ( .A(n41), .B(n66), .C(n43), .D(sfrdatai[1]), .Y(n109) );
  OAI21X1 U90 ( .B(iex2), .C(iex2_set), .A(n78), .Y(n66) );
  AO33X1 U91 ( .A(int1_ff1), .B(n9), .C(n82), .D(int1_fall), .E(n77), .F(n53), 
        .Y(n112) );
  AO33X1 U92 ( .A(int0_ff1), .B(n9), .C(n83), .D(int0_fall), .E(n32), .F(n53), 
        .Y(n116) );
  OAI32X1 U93 ( .A(n24), .B(iex8ack), .C(n18), .D(int8_ff1), .E(n40), .Y(n97)
         );
  INVX1 U94 ( .A(iex8_set), .Y(n24) );
  OAI32X1 U95 ( .A(n23), .B(iex7ack), .C(n18), .D(int7_ff1), .E(n37), .Y(n99)
         );
  INVX1 U96 ( .A(iex7_set), .Y(n23) );
  OAI32X1 U97 ( .A(n22), .B(iex6ack), .C(n18), .D(int6_ff1), .E(n36), .Y(n101)
         );
  INVX1 U98 ( .A(iex6_set), .Y(n22) );
  OAI31XL U99 ( .A(n27), .B(i3fr), .C(N90), .D(n69), .Y(n107) );
  INVX1 U100 ( .A(int3_ff1), .Y(n27) );
  AOI33X1 U101 ( .A(int3ff), .B(i3fr), .C(n70), .D(n53), .E(n79), .F(iex3_set), 
        .Y(n69) );
  NOR2X1 U102 ( .A(n7), .B(int3_ff1), .Y(n70) );
  OAI31XL U103 ( .A(n26), .B(i2fr), .C(N71), .D(n64), .Y(n110) );
  INVX1 U104 ( .A(int2_ff1), .Y(n26) );
  AOI33X1 U105 ( .A(int2ff), .B(i2fr), .C(n65), .D(n53), .E(n78), .F(iex2_set), 
        .Y(n64) );
  NOR2X1 U106 ( .A(n7), .B(int2_ff1), .Y(n65) );
  NAND2X1 U107 ( .A(int6ff), .B(n9), .Y(n36) );
  INVX1 U111 ( .A(int1ff), .Y(n82) );
  INVX1 U112 ( .A(int0ff), .Y(n83) );
  NOR2X1 U113 ( .A(ie1), .B(int1_fall), .Y(n62) );
  NOR2X1 U114 ( .A(ie0), .B(int0_fall), .Y(n57) );
  INVX1 U115 ( .A(it1), .Y(n30) );
  INVX1 U116 ( .A(it0), .Y(n31) );
  INVX1 U117 ( .A(int1_clr), .Y(n29) );
  INVX1 U118 ( .A(int0_clr), .Y(n28) );
endmodule


module isr_a0 ( clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, 
        t0ff, int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff, 
        int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b, 
        int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, int_vect_ab, irq, intvect, int_ack_03, int_ack_0b, 
        int_ack_13, int_ack_1b, int_ack_43, int_ack_4b, int_ack_53, int_ack_5b, 
        int_ack_63, int_ack_6b, int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, 
        int_ack_ab, is_reg, ip0, ip1, ien0, ien1, ien2, isr_tm, sfraddr, 
        sfrdatai, sfrwe, test_si, test_se );
  output [4:0] intvect;
  output [3:0] is_reg;
  output [5:0] ip0;
  output [5:0] ip1;
  output [7:0] ien0;
  output [5:0] ien1;
  output [5:0] ien2;
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, t0ff,
         int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff,
         int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b,
         int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b,
         int_vect_a3, int_vect_ab, sfrwe, test_si, test_se;
  output irq, int_ack_03, int_ack_0b, int_ack_13, int_ack_1b, int_ack_43,
         int_ack_4b, int_ack_53, int_ack_5b, int_ack_63, int_ack_6b,
         int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, int_ack_ab, isr_tm;
  wire   N38, N39, N40, N41, N42, N43, N44, N45, N49, N50, N51, N52, N53, N54,
         N55, N58, N59, N60, N61, N62, N63, N64, N67, N68, N69, N70, N71, N72,
         N73, N76, N77, N78, N79, N80, N81, N82, irq_r, N200, N207, N208, N209,
         N210, N211, N212, net12106, net12112, net12117, net12122, net12127,
         net12132, n196, n197, n198, n199, n200, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n201, n202, n203, n204, n205, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n206, n207, n208;

  SNPS_CLOCK_GATE_HIGH_isr_a0_0 clk_gate_ien0_reg_reg ( .CLK(clkper), .EN(N38), 
        .ENCLK(net12106), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_5 clk_gate_ien1_reg_reg ( .CLK(clkper), .EN(N49), 
        .ENCLK(net12112), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_4 clk_gate_ien2_reg_reg ( .CLK(clkper), .EN(N58), 
        .ENCLK(net12117), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_3 clk_gate_ip0_reg_reg ( .CLK(clkper), .EN(N67), 
        .ENCLK(net12122), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_2 clk_gate_ip1_reg_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12127), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_1 clk_gate_intvect_reg_reg ( .CLK(clkper), .EN(
        N207), .ENCLK(net12132), .TE(test_se) );
  SDFFQX1 intvect_reg_reg_0_ ( .D(N208), .SIN(ien2[5]), .SMC(test_se), .C(
        net12132), .Q(intvect[0]) );
  SDFFQX1 intvect_reg_reg_1_ ( .D(N209), .SIN(intvect[0]), .SMC(test_se), .C(
        net12132), .Q(intvect[1]) );
  SDFFQX1 intvect_reg_reg_4_ ( .D(N212), .SIN(intvect[3]), .SMC(test_se), .C(
        net12132), .Q(intvect[4]) );
  SDFFQX1 intvect_reg_reg_3_ ( .D(N211), .SIN(intvect[2]), .SMC(test_se), .C(
        net12132), .Q(intvect[3]) );
  SDFFQX1 intvect_reg_reg_2_ ( .D(N210), .SIN(intvect[1]), .SMC(test_se), .C(
        net12132), .Q(intvect[2]) );
  SDFFQX1 is_reg_s_reg_0_ ( .D(n199), .SIN(irq_r), .SMC(test_se), .C(clkper), 
        .Q(is_reg[0]) );
  SDFFQX1 is_reg_s_reg_1_ ( .D(n196), .SIN(is_reg[0]), .SMC(test_se), .C(
        clkper), .Q(is_reg[1]) );
  SDFFQX1 is_reg_s_reg_2_ ( .D(n197), .SIN(is_reg[1]), .SMC(test_se), .C(
        clkper), .Q(is_reg[2]) );
  SDFFQX1 is_reg_s_reg_3_ ( .D(n198), .SIN(is_reg[2]), .SMC(test_se), .C(
        clkper), .Q(is_reg[3]) );
  SDFFQX1 irq_r_reg ( .D(N200), .SIN(ip1[5]), .SMC(test_se), .C(clkper), .Q(
        irq_r) );
  SDFFQX1 ien2_reg_reg_5_ ( .D(N64), .SIN(ien2[4]), .SMC(test_se), .C(net12117), .Q(ien2[5]) );
  SDFFQX1 ien0_reg_reg_1_ ( .D(N40), .SIN(ien0[0]), .SMC(test_se), .C(net12106), .Q(ien0[1]) );
  SDFFQX1 ien2_reg_reg_4_ ( .D(N63), .SIN(ien2[3]), .SMC(test_se), .C(net12117), .Q(ien2[4]) );
  SDFFQX1 ien2_reg_reg_1_ ( .D(N60), .SIN(ien2[0]), .SMC(test_se), .C(net12117), .Q(ien2[1]) );
  SDFFQX1 ip0_reg_reg_3_ ( .D(N71), .SIN(ip0[2]), .SMC(test_se), .C(net12122), 
        .Q(ip0[3]) );
  SDFFQX1 ien1_reg_reg_1_ ( .D(N51), .SIN(ien1[0]), .SMC(test_se), .C(net12112), .Q(ien1[1]) );
  SDFFQX1 ip0_reg_reg_1_ ( .D(N69), .SIN(ip0[0]), .SMC(test_se), .C(net12122), 
        .Q(ip0[1]) );
  SDFFQX1 ip0_reg_reg_2_ ( .D(N70), .SIN(ip0[1]), .SMC(test_se), .C(net12122), 
        .Q(ip0[2]) );
  SDFFQX1 ip1_reg_reg_1_ ( .D(N78), .SIN(ip1[0]), .SMC(test_se), .C(net12127), 
        .Q(ip1[1]) );
  SDFFQX1 ien2_reg_reg_0_ ( .D(N59), .SIN(ien1[5]), .SMC(test_se), .C(net12117), .Q(ien2[0]) );
  SDFFQX1 ien0_reg_reg_3_ ( .D(N42), .SIN(ien0[2]), .SMC(test_se), .C(net12106), .Q(ien0[3]) );
  SDFFQX1 ien1_reg_reg_0_ ( .D(N50), .SIN(ien0[7]), .SMC(test_se), .C(net12112), .Q(ien1[0]) );
  SDFFQX1 ien1_reg_reg_2_ ( .D(N52), .SIN(ien1[1]), .SMC(test_se), .C(net12112), .Q(ien1[2]) );
  SDFFQX1 ien1_reg_reg_3_ ( .D(N53), .SIN(ien1[2]), .SMC(test_se), .C(net12112), .Q(ien1[3]) );
  SDFFQX1 ien1_reg_reg_5_ ( .D(N55), .SIN(ien1[4]), .SMC(test_se), .C(net12112), .Q(ien1[5]) );
  SDFFQX1 ien0_reg_reg_4_ ( .D(N43), .SIN(ien0[3]), .SMC(test_se), .C(net12106), .Q(ien0[4]) );
  SDFFQX1 ien2_reg_reg_3_ ( .D(N62), .SIN(ien2[2]), .SMC(test_se), .C(net12117), .Q(ien2[3]) );
  SDFFQX1 ien0_reg_reg_5_ ( .D(N44), .SIN(ien0[4]), .SMC(test_se), .C(net12106), .Q(ien0[5]) );
  SDFFQX1 ien2_reg_reg_2_ ( .D(N61), .SIN(ien2[1]), .SMC(test_se), .C(net12117), .Q(ien2[2]) );
  SDFFQX1 ien1_reg_reg_4_ ( .D(N54), .SIN(ien1[3]), .SMC(test_se), .C(net12112), .Q(ien1[4]) );
  SDFFQX1 ien0_reg_reg_6_ ( .D(N45), .SIN(ien0[5]), .SMC(test_se), .C(net12106), .Q(ien0[7]) );
  SDFFQX1 ien0_reg_reg_2_ ( .D(N41), .SIN(ien0[1]), .SMC(test_se), .C(net12106), .Q(ien0[2]) );
  SDFFQX1 ien0_reg_reg_0_ ( .D(N39), .SIN(test_si), .SMC(test_se), .C(net12106), .Q(ien0[0]) );
  SDFFQX1 ip1_reg_reg_5_ ( .D(N82), .SIN(ip1[4]), .SMC(test_se), .C(net12127), 
        .Q(ip1[5]) );
  SDFFQX1 ip0_reg_reg_0_ ( .D(N68), .SIN(intvect[4]), .SMC(test_se), .C(
        net12122), .Q(ip0[0]) );
  SDFFQX1 ip1_reg_reg_4_ ( .D(N81), .SIN(ip1[3]), .SMC(test_se), .C(net12127), 
        .Q(ip1[4]) );
  SDFFQX1 ip1_reg_reg_0_ ( .D(N77), .SIN(ip0[5]), .SMC(test_se), .C(net12127), 
        .Q(ip1[0]) );
  SDFFQX1 ip1_reg_reg_3_ ( .D(N80), .SIN(ip1[2]), .SMC(test_se), .C(net12127), 
        .Q(ip1[3]) );
  SDFFQX1 ip1_reg_reg_2_ ( .D(N79), .SIN(ip1[1]), .SMC(test_se), .C(net12127), 
        .Q(ip1[2]) );
  SDFFQX1 ip0_reg_reg_4_ ( .D(N72), .SIN(ip0[3]), .SMC(test_se), .C(net12122), 
        .Q(ip0[4]) );
  SDFFQX1 ip0_reg_reg_5_ ( .D(N73), .SIN(ip0[4]), .SMC(test_se), .C(net12122), 
        .Q(ip0[5]) );
  SDFFQX1 isr_tm_reg_reg ( .D(n200), .SIN(is_reg[3]), .SMC(test_se), .C(clkper), .Q(isr_tm) );
  INVX1 U3 ( .A(1'b1), .Y(ien0[6]) );
  NOR2XL U5 ( .A(n4), .B(sfraddr[3]), .Y(n59) );
  AND4XL U6 ( .A(sfraddr[3]), .B(sfrwe), .C(sfraddr[5]), .D(n98), .Y(n91) );
  NAND4XL U7 ( .A(sfraddr[2]), .B(sfraddr[0]), .C(n59), .D(n60), .Y(n58) );
  AOI221XL U8 ( .A(n204), .B(ien0[4]), .C(ien1[4]), .D(int_vect_63), .E(n47), 
        .Y(n172) );
  OAI222XL U9 ( .A(n25), .B(n176), .C(n177), .D(n46), .E(n206), .F(n178), .Y(
        n128) );
  OAI222XL U10 ( .A(n24), .B(n31), .C(n185), .D(n56), .E(n55), .F(n175), .Y(
        n130) );
  NAND3X1 U11 ( .A(n3), .B(n5), .C(n91), .Y(n97) );
  NAND3X1 U12 ( .A(sfraddr[0]), .B(n5), .C(n91), .Y(n92) );
  NOR2X1 U13 ( .A(n10), .B(n93), .Y(N63) );
  NOR2X1 U14 ( .A(n11), .B(n93), .Y(N64) );
  NOR2X1 U15 ( .A(n6), .B(n93), .Y(N59) );
  NOR2X1 U16 ( .A(n7), .B(n93), .Y(N60) );
  NOR2X1 U17 ( .A(n9), .B(n93), .Y(N62) );
  NOR2X1 U18 ( .A(n8), .B(n93), .Y(N61) );
  NOR2X1 U19 ( .A(n8), .B(n92), .Y(N70) );
  NOR2X1 U20 ( .A(n6), .B(n92), .Y(N68) );
  NOR2X1 U21 ( .A(n10), .B(n92), .Y(N72) );
  NOR2X1 U22 ( .A(n9), .B(n92), .Y(N71) );
  NOR2X1 U23 ( .A(n11), .B(n92), .Y(N73) );
  NOR2X1 U24 ( .A(n7), .B(n92), .Y(N69) );
  NOR2X1 U25 ( .A(n6), .B(n97), .Y(N39) );
  NOR2X1 U26 ( .A(n8), .B(n97), .Y(N41) );
  NOR2X1 U27 ( .A(n11), .B(n97), .Y(N44) );
  NOR2X1 U28 ( .A(n7), .B(n97), .Y(N40) );
  NOR2X1 U29 ( .A(n9), .B(n97), .Y(N42) );
  NOR2X1 U30 ( .A(n10), .B(n97), .Y(N43) );
  NAND2X1 U31 ( .A(n12), .B(n93), .Y(N58) );
  NAND3X1 U32 ( .A(n91), .B(n3), .C(n4), .Y(n96) );
  NAND3X1 U33 ( .A(n91), .B(sfraddr[0]), .C(n4), .Y(n90) );
  INVX1 U34 ( .A(sfraddr[0]), .Y(n3) );
  NOR2X1 U35 ( .A(n90), .B(n6), .Y(N77) );
  NOR2X1 U36 ( .A(n90), .B(n10), .Y(N81) );
  NOR2X1 U37 ( .A(n90), .B(n9), .Y(N80) );
  NOR2X1 U38 ( .A(n90), .B(n7), .Y(N78) );
  NOR2X1 U39 ( .A(n90), .B(n8), .Y(N79) );
  NOR2X1 U40 ( .A(n11), .B(n90), .Y(N82) );
  NOR2X1 U41 ( .A(n7), .B(n96), .Y(N51) );
  NOR2X1 U42 ( .A(n11), .B(n96), .Y(N55) );
  NOR2X1 U43 ( .A(n10), .B(n96), .Y(N54) );
  NOR2X1 U44 ( .A(n9), .B(n96), .Y(N53) );
  NOR2X1 U45 ( .A(n6), .B(n96), .Y(N50) );
  NOR2X1 U46 ( .A(n8), .B(n96), .Y(N52) );
  NAND2X1 U47 ( .A(n12), .B(n90), .Y(N76) );
  NAND2X1 U48 ( .A(n12), .B(n92), .Y(N67) );
  NAND2X1 U49 ( .A(n12), .B(n96), .Y(N49) );
  NAND2X1 U50 ( .A(n12), .B(n97), .Y(N38) );
  INVX1 U51 ( .A(n5), .Y(n4) );
  INVX1 U52 ( .A(n171), .Y(n24) );
  INVX1 U53 ( .A(n70), .Y(n34) );
  NAND2X1 U54 ( .A(n12), .B(n208), .Y(n66) );
  NOR4XL U55 ( .A(sfraddr[6]), .B(sfraddr[2]), .C(sfraddr[1]), .D(rst), .Y(n98) );
  NOR42XL U56 ( .C(n12), .D(n95), .A(sfraddr[5]), .B(sfraddr[6]), .Y(n60) );
  AND2X1 U57 ( .A(sfraddr[1]), .B(sfrwe), .Y(n95) );
  NAND4X1 U58 ( .A(n4), .B(sfraddr[3]), .C(n94), .D(n60), .Y(n93) );
  NOR2X1 U59 ( .A(sfraddr[2]), .B(sfraddr[0]), .Y(n94) );
  NOR21XL U60 ( .B(sfrdatai[7]), .A(n97), .Y(N45) );
  INVX1 U61 ( .A(sfraddr[4]), .Y(n5) );
  NAND4X1 U62 ( .A(n119), .B(n12), .C(n124), .D(n125), .Y(N207) );
  NOR21XL U63 ( .B(n100), .A(n99), .Y(n125) );
  NOR21XL U64 ( .B(n99), .A(rst), .Y(N212) );
  NOR3XL U65 ( .A(n176), .B(n25), .C(n188), .Y(n171) );
  NAND3X1 U66 ( .A(n118), .B(n119), .C(n120), .Y(n106) );
  NAND4X1 U67 ( .A(n118), .B(n123), .C(n102), .D(n126), .Y(n99) );
  AOI21AX1 U68 ( .B(n115), .C(n15), .A(n109), .Y(n126) );
  INVX1 U69 ( .A(n168), .Y(n27) );
  INVX1 U70 ( .A(n108), .Y(n17) );
  INVX1 U71 ( .A(n145), .Y(n15) );
  INVX1 U72 ( .A(n170), .Y(n31) );
  INVX1 U73 ( .A(n165), .Y(n25) );
  INVX1 U74 ( .A(sfrdatai[5]), .Y(n11) );
  INVX1 U75 ( .A(sfrdatai[0]), .Y(n6) );
  INVX1 U76 ( .A(sfrdatai[2]), .Y(n8) );
  INVX1 U77 ( .A(sfrdatai[1]), .Y(n7) );
  INVX1 U78 ( .A(sfrdatai[3]), .Y(n9) );
  INVX1 U79 ( .A(sfrdatai[4]), .Y(n10) );
  AOI31X1 U80 ( .A(n16), .B(n14), .C(n114), .D(rst), .Y(N208) );
  INVX1 U81 ( .A(n113), .Y(n16) );
  AOI211X1 U82 ( .C(n115), .D(n15), .A(n116), .B(n117), .Y(n114) );
  INVX1 U83 ( .A(n106), .Y(n14) );
  AOI31X1 U84 ( .A(n109), .B(n110), .C(n111), .D(rst), .Y(N209) );
  NOR2X1 U85 ( .A(n112), .B(n113), .Y(n111) );
  NOR2X1 U86 ( .A(rst), .B(n100), .Y(N211) );
  INVX1 U87 ( .A(n193), .Y(n26) );
  NOR21XL U88 ( .B(n62), .A(n61), .Y(n70) );
  INVX1 U89 ( .A(intcall), .Y(n208) );
  NAND32X1 U90 ( .B(retiinstr), .C(rst), .A(n61), .Y(n67) );
  INVX1 U91 ( .A(rst), .Y(n12) );
  NAND2X1 U92 ( .A(intcall), .B(n12), .Y(n61) );
  OAI32X1 U93 ( .A(n51), .B(rst), .C(n13), .D(n58), .E(n11), .Y(n200) );
  INVX1 U94 ( .A(n58), .Y(n13) );
  NOR32XL U95 ( .B(n105), .C(n122), .A(n104), .Y(n124) );
  NAND31X1 U96 ( .C(n127), .A(n128), .B(n129), .Y(n109) );
  OAI21X1 U97 ( .B(n172), .C(n56), .A(n186), .Y(n168) );
  NOR3XL U98 ( .A(n45), .B(n161), .C(n150), .Y(n170) );
  AOI211X1 U99 ( .C(n135), .D(n144), .A(n115), .B(n145), .Y(n129) );
  NOR2X1 U100 ( .A(n194), .B(n54), .Y(n187) );
  NOR2X1 U101 ( .A(n189), .B(n158), .Y(n165) );
  NAND3X1 U102 ( .A(n146), .B(n143), .C(n124), .Y(n139) );
  NOR42XL U103 ( .C(n120), .D(n137), .A(n112), .B(n117), .Y(n100) );
  AOI22AXL U104 ( .A(n17), .B(n142), .D(n143), .C(n124), .Y(n137) );
  NAND2X1 U105 ( .A(n121), .B(n107), .Y(n142) );
  OAI21X1 U106 ( .B(n170), .C(n54), .A(n182), .Y(n175) );
  NAND3X1 U107 ( .A(n121), .B(n107), .C(n17), .Y(n145) );
  NAND3X1 U108 ( .A(n162), .B(n152), .C(n138), .Y(n176) );
  AND2X1 U109 ( .A(n184), .B(n194), .Y(n186) );
  AOI31X1 U110 ( .A(n101), .B(n102), .C(n103), .D(rst), .Y(N210) );
  OR2X1 U111 ( .A(n107), .B(n108), .Y(n101) );
  AOI21X1 U112 ( .B(n104), .C(n105), .A(n106), .Y(n103) );
  NAND3X1 U113 ( .A(n144), .B(n135), .C(n15), .Y(n120) );
  INVX1 U114 ( .A(n130), .Y(n23) );
  OAI221X1 U115 ( .A(n21), .B(n141), .C(n140), .D(n138), .E(n18), .Y(n108) );
  INVX1 U116 ( .A(n139), .Y(n18) );
  NAND31X1 U117 ( .C(n153), .A(n141), .B(n127), .Y(n188) );
  OAI221X1 U118 ( .A(n108), .B(n121), .C(n19), .D(n122), .E(n123), .Y(n113) );
  INVX1 U119 ( .A(n105), .Y(n19) );
  OA21X1 U120 ( .B(n23), .C(n148), .A(n131), .Y(n134) );
  NAND2X1 U121 ( .A(n153), .B(n128), .Y(n110) );
  OAI21X1 U122 ( .B(n21), .C(n127), .A(n129), .Y(n132) );
  AOI21X1 U123 ( .B(n133), .C(n45), .A(n132), .Y(n131) );
  AOI21X1 U124 ( .B(n134), .C(n147), .A(n66), .Y(N200) );
  NAND2X1 U125 ( .A(n136), .B(n135), .Y(n147) );
  INVX1 U126 ( .A(n172), .Y(n29) );
  NOR2X1 U127 ( .A(n152), .B(n140), .Y(n116) );
  NAND2X1 U128 ( .A(n150), .B(n133), .Y(n122) );
  NAND21X1 U129 ( .B(n146), .A(n124), .Y(n119) );
  NOR2X1 U130 ( .A(n50), .B(n190), .Y(n193) );
  NOR3XL U131 ( .A(n139), .B(n21), .C(n141), .Y(n112) );
  NOR3XL U132 ( .A(n138), .B(n139), .C(n140), .Y(n117) );
  NAND2X1 U133 ( .A(n161), .B(n133), .Y(n121) );
  INVX1 U134 ( .A(n128), .Y(n21) );
  NAND2X1 U135 ( .A(n155), .B(n154), .Y(n143) );
  NOR2X1 U136 ( .A(n162), .B(n140), .Y(n115) );
  OAI21X1 U137 ( .B(n206), .C(n166), .A(n167), .Y(n180) );
  NAND2X1 U138 ( .A(n88), .B(n37), .Y(n89) );
  OAI22X1 U139 ( .A(n72), .B(n57), .C(n73), .D(n74), .Y(n62) );
  AOI22X1 U140 ( .A(n39), .B(n75), .C(n76), .D(n38), .Y(n74) );
  OAI22X1 U141 ( .A(n40), .B(n56), .C(n79), .D(n50), .Y(n75) );
  OAI222XL U142 ( .A(n77), .B(n49), .C(n78), .D(n46), .E(n79), .F(n48), .Y(n76) );
  OAI32X1 U143 ( .A(n61), .B(n33), .C(n62), .D(n71), .E(n42), .Y(n196) );
  AOI21BBXL U144 ( .B(n66), .C(n65), .A(n70), .Y(n71) );
  AOI211X1 U145 ( .C(n83), .D(n84), .A(int_ack_03), .B(int_ack_43), .Y(n72) );
  OAI22X1 U146 ( .A(n67), .B(n44), .C(n33), .D(n34), .Y(n198) );
  OAI22X1 U147 ( .A(n63), .B(n34), .C(n68), .D(n43), .Y(n197) );
  AOI21BX1 U148 ( .C(n66), .B(n69), .A(n70), .Y(n68) );
  NOR2X1 U149 ( .A(n87), .B(n40), .Y(int_ack_43) );
  INVX1 U150 ( .A(n63), .Y(n33) );
  INVX1 U151 ( .A(n86), .Y(n39) );
  NOR2X1 U152 ( .A(n77), .B(n89), .Y(int_ack_1b) );
  OAI31XL U153 ( .A(n61), .B(n62), .C(n63), .D(n64), .Y(n199) );
  GEN2XL U154 ( .D(n65), .E(n42), .C(n66), .B(n61), .A(n41), .Y(n64) );
  NAND2X1 U155 ( .A(n44), .B(n67), .Y(n69) );
  NOR2X1 U156 ( .A(n78), .B(n89), .Y(int_ack_13) );
  NOR2X1 U157 ( .A(n78), .B(n87), .Y(int_ack_53) );
  NOR2X1 U158 ( .A(n79), .B(n87), .Y(int_ack_4b) );
  NOR2X1 U159 ( .A(n78), .B(n36), .Y(int_ack_93) );
  NOR2X1 U160 ( .A(n79), .B(n36), .Y(int_ack_8b) );
  INVX1 U161 ( .A(n83), .Y(n40) );
  INVX1 U162 ( .A(n84), .Y(n36) );
  NOR2X1 U163 ( .A(n77), .B(n87), .Y(int_ack_5b) );
  NOR2X1 U164 ( .A(n79), .B(n89), .Y(int_ack_0b) );
  NAND31X1 U165 ( .C(n132), .A(n45), .B(n133), .Y(n123) );
  NAND3X1 U166 ( .A(n47), .B(n130), .C(n131), .Y(n102) );
  NAND3X1 U167 ( .A(n134), .B(n135), .C(n136), .Y(n118) );
  NOR3XL U168 ( .A(n85), .B(n40), .C(n86), .Y(int_ack_a3) );
  NOR3XL U169 ( .A(n85), .B(n79), .C(n86), .Y(int_ack_ab) );
  INVX1 U170 ( .A(n203), .Y(n45) );
  NOR2X1 U171 ( .A(n77), .B(n36), .Y(int_ack_9b) );
  INVX1 U172 ( .A(n148), .Y(n47) );
  AND2X1 U173 ( .A(irq_r), .B(ien0[7]), .Y(irq) );
  NOR21XL U174 ( .B(n202), .A(n166), .Y(n183) );
  AOI33X1 U175 ( .A(ip0[1]), .B(n176), .C(ip1[1]), .D(ip0[2]), .E(n188), .F(
        ip1[2]), .Y(n202) );
  NOR21XL U176 ( .B(ien1[0]), .A(n205), .Y(n155) );
  AOI22X1 U177 ( .A(int_vect_43), .B(n51), .C(sdaiff), .D(isr_tm), .Y(n205) );
  OAI211X1 U178 ( .C(n57), .D(n192), .A(n44), .B(ien0[7]), .Y(n166) );
  NOR43XL U179 ( .B(n27), .C(n192), .D(n26), .A(is_reg[1]), .Y(n164) );
  AOI31X1 U180 ( .A(ip0[4]), .B(n30), .C(n183), .D(n186), .Y(n185) );
  INVX1 U181 ( .A(n187), .Y(n30) );
  AO21X1 U182 ( .B(ien0[0]), .C(int_vect_03), .A(n155), .Y(n189) );
  AOI21X1 U183 ( .B(n188), .C(ip0[2]), .A(n178), .Y(n182) );
  OAI21X1 U184 ( .B(n50), .C(n168), .A(n169), .Y(n135) );
  AOI32X1 U185 ( .A(n170), .B(n171), .C(n172), .D(ip0[5]), .E(n173), .Y(n169)
         );
  OAI22X1 U186 ( .A(n50), .B(n160), .C(n174), .D(n175), .Y(n173) );
  NOR2X1 U187 ( .A(n172), .B(n55), .Y(n174) );
  AND3X1 U188 ( .A(ien0[3]), .B(int_vect_1b), .C(n51), .Y(n150) );
  AOI211X1 U189 ( .C(n51), .D(n207), .A(n23), .B(n149), .Y(n104) );
  OAI21X1 U190 ( .B(n51), .C(rxd0ff), .A(ien0[4]), .Y(n149) );
  NAND2X1 U191 ( .A(n201), .B(n183), .Y(n160) );
  AOI31X1 U192 ( .A(ip0[4]), .B(n29), .C(ip1[4]), .D(n187), .Y(n201) );
  OAI211X1 U193 ( .C(n190), .D(n53), .A(n41), .B(n191), .Y(n158) );
  AOI21X1 U194 ( .B(ip0[4]), .C(n29), .A(n175), .Y(n191) );
  AOI221XL U195 ( .A(n176), .B(ip1[1]), .C(n188), .D(ip1[2]), .E(n167), .Y(
        n184) );
  INVX1 U196 ( .A(isr_tm), .Y(n51) );
  NAND2X1 U197 ( .A(int_vect_8b), .B(ien2[1]), .Y(n162) );
  OAI21BBX1 U198 ( .A(n176), .B(ip0[1]), .C(n164), .Y(n178) );
  NAND4X1 U199 ( .A(int_vect_4b), .B(ien1[1]), .C(n162), .D(n51), .Y(n138) );
  NAND3X1 U200 ( .A(n159), .B(n43), .C(n195), .Y(n167) );
  AOI21X1 U201 ( .B(ip1[0]), .C(n189), .A(n160), .Y(n195) );
  NAND2X1 U202 ( .A(ip1[3]), .B(n31), .Y(n194) );
  NAND3X1 U203 ( .A(i2c_int), .B(n135), .C(ien0[5]), .Y(n146) );
  NAND2X1 U204 ( .A(ip0[0]), .B(n189), .Y(n192) );
  AOI32X1 U205 ( .A(ip0[2]), .B(n52), .C(n32), .D(n179), .E(n180), .Y(n177) );
  NAND2X1 U206 ( .A(ip1[1]), .B(n176), .Y(n179) );
  INVX1 U207 ( .A(n166), .Y(n32) );
  ENOX1 U208 ( .A(n207), .B(isr_tm), .C(rxd0ff), .D(isr_tm), .Y(n204) );
  OAI221X1 U209 ( .A(n181), .B(n49), .C(n54), .D(n20), .E(n24), .Y(n133) );
  AOI21X1 U210 ( .B(n183), .C(ip0[3]), .A(n184), .Y(n181) );
  INVX1 U211 ( .A(n182), .Y(n20) );
  AOI221XL U212 ( .A(n163), .B(ip1[1]), .C(ip0[1]), .D(n164), .E(n165), .Y(
        n140) );
  OAI21X1 U213 ( .B(n166), .C(n52), .A(n167), .Y(n163) );
  AND3X1 U214 ( .A(ien1[3]), .B(int_vect_5b), .C(n203), .Y(n161) );
  OAI211X1 U215 ( .C(n156), .D(n57), .A(n157), .B(n158), .Y(n154) );
  AOI33X1 U216 ( .A(n159), .B(n43), .C(n28), .D(ip0[0]), .E(n44), .F(ien0[7]), 
        .Y(n156) );
  NAND4X1 U217 ( .A(n27), .B(ip0[0]), .C(n26), .D(n42), .Y(n157) );
  INVX1 U218 ( .A(n160), .Y(n28) );
  AND2X1 U219 ( .A(int_vect_13), .B(ien0[2]), .Y(n153) );
  NAND2X1 U220 ( .A(int_vect_93), .B(ien2[2]), .Y(n127) );
  NAND3X1 U221 ( .A(ien1[2]), .B(n127), .C(int_vect_53), .Y(n141) );
  NAND3X1 U222 ( .A(ien0[1]), .B(n51), .C(int_vect_0b), .Y(n152) );
  INVX1 U223 ( .A(int_vect_23), .Y(n207) );
  AOI211X1 U224 ( .C(int_vect_03), .D(n151), .A(n22), .B(n116), .Y(n105) );
  AND2X1 U225 ( .A(ien0[0]), .B(n154), .Y(n151) );
  INVX1 U226 ( .A(n110), .Y(n22) );
  NOR32XL U227 ( .B(ien1[5]), .C(int_vect_6b), .A(n136), .Y(n144) );
  AOI211X1 U228 ( .C(i2c_int), .D(ien0[5]), .A(n144), .B(n136), .Y(n190) );
  NAND4X1 U229 ( .A(int_vect_63), .B(ien1[4]), .C(n130), .D(n148), .Y(n107) );
  INVX1 U230 ( .A(is_reg[3]), .Y(n44) );
  INVX1 U231 ( .A(ip0[3]), .Y(n54) );
  NAND2X1 U232 ( .A(n193), .B(ip0[5]), .Y(n159) );
  INVX1 U233 ( .A(ip1[0]), .Y(n57) );
  INVX1 U234 ( .A(ip1[5]), .Y(n50) );
  INVX1 U235 ( .A(is_reg[2]), .Y(n43) );
  INVX1 U236 ( .A(ip1[4]), .Y(n56) );
  INVX1 U237 ( .A(ip0[2]), .Y(n206) );
  INVX1 U238 ( .A(ip0[5]), .Y(n53) );
  INVX1 U239 ( .A(is_reg[1]), .Y(n42) );
  INVX1 U240 ( .A(ip0[4]), .Y(n55) );
  INVX1 U241 ( .A(ip0[1]), .Y(n52) );
  INVX1 U242 ( .A(ip1[2]), .Y(n46) );
  INVX1 U243 ( .A(is_reg[0]), .Y(n41) );
  INVX1 U244 ( .A(ip1[3]), .Y(n49) );
  AO222X1 U245 ( .A(intcall), .B(n73), .C(n39), .D(intvect[1]), .E(n83), .F(
        n35), .Y(int_ack_03) );
  INVX1 U246 ( .A(n89), .Y(n35) );
  OAI22AX1 U247 ( .D(ip0[0]), .C(n72), .A(n73), .B(n80), .Y(n63) );
  AOI22X1 U248 ( .A(n39), .B(n81), .C(n82), .D(n38), .Y(n80) );
  OAI22X1 U249 ( .A(n40), .B(n55), .C(n79), .D(n53), .Y(n81) );
  OAI222XL U250 ( .A(n77), .B(n54), .C(n78), .D(n206), .E(n79), .F(n52), .Y(
        n82) );
  NAND2X1 U251 ( .A(intvect[2]), .B(intcall), .Y(n86) );
  NOR3XL U252 ( .A(intvect[2]), .B(intvect[4]), .C(n208), .Y(n88) );
  NAND2X1 U253 ( .A(n88), .B(intvect[3]), .Y(n87) );
  NOR3XL U254 ( .A(n208), .B(intvect[2]), .C(n85), .Y(n84) );
  INVX1 U255 ( .A(intvect[3]), .Y(n37) );
  NOR2X1 U256 ( .A(n69), .B(is_reg[2]), .Y(n65) );
  NAND21X1 U257 ( .B(intvect[1]), .A(intvect[0]), .Y(n79) );
  NAND21X1 U258 ( .B(intvect[0]), .A(intvect[1]), .Y(n78) );
  NOR2X1 U259 ( .A(intvect[0]), .B(intvect[1]), .Y(n83) );
  AND2X1 U260 ( .A(intvect[4]), .B(intvect[3]), .Y(n73) );
  NAND2X1 U261 ( .A(intvect[1]), .B(intvect[0]), .Y(n77) );
  NOR4XL U262 ( .A(intvect[4]), .B(n37), .C(n79), .D(n86), .Y(int_ack_6b) );
  NOR4XL U263 ( .A(intvect[4]), .B(n37), .C(n40), .D(n86), .Y(int_ack_63) );
  NAND2X1 U264 ( .A(intvect[4]), .B(n37), .Y(n85) );
  INVX1 U265 ( .A(ip1[1]), .Y(n48) );
  INVX1 U266 ( .A(intvect[2]), .Y(n38) );
  AND2X1 U268 ( .A(int_vect_ab), .B(ien2[5]), .Y(n136) );
  NAND2X1 U269 ( .A(int_vect_a3), .B(ien2[4]), .Y(n148) );
  NAND2X1 U270 ( .A(int_vect_9b), .B(ien2[3]), .Y(n203) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module watchdog_a0 ( wdt_slow, clkwdt, clkper, resetff, newinstr, wdts_s, wdts, 
        ip0wdts, wdt_tm, sfrdatai, sfraddr, sfrwe, wdtrel, test_si, test_se );
  output [1:0] wdts_s;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] wdtrel;
  input wdt_slow, clkwdt, clkper, resetff, newinstr, sfrwe, test_si, test_se;
  output wdts, ip0wdts, wdt_tm;
  wire   wdt_tm_sync, wdt_act_sync, wdt_act, wdtrefresh_sync, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N67, N68, N69, N70, N71, pres_2, N112,
         N113, N114, N115, N116, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, wdt_normal, wdt_normal_ff, N212, net12155, net12161,
         net12166, net12171, net12176, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n117, n118;
  wire   [1:0] pres_8;
  wire   [3:0] cycles_reg;
  wire   [3:0] pres_16;
  wire   [6:0] wdth;
  wire   [7:0] wdtl;

  SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 clk_gate_wdtrel_s_reg ( .CLK(clkper), 
        .EN(N26), .ENCLK(net12155), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 clk_gate_cycles_reg_reg ( .CLK(clkwdt), 
        .EN(N67), .ENCLK(net12161), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 clk_gate_pres_16_reg ( .CLK(clkwdt), .EN(
        N112), .ENCLK(net12166), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 clk_gate_wdth_reg ( .CLK(clkwdt), .EN(
        N165), .ENCLK(net12171), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 clk_gate_wdtl_reg ( .CLK(clkwdt), .EN(
        n116), .ENCLK(net12176), .TE(test_se) );
  watchdog_a0_DW01_inc_0 add_278 ( .A(wdtl), .SUM({N144, N143, N142, N141, 
        N140, N139, N138, N137}) );
  watchdog_a0_DW01_inc_1 add_272 ( .A(wdth), .SUM({N136, N135, N134, N133, 
        N132, N131, N130}) );
  SDFFQX1 wdt_act_reg ( .D(n130), .SIN(pres_16[3]), .SMC(test_se), .C(clkper), 
        .Q(wdt_act) );
  SDFFQX1 wdts_reg ( .D(wdts_s[0]), .SIN(wdtrel[7]), .SMC(test_se), .C(clkper), 
        .Q(wdts) );
  SDFFQX1 wdts_s_reg_1_ ( .D(n126), .SIN(wdts_s[0]), .SMC(test_se), .C(
        net12176), .Q(wdts_s[1]) );
  SDFFQX1 wdts_s_reg_0_ ( .D(n132), .SIN(wdts), .SMC(test_se), .C(net12176), 
        .Q(wdts_s[0]) );
  SDFFQX1 wdt_normal_ff_reg ( .D(n115), .SIN(wdt_act_sync), .SMC(test_se), .C(
        clkper), .Q(wdt_normal_ff) );
  SDFFQX1 wdt_normal_reg ( .D(n133), .SIN(wdt_normal_ff), .SMC(test_se), .C(
        clkper), .Q(wdt_normal) );
  SDFFQX1 wdt_act_sync_reg ( .D(wdt_act), .SIN(wdt_act), .SMC(test_se), .C(
        clkwdt), .Q(wdt_act_sync) );
  SDFFQX1 pres_16_reg_3_ ( .D(N116), .SIN(pres_16[2]), .SMC(test_se), .C(
        net12166), .Q(pres_16[3]) );
  SDFFQX1 wdth_reg_6_ ( .D(N172), .SIN(wdth[5]), .SMC(test_se), .C(net12171), 
        .Q(wdth[6]) );
  SDFFQX1 pres_8_reg_1_ ( .D(n128), .SIN(pres_8[0]), .SMC(test_se), .C(
        net12161), .Q(pres_8[1]) );
  SDFFQX1 pres_16_reg_2_ ( .D(N115), .SIN(pres_16[1]), .SMC(test_se), .C(
        net12166), .Q(pres_16[2]) );
  SDFFQX1 pres_2_reg ( .D(n127), .SIN(ip0wdts), .SMC(test_se), .C(net12161), 
        .Q(pres_2) );
  SDFFQX1 pres_8_reg_0_ ( .D(n129), .SIN(pres_2), .SMC(test_se), .C(net12161), 
        .Q(pres_8[0]) );
  SDFFQX1 wdt_tm_sync_reg ( .D(wdt_tm), .SIN(wdt_tm), .SMC(test_se), .C(clkwdt), .Q(wdt_tm_sync) );
  SDFFQX1 pres_16_reg_1_ ( .D(N114), .SIN(pres_16[0]), .SMC(test_se), .C(
        net12166), .Q(pres_16[1]) );
  SDFFQX1 cycles_reg_reg_2_ ( .D(N70), .SIN(cycles_reg[1]), .SMC(test_se), .C(
        net12161), .Q(cycles_reg[2]) );
  SDFFQX1 pres_16_reg_0_ ( .D(N113), .SIN(pres_8[1]), .SMC(test_se), .C(
        net12166), .Q(pres_16[0]) );
  SDFFQX1 wdth_reg_4_ ( .D(N170), .SIN(wdth[3]), .SMC(test_se), .C(net12171), 
        .Q(wdth[4]) );
  SDFFQX1 wdtl_reg_2_ ( .D(N175), .SIN(wdtl[1]), .SMC(test_se), .C(net12176), 
        .Q(wdtl[2]) );
  SDFFQX1 cycles_reg_reg_3_ ( .D(N71), .SIN(cycles_reg[2]), .SMC(test_se), .C(
        net12161), .Q(cycles_reg[3]) );
  SDFFQX1 wdtl_reg_4_ ( .D(N177), .SIN(wdtl[3]), .SMC(test_se), .C(net12176), 
        .Q(wdtl[4]) );
  SDFFQX1 wdtrefresh_reg ( .D(N212), .SIN(wdtl[7]), .SMC(test_se), .C(clkper), 
        .Q(wdtrefresh_sync) );
  SDFFQX1 cycles_reg_reg_1_ ( .D(N69), .SIN(cycles_reg[0]), .SMC(test_se), .C(
        net12161), .Q(cycles_reg[1]) );
  SDFFQX1 cycles_reg_reg_0_ ( .D(N68), .SIN(test_si), .SMC(test_se), .C(
        net12161), .Q(cycles_reg[0]) );
  SDFFQX1 wdth_reg_1_ ( .D(N167), .SIN(wdth[0]), .SMC(test_se), .C(net12171), 
        .Q(wdth[1]) );
  SDFFQX1 wdth_reg_3_ ( .D(N169), .SIN(wdth[2]), .SMC(test_se), .C(net12171), 
        .Q(wdth[3]) );
  SDFFQX1 wdth_reg_2_ ( .D(N168), .SIN(wdth[1]), .SMC(test_se), .C(net12171), 
        .Q(wdth[2]) );
  SDFFQX1 wdtl_reg_6_ ( .D(N179), .SIN(wdtl[5]), .SMC(test_se), .C(net12176), 
        .Q(wdtl[6]) );
  SDFFQX1 wdtl_reg_5_ ( .D(N178), .SIN(wdtl[4]), .SMC(test_se), .C(net12176), 
        .Q(wdtl[5]) );
  SDFFQX1 wdtl_reg_7_ ( .D(N180), .SIN(wdtl[6]), .SMC(test_se), .C(net12176), 
        .Q(wdtl[7]) );
  SDFFQX1 wdth_reg_5_ ( .D(N171), .SIN(wdth[4]), .SMC(test_se), .C(net12171), 
        .Q(wdth[5]) );
  SDFFQX1 wdtl_reg_1_ ( .D(N174), .SIN(wdtl[0]), .SMC(test_se), .C(net12176), 
        .Q(wdtl[1]) );
  SDFFQX1 wdtl_reg_3_ ( .D(N176), .SIN(wdtl[2]), .SMC(test_se), .C(net12176), 
        .Q(wdtl[3]) );
  SDFFQX1 wdth_reg_0_ ( .D(N166), .SIN(wdt_tm_sync), .SMC(test_se), .C(
        net12171), .Q(wdth[0]) );
  SDFFQX1 wdtl_reg_0_ ( .D(N173), .SIN(wdth[6]), .SMC(test_se), .C(net12176), 
        .Q(wdtl[0]) );
  SDFFQX1 wdtrel_s_reg_1_ ( .D(N28), .SIN(wdtrel[0]), .SMC(test_se), .C(
        net12155), .Q(wdtrel[1]) );
  SDFFQX1 wdtrel_s_reg_3_ ( .D(N30), .SIN(wdtrel[2]), .SMC(test_se), .C(
        net12155), .Q(wdtrel[3]) );
  SDFFQX1 wdtrel_s_reg_2_ ( .D(N29), .SIN(wdtrel[1]), .SMC(test_se), .C(
        net12155), .Q(wdtrel[2]) );
  SDFFQX1 ip0wdts_reg ( .D(n131), .SIN(cycles_reg[3]), .SMC(test_se), .C(
        clkper), .Q(ip0wdts) );
  SDFFQX1 wdtrel_s_reg_7_ ( .D(N34), .SIN(wdtrel[6]), .SMC(test_se), .C(
        net12155), .Q(wdtrel[7]) );
  SDFFQX1 wdt_tm_s_reg ( .D(n134), .SIN(wdt_normal), .SMC(test_se), .C(clkper), 
        .Q(wdt_tm) );
  SDFFQX1 wdtrel_s_reg_6_ ( .D(N33), .SIN(wdtrel[5]), .SMC(test_se), .C(
        net12155), .Q(wdtrel[6]) );
  SDFFQX1 wdtrel_s_reg_4_ ( .D(N31), .SIN(wdtrel[3]), .SMC(test_se), .C(
        net12155), .Q(wdtrel[4]) );
  SDFFQX1 wdtrel_s_reg_0_ ( .D(N27), .SIN(wdtrefresh_sync), .SMC(test_se), .C(
        net12155), .Q(wdtrel[0]) );
  SDFFQX1 wdtrel_s_reg_5_ ( .D(N32), .SIN(wdtrel[4]), .SMC(test_se), .C(
        net12155), .Q(wdtrel[5]) );
  NOR2X1 U3 ( .A(n58), .B(wdtrefresh_sync), .Y(n1) );
  NAND2X1 U4 ( .A(n33), .B(n2), .Y(n32) );
  INVX1 U5 ( .A(sfraddr[0]), .Y(n2) );
  INVX1 U6 ( .A(n4), .Y(n3) );
  INVX1 U7 ( .A(n110), .Y(n11) );
  AND4X1 U8 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(n48), .D(n49), .Y(n33) );
  NOR2X1 U9 ( .A(sfraddr[2]), .B(sfraddr[1]), .Y(n48) );
  NOR31X1 U10 ( .C(sfrwe), .A(sfraddr[4]), .B(sfraddr[6]), .Y(n49) );
  INVX1 U11 ( .A(n25), .Y(n5) );
  NOR21XL U12 ( .B(sfrdatai[4]), .A(n97), .Y(N31) );
  NOR21XL U13 ( .B(sfrdatai[5]), .A(n97), .Y(N32) );
  NOR21XL U14 ( .B(sfrdatai[2]), .A(n97), .Y(N29) );
  NOR21XL U15 ( .B(sfrdatai[0]), .A(n97), .Y(N27) );
  NOR21XL U16 ( .B(sfrdatai[1]), .A(n97), .Y(N28) );
  NOR21XL U17 ( .B(sfrdatai[3]), .A(n97), .Y(N30) );
  NOR21XL U18 ( .B(sfrdatai[7]), .A(n97), .Y(N34) );
  NOR2X1 U19 ( .A(n4), .B(n97), .Y(N33) );
  NAND4X1 U20 ( .A(sfrwe), .B(n2), .C(n99), .D(n100), .Y(n50) );
  AND4X1 U21 ( .A(sfraddr[3]), .B(sfraddr[5]), .C(sfraddr[4]), .D(n3), .Y(n100) );
  NOR3XL U22 ( .A(sfraddr[1]), .B(sfraddr[6]), .C(sfraddr[2]), .Y(n99) );
  INVX1 U23 ( .A(sfrdatai[6]), .Y(n4) );
  NAND2X1 U24 ( .A(n61), .B(n12), .Y(n110) );
  NOR32XL U25 ( .B(n117), .C(n32), .A(newinstr), .Y(n25) );
  NAND2X1 U26 ( .A(n31), .B(n2), .Y(n97) );
  NAND2X1 U27 ( .A(n117), .B(n97), .Y(N26) );
  NOR32XL U28 ( .B(n39), .C(n9), .A(n61), .Y(n60) );
  NOR3XL U29 ( .A(n14), .B(n13), .C(n15), .Y(n61) );
  NAND3X1 U30 ( .A(n66), .B(n67), .C(n68), .Y(n64) );
  AOI211X1 U31 ( .C(n80), .D(n81), .A(n82), .B(n83), .Y(n67) );
  AOI211X1 U32 ( .C(n87), .D(n118), .A(n88), .B(n89), .Y(n66) );
  NOR4XL U33 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(n68) );
  INVX1 U34 ( .A(n57), .Y(n15) );
  NAND2X1 U35 ( .A(n73), .B(n23), .Y(n85) );
  INVX1 U36 ( .A(n102), .Y(n16) );
  NAND2X1 U37 ( .A(n26), .B(n38), .Y(n35) );
  NOR21XL U38 ( .B(N143), .A(n35), .Y(N179) );
  NOR21XL U39 ( .B(N142), .A(n35), .Y(N178) );
  NOR21XL U40 ( .B(N141), .A(n35), .Y(N177) );
  NOR21XL U41 ( .B(N140), .A(n35), .Y(N176) );
  NOR21XL U42 ( .B(N138), .A(n35), .Y(N174) );
  NOR21XL U43 ( .B(N139), .A(n35), .Y(N175) );
  OAI21X1 U44 ( .B(n112), .C(n110), .A(n53), .Y(N115) );
  XNOR2XL U45 ( .A(n111), .B(n20), .Y(n112) );
  ENOX1 U46 ( .A(n22), .B(n28), .C(N135), .D(n26), .Y(N171) );
  ENOX1 U47 ( .A(n23), .B(n28), .C(N134), .D(n1), .Y(N170) );
  NAND2X1 U48 ( .A(n1), .B(n16), .Y(n93) );
  NOR2X1 U49 ( .A(n20), .B(n111), .Y(n105) );
  OAI211X1 U50 ( .C(n38), .D(n101), .A(n28), .B(n117), .Y(N165) );
  NAND21X1 U51 ( .B(n27), .A(n26), .Y(n101) );
  INVX1 U52 ( .A(n58), .Y(n12) );
  OAI2B11X1 U53 ( .D(n1), .C(n27), .A(n28), .B(n117), .Y(n116) );
  INVX1 U54 ( .A(n94), .Y(n17) );
  NAND2X1 U55 ( .A(n117), .B(n58), .Y(N67) );
  OAI32X1 U56 ( .A(n32), .B(resetff), .C(n4), .D(n10), .E(n5), .Y(n133) );
  OAI32X1 U57 ( .A(n10), .B(resetff), .C(n25), .D(n5), .E(n6), .Y(n115) );
  AND4X1 U58 ( .A(sfraddr[1]), .B(n49), .C(sfraddr[2]), .D(n98), .Y(n31) );
  NOR3XL U59 ( .A(resetff), .B(sfraddr[5]), .C(sfraddr[3]), .Y(n98) );
  OAI21X1 U60 ( .B(n29), .C(n4), .A(n30), .Y(n134) );
  NAND3X1 U61 ( .A(n29), .B(n117), .C(wdt_tm), .Y(n30) );
  NAND2X1 U62 ( .A(sfraddr[0]), .B(n31), .Y(n29) );
  AOI21X1 U63 ( .B(n45), .C(n46), .A(resetff), .Y(n131) );
  NAND21X1 U64 ( .B(n47), .A(n3), .Y(n45) );
  OAI21X1 U65 ( .B(ip0wdts), .C(wdts_s[0]), .A(n47), .Y(n46) );
  NAND2X1 U66 ( .A(sfraddr[0]), .B(n33), .Y(n47) );
  OAI31XL U67 ( .A(n50), .B(wdts_s[0]), .C(resetff), .D(n51), .Y(n130) );
  OAI21X1 U68 ( .B(wdts_s[0]), .C(n117), .A(wdt_act), .Y(n51) );
  NOR3XL U69 ( .A(n50), .B(resetff), .C(n6), .Y(N212) );
  NOR21XL U70 ( .B(n75), .A(wdtrel[3]), .Y(n73) );
  NOR21XL U71 ( .B(n77), .A(wdtrel[2]), .Y(n75) );
  XNOR2XL U72 ( .A(wdtrel[1]), .B(wdth[0]), .Y(n80) );
  XNOR2XL U73 ( .A(wdtrel[6]), .B(wdth[5]), .Y(n86) );
  XNOR2XL U74 ( .A(n75), .B(n76), .Y(n71) );
  XNOR2XL U75 ( .A(wdtrel[3]), .B(wdth[2]), .Y(n76) );
  XNOR2XL U76 ( .A(n73), .B(n74), .Y(n72) );
  XNOR2XL U77 ( .A(wdtrel[4]), .B(wdth[3]), .Y(n74) );
  XNOR2XL U78 ( .A(n77), .B(n78), .Y(n70) );
  XNOR2XL U79 ( .A(wdtrel[2]), .B(wdth[1]), .Y(n78) );
  XNOR2XL U80 ( .A(wdtl[7]), .B(wdt_slow), .Y(n44) );
  NOR3XL U81 ( .A(n94), .B(cycles_reg[2]), .C(n21), .Y(n102) );
  OAI22BX1 U82 ( .B(n34), .A(n35), .D(wdts_s[0]), .C(n34), .Y(n132) );
  OAI211X1 U83 ( .C(n36), .D(n37), .A(n38), .B(n39), .Y(n34) );
  NAND4X1 U84 ( .A(wdth[6]), .B(wdth[5]), .C(n40), .D(wdth[4]), .Y(n37) );
  NAND41X1 U85 ( .D(n41), .A(wdth[0]), .B(wdth[1]), .C(n42), .Y(n36) );
  NOR2X1 U86 ( .A(n16), .B(wdtrefresh_sync), .Y(n57) );
  NAND2X1 U87 ( .A(cycles_reg[1]), .B(cycles_reg[0]), .Y(n94) );
  OAI32X1 U88 ( .A(n59), .B(resetff), .C(n60), .D(n7), .E(n8), .Y(n127) );
  INVX1 U89 ( .A(pres_2), .Y(n7) );
  AOI21BBXL U90 ( .B(pres_2), .C(wdtrefresh_sync), .A(wdt_tm_sync), .Y(n59) );
  INVX1 U91 ( .A(n60), .Y(n8) );
  OAI21X1 U92 ( .B(n84), .C(n85), .A(n18), .Y(n82) );
  AOI22X1 U93 ( .A(n86), .B(n22), .C(wdtrel[5]), .D(wdth[4]), .Y(n84) );
  OAI22X1 U94 ( .A(n62), .B(n63), .C(n35), .D(n64), .Y(n126) );
  NAND2X1 U95 ( .A(wdts_s[1]), .B(n39), .Y(n63) );
  OAI2B11X1 U96 ( .D(wdtl[2]), .C(n65), .A(n64), .B(n38), .Y(n62) );
  NAND21X1 U97 ( .B(n43), .A(n41), .Y(n65) );
  NAND4X1 U98 ( .A(n106), .B(n107), .C(wdtl[0]), .D(n108), .Y(n43) );
  XNOR2XL U99 ( .A(n118), .B(wdtl[5]), .Y(n106) );
  NOR2X1 U100 ( .A(n18), .B(n19), .Y(n108) );
  XNOR2XL U101 ( .A(n118), .B(wdtl[6]), .Y(n107) );
  NOR3XL U102 ( .A(n43), .B(wdtl[2]), .C(n44), .Y(n42) );
  AOI21AX1 U103 ( .B(n90), .C(n86), .A(n85), .Y(n89) );
  XNOR2XL U104 ( .A(wdtrel[5]), .B(wdth[4]), .Y(n90) );
  OAI211X1 U105 ( .C(wdtl[7]), .D(n80), .A(wdtl[6]), .B(wdtl[4]), .Y(n87) );
  NOR2X1 U106 ( .A(wdtrel[1]), .B(wdtrel[0]), .Y(n77) );
  NAND3X1 U107 ( .A(wdtl[2]), .B(wdtl[0]), .C(n79), .Y(n69) );
  AOI22AXL U108 ( .A(wdtl[3]), .B(wdtl[5]), .D(wdtl[5]), .C(wdtl[6]), .Y(n79)
         );
  INVX1 U109 ( .A(wdtl[3]), .Y(n19) );
  INVX1 U110 ( .A(wdtl[1]), .Y(n18) );
  NAND2X1 U111 ( .A(n53), .B(n113), .Y(N114) );
  OAI211X1 U112 ( .C(pres_16[1]), .D(pres_16[0]), .A(n111), .B(n11), .Y(n113)
         );
  NAND3X1 U113 ( .A(n53), .B(n117), .C(n114), .Y(N112) );
  AOI22X1 U114 ( .A(n11), .B(pres_2), .C(n12), .D(wdtrefresh_sync), .Y(n114)
         );
  NAND42X1 U115 ( .C(n44), .D(n43), .A(wdtl[2]), .B(wdtl[4]), .Y(n38) );
  NAND31X1 U116 ( .C(n52), .A(n53), .B(n54), .Y(n129) );
  NAND4X1 U117 ( .A(n39), .B(pres_8[0]), .C(n15), .D(n9), .Y(n54) );
  XNOR2XL U118 ( .A(wdtl[4]), .B(n118), .Y(n41) );
  NOR21XL U119 ( .B(N137), .A(n35), .Y(N173) );
  NOR21XL U120 ( .B(N144), .A(n35), .Y(N180) );
  NOR2X1 U121 ( .A(n58), .B(wdtrefresh_sync), .Y(n26) );
  AO22AXL U122 ( .A(N136), .B(n1), .C(wdtrel[6]), .D(n28), .Y(N172) );
  INVX1 U123 ( .A(resetff), .Y(n117) );
  NAND2X1 U124 ( .A(wdt_act_sync), .B(n117), .Y(n58) );
  AND2X1 U125 ( .A(wdth[2]), .B(wdth[3]), .Y(n40) );
  NOR3XL U126 ( .A(n58), .B(pres_8[0]), .C(n15), .Y(n52) );
  OAI22X1 U127 ( .A(wdth[4]), .B(n86), .C(n91), .D(n118), .Y(n88) );
  AOI211X1 U128 ( .C(n80), .D(wdtl[4]), .A(n19), .B(wdtl[7]), .Y(n91) );
  OAI21X1 U129 ( .B(pres_16[0]), .C(n110), .A(n53), .Y(N113) );
  OAI21X1 U130 ( .B(n109), .C(n110), .A(n53), .Y(N116) );
  XNOR2XL U131 ( .A(pres_16[3]), .B(n105), .Y(n109) );
  OAI21X1 U132 ( .B(n92), .C(n93), .A(n53), .Y(N71) );
  AOI32X1 U133 ( .A(n17), .B(n21), .C(cycles_reg[2]), .D(cycles_reg[3]), .E(
        n94), .Y(n92) );
  OAI21X1 U134 ( .B(cycles_reg[0]), .C(n93), .A(n53), .Y(N68) );
  NAND2X1 U135 ( .A(pres_16[1]), .B(pres_16[0]), .Y(n111) );
  AOI21X1 U136 ( .B(wdtl[4]), .C(n24), .A(n80), .Y(n83) );
  OAI211X1 U137 ( .C(n55), .D(n14), .A(n56), .B(n53), .Y(n128) );
  NAND4X1 U138 ( .A(n57), .B(n12), .C(pres_8[0]), .D(n14), .Y(n56) );
  AOI31X1 U139 ( .A(n15), .B(n9), .C(n39), .D(n52), .Y(n55) );
  NAND4X1 U140 ( .A(n102), .B(n103), .C(pres_2), .D(n104), .Y(n27) );
  NOR2X1 U141 ( .A(n13), .B(n14), .Y(n104) );
  OAI21BBX1 U142 ( .A(n105), .B(pres_16[3]), .C(wdtrel[7]), .Y(n103) );
  INVX1 U143 ( .A(wdtrel[4]), .Y(n23) );
  INVX1 U144 ( .A(wdtrel[0]), .Y(n24) );
  INVX1 U145 ( .A(wdtrel[5]), .Y(n22) );
  OR2X1 U146 ( .A(wdtl[7]), .B(n24), .Y(n81) );
  INVX1 U147 ( .A(cycles_reg[3]), .Y(n21) );
  AO22AXL U148 ( .A(N132), .B(n26), .C(wdtrel[2]), .D(n28), .Y(N168) );
  AO22AXL U149 ( .A(N133), .B(n1), .C(wdtrel[3]), .D(n28), .Y(N169) );
  AO22AXL U150 ( .A(N131), .B(n26), .C(wdtrel[1]), .D(n28), .Y(N167) );
  NAND2X1 U151 ( .A(wdt_tm_sync), .B(n12), .Y(n53) );
  NOR2X1 U152 ( .A(wdtrefresh_sync), .B(resetff), .Y(n39) );
  NAND2X1 U153 ( .A(wdtrefresh_sync), .B(n117), .Y(n28) );
  OAI21X1 U154 ( .B(n93), .C(n96), .A(n53), .Y(N69) );
  OAI21X1 U155 ( .B(cycles_reg[1]), .C(cycles_reg[0]), .A(n94), .Y(n96) );
  INVX1 U156 ( .A(wdt_tm_sync), .Y(n9) );
  NOR3XL U157 ( .A(n93), .B(wdt_tm_sync), .C(n95), .Y(N70) );
  XNOR2XL U158 ( .A(n17), .B(cycles_reg[2]), .Y(n95) );
  INVX1 U159 ( .A(pres_8[1]), .Y(n14) );
  ENOX1 U160 ( .A(n24), .B(n28), .C(N130), .D(n26), .Y(N166) );
  INVX1 U161 ( .A(pres_8[0]), .Y(n13) );
  INVX1 U162 ( .A(pres_16[2]), .Y(n20) );
  INVX1 U163 ( .A(wdt_normal), .Y(n10) );
  INVX1 U164 ( .A(wdt_normal_ff), .Y(n6) );
  INVX1 U165 ( .A(wdt_slow), .Y(n118) );
endmodule


module watchdog_a0_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module watchdog_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer1_a0 ( clkper, rst, newinstr, t1ff, t1ack, int1ff, t1_tf1, t1ov, 
        sfrdatai, sfraddr, sfrwe, t1_tmod, t1_tr1, tl1, th1, test_si, test_se
 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t1_tmod;
  output [7:0] tl1;
  output [7:0] th1;
  input clkper, rst, newinstr, t1ff, t1ack, int1ff, sfrwe, test_si, test_se;
  output t1_tf1, t1ov, t1_tr1;
  wire   t1clr, th1_ov_ff, tl1_ov_ff, N31, N32, N33, N34, N35, N36, N37, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N95, N97, N98, clk_ov12, N100, net12193,
         net12199, net12204, n54, n55, n56, n57, n58, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n59, n60, n61, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19;
  wire   [1:0] t0_mode;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer1_a0_0 clk_gate_t1_mode_reg ( .CLK(clkper), .EN(
        N31), .ENCLK(net12193), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_2 clk_gate_tl1_s_reg ( .CLK(clkper), .EN(N50), 
        .ENCLK(net12199), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_1 clk_gate_th1_s_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12204), .TE(test_se) );
  timer1_a0_DW01_inc_0 add_278 ( .A(th1), .SUM({N75, N74, N73, N72, N71, N70, 
        N69, N68}) );
  timer1_a0_DW01_inc_1 add_244 ( .A(tl1), .SUM({N49, N48, N47, N46, N45, N44, 
        N43, N42}) );
  SDFFQX1 th1_ov_ff_reg ( .D(n55), .SIN(t1clr), .SMC(test_se), .C(clkper), .Q(
        th1_ov_ff) );
  SDFFQX1 tl1_ov_ff_reg ( .D(n56), .SIN(th1[7]), .SMC(test_se), .C(clkper), 
        .Q(tl1_ov_ff) );
  SDFFQX1 clk_count_reg_3_ ( .D(N98), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 clk_count_reg_2_ ( .D(N97), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 t1clr_reg ( .D(n57), .SIN(t1_tr1), .SMC(test_se), .C(clkper), .Q(
        t1clr) );
  SDFFQX1 clk_count_reg_1_ ( .D(n10), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 clk_count_reg_0_ ( .D(N95), .SIN(test_si), .SMC(test_se), .C(clkper), 
        .Q(clk_count[0]) );
  SDFFQX1 clk_ov12_reg ( .D(N100), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 t0_mode_reg_1_ ( .D(N37), .SIN(t0_mode[0]), .SMC(test_se), .C(
        net12193), .Q(t0_mode[1]) );
  SDFFQX1 t0_mode_reg_0_ ( .D(N36), .SIN(clk_ov12), .SMC(test_se), .C(net12193), .Q(t0_mode[0]) );
  SDFFQX1 t1_gate_reg ( .D(N32), .SIN(t1_tmod[2]), .SMC(test_se), .C(net12193), 
        .Q(t1_tmod[3]) );
  SDFFQX1 t1_ct_reg ( .D(N33), .SIN(t0_mode[1]), .SMC(test_se), .C(net12193), 
        .Q(t1_tmod[2]) );
  SDFFQX1 tl1_s_reg_7_ ( .D(N58), .SIN(tl1[6]), .SMC(test_se), .C(net12199), 
        .Q(tl1[7]) );
  SDFFQX1 tl1_s_reg_5_ ( .D(N56), .SIN(tl1[4]), .SMC(test_se), .C(net12199), 
        .Q(tl1[5]) );
  SDFFQX1 tl1_s_reg_4_ ( .D(N55), .SIN(tl1[3]), .SMC(test_se), .C(net12199), 
        .Q(tl1[4]) );
  SDFFQX1 th1_s_reg_1_ ( .D(N78), .SIN(th1[0]), .SMC(test_se), .C(net12204), 
        .Q(th1[1]) );
  SDFFQX1 tl1_s_reg_1_ ( .D(N52), .SIN(tl1[0]), .SMC(test_se), .C(net12199), 
        .Q(tl1[1]) );
  SDFFQX1 t1_tf1_s_reg ( .D(n54), .SIN(t1_tmod[1]), .SMC(test_se), .C(clkper), 
        .Q(t1_tf1) );
  SDFFQX1 t1_tr1_s_reg ( .D(n58), .SIN(t1_tf1), .SMC(test_se), .C(clkper), .Q(
        t1_tr1) );
  SDFFQX1 th1_s_reg_7_ ( .D(N84), .SIN(th1[6]), .SMC(test_se), .C(net12204), 
        .Q(th1[7]) );
  SDFFQX1 tl1_s_reg_6_ ( .D(N57), .SIN(tl1[5]), .SMC(test_se), .C(net12199), 
        .Q(tl1[6]) );
  SDFFQX1 th1_s_reg_3_ ( .D(N80), .SIN(th1[2]), .SMC(test_se), .C(net12204), 
        .Q(th1[3]) );
  SDFFQX1 th1_s_reg_6_ ( .D(N83), .SIN(th1[5]), .SMC(test_se), .C(net12204), 
        .Q(th1[6]) );
  SDFFQX1 th1_s_reg_5_ ( .D(N82), .SIN(th1[4]), .SMC(test_se), .C(net12204), 
        .Q(th1[5]) );
  SDFFQX1 th1_s_reg_4_ ( .D(N81), .SIN(th1[3]), .SMC(test_se), .C(net12204), 
        .Q(th1[4]) );
  SDFFQX1 tl1_s_reg_3_ ( .D(N54), .SIN(tl1[2]), .SMC(test_se), .C(net12199), 
        .Q(tl1[3]) );
  SDFFQX1 tl1_s_reg_2_ ( .D(N53), .SIN(tl1[1]), .SMC(test_se), .C(net12199), 
        .Q(tl1[2]) );
  SDFFQX1 tl1_s_reg_0_ ( .D(N51), .SIN(tl1_ov_ff), .SMC(test_se), .C(net12199), 
        .Q(tl1[0]) );
  SDFFQX1 th1_s_reg_0_ ( .D(N77), .SIN(th1_ov_ff), .SMC(test_se), .C(net12204), 
        .Q(th1[0]) );
  SDFFQX1 th1_s_reg_2_ ( .D(N79), .SIN(th1[1]), .SMC(test_se), .C(net12204), 
        .Q(th1[2]) );
  SDFFQX1 t1_mode_reg_0_ ( .D(N34), .SIN(t1_tmod[3]), .SMC(test_se), .C(
        net12193), .Q(t1_tmod[0]) );
  SDFFQX1 t1_mode_reg_1_ ( .D(N35), .SIN(t1_tmod[0]), .SMC(test_se), .C(
        net12193), .Q(t1_tmod[1]) );
  NAND3XL U3 ( .A(sfraddr[0]), .B(n29), .C(sfraddr[1]), .Y(n49) );
  NAND32XL U4 ( .B(sfraddr[0]), .C(sfraddr[1]), .A(n29), .Y(n21) );
  NAND42XL U5 ( .C(sfraddr[1]), .D(rst), .A(sfraddr[0]), .B(n29), .Y(n60) );
  INVX1 U6 ( .A(n21), .Y(n8) );
  NAND21X1 U7 ( .B(n43), .A(n7), .Y(n41) );
  NOR2X1 U8 ( .A(n4), .B(n60), .Y(N35) );
  NOR2X1 U9 ( .A(n3), .B(n60), .Y(N34) );
  NOR2X1 U10 ( .A(n6), .B(n60), .Y(N32) );
  NOR2X1 U11 ( .A(n5), .B(n60), .Y(N33) );
  NOR2X1 U12 ( .A(n1), .B(n60), .Y(N36) );
  NOR2X1 U13 ( .A(n2), .B(n60), .Y(N37) );
  NAND2X1 U14 ( .A(n7), .B(n60), .Y(N31) );
  NOR43XL U15 ( .B(sfraddr[3]), .C(n61), .D(sfrwe), .A(sfraddr[2]), .Y(n29) );
  NOR3XL U16 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n61) );
  NOR2X1 U17 ( .A(n49), .B(rst), .Y(n47) );
  OR4X1 U18 ( .A(n47), .B(n46), .C(n48), .D(rst), .Y(N50) );
  NAND4X1 U19 ( .A(sfraddr[2]), .B(sfraddr[0]), .C(n44), .D(n45), .Y(n43) );
  NOR4XL U20 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[4]), .D(sfraddr[1]), 
        .Y(n45) );
  AND2X1 U21 ( .A(sfraddr[3]), .B(sfrwe), .Y(n44) );
  INVX1 U22 ( .A(n42), .Y(n9) );
  NAND3X1 U23 ( .A(n41), .B(n7), .C(n42), .Y(N76) );
  INVX1 U24 ( .A(sfrdatai[4]), .Y(n3) );
  INVX1 U25 ( .A(sfrdatai[5]), .Y(n4) );
  INVX1 U26 ( .A(sfrdatai[0]), .Y(n1) );
  INVX1 U27 ( .A(sfrdatai[1]), .Y(n2) );
  INVX1 U28 ( .A(sfrdatai[7]), .Y(n6) );
  INVX1 U29 ( .A(sfrdatai[6]), .Y(n5) );
  INVX1 U30 ( .A(rst), .Y(n7) );
  INVX1 U31 ( .A(n37), .Y(n11) );
  NOR42XL U32 ( .C(n31), .D(n49), .A(rst), .B(n50), .Y(n48) );
  NOR32XL U33 ( .B(n49), .C(n7), .A(n31), .Y(n46) );
  AO22AXL U34 ( .A(N70), .B(n9), .C(sfrdatai[2]), .D(n41), .Y(N79) );
  AO22AXL U35 ( .A(N71), .B(n9), .C(sfrdatai[3]), .D(n41), .Y(N80) );
  NAND4X1 U36 ( .A(n16), .B(n43), .C(n7), .D(n18), .Y(n42) );
  ENOX1 U37 ( .A(n41), .B(n3), .C(N72), .D(n9), .Y(N81) );
  ENOX1 U38 ( .A(n41), .B(n4), .C(N73), .D(n9), .Y(N82) );
  ENOX1 U39 ( .A(n41), .B(n2), .C(N69), .D(n9), .Y(N78) );
  ENOX1 U40 ( .A(n5), .B(n41), .C(N74), .D(n9), .Y(N83) );
  NAND21X1 U41 ( .B(newinstr), .A(n7), .Y(n22) );
  NAND2X1 U42 ( .A(n24), .B(n31), .Y(t1ov) );
  INVX1 U43 ( .A(n23), .Y(n16) );
  NAND2X1 U44 ( .A(n7), .B(n40), .Y(n37) );
  NAND2X1 U45 ( .A(n11), .B(n38), .Y(n35) );
  INVX1 U46 ( .A(n38), .Y(n12) );
  NOR2X1 U47 ( .A(rst), .B(n40), .Y(N100) );
  OR4X1 U48 ( .A(t1ack), .B(t1clr), .C(n8), .D(rst), .Y(n28) );
  OAI22BX1 U49 ( .B(n25), .A(n26), .D(t1_tf1), .C(n25), .Y(n54) );
  AOI31X1 U50 ( .A(n8), .B(n7), .C(sfrdatai[7]), .D(n27), .Y(n26) );
  GEN2XL U51 ( .D(th1_ov_ff), .E(n18), .C(n15), .B(n27), .A(n28), .Y(n25) );
  AOI21X1 U52 ( .B(t0_mode[0]), .C(t0_mode[1]), .A(n28), .Y(n27) );
  AO222X1 U53 ( .A(n46), .B(th1[0]), .C(n47), .D(sfrdatai[0]), .E(N42), .F(n48), .Y(N51) );
  AO222X1 U54 ( .A(n46), .B(th1[4]), .C(n47), .D(sfrdatai[4]), .E(N46), .F(n48), .Y(N55) );
  AO222X1 U55 ( .A(n46), .B(th1[2]), .C(n47), .D(sfrdatai[2]), .E(N44), .F(n48), .Y(N53) );
  AO222X1 U56 ( .A(n46), .B(th1[3]), .C(n47), .D(sfrdatai[3]), .E(N45), .F(n48), .Y(N54) );
  AO222X1 U57 ( .A(n46), .B(th1[1]), .C(n47), .D(sfrdatai[1]), .E(N43), .F(n48), .Y(N52) );
  AO222X1 U58 ( .A(n46), .B(th1[6]), .C(n47), .D(sfrdatai[6]), .E(N48), .F(n48), .Y(N57) );
  AO222X1 U59 ( .A(n46), .B(th1[5]), .C(n47), .D(sfrdatai[5]), .E(N47), .F(n48), .Y(N56) );
  AO222X1 U60 ( .A(n46), .B(th1[7]), .C(n47), .D(sfrdatai[7]), .E(N49), .F(n48), .Y(N58) );
  ENOX1 U61 ( .A(n41), .B(n1), .C(N68), .D(n9), .Y(N77) );
  ENOX1 U62 ( .A(n6), .B(n41), .C(N75), .D(n9), .Y(N84) );
  NOR2X1 U63 ( .A(rst), .B(n20), .Y(n58) );
  AOI22X1 U64 ( .A(sfrdatai[6]), .B(n8), .C(t1_tr1), .D(n21), .Y(n20) );
  AO22AXL U65 ( .A(t1ack), .B(n7), .C(t1clr), .D(n22), .Y(n57) );
  OAI22AX1 U66 ( .D(tl1_ov_ff), .C(n22), .A(rst), .B(n23), .Y(n56) );
  OAI22AX1 U67 ( .D(th1_ov_ff), .C(n22), .A(rst), .B(n24), .Y(n55) );
  NAND4X1 U68 ( .A(tl1[3]), .B(tl1[2]), .C(tl1[4]), .D(n51), .Y(n23) );
  NOR42XL U69 ( .C(tl1[1]), .D(tl1[0]), .A(n50), .B(n52), .Y(n51) );
  AOI32X1 U70 ( .A(tl1[6]), .B(tl1[5]), .C(tl1[7]), .D(n18), .E(n17), .Y(n52)
         );
  NAND2X1 U71 ( .A(n16), .B(t1_tmod[1]), .Y(n31) );
  OAI211X1 U72 ( .C(n17), .D(n18), .A(clk_ov12), .B(n53), .Y(n50) );
  AOI211X1 U73 ( .C(t1_tmod[3]), .D(n19), .A(t1_tmod[2]), .B(n59), .Y(n53) );
  INVX1 U74 ( .A(int1ff), .Y(n19) );
  AOI21X1 U75 ( .B(t0_mode[1]), .C(t0_mode[0]), .A(t1_tr1), .Y(n59) );
  NAND4X1 U76 ( .A(th1[2]), .B(th1[1]), .C(n32), .D(n33), .Y(n24) );
  NOR32XL U77 ( .B(th1[7]), .C(th1[6]), .A(n34), .Y(n33) );
  AND3X1 U78 ( .A(th1[0]), .B(n18), .C(n16), .Y(n32) );
  NAND3X1 U79 ( .A(th1[4]), .B(th1[3]), .C(th1[5]), .Y(n34) );
  INVX1 U80 ( .A(n30), .Y(n15) );
  AOI31X1 U81 ( .A(tl1_ov_ff), .B(n17), .C(t1_tmod[1]), .D(t1ov), .Y(n30) );
  INVX1 U82 ( .A(t1_tmod[1]), .Y(n18) );
  INVX1 U83 ( .A(t1_tmod[0]), .Y(n17) );
  NAND2X1 U84 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n38) );
  OAI32X1 U85 ( .A(n37), .B(clk_count[2]), .C(n38), .D(n13), .E(n35), .Y(N97)
         );
  OAI21X1 U86 ( .B(n14), .C(n35), .A(n36), .Y(N98) );
  NAND4X1 U87 ( .A(clk_count[2]), .B(n11), .C(n12), .D(n14), .Y(n36) );
  INVX1 U88 ( .A(clk_count[3]), .Y(n14) );
  NAND3X1 U89 ( .A(n12), .B(n13), .C(clk_count[3]), .Y(n40) );
  INVX1 U90 ( .A(clk_count[2]), .Y(n13) );
  NOR2X1 U91 ( .A(clk_count[0]), .B(n37), .Y(N95) );
  INVX1 U92 ( .A(n39), .Y(n10) );
  OAI211X1 U93 ( .C(clk_count[0]), .D(clk_count[1]), .A(n11), .B(n38), .Y(n39)
         );
endmodule


module timer1_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module timer1_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer0_a0 ( clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, t0_tf0, 
        t0_tf1, sfrdatai, sfraddr, sfrwe, t0_tmod, t0_tr0, t0_tr1, tl0, th0, 
        test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t0_tmod;
  output [7:0] tl0;
  output [7:0] th0;
  input clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, sfrwe, test_si,
         test_se;
  output t0_tf0, t0_tf1, t0_tr0, t0_tr1;
  wire   t0clr, th0_ov_ff, tl0_ov_ff, t1clr, N39, N40, N41, N42, N43, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N101, N103, N104, clk_ov12, N106, net12221,
         net12227, net12232, n60, n61, n62, n63, n64, n65, n66, n67, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n68, n69, n70, n71, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n72, n73;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer0_a0_0 clk_gate_t0_ct_reg ( .CLK(clkper), .EN(N39), 
        .ENCLK(net12221), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_2 clk_gate_th0_s_reg ( .CLK(clkper), .EN(N55), 
        .ENCLK(net12227), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_1 clk_gate_tl0_s_reg ( .CLK(clkper), .EN(N79), 
        .ENCLK(net12232), .TE(test_se) );
  timer0_a0_DW01_inc_0 add_347 ( .A(tl0), .SUM({N78, N77, N76, N75, N74, N73, 
        N72, N71}) );
  timer0_a0_DW01_inc_1 add_309 ( .A(th0), .SUM({N54, N53, N52, N51, N50, N49, 
        N48, N47}) );
  SDFFQX1 th0_ov_ff_reg ( .D(n61), .SIN(t1clr), .SMC(test_se), .C(clkper), .Q(
        th0_ov_ff) );
  SDFFQX1 t1clr_reg ( .D(n63), .SIN(t0clr), .SMC(test_se), .C(clkper), .Q(
        t1clr) );
  SDFFQX1 tl0_ov_ff_reg ( .D(n64), .SIN(th0[7]), .SMC(test_se), .C(clkper), 
        .Q(tl0_ov_ff) );
  SDFFQX1 t0clr_reg ( .D(n65), .SIN(t0_tr1), .SMC(test_se), .C(clkper), .Q(
        t0clr) );
  SDFFQX1 clk_count_reg_3_ ( .D(N104), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 clk_count_reg_2_ ( .D(N103), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 clk_count_reg_1_ ( .D(n16), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 clk_count_reg_0_ ( .D(N101), .SIN(test_si), .SMC(test_se), .C(clkper), .Q(clk_count[0]) );
  SDFFQX1 clk_ov12_reg ( .D(N106), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 tl0_s_reg_7_ ( .D(N87), .SIN(tl0[6]), .SMC(test_se), .C(net12232), 
        .Q(tl0[7]) );
  SDFFQX1 tl0_s_reg_5_ ( .D(N85), .SIN(tl0[4]), .SMC(test_se), .C(net12232), 
        .Q(tl0[5]) );
  SDFFQX1 tl0_s_reg_6_ ( .D(N86), .SIN(tl0[5]), .SMC(test_se), .C(net12232), 
        .Q(tl0[6]) );
  SDFFQX1 tl0_s_reg_4_ ( .D(N84), .SIN(tl0[3]), .SMC(test_se), .C(net12232), 
        .Q(tl0[4]) );
  SDFFQX1 th0_s_reg_1_ ( .D(N57), .SIN(th0[0]), .SMC(test_se), .C(net12227), 
        .Q(th0[1]) );
  SDFFQX1 t0_tf1_s_reg ( .D(n62), .SIN(t0_tf0), .SMC(test_se), .C(clkper), .Q(
        t0_tf1) );
  SDFFQX1 th0_s_reg_7_ ( .D(N63), .SIN(th0[6]), .SMC(test_se), .C(net12227), 
        .Q(th0[7]) );
  SDFFQX1 t0_ct_reg ( .D(N41), .SIN(clk_ov12), .SMC(test_se), .C(net12221), 
        .Q(t0_tmod[2]) );
  SDFFQX1 t0_gate_reg ( .D(N40), .SIN(t0_tmod[2]), .SMC(test_se), .C(net12221), 
        .Q(t0_tmod[3]) );
  SDFFQX1 tl0_s_reg_1_ ( .D(N81), .SIN(tl0[0]), .SMC(test_se), .C(net12232), 
        .Q(tl0[1]) );
  SDFFQX1 t0_tr1_s_reg ( .D(n66), .SIN(t0_tr0), .SMC(test_se), .C(clkper), .Q(
        t0_tr1) );
  SDFFQX1 th0_s_reg_6_ ( .D(N62), .SIN(th0[5]), .SMC(test_se), .C(net12227), 
        .Q(th0[6]) );
  SDFFQX1 th0_s_reg_5_ ( .D(N61), .SIN(th0[4]), .SMC(test_se), .C(net12227), 
        .Q(th0[5]) );
  SDFFQX1 th0_s_reg_4_ ( .D(N60), .SIN(th0[3]), .SMC(test_se), .C(net12227), 
        .Q(th0[4]) );
  SDFFQX1 tl0_s_reg_3_ ( .D(N83), .SIN(tl0[2]), .SMC(test_se), .C(net12232), 
        .Q(tl0[3]) );
  SDFFQX1 tl0_s_reg_2_ ( .D(N82), .SIN(tl0[1]), .SMC(test_se), .C(net12232), 
        .Q(tl0[2]) );
  SDFFQX1 th0_s_reg_3_ ( .D(N59), .SIN(th0[2]), .SMC(test_se), .C(net12227), 
        .Q(th0[3]) );
  SDFFQX1 t0_tf0_s_reg ( .D(n60), .SIN(t0_tmod[1]), .SMC(test_se), .C(clkper), 
        .Q(t0_tf0) );
  SDFFQX1 th0_s_reg_2_ ( .D(N58), .SIN(th0[1]), .SMC(test_se), .C(net12227), 
        .Q(th0[2]) );
  SDFFQX1 t0_mode_reg_0_ ( .D(N42), .SIN(t0_tmod[3]), .SMC(test_se), .C(
        net12221), .Q(t0_tmod[0]) );
  SDFFQX1 t0_tr0_s_reg ( .D(n67), .SIN(t0_tf1), .SMC(test_se), .C(clkper), .Q(
        t0_tr0) );
  SDFFQX1 tl0_s_reg_0_ ( .D(N80), .SIN(tl0_ov_ff), .SMC(test_se), .C(net12232), 
        .Q(tl0[0]) );
  SDFFQX1 th0_s_reg_0_ ( .D(N56), .SIN(th0_ov_ff), .SMC(test_se), .C(net12227), 
        .Q(th0[0]) );
  SDFFQX1 t0_mode_reg_1_ ( .D(N43), .SIN(t0_tmod[0]), .SMC(test_se), .C(
        net12221), .Q(t0_tmod[1]) );
  NAND3XL U3 ( .A(n40), .B(n1), .C(sfraddr[1]), .Y(n46) );
  INVX1 U4 ( .A(n31), .Y(n13) );
  NOR2X1 U5 ( .A(n29), .B(n10), .Y(n31) );
  NOR2X1 U6 ( .A(n46), .B(n10), .Y(n43) );
  NOR2X1 U7 ( .A(n31), .B(n10), .Y(n24) );
  INVX1 U8 ( .A(sfraddr[1]), .Y(n2) );
  NAND3X1 U9 ( .A(n1), .B(n2), .C(n40), .Y(n29) );
  NAND4X1 U10 ( .A(sfraddr[0]), .B(n40), .C(n12), .D(n2), .Y(n56) );
  OR2X1 U11 ( .A(n49), .B(n11), .Y(n48) );
  NOR2X1 U12 ( .A(n3), .B(n56), .Y(N42) );
  NOR2X1 U13 ( .A(n4), .B(n56), .Y(N43) );
  NOR2X1 U14 ( .A(n5), .B(n56), .Y(N41) );
  NOR2X1 U15 ( .A(n6), .B(n56), .Y(N40) );
  INVX1 U16 ( .A(sfraddr[0]), .Y(n1) );
  NAND2X1 U17 ( .A(n12), .B(n56), .Y(N39) );
  INVX1 U18 ( .A(n12), .Y(n10) );
  INVX1 U19 ( .A(n12), .Y(n11) );
  NOR43XL U20 ( .B(sfraddr[3]), .C(n57), .D(sfrwe), .A(sfraddr[2]), .Y(n40) );
  NOR3XL U21 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n57) );
  OR4X1 U22 ( .A(n43), .B(n41), .C(n42), .D(n10), .Y(N79) );
  NAND4X1 U23 ( .A(sfraddr[2]), .B(sfrwe), .C(n50), .D(n51), .Y(n49) );
  NOR4XL U24 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[4]), .D(sfraddr[1]), 
        .Y(n51) );
  NOR21XL U25 ( .B(sfraddr[3]), .A(sfraddr[0]), .Y(n50) );
  INVX1 U26 ( .A(n47), .Y(n14) );
  NAND3X1 U27 ( .A(n47), .B(n12), .C(n48), .Y(N55) );
  INVX1 U28 ( .A(sfrdatai[0]), .Y(n3) );
  INVX1 U29 ( .A(sfrdatai[1]), .Y(n4) );
  INVX1 U30 ( .A(sfrdatai[2]), .Y(n5) );
  INVX1 U31 ( .A(sfrdatai[3]), .Y(n6) );
  INVX1 U32 ( .A(sfrdatai[4]), .Y(n7) );
  INVX1 U33 ( .A(sfrdatai[6]), .Y(n9) );
  INVX1 U34 ( .A(sfrdatai[5]), .Y(n8) );
  INVX1 U35 ( .A(rst), .Y(n12) );
  INVX1 U36 ( .A(n69), .Y(n17) );
  NOR43XL U37 ( .B(n44), .C(n45), .D(n46), .A(n10), .Y(n42) );
  NOR32XL U38 ( .B(n46), .C(n12), .A(n45), .Y(n41) );
  NAND3X1 U39 ( .A(n39), .B(n12), .C(n49), .Y(n47) );
  ENOX1 U40 ( .A(n6), .B(n48), .C(N50), .D(n14), .Y(N59) );
  ENOX1 U41 ( .A(n4), .B(n48), .C(N48), .D(n14), .Y(N57) );
  ENOX1 U42 ( .A(n9), .B(n48), .C(N53), .D(n14), .Y(N62) );
  ENOX1 U43 ( .A(n7), .B(n48), .C(N51), .D(n14), .Y(N60) );
  ENOX1 U44 ( .A(n8), .B(n48), .C(N52), .D(n14), .Y(N61) );
  ENOX1 U45 ( .A(n5), .B(n48), .C(N49), .D(n14), .Y(N58) );
  OAI22X1 U46 ( .A(n10), .B(n15), .C(n25), .D(n21), .Y(n65) );
  OAI22X1 U47 ( .A(n10), .B(n26), .C(n25), .D(n19), .Y(n64) );
  OR2X1 U48 ( .A(newinstr), .B(n11), .Y(n25) );
  INVX1 U49 ( .A(t0ack), .Y(n15) );
  NAND2X1 U50 ( .A(n12), .B(n58), .Y(n69) );
  NAND2X1 U51 ( .A(n17), .B(n70), .Y(n59) );
  INVX1 U52 ( .A(n70), .Y(n18) );
  NOR2X1 U53 ( .A(n10), .B(n58), .Y(N106) );
  AO222X1 U54 ( .A(n41), .B(th0[0]), .C(N71), .D(n42), .E(sfrdatai[0]), .F(n43), .Y(N80) );
  AO222X1 U55 ( .A(n41), .B(th0[4]), .C(N75), .D(n42), .E(n43), .F(sfrdatai[4]), .Y(N84) );
  AO222X1 U56 ( .A(n41), .B(th0[6]), .C(N77), .D(n42), .E(n43), .F(sfrdatai[6]), .Y(N86) );
  AO222X1 U57 ( .A(n41), .B(th0[5]), .C(N76), .D(n42), .E(n43), .F(sfrdatai[5]), .Y(N85) );
  AO222X1 U58 ( .A(n41), .B(th0[2]), .C(N73), .D(n42), .E(sfrdatai[2]), .F(n43), .Y(N82) );
  AO222X1 U59 ( .A(n41), .B(th0[3]), .C(N74), .D(n42), .E(sfrdatai[3]), .F(n43), .Y(N83) );
  AO222X1 U60 ( .A(n41), .B(th0[1]), .C(N72), .D(n42), .E(sfrdatai[1]), .F(n43), .Y(N81) );
  AO222X1 U61 ( .A(n41), .B(th0[7]), .C(N78), .D(n42), .E(n43), .F(sfrdatai[7]), .Y(N87) );
  OAI22BX1 U62 ( .B(n27), .A(n28), .D(t0_tf1), .C(n27), .Y(n62) );
  AOI32X1 U63 ( .A(n29), .B(n12), .C(n30), .D(sfrdatai[7]), .E(n31), .Y(n28)
         );
  OAI211X1 U64 ( .C(n72), .D(n32), .A(n24), .B(n30), .Y(n27) );
  NOR2X1 U65 ( .A(t1clr), .B(t1ack), .Y(n30) );
  OAI31XL U66 ( .A(n23), .B(th0_ov_ff), .C(t0_tmod[1]), .D(n29), .Y(n36) );
  INVX1 U67 ( .A(n32), .Y(n23) );
  OAI211X1 U68 ( .C(n13), .D(n8), .A(n33), .B(n34), .Y(n60) );
  NAND4X1 U69 ( .A(t0_tf0), .B(n24), .C(n15), .D(n21), .Y(n33) );
  NAND4X1 U70 ( .A(n15), .B(n21), .C(n12), .D(n35), .Y(n34) );
  AOI31X1 U71 ( .A(n26), .B(n19), .C(t0_tmod[1]), .D(n36), .Y(n35) );
  OAI22BX1 U72 ( .B(N54), .A(n47), .D(sfrdatai[7]), .C(n48), .Y(N63) );
  ENOX1 U73 ( .A(n13), .B(n7), .C(n24), .D(t0_tr0), .Y(n67) );
  ENOX1 U74 ( .A(n13), .B(n9), .C(n24), .D(t0_tr1), .Y(n66) );
  ENOX1 U75 ( .A(n3), .B(n48), .C(N47), .D(n14), .Y(N56) );
  OAI22BX1 U76 ( .B(t1ack), .A(n10), .D(t1clr), .C(n25), .Y(n63) );
  OAI22AX1 U77 ( .D(th0_ov_ff), .C(n25), .A(n10), .B(n32), .Y(n61) );
  NOR43XL U78 ( .B(t0_tr0), .C(n55), .D(clk_ov12), .A(t0_tmod[2]), .Y(n44) );
  NAND21X1 U79 ( .B(int0ff), .A(t0_tmod[3]), .Y(n55) );
  NAND4X1 U80 ( .A(th0[3]), .B(th0[2]), .C(n37), .D(n38), .Y(n32) );
  AND4X1 U81 ( .A(th0[4]), .B(th0[5]), .C(th0[6]), .D(th0[7]), .Y(n38) );
  AND3X1 U82 ( .A(th0[1]), .B(n39), .C(th0[0]), .Y(n37) );
  OAI21X1 U83 ( .B(t0_tmod[1]), .C(n26), .A(n52), .Y(n39) );
  NAND4X1 U84 ( .A(t0_tmod[1]), .B(t0_tmod[0]), .C(clk_ov12), .D(t0_tr1), .Y(
        n52) );
  NAND4X1 U85 ( .A(tl0[3]), .B(tl0[2]), .C(tl0[4]), .D(n53), .Y(n26) );
  NOR43XL U86 ( .B(tl0[1]), .C(tl0[0]), .D(n44), .A(n54), .Y(n53) );
  AOI32X1 U87 ( .A(tl0[6]), .B(tl0[5]), .C(tl0[7]), .D(n72), .E(n73), .Y(n54)
         );
  INVX1 U88 ( .A(t0_tmod[1]), .Y(n72) );
  INVX1 U89 ( .A(t0_tmod[0]), .Y(n73) );
  NAND31X1 U90 ( .C(n26), .A(n73), .B(t0_tmod[1]), .Y(n45) );
  NAND2X1 U91 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n70) );
  OAI32X1 U92 ( .A(n69), .B(clk_count[2]), .C(n70), .D(n20), .E(n59), .Y(N103)
         );
  NAND3X1 U93 ( .A(n18), .B(n20), .C(clk_count[3]), .Y(n58) );
  OAI21X1 U94 ( .B(n22), .C(n59), .A(n68), .Y(N104) );
  NAND4X1 U95 ( .A(clk_count[2]), .B(n17), .C(n18), .D(n22), .Y(n68) );
  INVX1 U96 ( .A(clk_count[3]), .Y(n22) );
  INVX1 U97 ( .A(t0clr), .Y(n21) );
  INVX1 U98 ( .A(clk_count[2]), .Y(n20) );
  NOR2X1 U99 ( .A(clk_count[0]), .B(n69), .Y(N101) );
  INVX1 U100 ( .A(n71), .Y(n16) );
  OAI211X1 U101 ( .C(clk_count[0]), .D(clk_count[1]), .A(n17), .B(n70), .Y(n71) );
  INVX1 U102 ( .A(tl0_ov_ff), .Y(n19) );
endmodule


module timer0_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module timer0_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module serial0_a0 ( t_shift_clk, r_shift_clk, clkper, rst, newinstr, rxd0ff, 
        t1ov, rxd0o, rxd0oe, txd0, sfrdatai, sfraddr, sfrwe, s0con, s0buf, 
        s0rell, s0relh, smod, bd, test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] s0con;
  output [7:0] s0buf;
  output [7:0] s0rell;
  output [7:0] s0relh;
  input clkper, rst, newinstr, rxd0ff, t1ov, sfrwe, test_si, test_se;
  output t_shift_clk, r_shift_clk, rxd0o, rxd0oe, txd0, smod, bd;
  wire   r_clk_ov2, t1ov_ff, N59, ri_tmp, rxd0_val, s0con2_val, s0con2_tmp,
         ti_tmp, N108, N109, N110, N111, N112, N113, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, baud_rate_ov, N142, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N166, N169, N170, N185, N186, N187,
         N188, N190, clk_ov12, N191, r_start, baud_r_count, baud_r2_clk, N207,
         t_baud_ov, t_start, N223, N224, N225, N226, N227, N230, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N281,
         N282, N283, N284, N303, rxd0_fall, rxd0_ff, rxd0_fall_fl,
         receive_11_bits, N306, N307, N324, N325, N326, N327, N333, ri0_fall,
         ri0_ff, N348, N360, N361, N362, N363, N364, N375, N376, N377, N378,
         N379, N380, N381, N382, N424, N425, N426, N427, N428, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, net12260, net12266,
         net12271, net12276, net12281, net12286, net12291, net12296, net12301,
         net12306, net12311, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n245, n27, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228;
  wire   [3:0] r_baud_count;
  wire   [3:0] r_shift_count;
  wire   [3:0] t_shift_count;
  wire   [9:0] tim_baud;
  wire   [3:0] clk_count;
  wire   [3:0] t_baud_count;
  wire   [10:0] t_shift_reg;
  wire   [1:0] fluctuation_conter;
  wire   [2:0] rxd0_vec;
  wire   [7:0] r_shift_reg;

  MAJ3X1 U329 ( .A(rxd0_vec[1]), .B(rxd0_vec[0]), .C(rxd0_vec[2]), .Y(n173) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_0 clk_gate_s0con_s_reg ( .CLK(clkper), .EN(
        N108), .ENCLK(net12260), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_10 clk_gate_s0rell_s_reg ( .CLK(clkper), 
        .EN(N117), .ENCLK(net12266), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_9 clk_gate_s0relh_s_reg ( .CLK(clkper), .EN(
        N128), .ENCLK(net12271), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_8 clk_gate_tim_baud_reg ( .CLK(clkper), .EN(
        N166), .ENCLK(net12276), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_7 clk_gate_t_baud_count_reg ( .CLK(clkper), 
        .EN(N223), .ENCLK(net12281), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_6 clk_gate_t_shift_reg_reg ( .CLK(clkper), 
        .EN(N257), .ENCLK(net12286), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_5 clk_gate_rxd0_vec_reg ( .CLK(clkper), .EN(
        N324), .ENCLK(net12291), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_4 clk_gate_r_baud_count_reg ( .CLK(clkper), 
        .EN(N360), .ENCLK(net12296), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_3 clk_gate_r_shift_reg_reg ( .CLK(clkper), 
        .EN(n27), .ENCLK(net12301), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_2 clk_gate_r_shift_count_reg ( .CLK(clkper), 
        .EN(N428), .ENCLK(net12306), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_1 clk_gate_s0buf_r_reg ( .CLK(clkper), .EN(
        N471), .ENCLK(net12311), .TE(test_se) );
  serial0_a0_DW01_inc_0 add_584 ( .A(tim_baud), .SUM({N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145}) );
  SDFFQX1 t_shift_reg_reg_10_ ( .D(N268), .SIN(t_shift_reg[9]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[10]) );
  SDFFQX1 r_shift_reg_reg_0_ ( .D(N375), .SIN(r_shift_count[3]), .SMC(test_se), 
        .C(net12301), .Q(r_shift_reg[0]) );
  SDFFQX1 t_shift_reg_reg_1_ ( .D(N259), .SIN(t_shift_reg[0]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[1]) );
  SDFFQX1 ti_tmp_reg ( .D(n242), .SIN(t_start), .SMC(test_se), .C(clkper), .Q(
        ti_tmp) );
  SDFFQX1 ri_tmp_reg ( .D(n238), .SIN(ri0_ff), .SMC(test_se), .C(clkper), .Q(
        ri_tmp) );
  SDFFQX1 t_shift_reg_reg_2_ ( .D(N260), .SIN(t_shift_reg[1]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[2]) );
  SDFFQX1 t_baud_count_reg_3_ ( .D(N227), .SIN(t_baud_count[2]), .SMC(test_se), 
        .C(net12281), .Q(t_baud_count[3]) );
  SDFFQX1 t_shift_reg_reg_0_ ( .D(N258), .SIN(t_shift_count[3]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[0]) );
  SDFFQX1 baud_r_count_reg ( .D(n245), .SIN(baud_r2_clk), .SMC(test_se), .C(
        clkper), .Q(baud_r_count) );
  SDFFQX1 r_shift_reg_reg_7_ ( .D(N382), .SIN(r_shift_reg[6]), .SMC(test_se), 
        .C(net12301), .Q(r_shift_reg[7]) );
  SDFFQX1 r_shift_reg_reg_6_ ( .D(N381), .SIN(r_shift_reg[5]), .SMC(test_se), 
        .C(net12301), .Q(r_shift_reg[6]) );
  SDFFQX1 r_shift_reg_reg_5_ ( .D(N380), .SIN(r_shift_reg[4]), .SMC(test_se), 
        .C(net12301), .Q(r_shift_reg[5]) );
  SDFFQX1 r_shift_reg_reg_4_ ( .D(N379), .SIN(r_shift_reg[3]), .SMC(test_se), 
        .C(net12301), .Q(r_shift_reg[4]) );
  SDFFQX1 r_shift_reg_reg_3_ ( .D(N378), .SIN(r_shift_reg[2]), .SMC(test_se), 
        .C(net12301), .Q(r_shift_reg[3]) );
  SDFFQX1 r_shift_reg_reg_2_ ( .D(N377), .SIN(r_shift_reg[1]), .SMC(test_se), 
        .C(net12301), .Q(r_shift_reg[2]) );
  SDFFQX1 r_shift_reg_reg_1_ ( .D(N376), .SIN(r_shift_reg[0]), .SMC(test_se), 
        .C(net12301), .Q(r_shift_reg[1]) );
  SDFFQX1 fluctuation_conter_reg_1_ ( .D(n233), .SIN(fluctuation_conter[0]), 
        .SMC(test_se), .C(clkper), .Q(fluctuation_conter[1]) );
  SDFFQX1 t_shift_reg_reg_9_ ( .D(N267), .SIN(t_shift_reg[8]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[9]) );
  SDFFQX1 t_shift_reg_reg_8_ ( .D(N266), .SIN(t_shift_reg[7]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[8]) );
  SDFFQX1 t_shift_reg_reg_7_ ( .D(N265), .SIN(t_shift_reg[6]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[7]) );
  SDFFQX1 t_shift_reg_reg_6_ ( .D(N264), .SIN(t_shift_reg[5]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[6]) );
  SDFFQX1 t_shift_reg_reg_5_ ( .D(N263), .SIN(t_shift_reg[4]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[5]) );
  SDFFQX1 t_shift_reg_reg_4_ ( .D(N262), .SIN(t_shift_reg[3]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[4]) );
  SDFFQX1 t_shift_reg_reg_3_ ( .D(N261), .SIN(t_shift_reg[2]), .SMC(test_se), 
        .C(net12286), .Q(t_shift_reg[3]) );
  SDFFQX1 rxd0_vec_reg_2_ ( .D(N327), .SIN(rxd0_vec[1]), .SMC(test_se), .C(
        net12291), .Q(rxd0_vec[2]) );
  SDFFQX1 rxd0_vec_reg_1_ ( .D(N326), .SIN(rxd0_vec[0]), .SMC(test_se), .C(
        net12291), .Q(rxd0_vec[1]) );
  SDFFQX1 rxd0_fall_fl_reg ( .D(n235), .SIN(ri_tmp), .SMC(test_se), .C(clkper), 
        .Q(rxd0_fall_fl) );
  SDFFQX1 rxd0_ff_reg ( .D(N307), .SIN(rxd0_fall), .SMC(test_se), .C(clkper), 
        .Q(rxd0_ff) );
  SDFFQX1 rxd0_vec_reg_0_ ( .D(N325), .SIN(rxd0_val), .SMC(test_se), .C(
        net12291), .Q(rxd0_vec[0]) );
  SDFFQX1 receive_11_bits_reg ( .D(n229), .SIN(r_start), .SMC(test_se), .C(
        clkper), .Q(receive_11_bits) );
  SDFFQX1 t_shift_count_reg_3_ ( .D(N284), .SIN(t_shift_count[2]), .SMC(
        test_se), .C(net12286), .Q(t_shift_count[3]) );
  SDFFQX1 fluctuation_conter_reg_0_ ( .D(n234), .SIN(clk_ov12), .SMC(test_se), 
        .C(clkper), .Q(fluctuation_conter[0]) );
  SDFFQX1 clk_count_reg_3_ ( .D(N188), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 s0con2_val_reg ( .D(n231), .SIN(s0con2_tmp), .SMC(test_se), .C(
        net12291), .Q(s0con2_val) );
  SDFFQX1 s0con2_tmp_reg ( .D(n232), .SIN(s0buf[7]), .SMC(test_se), .C(clkper), 
        .Q(s0con2_tmp) );
  SDFFQX1 clk_count_reg_2_ ( .D(N187), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 ri0_ff_reg ( .D(N348), .SIN(ri0_fall), .SMC(test_se), .C(clkper), 
        .Q(ri0_ff) );
  SDFFQX1 clk_ov12_reg ( .D(N191), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 t_baud_ov_reg ( .D(N230), .SIN(t_baud_count[3]), .SMC(test_se), .C(
        clkper), .Q(t_baud_ov) );
  SDFFQX1 tim_baud_reg_9_ ( .D(n67), .SIN(tim_baud[8]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[9]) );
  SDFFQX1 tim_baud_reg_8_ ( .D(n74), .SIN(tim_baud[7]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[8]) );
  SDFFQX1 tim_baud_reg_4_ ( .D(n70), .SIN(tim_baud[3]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[4]) );
  SDFFQX1 t_shift_count_reg_1_ ( .D(N282), .SIN(t_shift_count[0]), .SMC(
        test_se), .C(net12286), .Q(t_shift_count[1]) );
  SDFFQX1 t_shift_count_reg_2_ ( .D(N283), .SIN(t_shift_count[1]), .SMC(
        test_se), .C(net12286), .Q(t_shift_count[2]) );
  SDFFQX1 t_shift_count_reg_0_ ( .D(N281), .SIN(t_baud_ov), .SMC(test_se), .C(
        net12286), .Q(t_shift_count[0]) );
  SDFFQX1 ri0_fall_reg ( .D(n236), .SIN(receive_11_bits), .SMC(test_se), .C(
        clkper), .Q(ri0_fall) );
  SDFFQX1 rxd0_val_reg ( .D(N333), .SIN(rxd0_ff), .SMC(test_se), .C(clkper), 
        .Q(rxd0_val) );
  SDFFQX1 t_baud_count_reg_1_ ( .D(N225), .SIN(t_baud_count[0]), .SMC(test_se), 
        .C(net12281), .Q(t_baud_count[1]) );
  SDFFQX1 t_baud_count_reg_2_ ( .D(N226), .SIN(t_baud_count[1]), .SMC(test_se), 
        .C(net12281), .Q(t_baud_count[2]) );
  SDFFQX1 clk_count_reg_1_ ( .D(N186), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 t_baud_count_reg_0_ ( .D(N224), .SIN(t1ov_ff), .SMC(test_se), .C(
        net12281), .Q(t_baud_count[0]) );
  SDFFQX1 r_start_reg ( .D(n240), .SIN(r_shift_reg[7]), .SMC(test_se), .C(
        clkper), .Q(r_start) );
  SDFFQX1 clk_count_reg_0_ ( .D(N185), .SIN(bd), .SMC(test_se), .C(clkper), 
        .Q(clk_count[0]) );
  SDFFQX1 rxd0_fall_reg ( .D(N306), .SIN(rxd0_fall_fl), .SMC(test_se), .C(
        clkper), .Q(rxd0_fall) );
  SDFFQX1 baud_r2_clk_reg ( .D(N207), .SIN(test_si), .SMC(test_se), .C(clkper), 
        .Q(baud_r2_clk) );
  SDFFQX1 tim_baud_reg_2_ ( .D(N169), .SIN(tim_baud[1]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[2]) );
  SDFFQX1 tim_baud_reg_7_ ( .D(n73), .SIN(tim_baud[6]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[7]) );
  SDFFQX1 tim_baud_reg_5_ ( .D(n71), .SIN(tim_baud[4]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[5]) );
  SDFFQX1 tim_baud_reg_1_ ( .D(n69), .SIN(tim_baud[0]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[1]) );
  SDFFQX1 tim_baud_reg_6_ ( .D(n72), .SIN(tim_baud[5]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[6]) );
  SDFFQX1 tim_baud_reg_3_ ( .D(N170), .SIN(tim_baud[2]), .SMC(test_se), .C(
        net12276), .Q(tim_baud[3]) );
  SDFFQX1 r_shift_count_reg_1_ ( .D(N425), .SIN(r_shift_count[0]), .SMC(
        test_se), .C(net12306), .Q(r_shift_count[1]) );
  SDFFQX1 r_shift_count_reg_3_ ( .D(N427), .SIN(r_shift_count[2]), .SMC(
        test_se), .C(net12306), .Q(r_shift_count[3]) );
  SDFFQX1 r_baud_count_reg_1_ ( .D(N362), .SIN(r_baud_count[0]), .SMC(test_se), 
        .C(net12296), .Q(r_baud_count[1]) );
  SDFFQX1 r_shift_count_reg_2_ ( .D(N426), .SIN(r_shift_count[1]), .SMC(
        test_se), .C(net12306), .Q(r_shift_count[2]) );
  SDFFQX1 r_shift_count_reg_0_ ( .D(N424), .SIN(r_clk_ov2), .SMC(test_se), .C(
        net12306), .Q(r_shift_count[0]) );
  SDFFQX1 r_baud_count_reg_3_ ( .D(N364), .SIN(r_baud_count[2]), .SMC(test_se), 
        .C(net12296), .Q(r_baud_count[3]) );
  SDFFQX1 r_baud_count_reg_2_ ( .D(N363), .SIN(r_baud_count[1]), .SMC(test_se), 
        .C(net12296), .Q(r_baud_count[2]) );
  SDFFQX1 tim_baud_reg_0_ ( .D(n68), .SIN(ti_tmp), .SMC(test_se), .C(net12276), 
        .Q(tim_baud[0]) );
  SDFFQX1 r_baud_count_reg_0_ ( .D(N361), .SIN(fluctuation_conter[1]), .SMC(
        test_se), .C(net12296), .Q(r_baud_count[0]) );
  SDFFQX1 t1ov_ff_reg ( .D(N59), .SIN(smod), .SMC(test_se), .C(clkper), .Q(
        t1ov_ff) );
  SDFFQX1 baud_rate_ov_reg ( .D(N142), .SIN(baud_r_count), .SMC(test_se), .C(
        clkper), .Q(baud_rate_ov) );
  SDFFQX1 r_clk_ov2_reg ( .D(N190), .SIN(r_baud_count[3]), .SMC(test_se), .C(
        clkper), .Q(r_clk_ov2) );
  SDFFQX1 t_start_reg ( .D(n243), .SIN(t_shift_reg[10]), .SMC(test_se), .C(
        clkper), .Q(t_start) );
  SDFFQX1 rxd0o_reg ( .D(N303), .SIN(rxd0_vec[2]), .SMC(test_se), .C(clkper), 
        .Q(rxd0o) );
  SDFFQX1 txd0_reg ( .D(n239), .SIN(tim_baud[9]), .SMC(test_se), .C(clkper), 
        .Q(txd0) );
  SDFFQX1 s0buf_r_reg_7_ ( .D(N479), .SIN(s0buf[6]), .SMC(test_se), .C(
        net12311), .Q(s0buf[7]) );
  SDFFQX1 s0relh_s_reg_3_ ( .D(N132), .SIN(s0relh[2]), .SMC(test_se), .C(
        net12271), .Q(s0relh[3]) );
  SDFFQX1 s0rell_s_reg_3_ ( .D(N121), .SIN(s0rell[2]), .SMC(test_se), .C(
        net12266), .Q(s0rell[3]) );
  SDFFQX1 s0rell_s_reg_7_ ( .D(N125), .SIN(s0rell[6]), .SMC(test_se), .C(
        net12266), .Q(s0rell[7]) );
  SDFFQX1 s0rell_s_reg_6_ ( .D(N124), .SIN(s0rell[5]), .SMC(test_se), .C(
        net12266), .Q(s0rell[6]) );
  SDFFQX1 s0rell_s_reg_0_ ( .D(N118), .SIN(s0relh[7]), .SMC(test_se), .C(
        net12266), .Q(s0rell[0]) );
  SDFFQX1 s0relh_s_reg_0_ ( .D(N129), .SIN(s0con[7]), .SMC(test_se), .C(
        net12271), .Q(s0relh[0]) );
  SDFFQX1 bd_s_reg ( .D(n29), .SIN(baud_rate_ov), .SMC(test_se), .C(clkper), 
        .Q(bd) );
  SDFFQX1 s0relh_s_reg_1_ ( .D(N130), .SIN(s0relh[0]), .SMC(test_se), .C(
        net12271), .Q(s0relh[1]) );
  SDFFQX1 s0rell_s_reg_1_ ( .D(N119), .SIN(s0rell[0]), .SMC(test_se), .C(
        net12266), .Q(s0rell[1]) );
  SDFFQX1 s0con_s_reg_1_ ( .D(n241), .SIN(s0con[0]), .SMC(test_se), .C(clkper), 
        .Q(s0con[1]) );
  SDFFQX1 s0buf_r_reg_1_ ( .D(N473), .SIN(s0buf[0]), .SMC(test_se), .C(
        net12311), .Q(s0buf[1]) );
  SDFFQX1 s0buf_r_reg_3_ ( .D(N475), .SIN(s0buf[2]), .SMC(test_se), .C(
        net12311), .Q(s0buf[3]) );
  SDFFQX1 s0buf_r_reg_6_ ( .D(N478), .SIN(s0buf[5]), .SMC(test_se), .C(
        net12311), .Q(s0buf[6]) );
  SDFFQX1 s0buf_r_reg_0_ ( .D(N472), .SIN(rxd0o), .SMC(test_se), .C(net12311), 
        .Q(s0buf[0]) );
  SDFFQX1 s0buf_r_reg_2_ ( .D(N474), .SIN(s0buf[1]), .SMC(test_se), .C(
        net12311), .Q(s0buf[2]) );
  SDFFQX1 s0relh_s_reg_4_ ( .D(N133), .SIN(s0relh[3]), .SMC(test_se), .C(
        net12271), .Q(s0relh[4]) );
  SDFFQX1 s0relh_s_reg_2_ ( .D(N131), .SIN(s0relh[1]), .SMC(test_se), .C(
        net12271), .Q(s0relh[2]) );
  SDFFQX1 s0relh_s_reg_5_ ( .D(N134), .SIN(s0relh[4]), .SMC(test_se), .C(
        net12271), .Q(s0relh[5]) );
  SDFFQX1 s0buf_r_reg_5_ ( .D(N477), .SIN(s0buf[4]), .SMC(test_se), .C(
        net12311), .Q(s0buf[5]) );
  SDFFQX1 s0buf_r_reg_4_ ( .D(N476), .SIN(s0buf[3]), .SMC(test_se), .C(
        net12311), .Q(s0buf[4]) );
  SDFFQX1 s0con_s_reg_3_ ( .D(N109), .SIN(s0con[2]), .SMC(test_se), .C(
        net12260), .Q(s0con[3]) );
  SDFFQX1 s0rell_s_reg_2_ ( .D(N120), .SIN(s0rell[1]), .SMC(test_se), .C(
        net12266), .Q(s0rell[2]) );
  SDFFQX1 s0rell_s_reg_4_ ( .D(N122), .SIN(s0rell[3]), .SMC(test_se), .C(
        net12266), .Q(s0rell[4]) );
  SDFFQX1 s0rell_s_reg_5_ ( .D(N123), .SIN(s0rell[4]), .SMC(test_se), .C(
        net12266), .Q(s0rell[5]) );
  SDFFQX1 s0con_s_reg_5_ ( .D(N111), .SIN(s0con[4]), .SMC(test_se), .C(
        net12260), .Q(s0con[5]) );
  SDFFQX1 smod_s_reg ( .D(n28), .SIN(s0rell[7]), .SMC(test_se), .C(clkper), 
        .Q(smod) );
  SDFFQX1 s0con_s_reg_0_ ( .D(n237), .SIN(s0con2_val), .SMC(test_se), .C(
        clkper), .Q(s0con[0]) );
  SDFFQX1 s0con_s_reg_6_ ( .D(N112), .SIN(s0con[5]), .SMC(test_se), .C(
        net12260), .Q(s0con[6]) );
  SDFFQX1 s0con_s_reg_4_ ( .D(N110), .SIN(s0con[3]), .SMC(test_se), .C(
        net12260), .Q(s0con[4]) );
  SDFFQX1 s0relh_s_reg_7_ ( .D(N136), .SIN(s0relh[6]), .SMC(test_se), .C(
        net12271), .Q(s0relh[7]) );
  SDFFQX1 s0relh_s_reg_6_ ( .D(N135), .SIN(s0relh[5]), .SMC(test_se), .C(
        net12271), .Q(s0relh[6]) );
  SDFFQX1 s0con_s_reg_7_ ( .D(N113), .SIN(s0con[6]), .SMC(test_se), .C(
        net12260), .Q(s0con[7]) );
  SDFFQX1 s0con_s_reg_2_ ( .D(n230), .SIN(s0con[1]), .SMC(test_se), .C(clkper), 
        .Q(s0con[2]) );
  BUFX3 U3 ( .A(n84), .Y(n1) );
  BUFX3 U4 ( .A(n83), .Y(n2) );
  NAND2X1 U5 ( .A(n227), .B(n226), .Y(n3) );
  AOI221XL U6 ( .A(r_start), .B(n114), .C(n3), .D(r_shift_clk), .E(n20), .Y(
        n81) );
  INVX1 U7 ( .A(N108), .Y(n32) );
  NAND2X1 U8 ( .A(n15), .B(n131), .Y(N108) );
  INVX1 U9 ( .A(n181), .Y(n35) );
  INVX1 U10 ( .A(n131), .Y(n31) );
  NAND2X1 U11 ( .A(n26), .B(n212), .Y(N128) );
  NAND4X1 U12 ( .A(n94), .B(n95), .C(n15), .D(n6), .Y(n131) );
  NOR2X1 U13 ( .A(n193), .B(n19), .Y(n181) );
  INVX1 U14 ( .A(n183), .Y(n36) );
  NAND2X1 U15 ( .A(n213), .B(sfraddr[4]), .Y(n212) );
  AOI31X1 U16 ( .A(n94), .B(n6), .C(n95), .D(n22), .Y(n107) );
  NAND2X1 U17 ( .A(n15), .B(n214), .Y(N117) );
  NOR32XL U18 ( .B(n16), .C(sfraddr[1]), .A(sfraddr[6]), .Y(n100) );
  INVX1 U19 ( .A(n21), .Y(n16) );
  INVX1 U20 ( .A(n21), .Y(n15) );
  INVX1 U21 ( .A(n20), .Y(n18) );
  INVX1 U22 ( .A(n21), .Y(n17) );
  NOR4XL U23 ( .A(n34), .B(n4), .C(sfraddr[0]), .D(sfraddr[2]), .Y(n94) );
  NAND2X1 U24 ( .A(n181), .B(n225), .Y(n183) );
  NAND4X1 U25 ( .A(n95), .B(sfrwe), .C(sfraddr[0]), .D(n194), .Y(n193) );
  NOR3XL U26 ( .A(n4), .B(sfraddr[6]), .C(sfraddr[2]), .Y(n194) );
  INVX1 U27 ( .A(sfrwe), .Y(n34) );
  AND3X1 U28 ( .A(n100), .B(n94), .C(sfraddr[5]), .Y(n213) );
  NAND2X1 U29 ( .A(n213), .B(n5), .Y(n214) );
  INVX1 U30 ( .A(n176), .Y(n38) );
  OAI21X1 U31 ( .B(n131), .C(n13), .A(n18), .Y(N112) );
  OAI21X1 U32 ( .B(n13), .C(n214), .A(n18), .Y(N124) );
  OAI21X1 U33 ( .B(n7), .C(n214), .A(n24), .Y(N118) );
  OAI21X1 U34 ( .B(n11), .C(n214), .A(n18), .Y(N122) );
  OAI21X1 U35 ( .B(n14), .C(n214), .A(n18), .Y(N125) );
  OAI21X1 U36 ( .B(n10), .C(n214), .A(n24), .Y(N121) );
  OAI21X1 U37 ( .B(n7), .C(n212), .A(n18), .Y(N129) );
  OAI21X1 U38 ( .B(n8), .C(n212), .A(n18), .Y(N130) );
  NOR2X1 U39 ( .A(n12), .B(n214), .Y(N123) );
  NOR2X1 U40 ( .A(n8), .B(n214), .Y(N119) );
  NOR2X1 U41 ( .A(n9), .B(n214), .Y(N120) );
  NOR2X1 U42 ( .A(n13), .B(n212), .Y(N135) );
  NOR2X1 U43 ( .A(n14), .B(n212), .Y(N136) );
  NOR2X1 U44 ( .A(n9), .B(n212), .Y(N131) );
  NOR2X1 U45 ( .A(n10), .B(n212), .Y(N132) );
  NOR2X1 U46 ( .A(n11), .B(n212), .Y(N133) );
  NOR2X1 U47 ( .A(n12), .B(n212), .Y(N134) );
  NOR2X1 U48 ( .A(n14), .B(n131), .Y(N113) );
  NOR3XL U49 ( .A(sfraddr[1]), .B(sfraddr[5]), .C(n5), .Y(n95) );
  INVX1 U50 ( .A(sfraddr[6]), .Y(n6) );
  NOR2X1 U51 ( .A(n131), .B(n11), .Y(N110) );
  NOR2X1 U52 ( .A(n131), .B(n10), .Y(N109) );
  NOR2X1 U53 ( .A(n131), .B(n12), .Y(N111) );
  NAND3X1 U54 ( .A(n35), .B(n17), .C(n176), .Y(N257) );
  NAND21X1 U55 ( .B(n130), .A(n15), .Y(n127) );
  INVX1 U56 ( .A(n25), .Y(n21) );
  INVX1 U57 ( .A(n24), .Y(n23) );
  INVX1 U58 ( .A(n26), .Y(n19) );
  INVX1 U59 ( .A(n25), .Y(n22) );
  INVX1 U60 ( .A(n26), .Y(n20) );
  NAND3X1 U61 ( .A(n193), .B(n16), .C(t_shift_clk), .Y(n176) );
  NAND2X1 U62 ( .A(n181), .B(n80), .Y(n179) );
  NOR4XL U63 ( .A(sfraddr[5]), .B(sfraddr[4]), .C(sfraddr[3]), .D(n34), .Y(
        n101) );
  INVX1 U64 ( .A(sfraddr[4]), .Y(n5) );
  INVX1 U65 ( .A(sfraddr[3]), .Y(n4) );
  INVX1 U66 ( .A(sfrdatai[5]), .Y(n12) );
  INVX1 U67 ( .A(sfrdatai[3]), .Y(n10) );
  INVX1 U68 ( .A(sfrdatai[4]), .Y(n11) );
  INVX1 U69 ( .A(sfrdatai[2]), .Y(n9) );
  INVX1 U70 ( .A(sfrdatai[6]), .Y(n13) );
  INVX1 U71 ( .A(sfrdatai[7]), .Y(n14) );
  INVX1 U72 ( .A(sfrdatai[0]), .Y(n7) );
  INVX1 U73 ( .A(sfrdatai[1]), .Y(n8) );
  INVX1 U74 ( .A(n3), .Y(n225) );
  NAND2X1 U75 ( .A(n145), .B(n3), .Y(n130) );
  NAND32X1 U76 ( .B(n114), .C(n23), .A(n145), .Y(n153) );
  NOR21XL U77 ( .B(t1ov), .A(n19), .Y(N59) );
  OAI211X1 U78 ( .C(n59), .D(n153), .A(n129), .B(n24), .Y(N471) );
  INVX1 U79 ( .A(rst), .Y(n25) );
  NOR3XL U80 ( .A(n120), .B(n22), .C(n3), .Y(n166) );
  INVX1 U81 ( .A(rst), .Y(n24) );
  INVX1 U82 ( .A(rst), .Y(n26) );
  NOR2X1 U83 ( .A(n21), .B(n114), .Y(n134) );
  INVX1 U84 ( .A(n140), .Y(n54) );
  NAND3X1 U85 ( .A(n114), .B(n16), .C(n76), .Y(n129) );
  NOR2X1 U86 ( .A(n22), .B(newinstr), .Y(n104) );
  NAND2X1 U87 ( .A(n227), .B(n226), .Y(n80) );
  NOR2X1 U88 ( .A(n80), .B(n220), .Y(rxd0oe) );
  NOR32XL U89 ( .B(r_shift_clk), .C(n224), .A(n138), .Y(n145) );
  AOI21X1 U90 ( .B(n77), .C(n196), .A(N224), .Y(n199) );
  INVX1 U91 ( .A(n117), .Y(n66) );
  NOR3XL U92 ( .A(n115), .B(n117), .C(n216), .Y(r_shift_clk) );
  INVX1 U93 ( .A(n196), .Y(n65) );
  OAI22X1 U94 ( .A(n153), .B(n47), .C(n129), .D(n46), .Y(N473) );
  OAI22X1 U95 ( .A(n153), .B(n45), .C(n129), .D(n44), .Y(N475) );
  OAI22X1 U96 ( .A(n153), .B(n42), .C(n129), .D(n41), .Y(N478) );
  OAI22X1 U97 ( .A(n153), .B(n44), .C(n129), .D(n43), .Y(N476) );
  OAI22X1 U98 ( .A(n153), .B(n43), .C(n129), .D(n42), .Y(N477) );
  OAI22X1 U99 ( .A(n153), .B(n46), .C(n129), .D(n45), .Y(N474) );
  OAI22X1 U100 ( .A(n153), .B(n41), .C(n60), .D(n129), .Y(N479) );
  AOI211X1 U101 ( .C(n79), .D(n77), .A(n65), .B(n78), .Y(N225) );
  OAI21X1 U102 ( .B(n216), .C(n108), .A(n109), .Y(n240) );
  OAI211X1 U103 ( .C(n110), .D(n111), .A(n108), .B(n24), .Y(n109) );
  NAND32X1 U104 ( .B(n110), .C(n23), .A(n112), .Y(n108) );
  AND3X1 U105 ( .A(n225), .B(n120), .C(n216), .Y(n110) );
  NAND2X1 U106 ( .A(n154), .B(n81), .Y(N428) );
  OAI21X1 U107 ( .B(n61), .C(n126), .A(n18), .Y(n204) );
  NAND21X1 U108 ( .B(n204), .A(n126), .Y(n205) );
  INVX1 U109 ( .A(n138), .Y(n76) );
  AOI22AXL U110 ( .A(n225), .B(n120), .D(n159), .C(n3), .Y(n154) );
  NAND2X1 U111 ( .A(n55), .B(n117), .Y(n140) );
  OAI21AX1 U112 ( .B(n166), .C(n159), .A(n164), .Y(n162) );
  OAI32X1 U113 ( .A(n62), .B(n126), .C(n204), .D(n61), .E(n205), .Y(N188) );
  NOR2X1 U114 ( .A(n156), .B(n80), .Y(n114) );
  NOR3XL U115 ( .A(n52), .B(n156), .C(n223), .Y(n120) );
  OAI21X1 U116 ( .B(n117), .C(n228), .A(n18), .Y(N325) );
  AOI211X1 U117 ( .C(n152), .D(n217), .A(n169), .B(n170), .Y(N363) );
  NOR2X1 U118 ( .A(n220), .B(n156), .Y(t_shift_clk) );
  INVX1 U119 ( .A(n139), .Y(n55) );
  INVX1 U120 ( .A(n81), .Y(n27) );
  NAND2X1 U121 ( .A(n25), .B(n200), .Y(N223) );
  NAND3X1 U122 ( .A(n16), .B(n63), .C(n169), .Y(N360) );
  NOR43XL U123 ( .B(n62), .C(n56), .D(N190), .A(n61), .Y(N191) );
  NAND32X1 U124 ( .B(n1), .C(n2), .A(n15), .Y(N166) );
  AOI21AX1 U125 ( .B(n220), .C(n216), .A(n24), .Y(n122) );
  AOI211X1 U126 ( .C(n58), .D(n56), .A(n204), .B(n57), .Y(N186) );
  INVX1 U127 ( .A(n126), .Y(n57) );
  NOR3XL U128 ( .A(n97), .B(n22), .C(n40), .Y(N207) );
  NOR2X1 U129 ( .A(n58), .B(n20), .Y(N190) );
  NOR2X1 U130 ( .A(n224), .B(n20), .Y(N348) );
  NAND2X1 U131 ( .A(n60), .B(n15), .Y(N382) );
  NOR2X1 U132 ( .A(n22), .B(n96), .Y(n245) );
  XNOR2XL U133 ( .A(n40), .B(n97), .Y(n96) );
  NAND3X1 U134 ( .A(n225), .B(n39), .C(n122), .Y(N303) );
  NAND2X1 U135 ( .A(n26), .B(n117), .Y(N324) );
  INVX1 U136 ( .A(n198), .Y(n78) );
  NOR3XL U137 ( .A(n208), .B(n22), .C(n203), .Y(N142) );
  NOR2X1 U138 ( .A(n152), .B(n217), .Y(n170) );
  NAND2X1 U139 ( .A(n24), .B(n46), .Y(N376) );
  NAND2X1 U140 ( .A(n26), .B(n45), .Y(N377) );
  NAND2X1 U141 ( .A(n26), .B(n44), .Y(N378) );
  NAND2X1 U142 ( .A(n26), .B(n43), .Y(N379) );
  NAND2X1 U143 ( .A(n26), .B(n42), .Y(N380) );
  NAND2X1 U144 ( .A(n26), .B(n41), .Y(N381) );
  NAND2X1 U145 ( .A(n26), .B(n47), .Y(N375) );
  NOR2X1 U146 ( .A(n22), .B(n228), .Y(N307) );
  INVX1 U147 ( .A(n143), .Y(n59) );
  AO222X1 U148 ( .A(sfrdatai[1]), .B(n31), .C(n107), .D(ti_tmp), .E(s0con[1]), 
        .F(n32), .Y(n241) );
  OAI211X1 U149 ( .C(n7), .D(n179), .A(n18), .B(n191), .Y(N260) );
  AOI22X1 U150 ( .A(n36), .B(sfrdatai[1]), .C(t_shift_reg[3]), .D(n38), .Y(
        n191) );
  OAI211X1 U151 ( .C(n8), .D(n179), .A(n17), .B(n190), .Y(N261) );
  AOI22X1 U152 ( .A(n36), .B(sfrdatai[2]), .C(t_shift_reg[4]), .D(n38), .Y(
        n190) );
  OAI211X1 U153 ( .C(n179), .D(n12), .A(n17), .B(n186), .Y(N265) );
  AOI22X1 U154 ( .A(n36), .B(sfrdatai[6]), .C(t_shift_reg[8]), .D(n38), .Y(
        n186) );
  OAI211X1 U155 ( .C(n9), .D(n179), .A(n18), .B(n189), .Y(N262) );
  AOI22X1 U156 ( .A(sfrdatai[3]), .B(n36), .C(t_shift_reg[5]), .D(n38), .Y(
        n189) );
  OAI211X1 U157 ( .C(n179), .D(n10), .A(n17), .B(n188), .Y(N263) );
  AOI22X1 U158 ( .A(sfrdatai[4]), .B(n36), .C(t_shift_reg[6]), .D(n38), .Y(
        n188) );
  OAI211X1 U159 ( .C(n179), .D(n11), .A(n17), .B(n187), .Y(N264) );
  AOI22X1 U160 ( .A(sfrdatai[5]), .B(n36), .C(t_shift_reg[7]), .D(n38), .Y(
        n187) );
  OAI211X1 U161 ( .C(n179), .D(n13), .A(n17), .B(n185), .Y(N266) );
  AOI22X1 U162 ( .A(n36), .B(sfrdatai[7]), .C(t_shift_reg[9]), .D(n38), .Y(
        n185) );
  AO222X1 U163 ( .A(n131), .B(N348), .C(n107), .D(ri_tmp), .E(n31), .F(
        sfrdatai[0]), .Y(n237) );
  GEN2XL U164 ( .D(t_shift_count[1]), .E(t_shift_count[0]), .C(n178), .B(n38), 
        .A(n37), .Y(N282) );
  INVX1 U165 ( .A(n179), .Y(n37) );
  NAND3X1 U166 ( .A(n176), .B(n17), .C(n182), .Y(N268) );
  OAI21X1 U167 ( .B(s0con[3]), .C(n227), .A(n181), .Y(n182) );
  OAI21X1 U168 ( .B(n131), .C(n9), .A(n147), .Y(n230) );
  AOI33X1 U169 ( .A(s0con2_tmp), .B(n107), .C(s0con2_val), .D(n32), .E(n50), 
        .F(s0con[2]), .Y(n147) );
  INVX1 U170 ( .A(s0con2_tmp), .Y(n50) );
  OAI21X1 U171 ( .B(t_shift_count[0]), .C(n176), .A(n180), .Y(N281) );
  OAI21X1 U172 ( .B(s0con[7]), .C(n226), .A(n181), .Y(n180) );
  OAI21X1 U173 ( .B(n175), .C(n176), .A(n35), .Y(N284) );
  XOR2X1 U174 ( .A(n103), .B(t_shift_count[3]), .Y(n175) );
  NAND3X1 U175 ( .A(n183), .B(n16), .C(n184), .Y(N267) );
  AOI22X1 U176 ( .A(t_shift_reg[10]), .B(n38), .C(n181), .D(sfrdatai[7]), .Y(
        n184) );
  OAI2B11X1 U177 ( .D(t_shift_reg[1]), .C(n176), .A(n35), .B(n17), .Y(N258) );
  OAI211X1 U178 ( .C(n7), .D(n183), .A(n17), .B(n192), .Y(N259) );
  NAND2X1 U179 ( .A(t_shift_reg[2]), .B(n38), .Y(n192) );
  INVX1 U180 ( .A(n98), .Y(n28) );
  AOI32X1 U181 ( .A(smod), .B(n16), .C(n99), .D(sfrdatai[7]), .E(n30), .Y(n98)
         );
  INVX1 U182 ( .A(n99), .Y(n30) );
  NAND4X1 U183 ( .A(sfraddr[0]), .B(n100), .C(sfraddr[2]), .D(n101), .Y(n99)
         );
  INVX1 U184 ( .A(n92), .Y(n29) );
  AOI32X1 U185 ( .A(bd), .B(n16), .C(n93), .D(n33), .E(sfrdatai[7]), .Y(n92)
         );
  INVX1 U186 ( .A(n93), .Y(n33) );
  NAND4X1 U187 ( .A(sfraddr[6]), .B(n94), .C(n95), .D(n15), .Y(n93) );
  AOI21X1 U188 ( .B(n103), .C(n177), .A(n176), .Y(N283) );
  NAND21X1 U189 ( .B(n178), .A(t_shift_count[2]), .Y(n177) );
  NAND2X1 U190 ( .A(n35), .B(n102), .Y(n243) );
  OAI211X1 U191 ( .C(t_shift_count[3]), .D(n103), .A(n17), .B(t_start), .Y(
        n102) );
  ENOX1 U192 ( .A(n127), .B(n142), .C(n142), .D(s0con2_tmp), .Y(n232) );
  ENOX1 U193 ( .A(n127), .B(n143), .C(n130), .D(n104), .Y(n142) );
  OAI211X1 U194 ( .C(n59), .D(n127), .A(n128), .B(n129), .Y(n238) );
  NAND3X1 U195 ( .A(n104), .B(n130), .C(ri_tmp), .Y(n128) );
  OAI21BBX1 U196 ( .A(n104), .B(ti_tmp), .C(n105), .Y(n242) );
  NAND4X1 U197 ( .A(t_shift_clk), .B(n16), .C(t_shift_count[0]), .D(n106), .Y(
        n105) );
  NOR3XL U198 ( .A(t_shift_count[1]), .B(t_shift_count[3]), .C(
        t_shift_count[2]), .Y(n106) );
  INVX1 U199 ( .A(s0con[6]), .Y(n226) );
  INVX1 U200 ( .A(s0con[7]), .Y(n227) );
  INVX1 U201 ( .A(t_start), .Y(n220) );
  ENOX1 U202 ( .A(smod), .B(baud_r2_clk), .C(n97), .D(smod), .Y(n117) );
  AOI31X1 U203 ( .A(t_baud_count[2]), .B(s0relh[6]), .C(n78), .D(n200), .Y(
        n196) );
  OAI32X1 U204 ( .A(n65), .B(t_baud_count[2]), .C(n198), .D(n199), .E(n215), 
        .Y(N226) );
  OAI32X1 U205 ( .A(n49), .B(n23), .C(n144), .D(n60), .E(n127), .Y(n231) );
  INVX1 U206 ( .A(s0con2_val), .Y(n49) );
  NOR4XL U207 ( .A(n146), .B(n138), .C(n115), .D(n216), .Y(n144) );
  NAND3X1 U208 ( .A(n3), .B(n224), .C(n143), .Y(n146) );
  OAI22AX1 U209 ( .D(n201), .C(t1ov_ff), .A(n202), .B(n201), .Y(n97) );
  NOR2X1 U210 ( .A(n226), .B(bd), .Y(n201) );
  AOI221XL U211 ( .A(s0con[6]), .B(n219), .C(n203), .D(n226), .E(n225), .Y(
        n202) );
  NAND3X1 U212 ( .A(t_start), .B(n16), .C(n66), .Y(n200) );
  NOR2X1 U213 ( .A(s0relh[7]), .B(r_clk_ov2), .Y(n203) );
  NOR2X1 U214 ( .A(n65), .B(t_baud_count[0]), .Y(N224) );
  GEN2XL U215 ( .D(n196), .E(n215), .C(n64), .B(t_baud_count[3]), .A(n197), 
        .Y(N227) );
  NOR4XL U216 ( .A(t_baud_count[3]), .B(n198), .C(n215), .D(n65), .Y(n197) );
  INVX1 U217 ( .A(n199), .Y(n64) );
  AOI22X1 U218 ( .A(n113), .B(n80), .C(n76), .D(n114), .Y(n112) );
  OAI32X1 U219 ( .A(n115), .B(n116), .C(n117), .D(n223), .E(n118), .Y(n113) );
  AOI21X1 U220 ( .B(rxd0_val), .C(n119), .A(n76), .Y(n116) );
  OAI22AX1 U221 ( .D(r_shift_reg[0]), .C(n153), .A(n129), .B(n47), .Y(N472) );
  INVX1 U222 ( .A(baud_rate_ov), .Y(n219) );
  NAND43X1 U223 ( .B(r_shift_count[3]), .C(r_shift_count[1]), .D(
        r_shift_count[2]), .A(r_shift_count[0]), .Y(n138) );
  AOI22X1 U224 ( .A(n221), .B(n219), .C(n208), .D(s0relh[7]), .Y(n83) );
  AOI21X1 U225 ( .B(n221), .C(r_clk_ov2), .A(n83), .Y(n84) );
  GEN2XL U226 ( .D(n55), .E(n48), .C(n54), .B(fluctuation_conter[1]), .A(n141), 
        .Y(n233) );
  NOR4XL U227 ( .A(fluctuation_conter[1]), .B(n54), .C(n139), .D(n48), .Y(n141) );
  INVX1 U228 ( .A(n85), .Y(n74) );
  AOI221XL U229 ( .A(s0relh[0]), .B(n83), .C(N153), .D(n84), .E(n21), .Y(n85)
         );
  NAND21X1 U230 ( .B(r_shift_count[2]), .A(n163), .Y(n160) );
  OAI22X1 U231 ( .A(t_baud_ov), .B(n225), .C(clk_ov12), .D(n80), .Y(n156) );
  NAND2X1 U232 ( .A(rxd0_fall_fl), .B(n15), .Y(n139) );
  NOR42XL U233 ( .C(r_shift_count[3]), .D(r_shift_count[1]), .A(
        r_shift_count[0]), .B(r_shift_count[2]), .Y(n119) );
  OAI32X1 U234 ( .A(n204), .B(clk_count[2]), .C(n126), .D(n62), .E(n205), .Y(
        N187) );
  OAI32X1 U235 ( .A(n139), .B(fluctuation_conter[0]), .C(n54), .D(n140), .E(
        n48), .Y(n234) );
  OAI32X1 U236 ( .A(n48), .B(n63), .C(n139), .D(r_baud_count[0]), .E(n169), 
        .Y(N361) );
  OAI32X1 U237 ( .A(n51), .B(n63), .C(n139), .D(n171), .E(n169), .Y(N362) );
  INVX1 U238 ( .A(fluctuation_conter[1]), .Y(n51) );
  AOI21X1 U239 ( .B(r_baud_count[1]), .C(n218), .A(n151), .Y(n171) );
  OAI32X1 U240 ( .A(n159), .B(n22), .C(n225), .D(n164), .E(n165), .Y(N425) );
  AOI21X1 U241 ( .B(r_shift_count[0]), .C(r_shift_count[1]), .A(n163), .Y(n165) );
  NAND4X1 U242 ( .A(r_start), .B(n66), .C(n15), .D(n63), .Y(n169) );
  NOR2X1 U243 ( .A(r_shift_count[0]), .B(r_shift_count[1]), .Y(n163) );
  NAND41X1 U244 ( .D(n209), .A(n210), .B(tim_baud[8]), .C(tim_baud[9]), .Y(
        n208) );
  NAND3X1 U245 ( .A(tim_baud[6]), .B(tim_baud[5]), .C(tim_baud[7]), .Y(n209)
         );
  NOR32XL U246 ( .B(tim_baud[4]), .C(tim_baud[3]), .A(n211), .Y(n210) );
  NAND3X1 U247 ( .A(tim_baud[1]), .B(tim_baud[0]), .C(tim_baud[2]), .Y(n211)
         );
  INVX1 U248 ( .A(r_baud_count[2]), .Y(n217) );
  NOR4XL U249 ( .A(rxd0_fall), .B(receive_11_bits), .C(r_start), .D(n174), .Y(
        N306) );
  AOI31X1 U250 ( .A(n16), .B(n228), .C(rxd0_ff), .D(n55), .Y(n174) );
  NOR2X1 U251 ( .A(n218), .B(r_baud_count[1]), .Y(n151) );
  NOR2X1 U252 ( .A(n160), .B(r_shift_count[3]), .Y(n111) );
  OAI21X1 U253 ( .B(N382), .C(n157), .A(n158), .Y(N427) );
  GEN2XL U254 ( .D(n119), .E(n80), .C(n157), .B(n154), .A(n23), .Y(n158) );
  AOI21X1 U255 ( .B(n160), .C(r_shift_count[3]), .A(n111), .Y(n157) );
  OAI21X1 U256 ( .B(n52), .C(n132), .A(n133), .Y(n236) );
  NAND4X1 U257 ( .A(ri0_ff), .B(n132), .C(n15), .D(n224), .Y(n133) );
  OAI31XL U258 ( .A(n53), .B(s0con[0]), .C(n80), .D(n134), .Y(n132) );
  INVX1 U259 ( .A(ri0_ff), .Y(n53) );
  AOI221XL U260 ( .A(s0relh[6]), .B(n217), .C(n75), .D(n222), .E(n135), .Y(
        n235) );
  AOI22X1 U261 ( .A(n136), .B(n137), .C(n55), .D(n118), .Y(n135) );
  NOR32XL U262 ( .B(rxd0_ff), .C(s0con[6]), .A(n138), .Y(n136) );
  NOR3XL U263 ( .A(n22), .B(s0con[7]), .C(rxd0ff), .Y(n137) );
  NAND2X1 U264 ( .A(n151), .B(n155), .Y(n115) );
  OAI32X1 U265 ( .A(n75), .B(s0relh[6]), .C(r_baud_count[2]), .D(n217), .E(
        n222), .Y(n155) );
  NOR4XL U266 ( .A(n195), .B(n79), .C(n19), .D(n117), .Y(N230) );
  NAND32X1 U267 ( .B(t_baud_count[3]), .C(t_baud_count[2]), .A(n77), .Y(n195)
         );
  AOI21X1 U268 ( .B(n160), .C(n161), .A(n162), .Y(N426) );
  NAND21X1 U269 ( .B(n163), .A(r_shift_count[2]), .Y(n161) );
  INVX1 U270 ( .A(s0relh[6]), .Y(n222) );
  OAI21BBX1 U271 ( .A(n66), .B(rxd0_vec[0]), .C(n24), .Y(N326) );
  OAI21BBX1 U272 ( .A(n66), .B(rxd0_vec[1]), .C(n24), .Y(N327) );
  NOR2X1 U273 ( .A(n167), .B(n166), .Y(n164) );
  AOI211X1 U274 ( .C(n119), .D(rxd0_val), .A(n225), .B(n23), .Y(n167) );
  NAND2X1 U275 ( .A(rxd0_fall), .B(n111), .Y(n118) );
  INVX1 U276 ( .A(r_baud_count[0]), .Y(n218) );
  INVX1 U277 ( .A(r_baud_count[3]), .Y(n75) );
  NOR2X1 U278 ( .A(n168), .B(n169), .Y(N364) );
  XNOR2XL U279 ( .A(r_baud_count[3]), .B(n170), .Y(n168) );
  NOR2X1 U280 ( .A(n22), .B(n207), .Y(N169) );
  AOI22X1 U281 ( .A(N147), .B(n84), .C(s0rell[2]), .D(n2), .Y(n207) );
  NOR2X1 U282 ( .A(n20), .B(n206), .Y(N170) );
  AOI22X1 U283 ( .A(N148), .B(n1), .C(s0rell[3]), .D(n2), .Y(n206) );
  NOR2X1 U284 ( .A(r_shift_count[0]), .B(n162), .Y(N424) );
  INVX1 U285 ( .A(n87), .Y(n72) );
  AOI221XL U286 ( .A(s0rell[6]), .B(n83), .C(N151), .D(n84), .E(n23), .Y(n87)
         );
  INVX1 U287 ( .A(n90), .Y(n69) );
  AOI221XL U288 ( .A(s0rell[1]), .B(n83), .C(N146), .D(n84), .E(n23), .Y(n90)
         );
  INVX1 U289 ( .A(n88), .Y(n71) );
  AOI221XL U290 ( .A(s0rell[5]), .B(n83), .C(N150), .D(n84), .E(n23), .Y(n88)
         );
  INVX1 U291 ( .A(n86), .Y(n73) );
  AOI221XL U292 ( .A(s0rell[7]), .B(n83), .C(N152), .D(n84), .E(n23), .Y(n86)
         );
  INVX1 U293 ( .A(n89), .Y(n70) );
  AOI221XL U294 ( .A(s0rell[4]), .B(n83), .C(N149), .D(n84), .E(n23), .Y(n89)
         );
  INVX1 U295 ( .A(n82), .Y(n67) );
  AOI221XL U296 ( .A(s0relh[1]), .B(n83), .C(N154), .D(n84), .E(n20), .Y(n82)
         );
  INVX1 U297 ( .A(n91), .Y(n68) );
  AOI221XL U298 ( .A(s0rell[0]), .B(n83), .C(N145), .D(n84), .E(n20), .Y(n91)
         );
  NAND2X1 U299 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n126) );
  NAND2X1 U300 ( .A(t_baud_count[1]), .B(t_baud_count[0]), .Y(n198) );
  NAND2X1 U301 ( .A(s0con[5]), .B(n60), .Y(n143) );
  NOR31X1 U302 ( .C(t_shift_count[0]), .A(t_shift_count[2]), .B(
        t_shift_count[1]), .Y(n125) );
  OAI21X1 U303 ( .B(n80), .C(n228), .A(n172), .Y(N333) );
  AOI21X1 U304 ( .B(n173), .C(n3), .A(n20), .Y(n172) );
  AND2X1 U305 ( .A(n148), .B(s0con[7]), .Y(n229) );
  OAI33XL U306 ( .A(n149), .B(n19), .C(n150), .D(n138), .E(n20), .F(n115), .Y(
        n148) );
  OAI31XL U307 ( .A(n152), .B(r_baud_count[2]), .C(n222), .D(receive_11_bits), 
        .Y(n149) );
  NOR43XL U308 ( .B(n222), .C(n75), .D(n151), .A(n217), .Y(n150) );
  INVX1 U309 ( .A(s0con[0]), .Y(n224) );
  INVX1 U310 ( .A(r_start), .Y(n216) );
  INVX1 U311 ( .A(rxd0_val), .Y(n60) );
  OAI211X1 U312 ( .C(n225), .D(n39), .A(n121), .B(n122), .Y(n239) );
  OAI21BBX1 U313 ( .A(n123), .B(n124), .C(n225), .Y(n121) );
  OAI31XL U314 ( .A(clk_count[0]), .B(clk_count[2]), .C(clk_count[1]), .D(
        clk_count[3]), .Y(n124) );
  AOI33X1 U315 ( .A(txd0), .B(t_shift_count[3]), .C(n125), .D(n62), .E(n61), 
        .F(n126), .Y(n123) );
  NAND2X1 U316 ( .A(rxd0_fall), .B(s0con[4]), .Y(n159) );
  INVX1 U317 ( .A(s0con[4]), .Y(n223) );
  NOR2X1 U318 ( .A(clk_count[0]), .B(n204), .Y(N185) );
  INVX1 U319 ( .A(s0relh[7]), .Y(n221) );
  INVX1 U320 ( .A(ri0_fall), .Y(n52) );
  NAND21X1 U321 ( .B(t_shift_count[2]), .A(n178), .Y(n103) );
  NOR2X1 U322 ( .A(t_shift_count[1]), .B(t_shift_count[0]), .Y(n178) );
  INVX1 U323 ( .A(rxd0_fall), .Y(n63) );
  INVX1 U324 ( .A(clk_count[3]), .Y(n61) );
  NAND2X1 U325 ( .A(r_baud_count[1]), .B(r_baud_count[0]), .Y(n152) );
  INVX1 U326 ( .A(t_baud_count[1]), .Y(n77) );
  INVX1 U327 ( .A(rxd0ff), .Y(n228) );
  INVX1 U328 ( .A(fluctuation_conter[0]), .Y(n48) );
  INVX1 U330 ( .A(clk_count[2]), .Y(n62) );
  INVX1 U331 ( .A(t_baud_count[2]), .Y(n215) );
  INVX1 U332 ( .A(clk_count[0]), .Y(n58) );
  INVX1 U333 ( .A(r_shift_reg[1]), .Y(n47) );
  INVX1 U334 ( .A(r_shift_reg[2]), .Y(n46) );
  INVX1 U335 ( .A(r_shift_reg[3]), .Y(n45) );
  INVX1 U336 ( .A(r_shift_reg[4]), .Y(n44) );
  INVX1 U337 ( .A(r_shift_reg[5]), .Y(n43) );
  INVX1 U338 ( .A(r_shift_reg[6]), .Y(n42) );
  INVX1 U339 ( .A(r_shift_reg[7]), .Y(n41) );
  INVX1 U340 ( .A(t_baud_count[0]), .Y(n79) );
  INVX1 U341 ( .A(clk_count[1]), .Y(n56) );
  INVX1 U342 ( .A(baud_r_count), .Y(n40) );
  INVX1 U343 ( .A(t_shift_reg[0]), .Y(n39) );
endmodule


module serial0_a0_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ports_a0 ( clkper, rst, port0, sfrdatai, sfraddr, sfrwe, test_si, 
        test_se );
  output [7:0] port0;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkper, rst, sfrwe, test_si, test_se;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, net12328, n2, n3, n4, n1;

  SNPS_CLOCK_GATE_HIGH_ports_a0 clk_gate_p0_reg ( .CLK(clkper), .EN(N2), 
        .ENCLK(net12328), .TE(test_se) );
  SDFFQX1 p0_reg_7_ ( .D(N10), .SIN(port0[6]), .SMC(test_se), .C(net12328), 
        .Q(port0[7]) );
  SDFFQX1 p0_reg_3_ ( .D(N6), .SIN(port0[2]), .SMC(test_se), .C(net12328), .Q(
        port0[3]) );
  SDFFQX1 p0_reg_1_ ( .D(N4), .SIN(port0[0]), .SMC(test_se), .C(net12328), .Q(
        port0[1]) );
  SDFFQX1 p0_reg_6_ ( .D(N9), .SIN(port0[5]), .SMC(test_se), .C(net12328), .Q(
        port0[6]) );
  SDFFQX1 p0_reg_5_ ( .D(N8), .SIN(port0[4]), .SMC(test_se), .C(net12328), .Q(
        port0[5]) );
  SDFFQX1 p0_reg_4_ ( .D(N7), .SIN(port0[3]), .SMC(test_se), .C(net12328), .Q(
        port0[4]) );
  SDFFQX1 p0_reg_2_ ( .D(N5), .SIN(port0[1]), .SMC(test_se), .C(net12328), .Q(
        port0[2]) );
  SDFFQX1 p0_reg_0_ ( .D(N3), .SIN(test_si), .SMC(test_se), .C(net12328), .Q(
        port0[0]) );
  NAND2X1 U2 ( .A(n1), .B(n2), .Y(N2) );
  NAND42XL U3 ( .C(sfraddr[3]), .D(sfraddr[2]), .A(n3), .B(n4), .Y(n2) );
  NOR3XL U4 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n3) );
  NOR42XL U5 ( .C(sfrwe), .D(n1), .A(sfraddr[1]), .B(sfraddr[0]), .Y(n4) );
  NOR21XL U6 ( .B(sfrdatai[0]), .A(n2), .Y(N3) );
  NOR21XL U7 ( .B(sfrdatai[3]), .A(n2), .Y(N6) );
  NOR21XL U8 ( .B(sfrdatai[1]), .A(n2), .Y(N4) );
  NOR21XL U9 ( .B(sfrdatai[4]), .A(n2), .Y(N7) );
  NOR21XL U10 ( .B(sfrdatai[5]), .A(n2), .Y(N8) );
  NOR21XL U11 ( .B(sfrdatai[6]), .A(n2), .Y(N9) );
  NOR21XL U12 ( .B(sfrdatai[7]), .A(n2), .Y(N10) );
  NOR21XL U13 ( .B(sfrdatai[2]), .A(n2), .Y(N5) );
  INVX1 U14 ( .A(rst), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ports_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mdu_a0 ( clkper, rst, mdubsy, sfrdatai, sfraddr, sfrwe, sfroe, arcon, 
        md0, md1, md2, md3, md4, md5, test_si, test_so, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] arcon;
  output [7:0] md0;
  output [7:0] md1;
  output [7:0] md2;
  output [7:0] md3;
  output [7:0] md4;
  output [7:0] md5;
  input clkper, rst, sfrwe, sfroe, test_si, test_se;
  output mdubsy, test_so;
  wire   N104, N105, N106, N107, N108, N109, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N332, N333, N334, N335, N336, N337, N338, N339, N340,
         N405, N406, N407, N408, N409, N410, N411, N412, N413, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N566, N567, N568, N569, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N610,
         N674, N675, N676, N677, N678, set_div16, set_div32, N802, N892, N893,
         N894, N895, net12346, net12352, net12357, net12362, net12367,
         net12372, net12377, n408, n409, n410, n411, n412, n413, n414, n137,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n1, n2, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n405, n406, n407, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2;
  wire   [3:0] oper_reg;
  wire   [4:1] counter_st;
  wire   [17:1] sum1;
  wire   [17:1] sum;
  wire   [15:0] norm_reg;
  wire   [1:0] mdu_op;
  wire   [17:1] arg_a;
  wire   [16:1] arg_b;
  wire   [17:0] arg_c;
  wire   [16:1] arg_d;

  SNPS_CLOCK_GATE_HIGH_mdu_a0_0 clk_gate_arcon_s_reg ( .CLK(clkper), .EN(N104), 
        .ENCLK(net12346), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_6 clk_gate_md0_s_reg ( .CLK(clkper), .EN(N190), 
        .ENCLK(net12352), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_5 clk_gate_md1_s_reg ( .CLK(clkper), .EN(N258), 
        .ENCLK(net12357), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_4 clk_gate_md2_s_reg ( .CLK(clkper), .EN(N332), 
        .ENCLK(net12362), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_3 clk_gate_md3_s_reg ( .CLK(clkper), .EN(N405), 
        .ENCLK(net12367), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_2 clk_gate_md4_s_reg ( .CLK(clkper), .EN(N453), 
        .ENCLK(net12372), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_1 clk_gate_md5_s_reg ( .CLK(clkper), .EN(N483), 
        .ENCLK(net12377), .TE(test_se) );
  mdu_a0_DW01_add_0 add_1040 ( .A(arg_c), .B({1'b0, arg_d, n404}), .CI(1'b0), 
        .SUM({sum, SYNOPSYS_UNCONNECTED_1}), .CO() );
  mdu_a0_DW01_add_1 add_961 ( .A({arg_a, n137}), .B({1'b0, arg_b, n404}), .CI(
        1'b0), .SUM({sum1, SYNOPSYS_UNCONNECTED_2}), .CO() );
  SDFFQX1 set_div16_reg ( .D(n414), .SIN(oper_reg[3]), .SMC(test_se), .C(
        clkper), .Q(set_div16) );
  SDFFQX1 setmdef_reg ( .D(N802), .SIN(set_div32), .SMC(test_se), .C(clkper), 
        .Q(test_so) );
  SDFFQX1 set_div32_reg ( .D(n413), .SIN(set_div16), .SMC(test_se), .C(clkper), 
        .Q(set_div32) );
  SDFFQX1 counter_st_reg_0_ ( .D(N674), .SIN(arcon[7]), .SMC(test_se), .C(
        clkper), .Q(N610) );
  SDFFQX1 counter_st_reg_1_ ( .D(N675), .SIN(N610), .SMC(test_se), .C(clkper), 
        .Q(counter_st[1]) );
  SDFFQX1 counter_st_reg_2_ ( .D(N676), .SIN(counter_st[1]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[2]) );
  SDFFQX1 counter_st_reg_4_ ( .D(N678), .SIN(counter_st[3]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[4]) );
  SDFFQX1 counter_st_reg_3_ ( .D(N677), .SIN(counter_st[2]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[3]) );
  SDFFQX1 oper_reg_reg_3_ ( .D(N895), .SIN(oper_reg[2]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[3]) );
  SDFFQX1 oper_reg_reg_0_ ( .D(N892), .SIN(norm_reg[15]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[0]) );
  SDFFQX1 oper_reg_reg_1_ ( .D(N893), .SIN(oper_reg[0]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[1]) );
  SDFFQX1 oper_reg_reg_2_ ( .D(N894), .SIN(oper_reg[1]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[2]) );
  SDFFQX1 norm_reg_reg_15_ ( .D(N581), .SIN(norm_reg[14]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[15]) );
  SDFFQX1 norm_reg_reg_14_ ( .D(N580), .SIN(norm_reg[13]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[14]) );
  SDFFQX1 norm_reg_reg_13_ ( .D(N579), .SIN(norm_reg[12]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[13]) );
  SDFFQX1 norm_reg_reg_12_ ( .D(N578), .SIN(norm_reg[11]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[12]) );
  SDFFQX1 norm_reg_reg_11_ ( .D(N577), .SIN(norm_reg[10]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[11]) );
  SDFFQX1 norm_reg_reg_10_ ( .D(N576), .SIN(norm_reg[9]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[10]) );
  SDFFQX1 norm_reg_reg_9_ ( .D(N575), .SIN(norm_reg[8]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[9]) );
  SDFFQX1 norm_reg_reg_8_ ( .D(N574), .SIN(norm_reg[7]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[8]) );
  SDFFQX1 norm_reg_reg_7_ ( .D(N573), .SIN(norm_reg[6]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[7]) );
  SDFFQX1 arcon_s_reg_6_ ( .D(n408), .SIN(arcon[5]), .SMC(test_se), .C(clkper), 
        .Q(arcon[6]) );
  SDFFQX1 arcon_s_reg_2_ ( .D(N107), .SIN(arcon[1]), .SMC(test_se), .C(
        net12346), .Q(arcon[2]) );
  SDFFQX1 arcon_s_reg_7_ ( .D(n410), .SIN(arcon[6]), .SMC(test_se), .C(clkper), 
        .Q(arcon[7]) );
  SDFFQX1 arcon_s_reg_3_ ( .D(N108), .SIN(arcon[2]), .SMC(test_se), .C(
        net12346), .Q(arcon[3]) );
  SDFFQX1 md1_s_reg_6_ ( .D(N265), .SIN(md1[5]), .SMC(test_se), .C(net12357), 
        .Q(md1[6]) );
  SDFFQX1 md1_s_reg_5_ ( .D(N264), .SIN(md1[4]), .SMC(test_se), .C(net12357), 
        .Q(md1[5]) );
  SDFFQX1 md0_s_reg_1_ ( .D(N192), .SIN(md0[0]), .SMC(test_se), .C(net12352), 
        .Q(md0[1]) );
  SDFFQX1 norm_reg_reg_6_ ( .D(N572), .SIN(norm_reg[5]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[6]) );
  SDFFQX1 arcon_s_reg_1_ ( .D(N106), .SIN(arcon[0]), .SMC(test_se), .C(
        net12346), .Q(arcon[1]) );
  SDFFQX1 md1_s_reg_4_ ( .D(N263), .SIN(md1[3]), .SMC(test_se), .C(net12357), 
        .Q(md1[4]) );
  SDFFQX1 md0_s_reg_6_ ( .D(N197), .SIN(md0[5]), .SMC(test_se), .C(net12352), 
        .Q(md0[6]) );
  SDFFQX1 md0_s_reg_7_ ( .D(N198), .SIN(md0[6]), .SMC(test_se), .C(net12352), 
        .Q(md0[7]) );
  SDFFQX1 md1_s_reg_1_ ( .D(N260), .SIN(md1[0]), .SMC(test_se), .C(net12357), 
        .Q(md1[1]) );
  SDFFQX1 md5_s_reg_3_ ( .D(N487), .SIN(md5[2]), .SMC(test_se), .C(net12377), 
        .Q(md5[3]) );
  SDFFQX1 md4_s_reg_7_ ( .D(N461), .SIN(md4[6]), .SMC(test_se), .C(net12372), 
        .Q(md4[7]) );
  SDFFQX1 md5_s_reg_2_ ( .D(N486), .SIN(md5[1]), .SMC(test_se), .C(net12377), 
        .Q(md5[2]) );
  SDFFQX1 md3_s_reg_6_ ( .D(N412), .SIN(md3[5]), .SMC(test_se), .C(net12367), 
        .Q(md3[6]) );
  SDFFQX1 md5_s_reg_1_ ( .D(N485), .SIN(md5[0]), .SMC(test_se), .C(net12377), 
        .Q(md5[1]) );
  SDFFQX1 arcon_s_reg_0_ ( .D(N105), .SIN(test_si), .SMC(test_se), .C(net12346), .Q(arcon[0]) );
  SDFFQX1 arcon_s_reg_4_ ( .D(N109), .SIN(arcon[3]), .SMC(test_se), .C(
        net12346), .Q(arcon[4]) );
  SDFFQX1 md0_s_reg_3_ ( .D(N194), .SIN(md0[2]), .SMC(test_se), .C(net12352), 
        .Q(md0[3]) );
  SDFFQX1 norm_reg_reg_5_ ( .D(N571), .SIN(norm_reg[4]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[5]) );
  SDFFQX1 norm_reg_reg_4_ ( .D(N570), .SIN(norm_reg[3]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[4]) );
  SDFFQX1 arcon_s_reg_5_ ( .D(n409), .SIN(arcon[4]), .SMC(test_se), .C(
        net12346), .Q(arcon[5]) );
  SDFFQX1 md2_s_reg_5_ ( .D(N338), .SIN(md2[4]), .SMC(test_se), .C(net12362), 
        .Q(md2[5]) );
  SDFFQX1 md0_s_reg_5_ ( .D(N196), .SIN(md0[4]), .SMC(test_se), .C(net12352), 
        .Q(md0[5]) );
  SDFFQX1 md5_s_reg_6_ ( .D(N490), .SIN(md5[5]), .SMC(test_se), .C(net12377), 
        .Q(md5[6]) );
  SDFFQX1 md5_s_reg_7_ ( .D(N491), .SIN(md5[6]), .SMC(test_se), .C(net12377), 
        .Q(md5[7]) );
  SDFFQX1 md1_s_reg_2_ ( .D(N261), .SIN(md1[1]), .SMC(test_se), .C(net12357), 
        .Q(md1[2]) );
  SDFFQX1 md1_s_reg_0_ ( .D(N259), .SIN(md0[7]), .SMC(test_se), .C(net12357), 
        .Q(md1[0]) );
  SDFFQX1 md1_s_reg_3_ ( .D(N262), .SIN(md1[2]), .SMC(test_se), .C(net12357), 
        .Q(md1[3]) );
  SDFFQX1 md5_s_reg_5_ ( .D(N489), .SIN(md5[4]), .SMC(test_se), .C(net12377), 
        .Q(md5[5]) );
  SDFFQX1 md0_s_reg_4_ ( .D(N195), .SIN(md0[3]), .SMC(test_se), .C(net12352), 
        .Q(md0[4]) );
  SDFFQX1 md5_s_reg_4_ ( .D(N488), .SIN(md5[3]), .SMC(test_se), .C(net12377), 
        .Q(md5[4]) );
  SDFFQX1 md3_s_reg_1_ ( .D(N407), .SIN(md3[0]), .SMC(test_se), .C(net12367), 
        .Q(md3[1]) );
  SDFFQX1 md4_s_reg_6_ ( .D(N460), .SIN(md4[5]), .SMC(test_se), .C(net12372), 
        .Q(md4[6]) );
  SDFFQX1 md2_s_reg_6_ ( .D(N339), .SIN(md2[5]), .SMC(test_se), .C(net12362), 
        .Q(md2[6]) );
  SDFFQX1 md2_s_reg_7_ ( .D(N340), .SIN(md2[6]), .SMC(test_se), .C(net12362), 
        .Q(md2[7]) );
  SDFFQX1 md3_s_reg_0_ ( .D(N406), .SIN(md2[7]), .SMC(test_se), .C(net12367), 
        .Q(md3[0]) );
  SDFFQX1 md3_s_reg_2_ ( .D(N408), .SIN(md3[1]), .SMC(test_se), .C(net12367), 
        .Q(md3[2]) );
  SDFFQX1 md3_s_reg_3_ ( .D(N409), .SIN(md3[2]), .SMC(test_se), .C(net12367), 
        .Q(md3[3]) );
  SDFFQX1 md5_s_reg_0_ ( .D(N484), .SIN(md4[7]), .SMC(test_se), .C(net12377), 
        .Q(md5[0]) );
  SDFFQX1 md0_s_reg_2_ ( .D(N193), .SIN(md0[1]), .SMC(test_se), .C(net12352), 
        .Q(md0[2]) );
  SDFFQX1 md3_s_reg_5_ ( .D(N411), .SIN(md3[4]), .SMC(test_se), .C(net12367), 
        .Q(md3[5]) );
  SDFFQX1 norm_reg_reg_3_ ( .D(N569), .SIN(norm_reg[2]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[3]) );
  SDFFQX1 md2_s_reg_4_ ( .D(N337), .SIN(md2[3]), .SMC(test_se), .C(net12362), 
        .Q(md2[4]) );
  SDFFQX1 md4_s_reg_5_ ( .D(N459), .SIN(md4[4]), .SMC(test_se), .C(net12372), 
        .Q(md4[5]) );
  SDFFQX1 md4_s_reg_4_ ( .D(N458), .SIN(md4[3]), .SMC(test_se), .C(net12372), 
        .Q(md4[4]) );
  SDFFQX1 md3_s_reg_4_ ( .D(N410), .SIN(md3[3]), .SMC(test_se), .C(net12367), 
        .Q(md3[4]) );
  SDFFQX1 norm_reg_reg_2_ ( .D(N568), .SIN(norm_reg[1]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[2]) );
  SDFFQX1 norm_reg_reg_1_ ( .D(N567), .SIN(norm_reg[0]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[1]) );
  SDFFQX1 md2_s_reg_3_ ( .D(N336), .SIN(md2[2]), .SMC(test_se), .C(net12362), 
        .Q(md2[3]) );
  SDFFQX1 md2_s_reg_2_ ( .D(N335), .SIN(md2[1]), .SMC(test_se), .C(net12362), 
        .Q(md2[2]) );
  SDFFQX1 md4_s_reg_2_ ( .D(N456), .SIN(md4[1]), .SMC(test_se), .C(net12372), 
        .Q(md4[2]) );
  SDFFQX1 md4_s_reg_3_ ( .D(N457), .SIN(md4[2]), .SMC(test_se), .C(net12372), 
        .Q(md4[3]) );
  SDFFQX1 norm_reg_reg_0_ ( .D(N566), .SIN(mdu_op[1]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[0]) );
  SDFFQX1 md2_s_reg_1_ ( .D(N334), .SIN(md2[0]), .SMC(test_se), .C(net12362), 
        .Q(md2[1]) );
  SDFFQX1 md4_s_reg_1_ ( .D(N455), .SIN(md4[0]), .SMC(test_se), .C(net12372), 
        .Q(md4[1]) );
  SDFFQX1 md0_s_reg_0_ ( .D(N191), .SIN(counter_st[4]), .SMC(test_se), .C(
        net12352), .Q(md0[0]) );
  SDFFQX1 md2_s_reg_0_ ( .D(N333), .SIN(md1[7]), .SMC(test_se), .C(net12362), 
        .Q(md2[0]) );
  SDFFQX1 md1_s_reg_7_ ( .D(N266), .SIN(md1[6]), .SMC(test_se), .C(net12357), 
        .Q(md1[7]) );
  SDFFQX1 md4_s_reg_0_ ( .D(N454), .SIN(md3[7]), .SMC(test_se), .C(net12372), 
        .Q(md4[0]) );
  SDFFQX1 md3_s_reg_7_ ( .D(N413), .SIN(md3[6]), .SMC(test_se), .C(net12367), 
        .Q(md3[7]) );
  SDFFQX1 mdu_op_reg_0_ ( .D(n411), .SIN(md5[7]), .SMC(test_se), .C(clkper), 
        .Q(mdu_op[0]) );
  SDFFQX1 mdu_op_reg_1_ ( .D(n412), .SIN(mdu_op[0]), .SMC(test_se), .C(clkper), 
        .Q(mdu_op[1]) );
  NAND41XL U5 ( .D(sfraddr[4]), .A(sfraddr[5]), .B(sfraddr[3]), .C(sfraddr[6]), 
        .Y(n243) );
  NAND2X1 U6 ( .A(n242), .B(n271), .Y(n1) );
  NAND2X1 U7 ( .A(n271), .B(n55), .Y(n2) );
  INVX1 U8 ( .A(n298), .Y(n5) );
  INVX1 U9 ( .A(n50), .Y(n6) );
  INVX1 U10 ( .A(n65), .Y(n7) );
  NAND2X1 U11 ( .A(n106), .B(arg_c[0]), .Y(n8) );
  NAND2X1 U12 ( .A(n27), .B(n260), .Y(n9) );
  INVX1 U13 ( .A(n66), .Y(n10) );
  INVX1 U14 ( .A(n22), .Y(n11) );
  NAND2X1 U15 ( .A(n259), .B(n260), .Y(n12) );
  BUFX3 U16 ( .A(n188), .Y(n13) );
  NOR2X1 U17 ( .A(sum1[17]), .B(n26), .Y(n14) );
  INVX1 U18 ( .A(n64), .Y(n15) );
  BUFX3 U19 ( .A(n254), .Y(n16) );
  NAND2X1 U20 ( .A(sum1[17]), .B(arg_c[0]), .Y(n17) );
  BUFX3 U21 ( .A(n194), .Y(n18) );
  INVX1 U22 ( .A(n75), .Y(n19) );
  NOR2X1 U23 ( .A(n106), .B(n26), .Y(n20) );
  INVX1 U24 ( .A(n49), .Y(n21) );
  BUFX3 U25 ( .A(n294), .Y(n22) );
  NOR2X1 U26 ( .A(n376), .B(n67), .Y(n23) );
  INVX1 U27 ( .A(n137), .Y(n24) );
  INVX1 U28 ( .A(sum[17]), .Y(n25) );
  INVX1 U29 ( .A(n25), .Y(n26) );
  INVX1 U30 ( .A(n25), .Y(n27) );
  NOR4XL U31 ( .A(n252), .B(n84), .C(n86), .D(n85), .Y(n380) );
  INVX1 U32 ( .A(n168), .Y(n49) );
  NAND2X1 U33 ( .A(n52), .B(n271), .Y(n166) );
  NAND2X1 U34 ( .A(n54), .B(n271), .Y(n168) );
  NAND2X1 U35 ( .A(n271), .B(n55), .Y(n162) );
  NAND2X1 U36 ( .A(n271), .B(n53), .Y(n237) );
  INVX1 U37 ( .A(n352), .Y(n53) );
  INVX1 U38 ( .A(n328), .Y(n55) );
  INVX1 U39 ( .A(n336), .Y(n76) );
  INVX1 U40 ( .A(n369), .Y(n78) );
  INVX1 U41 ( .A(n342), .Y(n66) );
  INVX1 U42 ( .A(n32), .Y(n30) );
  INVX1 U43 ( .A(n404), .Y(n35) );
  INVX1 U44 ( .A(n32), .Y(n31) );
  INVX1 U45 ( .A(n404), .Y(n34) );
  NOR2X1 U46 ( .A(n51), .B(n46), .Y(n271) );
  OAI21AX1 U47 ( .B(n164), .C(n228), .A(n229), .Y(n197) );
  NAND2X1 U48 ( .A(n242), .B(n271), .Y(n161) );
  NAND3X1 U49 ( .A(n272), .B(n37), .C(sfraddr[0]), .Y(n328) );
  NAND3X1 U50 ( .A(n36), .B(n37), .C(n272), .Y(n352) );
  NAND2X1 U51 ( .A(n165), .B(n271), .Y(n355) );
  OR2X1 U52 ( .A(n240), .B(n46), .Y(n159) );
  INVX1 U53 ( .A(n228), .Y(n54) );
  INVX1 U54 ( .A(n244), .Y(n52) );
  NAND2X1 U55 ( .A(n311), .B(n161), .Y(N405) );
  NAND2X1 U56 ( .A(n311), .B(n162), .Y(N332) );
  INVX1 U57 ( .A(n374), .Y(n77) );
  NOR2X1 U58 ( .A(n23), .B(n76), .Y(n342) );
  NAND2X1 U59 ( .A(n80), .B(n374), .Y(n369) );
  NAND2X1 U60 ( .A(n80), .B(n77), .Y(n336) );
  NAND2X1 U61 ( .A(n259), .B(n260), .Y(n253) );
  INVX1 U62 ( .A(n404), .Y(n33) );
  INVX1 U63 ( .A(n440), .Y(n32) );
  NAND42X1 U64 ( .C(n243), .D(sfraddr[1]), .A(sfraddr[0]), .B(n285), .Y(n240)
         );
  NOR2X1 U65 ( .A(n37), .B(n51), .Y(n285) );
  OAI21X1 U66 ( .B(n164), .C(n352), .A(n48), .Y(n158) );
  OAI21X1 U67 ( .B(n164), .C(n244), .A(n48), .Y(n229) );
  OAI21BX1 U68 ( .C(n242), .B(n164), .A(n48), .Y(n288) );
  OAI21BX1 U69 ( .C(n165), .B(n164), .A(n48), .Y(n357) );
  OAI21X1 U70 ( .B(n164), .C(n328), .A(n48), .Y(n313) );
  AOI21AX1 U71 ( .B(sfrwe), .C(n54), .A(n47), .Y(n403) );
  NAND3X1 U72 ( .A(n272), .B(n36), .C(sfraddr[2]), .Y(n244) );
  NOR4XL U73 ( .A(n36), .B(n243), .C(sfraddr[1]), .D(sfraddr[2]), .Y(n165) );
  NAND3X1 U74 ( .A(sfraddr[0]), .B(n272), .C(sfraddr[2]), .Y(n228) );
  NOR2X1 U75 ( .A(n46), .B(sfrwe), .Y(n164) );
  NOR4XL U76 ( .A(n37), .B(n243), .C(sfraddr[0]), .D(sfraddr[1]), .Y(n242) );
  OAI31XL U77 ( .A(n36), .B(sfraddr[1]), .C(n243), .D(n244), .Y(n241) );
  NAND2X1 U78 ( .A(n240), .B(n48), .Y(n274) );
  NAND2X1 U79 ( .A(n403), .B(n84), .Y(n379) );
  INVX1 U80 ( .A(sfraddr[2]), .Y(n37) );
  OAI31XL U81 ( .A(n52), .B(n54), .C(n165), .D(sfrwe), .Y(n239) );
  INVX1 U82 ( .A(sfrwe), .Y(n51) );
  NAND3X1 U83 ( .A(n74), .B(n48), .C(n159), .Y(N453) );
  NOR21XL U84 ( .B(sfraddr[1]), .A(n243), .Y(n272) );
  INVX1 U85 ( .A(sfraddr[0]), .Y(n36) );
  NAND2X1 U86 ( .A(n354), .B(n355), .Y(N190) );
  NAND2X1 U87 ( .A(n354), .B(n237), .Y(N258) );
  NAND3X1 U88 ( .A(n74), .B(n47), .C(n6), .Y(N483) );
  NOR2X1 U89 ( .A(n376), .B(n67), .Y(n299) );
  NAND2X1 U90 ( .A(n81), .B(n79), .Y(n374) );
  NAND2X1 U91 ( .A(n77), .B(n262), .Y(n376) );
  NAND2X1 U92 ( .A(n330), .B(n331), .Y(n289) );
  OR2X1 U93 ( .A(n375), .B(n67), .Y(n331) );
  INVX1 U94 ( .A(n262), .Y(n80) );
  INVX1 U95 ( .A(n372), .Y(n71) );
  NOR3XL U96 ( .A(n81), .B(n46), .C(n262), .Y(n260) );
  INVX1 U97 ( .A(n298), .Y(n68) );
  NOR32XL U98 ( .B(n330), .C(n332), .A(n76), .Y(n311) );
  NOR43XL U99 ( .B(n291), .C(n375), .D(n376), .A(n46), .Y(n332) );
  INVX1 U100 ( .A(n380), .Y(n83) );
  INVX1 U101 ( .A(n47), .Y(n46) );
  INVX1 U102 ( .A(n286), .Y(n74) );
  NOR2X1 U103 ( .A(n106), .B(n26), .Y(n259) );
  NAND2X1 U104 ( .A(n27), .B(n260), .Y(n255) );
  NAND2X1 U105 ( .A(n261), .B(n260), .Y(n254) );
  NAND2X1 U106 ( .A(n106), .B(arg_c[0]), .Y(n190) );
  INVX1 U107 ( .A(n195), .Y(n440) );
  INVX1 U108 ( .A(n404), .Y(n441) );
  INVX1 U109 ( .A(n195), .Y(n137) );
  AOI31X1 U110 ( .A(n1), .B(n2), .C(n234), .D(n235), .Y(N802) );
  AOI21AX1 U111 ( .B(n236), .C(n48), .A(n237), .Y(n234) );
  OAI2B11X1 U112 ( .D(sfroe), .C(n238), .A(n239), .B(n240), .Y(n236) );
  NOR4XL U113 ( .A(n241), .B(n242), .C(n53), .D(n55), .Y(n238) );
  NAND4X1 U114 ( .A(n377), .B(n379), .C(n168), .D(n48), .Y(N104) );
  INVX1 U115 ( .A(sfrdatai[3]), .Y(n41) );
  INVX1 U116 ( .A(sfrdatai[1]), .Y(n39) );
  INVX1 U117 ( .A(sfrdatai[2]), .Y(n40) );
  INVX1 U118 ( .A(sfrdatai[4]), .Y(n42) );
  INVX1 U119 ( .A(sfrdatai[0]), .Y(n38) );
  INVX1 U120 ( .A(sfrdatai[5]), .Y(n43) );
  INVX1 U121 ( .A(sfrdatai[7]), .Y(n45) );
  INVX1 U122 ( .A(sfrdatai[6]), .Y(n44) );
  NOR32XL U123 ( .B(n201), .C(n398), .A(n85), .Y(n396) );
  NAND2X1 U124 ( .A(n396), .B(n397), .Y(n262) );
  NOR3XL U125 ( .A(n333), .B(n79), .C(n262), .Y(n286) );
  AOI31X1 U126 ( .A(n80), .B(n333), .C(n79), .D(n286), .Y(n330) );
  INVX1 U127 ( .A(n257), .Y(n79) );
  INVX1 U128 ( .A(n388), .Y(n63) );
  INVX1 U129 ( .A(n294), .Y(n70) );
  NOR2X1 U130 ( .A(n383), .B(n375), .Y(n372) );
  NOR2X1 U131 ( .A(n383), .B(n376), .Y(n28) );
  INVX1 U132 ( .A(n333), .Y(n81) );
  NAND3X1 U133 ( .A(n257), .B(n262), .C(n81), .Y(n291) );
  NAND3X1 U134 ( .A(n262), .B(n333), .C(n79), .Y(n375) );
  NAND2X1 U135 ( .A(n207), .B(n205), .Y(n252) );
  INVX1 U136 ( .A(n392), .Y(n69) );
  NOR2X1 U137 ( .A(n383), .B(n376), .Y(n29) );
  NOR2X1 U138 ( .A(n383), .B(n376), .Y(n298) );
  INVX1 U139 ( .A(n397), .Y(n84) );
  NOR32XL U140 ( .B(n19), .C(n332), .A(n78), .Y(n354) );
  INVX1 U141 ( .A(n209), .Y(n86) );
  INVX1 U142 ( .A(n383), .Y(n67) );
  INVX1 U143 ( .A(rst), .Y(n47) );
  INVX1 U144 ( .A(n214), .Y(n82) );
  INVX1 U145 ( .A(rst), .Y(n48) );
  INVX1 U146 ( .A(n206), .Y(n60) );
  OAI21X1 U147 ( .B(n445), .C(n443), .A(n404), .Y(n195) );
  OAI22X1 U148 ( .A(n17), .B(n108), .C(n190), .D(n109), .Y(arg_c[17]) );
  NOR2X1 U149 ( .A(sum1[17]), .B(n26), .Y(n261) );
  INVX1 U150 ( .A(sum[15]), .Y(n93) );
  INVX1 U151 ( .A(sum[16]), .Y(n92) );
  NAND2X1 U152 ( .A(sum1[17]), .B(arg_c[0]), .Y(n189) );
  INVX1 U153 ( .A(sum1[17]), .Y(n106) );
  NAND2X1 U154 ( .A(n443), .B(n445), .Y(n404) );
  OAI222XL U155 ( .A(n427), .B(n12), .C(n428), .D(n254), .E(n255), .F(n104), 
        .Y(N569) );
  OAI222XL U156 ( .A(n431), .B(n253), .C(n432), .D(n254), .E(n9), .F(n105), 
        .Y(N568) );
  OAI222XL U157 ( .A(n420), .B(n12), .C(n421), .D(n254), .E(n255), .F(n103), 
        .Y(N570) );
  OAI222XL U158 ( .A(n419), .B(n253), .C(n422), .D(n254), .E(n9), .F(n102), 
        .Y(N571) );
  OAI222XL U159 ( .A(n407), .B(n12), .C(n415), .D(n254), .E(n255), .F(n101), 
        .Y(N572) );
  OAI222XL U160 ( .A(n139), .B(n253), .C(n140), .D(n254), .E(n9), .F(n100), 
        .Y(N573) );
  OAI222XL U161 ( .A(n122), .B(n12), .C(n123), .D(n254), .E(n255), .F(n98), 
        .Y(N575) );
  OAI222XL U162 ( .A(n136), .B(n253), .C(n138), .D(n254), .E(n9), .F(n99), .Y(
        N574) );
  OAI222XL U163 ( .A(n119), .B(n12), .C(n120), .D(n254), .E(n255), .F(n97), 
        .Y(N576) );
  OAI222XL U164 ( .A(n118), .B(n253), .C(n121), .D(n16), .E(n9), .F(n96), .Y(
        N577) );
  OAI222XL U165 ( .A(n116), .B(n12), .C(n117), .D(n16), .E(n255), .F(n95), .Y(
        N578) );
  OAI222XL U166 ( .A(n114), .B(n253), .C(n115), .D(n16), .E(n9), .F(n94), .Y(
        N579) );
  OAI222XL U167 ( .A(n112), .B(n12), .C(n113), .D(n16), .E(n255), .F(n93), .Y(
        N580) );
  OAI222XL U168 ( .A(n110), .B(n253), .C(n111), .D(n16), .E(n9), .F(n92), .Y(
        N581) );
  OAI22X1 U169 ( .A(n39), .B(n159), .C(n280), .D(n274), .Y(N455) );
  AOI222XL U170 ( .A(sum[2]), .B(n27), .C(n14), .D(n281), .E(n20), .F(sum1[1]), 
        .Y(n280) );
  OAI22X1 U171 ( .A(n192), .B(n439), .C(n442), .D(n438), .Y(n281) );
  OAI22X1 U172 ( .A(n38), .B(n159), .C(n282), .D(n274), .Y(N454) );
  AOI22X1 U173 ( .A(n283), .B(n284), .C(sum[1]), .D(n27), .Y(n282) );
  OAI22X1 U174 ( .A(n192), .B(n133), .C(n442), .D(n127), .Y(n284) );
  OR2X1 U175 ( .A(n259), .B(n261), .Y(n283) );
  OAI21X1 U176 ( .B(n9), .C(n126), .A(n258), .Y(N566) );
  AO222X1 U177 ( .A(n127), .B(n257), .C(n133), .D(n79), .E(n16), .F(n253), .Y(
        n258) );
  INVX1 U178 ( .A(n192), .Y(n442) );
  INVX1 U179 ( .A(n193), .Y(n444) );
  INVX1 U180 ( .A(sum[14]), .Y(n94) );
  INVX1 U181 ( .A(sum[13]), .Y(n95) );
  INVX1 U182 ( .A(sum[12]), .Y(n96) );
  INVX1 U183 ( .A(sum[11]), .Y(n97) );
  INVX1 U184 ( .A(sum[9]), .Y(n99) );
  INVX1 U185 ( .A(sum[10]), .Y(n98) );
  INVX1 U186 ( .A(sum[8]), .Y(n100) );
  INVX1 U187 ( .A(sum[6]), .Y(n102) );
  INVX1 U188 ( .A(sum[7]), .Y(n101) );
  INVX1 U189 ( .A(sum[5]), .Y(n103) );
  INVX1 U190 ( .A(sum[3]), .Y(n105) );
  INVX1 U191 ( .A(sum[4]), .Y(n104) );
  NAND21X1 U192 ( .B(n401), .A(n403), .Y(n377) );
  INVX1 U193 ( .A(sum1[2]), .Y(n431) );
  INVX1 U194 ( .A(sum1[3]), .Y(n427) );
  INVX1 U195 ( .A(sum1[4]), .Y(n420) );
  INVX1 U196 ( .A(sum1[5]), .Y(n419) );
  INVX1 U197 ( .A(sum1[6]), .Y(n407) );
  INVX1 U198 ( .A(sum1[7]), .Y(n139) );
  INVX1 U199 ( .A(sum1[8]), .Y(n136) );
  INVX1 U200 ( .A(sum1[9]), .Y(n122) );
  INVX1 U201 ( .A(sum1[10]), .Y(n119) );
  INVX1 U202 ( .A(sum1[11]), .Y(n118) );
  INVX1 U203 ( .A(sum1[12]), .Y(n116) );
  INVX1 U204 ( .A(sum1[13]), .Y(n114) );
  INVX1 U205 ( .A(sum1[14]), .Y(n112) );
  INVX1 U206 ( .A(sum1[15]), .Y(n110) );
  INVX1 U207 ( .A(sum[2]), .Y(n107) );
  INVX1 U208 ( .A(sum1[16]), .Y(n108) );
  OAI222XL U209 ( .A(n377), .B(n386), .C(n247), .D(n379), .E(n21), .F(n41), 
        .Y(N108) );
  OAI222XL U210 ( .A(n168), .B(n38), .C(n250), .D(n379), .E(n58), .F(n377), 
        .Y(N105) );
  OAI222XL U211 ( .A(n377), .B(n59), .C(n249), .D(n379), .E(n168), .F(n39), 
        .Y(N106) );
  INVX1 U212 ( .A(n391), .Y(n59) );
  OAI222XL U213 ( .A(n377), .B(n389), .C(n248), .D(n379), .E(n168), .F(n40), 
        .Y(N107) );
  OAI222XL U214 ( .A(n377), .B(n378), .C(n245), .D(n379), .E(n168), .F(n42), 
        .Y(N109) );
  OAI32X1 U215 ( .A(n124), .B(n46), .C(n49), .D(n168), .E(n43), .Y(n409) );
  OAI211X1 U216 ( .C(n196), .D(n197), .A(n166), .B(n168), .Y(N895) );
  AOI211X1 U217 ( .C(n85), .D(n198), .A(n199), .B(n200), .Y(n196) );
  OAI32X1 U218 ( .A(n201), .B(n439), .C(n202), .D(n404), .E(n203), .Y(n200) );
  OAI222XL U219 ( .A(n204), .B(n205), .C(n206), .D(n207), .E(n208), .F(n209), 
        .Y(n199) );
  OAI211X1 U220 ( .C(n160), .D(n56), .A(n161), .B(n162), .Y(n413) );
  NOR2X1 U221 ( .A(n163), .B(n164), .Y(n160) );
  NOR4XL U222 ( .A(n46), .B(n54), .C(n165), .D(n52), .Y(n163) );
  AOI31X1 U223 ( .A(n217), .B(n218), .C(n219), .D(n197), .Y(N893) );
  AOI22AXL U224 ( .A(n86), .B(n208), .D(n207), .C(n60), .Y(n218) );
  AOI21X1 U225 ( .B(n223), .C(n213), .A(n224), .Y(n217) );
  AOI221XL U226 ( .A(n82), .B(n124), .C(n88), .D(n444), .E(n220), .Y(n219) );
  INVX1 U227 ( .A(sum1[1]), .Y(n433) );
  NAND2X1 U228 ( .A(n192), .B(n193), .Y(arg_c[0]) );
  INVX1 U229 ( .A(sum[1]), .Y(n126) );
  NOR42XL U230 ( .C(n400), .D(n401), .A(n235), .B(n172), .Y(n398) );
  NOR21XL U231 ( .B(n178), .A(n88), .Y(n400) );
  NAND3X1 U232 ( .A(n205), .B(n182), .C(n396), .Y(n257) );
  AOI31X1 U233 ( .A(n394), .B(n331), .C(n262), .D(n380), .Y(n388) );
  AOI21X1 U234 ( .B(n133), .C(n257), .A(n299), .Y(n394) );
  INVX1 U235 ( .A(n203), .Y(n88) );
  OAI31XL U236 ( .A(n91), .B(n90), .C(n87), .D(mdubsy), .Y(n235) );
  NAND2X1 U237 ( .A(n172), .B(n90), .Y(mdubsy) );
  NAND42X1 U238 ( .C(n252), .D(n223), .A(n398), .B(n201), .Y(n333) );
  OAI21X1 U239 ( .B(n133), .C(n291), .A(n71), .Y(n294) );
  OAI31XL U240 ( .A(n393), .B(n28), .C(n372), .D(n83), .Y(n392) );
  NOR3XL U241 ( .A(n133), .B(n80), .C(n79), .Y(n393) );
  NAND2X1 U242 ( .A(n76), .B(n221), .Y(n292) );
  NAND3X1 U243 ( .A(n87), .B(n90), .C(n402), .Y(n201) );
  NAND2X1 U244 ( .A(n395), .B(n402), .Y(n205) );
  INVX1 U245 ( .A(n339), .Y(n64) );
  NAND2X1 U246 ( .A(n399), .B(n90), .Y(n207) );
  INVX1 U247 ( .A(n181), .Y(n85) );
  NOR2X1 U248 ( .A(n249), .B(n246), .Y(N675) );
  NOR2X1 U249 ( .A(n247), .B(n246), .Y(N677) );
  NOR2X1 U250 ( .A(n245), .B(n246), .Y(N678) );
  NOR2X1 U251 ( .A(n248), .B(n246), .Y(N676) );
  AOI21X1 U252 ( .B(n90), .C(n232), .A(n223), .Y(n397) );
  NOR2X1 U253 ( .A(n250), .B(n246), .Y(N674) );
  NAND2X1 U254 ( .A(n382), .B(n216), .Y(n383) );
  NAND3X1 U255 ( .A(n89), .B(n91), .C(n395), .Y(n209) );
  NAND21X1 U256 ( .B(n201), .A(n202), .Y(n214) );
  NAND2X1 U257 ( .A(n222), .B(n72), .Y(n206) );
  AOI31X1 U258 ( .A(n216), .B(n61), .C(n58), .D(n67), .Y(n213) );
  OAI31XL U259 ( .A(n251), .B(n84), .C(n252), .D(n48), .Y(n246) );
  NAND3X1 U260 ( .A(n201), .B(n181), .C(n209), .Y(n251) );
  OAI21X1 U261 ( .B(n231), .C(n61), .A(n384), .Y(n389) );
  NAND2X1 U262 ( .A(n382), .B(n58), .Y(n384) );
  NAND2X1 U263 ( .A(n205), .B(n221), .Y(n220) );
  INVX1 U264 ( .A(n208), .Y(n57) );
  OAI22X1 U265 ( .A(md4[1]), .B(n35), .C(n437), .D(n194), .Y(arg_b[2]) );
  OAI22X1 U266 ( .A(n432), .B(n195), .C(n30), .D(n435), .Y(arg_a[2]) );
  OAI22X1 U267 ( .A(md4[2]), .B(n35), .C(n429), .D(n194), .Y(arg_b[3]) );
  OAI22X1 U268 ( .A(n428), .B(n195), .C(n30), .D(n430), .Y(arg_a[3]) );
  OAI22X1 U269 ( .A(md4[3]), .B(n35), .C(n424), .D(n194), .Y(arg_b[4]) );
  OAI22X1 U270 ( .A(n421), .B(n195), .C(n30), .D(n426), .Y(arg_a[4]) );
  OAI22X1 U271 ( .A(md4[4]), .B(n35), .C(n423), .D(n194), .Y(arg_b[5]) );
  OAI22X1 U272 ( .A(n422), .B(n195), .C(n30), .D(n425), .Y(arg_a[5]) );
  OAI22X1 U273 ( .A(md4[5]), .B(n35), .C(n416), .D(n194), .Y(arg_b[6]) );
  OAI22X1 U274 ( .A(n415), .B(n195), .C(n31), .D(n417), .Y(arg_a[6]) );
  OAI22X1 U275 ( .A(md4[2]), .B(n33), .C(n188), .D(n429), .Y(arg_d[3]) );
  OAI222XL U276 ( .A(n17), .B(n431), .C(n190), .D(n432), .E(n137), .F(n420), 
        .Y(arg_c[3]) );
  OAI22X1 U277 ( .A(md4[6]), .B(n35), .C(n150), .D(n194), .Y(arg_b[7]) );
  OAI22X1 U278 ( .A(n140), .B(n195), .C(n31), .D(n418), .Y(arg_a[7]) );
  OAI22X1 U279 ( .A(md4[3]), .B(n33), .C(n188), .D(n424), .Y(arg_d[4]) );
  OAI222XL U280 ( .A(n189), .B(n427), .C(n8), .D(n428), .E(n137), .F(n419), 
        .Y(arg_c[4]) );
  OAI22X1 U281 ( .A(md4[7]), .B(n35), .C(n405), .D(n194), .Y(arg_b[8]) );
  OAI22X1 U282 ( .A(n138), .B(n195), .C(n440), .D(n154), .Y(arg_a[8]) );
  OAI22X1 U283 ( .A(md4[4]), .B(n33), .C(n188), .D(n423), .Y(arg_d[5]) );
  OAI222XL U284 ( .A(n17), .B(n420), .C(n190), .D(n421), .E(n137), .F(n407), 
        .Y(arg_c[5]) );
  OAI22X1 U285 ( .A(md5[0]), .B(n34), .C(n406), .D(n194), .Y(arg_b[9]) );
  OAI22X1 U286 ( .A(n123), .B(n195), .C(n440), .D(n153), .Y(arg_a[9]) );
  OAI22X1 U287 ( .A(md4[5]), .B(n33), .C(n188), .D(n416), .Y(arg_d[6]) );
  OAI222XL U288 ( .A(n189), .B(n419), .C(n8), .D(n422), .E(n137), .F(n139), 
        .Y(arg_c[6]) );
  OAI22X1 U289 ( .A(md5[1]), .B(n33), .C(n157), .D(n18), .Y(arg_b[10]) );
  OAI22X1 U290 ( .A(n120), .B(n24), .C(n30), .D(n152), .Y(arg_a[10]) );
  OAI22X1 U291 ( .A(md4[6]), .B(n34), .C(n188), .D(n150), .Y(arg_d[7]) );
  OAI222XL U292 ( .A(n17), .B(n407), .C(n190), .D(n415), .E(n137), .F(n136), 
        .Y(arg_c[7]) );
  OAI22X1 U293 ( .A(md5[2]), .B(n441), .C(n134), .D(n18), .Y(arg_b[11]) );
  OAI22X1 U294 ( .A(n121), .B(n24), .C(n30), .D(n131), .Y(arg_a[11]) );
  OAI22X1 U295 ( .A(md4[7]), .B(n33), .C(n188), .D(n405), .Y(arg_d[8]) );
  OAI222XL U296 ( .A(n189), .B(n139), .C(n8), .D(n140), .E(n137), .F(n122), 
        .Y(arg_c[8]) );
  OAI22X1 U297 ( .A(md5[3]), .B(n441), .C(n149), .D(n18), .Y(arg_b[12]) );
  OAI22X1 U298 ( .A(n117), .B(n24), .C(n30), .D(n156), .Y(arg_a[12]) );
  OAI22X1 U299 ( .A(md5[0]), .B(n34), .C(n188), .D(n406), .Y(arg_d[9]) );
  OAI222XL U300 ( .A(n17), .B(n136), .C(n190), .D(n138), .E(n440), .F(n119), 
        .Y(arg_c[9]) );
  OAI22X1 U301 ( .A(md5[4]), .B(n441), .C(n151), .D(n18), .Y(arg_b[13]) );
  OAI22X1 U302 ( .A(n115), .B(n24), .C(n30), .D(n142), .Y(arg_a[13]) );
  OAI22X1 U303 ( .A(md5[1]), .B(n34), .C(n13), .D(n157), .Y(arg_d[10]) );
  OAI222XL U304 ( .A(n189), .B(n122), .C(n8), .D(n123), .E(n440), .F(n118), 
        .Y(arg_c[10]) );
  ENOX1 U305 ( .A(n113), .B(n24), .C(n24), .D(md3[5]), .Y(arg_a[14]) );
  OAI22X1 U306 ( .A(md5[5]), .B(n441), .C(n155), .D(n18), .Y(arg_b[14]) );
  OAI22X1 U307 ( .A(md5[2]), .B(n34), .C(n13), .D(n134), .Y(arg_d[11]) );
  OAI222XL U308 ( .A(n17), .B(n119), .C(n190), .D(n120), .E(n440), .F(n116), 
        .Y(arg_c[11]) );
  OAI22X1 U309 ( .A(md5[6]), .B(n35), .C(n130), .D(n18), .Y(arg_b[15]) );
  OAI22X1 U310 ( .A(n111), .B(n24), .C(n30), .D(n133), .Y(arg_a[15]) );
  OAI22X1 U311 ( .A(md5[3]), .B(n34), .C(n13), .D(n149), .Y(arg_d[12]) );
  OAI222XL U312 ( .A(n189), .B(n118), .C(n8), .D(n121), .E(n440), .F(n114), 
        .Y(arg_c[12]) );
  OAI22X1 U313 ( .A(md5[4]), .B(n34), .C(n13), .D(n151), .Y(arg_d[13]) );
  OAI222XL U314 ( .A(n17), .B(n116), .C(n190), .D(n117), .E(n440), .F(n112), 
        .Y(arg_c[13]) );
  OAI22X1 U315 ( .A(md5[5]), .B(n34), .C(n13), .D(n155), .Y(arg_d[14]) );
  OAI222XL U316 ( .A(n189), .B(n114), .C(n8), .D(n115), .E(n440), .F(n110), 
        .Y(arg_c[14]) );
  OAI22X1 U317 ( .A(md5[6]), .B(n34), .C(n13), .D(n130), .Y(arg_d[15]) );
  OAI222XL U318 ( .A(n17), .B(n112), .C(n190), .D(n113), .E(n31), .F(n108), 
        .Y(arg_c[15]) );
  OAI22X1 U319 ( .A(md4[0]), .B(n35), .C(n436), .D(n194), .Y(arg_b[1]) );
  OAI21X1 U320 ( .B(n31), .C(n434), .A(n191), .Y(arg_a[1]) );
  NOR21XL U321 ( .B(norm_reg[15]), .A(n24), .Y(arg_a[17]) );
  OAI22X1 U322 ( .A(md5[7]), .B(n35), .C(n129), .D(n18), .Y(arg_b[16]) );
  OAI22X1 U323 ( .A(n109), .B(n24), .C(n30), .D(n439), .Y(arg_a[16]) );
  OAI22X1 U324 ( .A(md5[7]), .B(n34), .C(n13), .D(n129), .Y(arg_d[16]) );
  OAI222XL U325 ( .A(n189), .B(n110), .C(n8), .D(n111), .E(n31), .F(n106), .Y(
        arg_c[16]) );
  NAND2X1 U326 ( .A(md0[0]), .B(n33), .Y(n194) );
  NAND2X1 U327 ( .A(mdu_op[1]), .B(n443), .Y(n192) );
  OAI22X1 U328 ( .A(md4[1]), .B(n33), .C(n188), .D(n437), .Y(arg_d[2]) );
  OAI222XL U329 ( .A(n189), .B(n433), .C(sum1[17]), .D(n191), .E(n137), .F(
        n427), .Y(arg_c[2]) );
  NAND2X1 U330 ( .A(mdu_op[0]), .B(n445), .Y(n193) );
  OAI222XL U331 ( .A(n433), .B(n12), .C(n256), .D(n16), .E(n255), .F(n107), 
        .Y(N567) );
  AOI22X1 U332 ( .A(n79), .B(md3[7]), .C(md1[7]), .D(n257), .Y(n256) );
  AOI22X1 U333 ( .A(n442), .B(md3[7]), .C(n444), .D(md1[7]), .Y(n191) );
  OAI22X1 U334 ( .A(n38), .B(n355), .C(n373), .D(n357), .Y(N191) );
  AOI222XL U335 ( .A(n29), .B(md0[1]), .C(md0[2]), .D(n66), .E(n78), .F(
        sum[17]), .Y(n373) );
  OAI22X1 U336 ( .A(n40), .B(n159), .C(n279), .D(n274), .Y(N456) );
  AOI222XL U337 ( .A(sum[3]), .B(sum[17]), .C(n261), .D(norm_reg[0]), .E(n259), 
        .F(sum1[2]), .Y(n279) );
  OAI22X1 U338 ( .A(n41), .B(n159), .C(n278), .D(n274), .Y(N457) );
  AOI222XL U339 ( .A(sum[4]), .B(n27), .C(n14), .D(norm_reg[1]), .E(n20), .F(
        sum1[3]), .Y(n278) );
  OAI22X1 U340 ( .A(n42), .B(n159), .C(n277), .D(n274), .Y(N458) );
  AOI222XL U341 ( .A(sum[5]), .B(sum[17]), .C(n261), .D(norm_reg[2]), .E(n259), 
        .F(sum1[4]), .Y(n277) );
  OAI22X1 U342 ( .A(n43), .B(n159), .C(n276), .D(n274), .Y(N459) );
  AOI222XL U343 ( .A(sum[6]), .B(n27), .C(n14), .D(norm_reg[3]), .E(n20), .F(
        sum1[5]), .Y(n276) );
  OAI22X1 U344 ( .A(n166), .B(n38), .C(n270), .D(n229), .Y(N484) );
  AOI222XL U345 ( .A(sum[9]), .B(n27), .C(n14), .D(norm_reg[6]), .E(n20), .F(
        sum1[8]), .Y(n270) );
  OAI22X1 U346 ( .A(n45), .B(n159), .C(n273), .D(n274), .Y(N461) );
  AOI222XL U347 ( .A(sum[8]), .B(sum[17]), .C(n261), .D(norm_reg[5]), .E(n259), 
        .F(sum1[7]), .Y(n273) );
  OAI22X1 U348 ( .A(n166), .B(n39), .C(n269), .D(n229), .Y(N485) );
  AOI222XL U349 ( .A(sum[10]), .B(sum[17]), .C(n261), .D(norm_reg[7]), .E(n259), .F(sum1[9]), .Y(n269) );
  OAI22X1 U350 ( .A(n166), .B(n43), .C(n265), .D(n229), .Y(N489) );
  AOI222XL U351 ( .A(sum[14]), .B(n27), .C(n14), .D(norm_reg[11]), .E(n20), 
        .F(sum1[13]), .Y(n265) );
  OAI22X1 U352 ( .A(n166), .B(n42), .C(n266), .D(n229), .Y(N488) );
  AOI222XL U353 ( .A(sum[13]), .B(sum[17]), .C(n261), .D(norm_reg[10]), .E(
        n259), .F(sum1[12]), .Y(n266) );
  OAI22X1 U354 ( .A(n44), .B(n159), .C(n275), .D(n274), .Y(N460) );
  AOI222XL U355 ( .A(sum[7]), .B(sum[17]), .C(n14), .D(norm_reg[4]), .E(n20), 
        .F(sum1[6]), .Y(n275) );
  OAI22X1 U356 ( .A(n166), .B(n41), .C(n267), .D(n229), .Y(N487) );
  AOI222XL U357 ( .A(sum[12]), .B(n27), .C(n14), .D(norm_reg[9]), .E(n20), .F(
        sum1[11]), .Y(n267) );
  OAI22X1 U358 ( .A(n6), .B(n40), .C(n268), .D(n229), .Y(N486) );
  AOI222XL U359 ( .A(sum[11]), .B(sum[17]), .C(n261), .D(norm_reg[8]), .E(n259), .F(sum1[10]), .Y(n268) );
  OAI22X1 U360 ( .A(n6), .B(n44), .C(n264), .D(n229), .Y(N490) );
  AOI222XL U361 ( .A(sum[15]), .B(n27), .C(n14), .D(norm_reg[12]), .E(n20), 
        .F(sum1[14]), .Y(n264) );
  OAI22X1 U362 ( .A(n6), .B(n45), .C(n263), .D(n229), .Y(N491) );
  AOI222XL U363 ( .A(sum[16]), .B(sum[17]), .C(n261), .D(norm_reg[13]), .E(
        n259), .F(sum1[15]), .Y(n263) );
  OAI22X1 U364 ( .A(n43), .B(n161), .C(n297), .D(n288), .Y(N411) );
  AOI221XL U365 ( .A(n28), .B(md3[6]), .C(n299), .D(md3[7]), .E(n300), .Y(n297) );
  OAI222XL U366 ( .A(n296), .B(n156), .C(n70), .D(n142), .E(n93), .F(n292), 
        .Y(n300) );
  OAI22X1 U367 ( .A(n44), .B(n1), .C(n293), .D(n288), .Y(N412) );
  AOI221XL U368 ( .A(md3[5]), .B(n22), .C(md3[4]), .D(n65), .E(n295), .Y(n293)
         );
  INVX1 U369 ( .A(n296), .Y(n65) );
  OAI22X1 U370 ( .A(n439), .B(n68), .C(n92), .D(n19), .Y(n295) );
  INVX1 U371 ( .A(mdu_op[0]), .Y(n443) );
  OAI22X1 U372 ( .A(n45), .B(n161), .C(n287), .D(n288), .Y(N413) );
  AOI221XL U373 ( .A(md3[5]), .B(n289), .C(n75), .D(n26), .E(n290), .Y(n287)
         );
  INVX1 U374 ( .A(n292), .Y(n75) );
  OAI22X1 U375 ( .A(n179), .B(n291), .C(n133), .D(n71), .Y(n290) );
  INVX1 U376 ( .A(mdu_op[1]), .Y(n445) );
  OAI22X1 U377 ( .A(n42), .B(n1), .C(n301), .D(n288), .Y(N410) );
  AOI221XL U378 ( .A(n298), .B(md3[5]), .C(n23), .D(md3[6]), .E(n302), .Y(n301) );
  OAI222XL U379 ( .A(n296), .B(n131), .C(n70), .D(n156), .E(n94), .F(n292), 
        .Y(n302) );
  INVX1 U380 ( .A(md2[0]), .Y(n434) );
  INVX1 U381 ( .A(md4[0]), .Y(n436) );
  OAI22X1 U382 ( .A(n40), .B(n161), .C(n305), .D(n288), .Y(N408) );
  AOI221XL U383 ( .A(n28), .B(md3[3]), .C(n299), .D(md3[4]), .E(n306), .Y(n305) );
  OAI222XL U384 ( .A(n296), .B(n153), .C(n70), .D(n152), .E(n96), .F(n292), 
        .Y(n306) );
  OAI22X1 U385 ( .A(n41), .B(n1), .C(n303), .D(n288), .Y(N409) );
  AOI221XL U386 ( .A(n29), .B(md3[4]), .C(n23), .D(md3[5]), .E(n304), .Y(n303)
         );
  OAI222XL U387 ( .A(n296), .B(n152), .C(n70), .D(n131), .E(n95), .F(n292), 
        .Y(n304) );
  INVX1 U388 ( .A(md2[1]), .Y(n435) );
  INVX1 U389 ( .A(md4[1]), .Y(n437) );
  INVX1 U390 ( .A(norm_reg[0]), .Y(n432) );
  OAI22X1 U391 ( .A(n39), .B(n161), .C(n307), .D(n288), .Y(N407) );
  AOI221XL U392 ( .A(n29), .B(md3[2]), .C(n299), .D(md3[3]), .E(n308), .Y(n307) );
  OAI222XL U393 ( .A(n296), .B(n154), .C(n70), .D(n153), .E(n97), .F(n292), 
        .Y(n308) );
  INVX1 U394 ( .A(md2[3]), .Y(n426) );
  INVX1 U395 ( .A(md2[2]), .Y(n430) );
  INVX1 U396 ( .A(md4[3]), .Y(n424) );
  INVX1 U397 ( .A(md4[2]), .Y(n429) );
  INVX1 U398 ( .A(norm_reg[1]), .Y(n428) );
  INVX1 U399 ( .A(norm_reg[2]), .Y(n421) );
  OAI22X1 U400 ( .A(n45), .B(n162), .C(n312), .D(n313), .Y(N340) );
  AOI221XL U401 ( .A(n29), .B(md3[0]), .C(n299), .D(md3[1]), .E(n314), .Y(n312) );
  OAI222XL U402 ( .A(n296), .B(n417), .C(n70), .D(n418), .E(n99), .F(n292), 
        .Y(n314) );
  OAI22X1 U403 ( .A(n38), .B(n1), .C(n309), .D(n288), .Y(N406) );
  AOI221XL U404 ( .A(n28), .B(md3[1]), .C(n23), .D(md3[2]), .E(n310), .Y(n309)
         );
  OAI222XL U405 ( .A(n296), .B(n418), .C(n70), .D(n154), .E(n98), .F(n292), 
        .Y(n310) );
  INVX1 U406 ( .A(md2[4]), .Y(n425) );
  INVX1 U407 ( .A(md4[4]), .Y(n423) );
  INVX1 U408 ( .A(norm_reg[3]), .Y(n422) );
  OAI22X1 U409 ( .A(n44), .B(n2), .C(n315), .D(n313), .Y(N339) );
  AOI221XL U410 ( .A(n28), .B(md2[7]), .C(n23), .D(md3[0]), .E(n316), .Y(n315)
         );
  OAI222XL U411 ( .A(n296), .B(n425), .C(n70), .D(n417), .E(n100), .F(n292), 
        .Y(n316) );
  INVX1 U412 ( .A(md2[5]), .Y(n417) );
  INVX1 U413 ( .A(md2[6]), .Y(n418) );
  INVX1 U414 ( .A(md4[5]), .Y(n416) );
  INVX1 U415 ( .A(md4[6]), .Y(n150) );
  INVX1 U416 ( .A(norm_reg[4]), .Y(n415) );
  INVX1 U417 ( .A(norm_reg[5]), .Y(n140) );
  OAI22X1 U418 ( .A(n42), .B(n162), .C(n319), .D(n313), .Y(N337) );
  AOI221XL U419 ( .A(n28), .B(md2[5]), .C(n299), .D(md2[6]), .E(n320), .Y(n319) );
  OAI222XL U420 ( .A(n296), .B(n430), .C(n70), .D(n426), .E(n102), .F(n292), 
        .Y(n320) );
  OAI22X1 U421 ( .A(n43), .B(n2), .C(n317), .D(n313), .Y(N338) );
  AOI221XL U422 ( .A(n29), .B(md2[6]), .C(n23), .D(md2[7]), .E(n318), .Y(n317)
         );
  OAI222XL U423 ( .A(n7), .B(n426), .C(n70), .D(n425), .E(n101), .F(n19), .Y(
        n318) );
  INVX1 U424 ( .A(md2[7]), .Y(n154) );
  INVX1 U425 ( .A(md4[7]), .Y(n405) );
  INVX1 U426 ( .A(norm_reg[6]), .Y(n138) );
  OAI22X1 U427 ( .A(n41), .B(n162), .C(n321), .D(n313), .Y(N336) );
  AOI221XL U428 ( .A(n29), .B(md2[4]), .C(n299), .D(md2[5]), .E(n322), .Y(n321) );
  OAI222XL U429 ( .A(n7), .B(n435), .C(n11), .D(n430), .E(n103), .F(n19), .Y(
        n322) );
  INVX1 U430 ( .A(md3[0]), .Y(n153) );
  INVX1 U431 ( .A(md5[1]), .Y(n157) );
  INVX1 U432 ( .A(md3[1]), .Y(n152) );
  INVX1 U433 ( .A(md5[0]), .Y(n406) );
  INVX1 U434 ( .A(norm_reg[7]), .Y(n123) );
  INVX1 U435 ( .A(norm_reg[8]), .Y(n120) );
  OAI22X1 U436 ( .A(n39), .B(n2), .C(n325), .D(n313), .Y(N334) );
  AOI221XL U437 ( .A(n29), .B(md2[2]), .C(n23), .D(md2[3]), .E(n326), .Y(n325)
         );
  OAI222XL U438 ( .A(n7), .B(n438), .C(n11), .D(n434), .E(n105), .F(n19), .Y(
        n326) );
  OAI22X1 U439 ( .A(n40), .B(n162), .C(n323), .D(n313), .Y(N335) );
  AOI221XL U440 ( .A(n28), .B(md2[3]), .C(n299), .D(md2[4]), .E(n324), .Y(n323) );
  OAI222XL U441 ( .A(n7), .B(n434), .C(n11), .D(n435), .E(n104), .F(n19), .Y(
        n324) );
  INVX1 U442 ( .A(md3[2]), .Y(n131) );
  INVX1 U443 ( .A(md5[2]), .Y(n134) );
  INVX1 U444 ( .A(norm_reg[9]), .Y(n121) );
  OAI22X1 U445 ( .A(md4[0]), .B(n33), .C(n188), .D(n436), .Y(arg_d[1]) );
  OAI222XL U446 ( .A(n192), .B(n133), .C(n193), .D(n127), .E(n137), .F(n431), 
        .Y(arg_c[1]) );
  OAI22X1 U447 ( .A(n38), .B(n2), .C(n327), .D(n313), .Y(N333) );
  AOI221XL U448 ( .A(n28), .B(md2[1]), .C(n23), .D(md2[2]), .E(n329), .Y(n327)
         );
  OAI222XL U449 ( .A(n7), .B(n127), .C(n11), .D(n438), .E(n107), .F(n19), .Y(
        n329) );
  OAI22X1 U450 ( .A(n45), .B(n355), .C(n356), .D(n357), .Y(N198) );
  AOI221XL U451 ( .A(md0[6]), .B(n294), .C(md0[5]), .D(n339), .E(n358), .Y(
        n356) );
  OAI22X1 U452 ( .A(n68), .B(n141), .C(n342), .D(n143), .Y(n358) );
  OAI22X1 U453 ( .A(n44), .B(n355), .C(n359), .D(n357), .Y(N197) );
  AOI221XL U454 ( .A(md0[5]), .B(n294), .C(md0[4]), .D(n339), .E(n360), .Y(
        n359) );
  OAI22X1 U455 ( .A(n68), .B(n148), .C(n342), .D(n141), .Y(n360) );
  OAI22X1 U456 ( .A(n43), .B(n355), .C(n361), .D(n357), .Y(N196) );
  AOI221XL U457 ( .A(md0[4]), .B(n22), .C(md0[3]), .D(n339), .E(n362), .Y(n361) );
  OAI22X1 U458 ( .A(n68), .B(n147), .C(n342), .D(n148), .Y(n362) );
  OAI22X1 U459 ( .A(n42), .B(n355), .C(n363), .D(n357), .Y(N195) );
  AOI221XL U460 ( .A(md0[3]), .B(n22), .C(md0[2]), .D(n15), .E(n364), .Y(n363)
         );
  OAI22X1 U461 ( .A(n5), .B(n146), .C(n10), .D(n147), .Y(n364) );
  OAI22X1 U462 ( .A(n41), .B(n355), .C(n365), .D(n357), .Y(N194) );
  AOI221XL U463 ( .A(md0[2]), .B(n22), .C(md0[1]), .D(n15), .E(n366), .Y(n365)
         );
  OAI22X1 U464 ( .A(n5), .B(n145), .C(n10), .D(n146), .Y(n366) );
  OAI22X1 U465 ( .A(n39), .B(n355), .C(n370), .D(n357), .Y(N192) );
  AOI221XL U466 ( .A(md0[0]), .B(n22), .C(md0[3]), .D(n66), .E(n371), .Y(n370)
         );
  ENOX1 U467 ( .A(n106), .B(n369), .C(n29), .D(md0[2]), .Y(n371) );
  OAI22X1 U468 ( .A(n40), .B(n355), .C(n367), .D(n357), .Y(N193) );
  AOI221XL U469 ( .A(md0[1]), .B(n22), .C(md0[0]), .D(n15), .E(n368), .Y(n367)
         );
  ENOX1 U470 ( .A(n10), .B(n145), .C(n29), .D(md0[3]), .Y(n368) );
  OAI22X1 U471 ( .A(n45), .B(n237), .C(n334), .D(n158), .Y(N266) );
  AOI221XL U472 ( .A(n29), .B(md2[0]), .C(n299), .D(md2[1]), .E(n335), .Y(n334) );
  OAI222XL U473 ( .A(n64), .B(n125), .C(n11), .D(n127), .E(n126), .F(n336), 
        .Y(n335) );
  OAI22X1 U474 ( .A(n41), .B(n237), .C(n345), .D(n158), .Y(N262) );
  AOI221XL U475 ( .A(md1[2]), .B(n294), .C(md1[1]), .D(n339), .E(n346), .Y(
        n345) );
  OAI22X1 U476 ( .A(n68), .B(n128), .C(n342), .D(n125), .Y(n346) );
  OAI22X1 U477 ( .A(n39), .B(n237), .C(n349), .D(n158), .Y(N260) );
  AOI221XL U478 ( .A(md1[0]), .B(n294), .C(md0[7]), .D(n339), .E(n350), .Y(
        n349) );
  OAI22X1 U479 ( .A(n68), .B(n132), .C(n342), .D(n144), .Y(n350) );
  OAI22X1 U480 ( .A(n38), .B(n237), .C(n351), .D(n158), .Y(N259) );
  AOI221XL U481 ( .A(md0[7]), .B(n294), .C(md0[6]), .D(n339), .E(n353), .Y(
        n351) );
  OAI22X1 U482 ( .A(n68), .B(n143), .C(n342), .D(n132), .Y(n353) );
  OAI22X1 U483 ( .A(n40), .B(n237), .C(n347), .D(n158), .Y(N261) );
  AOI221XL U484 ( .A(md1[1]), .B(n294), .C(md1[0]), .D(n339), .E(n348), .Y(
        n347) );
  OAI22X1 U485 ( .A(n68), .B(n144), .C(n342), .D(n128), .Y(n348) );
  OAI22X1 U486 ( .A(n42), .B(n237), .C(n343), .D(n158), .Y(N263) );
  AOI221XL U487 ( .A(md1[3]), .B(n294), .C(md1[2]), .D(n339), .E(n344), .Y(
        n343) );
  OAI22X1 U488 ( .A(n68), .B(n125), .C(n342), .D(n127), .Y(n344) );
  OAI22X1 U489 ( .A(n44), .B(n237), .C(n337), .D(n158), .Y(N265) );
  AOI221XL U490 ( .A(n28), .B(md1[7]), .C(n23), .D(md2[0]), .E(n338), .Y(n337)
         );
  OAI222XL U491 ( .A(n64), .B(n128), .C(n11), .D(n125), .E(n433), .F(n336), 
        .Y(n338) );
  OAI22X1 U492 ( .A(n43), .B(n237), .C(n340), .D(n158), .Y(N264) );
  AOI221XL U493 ( .A(md1[4]), .B(n294), .C(md1[3]), .D(n339), .E(n341), .Y(
        n340) );
  OAI22X1 U494 ( .A(n127), .B(n68), .C(n342), .D(n438), .Y(n341) );
  OAI21BX1 U495 ( .C(set_div16), .B(n158), .A(n159), .Y(n414) );
  OAI31XL U496 ( .A(n443), .B(n46), .C(n50), .D(n169), .Y(n411) );
  AOI31X1 U497 ( .A(set_div16), .B(n56), .C(n50), .D(n49), .Y(n169) );
  INVX1 U498 ( .A(n166), .Y(n50) );
  OAI211X1 U499 ( .C(n56), .D(n166), .A(n167), .B(n168), .Y(n412) );
  NAND3X1 U500 ( .A(n166), .B(n47), .C(mdu_op[1]), .Y(n167) );
  OAI211X1 U501 ( .C(n210), .D(n197), .A(n166), .B(n168), .Y(N894) );
  AOI211X1 U502 ( .C(n88), .D(n443), .A(n211), .B(n212), .Y(n210) );
  OAI221X1 U503 ( .A(n181), .B(n198), .C(n60), .D(n207), .E(n214), .Y(n211) );
  ENOX1 U504 ( .A(md3[7]), .B(n201), .C(n84), .D(n213), .Y(n212) );
  AOI31X1 U505 ( .A(n225), .B(n226), .C(n227), .D(n197), .Y(N892) );
  NAND21X1 U506 ( .B(n205), .A(n204), .Y(n226) );
  AOI32X1 U507 ( .A(n232), .B(n90), .C(n213), .D(n82), .E(arcon[5]), .Y(n225)
         );
  AOI221XL U508 ( .A(n86), .B(n57), .C(n88), .D(n192), .E(n224), .Y(n227) );
  INVX1 U509 ( .A(md3[3]), .Y(n156) );
  INVX1 U510 ( .A(md3[4]), .Y(n142) );
  INVX1 U511 ( .A(norm_reg[10]), .Y(n117) );
  INVX1 U512 ( .A(norm_reg[11]), .Y(n115) );
  INVX1 U513 ( .A(md5[3]), .Y(n149) );
  INVX1 U514 ( .A(md5[4]), .Y(n151) );
  INVX1 U515 ( .A(md5[5]), .Y(n155) );
  INVX1 U516 ( .A(norm_reg[12]), .Y(n113) );
  INVX1 U517 ( .A(md3[6]), .Y(n133) );
  AOI211X1 U518 ( .C(sfroe), .D(n54), .A(n170), .B(n46), .Y(n410) );
  NOR2X1 U519 ( .A(arcon[7]), .B(test_so), .Y(n170) );
  INVX1 U520 ( .A(md3[7]), .Y(n439) );
  INVX1 U521 ( .A(md5[7]), .Y(n129) );
  INVX1 U522 ( .A(md5[6]), .Y(n130) );
  INVX1 U523 ( .A(norm_reg[13]), .Y(n111) );
  INVX1 U524 ( .A(norm_reg[14]), .Y(n109) );
  NAND2X1 U525 ( .A(md0[1]), .B(n33), .Y(n188) );
  INVX1 U526 ( .A(md1[6]), .Y(n127) );
  AOI21BBXL U527 ( .B(md3[6]), .C(n291), .A(n289), .Y(n296) );
  AOI221XL U528 ( .A(n378), .B(n69), .C(n380), .D(arcon[4]), .E(n62), .Y(n245)
         );
  INVX1 U529 ( .A(n381), .Y(n62) );
  GEN2XL U530 ( .D(n382), .E(n73), .C(n72), .B(n383), .A(n63), .Y(n381) );
  NAND2X1 U531 ( .A(n399), .B(oper_reg[3]), .Y(n203) );
  NOR3XL U532 ( .A(oper_reg[0]), .B(oper_reg[1]), .C(n91), .Y(n399) );
  NOR3XL U533 ( .A(oper_reg[1]), .B(oper_reg[2]), .C(oper_reg[0]), .Y(n172) );
  NOR2X1 U534 ( .A(n89), .B(oper_reg[2]), .Y(n402) );
  INVX1 U535 ( .A(oper_reg[0]), .Y(n89) );
  INVX1 U536 ( .A(oper_reg[2]), .Y(n91) );
  NAND3X1 U537 ( .A(oper_reg[3]), .B(n87), .C(n402), .Y(n178) );
  OAI211X1 U538 ( .C(md3[6]), .D(n291), .A(n331), .B(n369), .Y(n339) );
  OA222X1 U539 ( .A(counter_st[1]), .B(n63), .C(n391), .D(n392), .E(n83), .F(
        n135), .Y(n249) );
  NAND3X1 U540 ( .A(n395), .B(oper_reg[0]), .C(oper_reg[2]), .Y(n181) );
  AOI222XL U541 ( .A(n389), .B(n69), .C(n390), .D(n388), .E(n380), .F(arcon[2]), .Y(n248) );
  AO21X1 U542 ( .B(counter_st[2]), .C(counter_st[1]), .A(n382), .Y(n390) );
  AOI222XL U543 ( .A(n388), .B(N610), .C(n58), .D(n69), .E(n380), .F(arcon[0]), 
        .Y(n250) );
  AOI222XL U544 ( .A(n386), .B(n69), .C(n387), .D(n388), .E(n380), .F(arcon[3]), .Y(n247) );
  XNOR2XL U545 ( .A(n73), .B(n382), .Y(n387) );
  INVX1 U546 ( .A(oper_reg[3]), .Y(n90) );
  NOR2X1 U547 ( .A(n87), .B(oper_reg[3]), .Y(n395) );
  INVX1 U548 ( .A(oper_reg[1]), .Y(n87) );
  NAND3X1 U549 ( .A(n402), .B(oper_reg[3]), .C(oper_reg[1]), .Y(n401) );
  AND3X1 U550 ( .A(n395), .B(n89), .C(oper_reg[2]), .Y(n223) );
  NOR3XL U551 ( .A(n89), .B(oper_reg[1]), .C(n91), .Y(n232) );
  NAND3X1 U552 ( .A(n89), .B(n91), .C(oper_reg[3]), .Y(n182) );
  NOR2X1 U553 ( .A(counter_st[2]), .B(counter_st[1]), .Y(n382) );
  NOR2X1 U554 ( .A(counter_st[3]), .B(counter_st[4]), .Y(n216) );
  AND3X1 U555 ( .A(n231), .B(n73), .C(counter_st[2]), .Y(n222) );
  NAND2X1 U556 ( .A(n232), .B(oper_reg[3]), .Y(n221) );
  NOR2X1 U557 ( .A(counter_st[1]), .B(N610), .Y(n231) );
  NAND2X1 U558 ( .A(n179), .B(n215), .Y(n198) );
  NAND4X1 U559 ( .A(counter_st[1]), .B(n216), .C(n58), .D(n61), .Y(n215) );
  NAND42X1 U560 ( .C(arcon[0]), .D(arcon[2]), .A(n135), .B(n233), .Y(n202) );
  NOR2X1 U561 ( .A(arcon[4]), .B(arcon[3]), .Y(n233) );
  AOI21X1 U562 ( .B(counter_st[1]), .C(N610), .A(n231), .Y(n391) );
  XNOR2XL U563 ( .A(n384), .B(counter_st[3]), .Y(n386) );
  NAND4X1 U564 ( .A(counter_st[4]), .B(counter_st[1]), .C(n230), .D(n58), .Y(
        n208) );
  NOR2X1 U565 ( .A(counter_st[3]), .B(counter_st[2]), .Y(n230) );
  OAI22AX1 U566 ( .D(n216), .C(n384), .A(n385), .B(n72), .Y(n378) );
  NOR2X1 U567 ( .A(counter_st[3]), .B(n384), .Y(n385) );
  INVX1 U568 ( .A(N610), .Y(n58) );
  OAI31XL U569 ( .A(n201), .B(md3[7]), .C(n202), .D(n181), .Y(n224) );
  NOR2X1 U570 ( .A(md3[6]), .B(md3[5]), .Y(n179) );
  NOR42XL U571 ( .C(n434), .D(n179), .A(md2[1]), .B(n180), .Y(n177) );
  NAND4X1 U572 ( .A(n430), .B(n426), .C(n425), .D(n417), .Y(n180) );
  NOR4XL U573 ( .A(md3[1]), .B(md3[0]), .C(md2[7]), .D(md2[6]), .Y(n175) );
  NOR4XL U574 ( .A(md3[7]), .B(md3[4]), .C(md3[3]), .D(md3[2]), .Y(n176) );
  NOR4XL U575 ( .A(md4[2]), .B(md4[1]), .C(md4[0]), .D(n182), .Y(n183) );
  NAND2X1 U576 ( .A(counter_st[4]), .B(n222), .Y(n204) );
  NOR3XL U577 ( .A(n187), .B(md5[4]), .C(md5[3]), .Y(n186) );
  NAND3X1 U578 ( .A(n130), .B(n129), .C(n155), .Y(n187) );
  INVX1 U579 ( .A(counter_st[2]), .Y(n61) );
  INVX1 U580 ( .A(counter_st[4]), .Y(n72) );
  INVX1 U581 ( .A(counter_st[3]), .Y(n73) );
  INVX1 U582 ( .A(md1[7]), .Y(n438) );
  INVX1 U583 ( .A(arcon[1]), .Y(n135) );
  INVX1 U584 ( .A(md1[5]), .Y(n125) );
  INVX1 U585 ( .A(md1[4]), .Y(n128) );
  NOR2X1 U586 ( .A(n46), .B(n171), .Y(n408) );
  AOI211X1 U587 ( .C(n172), .D(oper_reg[3]), .A(n173), .B(n174), .Y(n171) );
  AO44X1 U588 ( .A(arcon[6]), .B(n181), .C(n182), .D(n178), .E(n183), .F(n184), 
        .G(n185), .H(n186), .Y(n173) );
  AOI31X1 U589 ( .A(n175), .B(n176), .C(n177), .D(n178), .Y(n174) );
  NOR4XL U590 ( .A(md5[2]), .B(md5[1]), .C(md5[0]), .D(md4[7]), .Y(n185) );
  NOR4XL U591 ( .A(md4[6]), .B(md4[5]), .C(md4[4]), .D(md4[3]), .Y(n184) );
  INVX1 U592 ( .A(set_div32), .Y(n56) );
  INVX1 U593 ( .A(md1[1]), .Y(n143) );
  INVX1 U594 ( .A(md0[4]), .Y(n145) );
  INVX1 U595 ( .A(md0[7]), .Y(n148) );
  INVX1 U596 ( .A(md0[6]), .Y(n147) );
  INVX1 U597 ( .A(md1[0]), .Y(n141) );
  INVX1 U598 ( .A(md1[2]), .Y(n132) );
  INVX1 U599 ( .A(md1[3]), .Y(n144) );
  INVX1 U600 ( .A(md0[5]), .Y(n146) );
  INVX1 U601 ( .A(arcon[5]), .Y(n124) );
endmodule


module mdu_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
endmodule


module mdu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module wakeupctrl_a0 ( irq, int0ff, int1ff, it0, it1, isreg, intprior0, 
        intprior1, eal, eint0, eint1, pmuintreq );
  input [3:0] isreg;
  input [1:0] intprior0;
  input [1:0] intprior1;
  input irq, int0ff, int1ff, it0, it1, eal, eint0, eint1;
  output pmuintreq;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n1;

  NAND42X1 U1 ( .C(it0), .D(int0ff), .A(eint0), .B(n9), .Y(n3) );
  OAI2B11X1 U2 ( .D(intprior0[0]), .C(n6), .A(n10), .B(n8), .Y(n9) );
  OAI21X1 U3 ( .B(intprior0[0]), .C(n1), .A(intprior1[0]), .Y(n10) );
  AO21X1 U4 ( .B(n2), .C(eal), .A(irq), .Y(pmuintreq) );
  AOI21X1 U5 ( .B(n3), .C(n4), .A(isreg[3]), .Y(n2) );
  NAND42X1 U6 ( .C(it1), .D(int1ff), .A(eint1), .B(n5), .Y(n4) );
  OAI2B11X1 U7 ( .D(intprior0[1]), .C(n6), .A(n7), .B(n8), .Y(n5) );
  OAI21X1 U8 ( .B(intprior0[1]), .C(n1), .A(intprior1[1]), .Y(n7) );
  OR2X1 U9 ( .A(isreg[1]), .B(isreg[2]), .Y(n6) );
  OR2X1 U10 ( .A(isreg[0]), .B(n6), .Y(n8) );
  INVX1 U11 ( .A(isreg[2]), .Y(n1) );
endmodule


module pmurstctrl_a0 ( resetff, wdts, srst, pmuintreq, stop, idle, clkcpu_en, 
        clkper_en, cpu_resume, rsttowdt, rsttosrst, rst );
  input resetff, wdts, srst, pmuintreq, stop, idle;
  output clkcpu_en, clkper_en, cpu_resume, rsttowdt, rsttosrst, rst;
  wire   n2;

  OAI21X1 U1 ( .B(stop), .C(idle), .A(n2), .Y(clkcpu_en) );
  NAND2X1 U2 ( .A(stop), .B(n2), .Y(clkper_en) );
  BUFX3 U3 ( .A(pmuintreq), .Y(cpu_resume) );
  INVX1 U4 ( .A(pmuintreq), .Y(n2) );
  OR2X1 U5 ( .A(srst), .B(resetff), .Y(rsttowdt) );
  OR2X1 U6 ( .A(wdts), .B(rsttowdt), .Y(rst) );
  OR2X1 U7 ( .A(resetff), .B(wdts), .Y(rsttosrst) );
endmodule


module sfrmux_a0 ( isfrwait, sfraddr, c, ac, f0, rs, ov, f1, p, acc, b, dpl, 
        dph, dps, dpc, p2, sp, smod, pmw, p2sel, gf0, stop, idle, ckcon, port0, 
        port0ff, rmwinstr, arcon, md0, md1, md2, md3, md4, md5, t0_tmod, 
        t0_tf0, t0_tf1, t0_tr0, t0_tr1, tl0, th0, t1_tmod, t1_tf1, t1_tr1, tl1, 
        th1, wdtrel, ip0wdts, wdt_tm, t2con, s0con, s0buf, s0rell, s0relh, bd, 
        ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9, 
        iex10, iex11, iex12, ien0, ien1, ien2, ip0, ip1, isr_tm, i2c_int, 
        i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o, sfrdatai, tf1_gate, riti0_gate, 
        iex7_gate, iex2_gate, srstflag, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, ext_sfr_sel, sfrdatao );
  input [6:0] sfraddr;
  input [1:0] rs;
  input [7:0] acc;
  input [7:0] b;
  input [7:0] dpl;
  input [7:0] dph;
  input [3:0] dps;
  input [5:0] dpc;
  input [7:0] p2;
  input [7:0] sp;
  input [7:0] ckcon;
  input [7:0] port0;
  input [7:0] port0ff;
  input [7:0] arcon;
  input [7:0] md0;
  input [7:0] md1;
  input [7:0] md2;
  input [7:0] md3;
  input [7:0] md4;
  input [7:0] md5;
  input [3:0] t0_tmod;
  input [7:0] tl0;
  input [7:0] th0;
  input [3:0] t1_tmod;
  input [7:0] tl1;
  input [7:0] th1;
  input [7:0] wdtrel;
  input [7:0] t2con;
  input [7:0] s0con;
  input [7:0] s0buf;
  input [7:0] s0rell;
  input [7:0] s0relh;
  input [7:0] ien0;
  input [5:0] ien1;
  input [5:0] ien2;
  input [5:0] ip0;
  input [5:0] ip1;
  input [7:0] i2cdat_o;
  input [7:0] i2cadr_o;
  input [7:0] i2ccon_o;
  input [7:0] i2csta_o;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  input isfrwait, c, ac, f0, ov, f1, p, smod, pmw, p2sel, gf0, stop, idle,
         rmwinstr, t0_tf0, t0_tf1, t0_tr0, t0_tr1, t1_tf1, t1_tr1, ip0wdts,
         wdt_tm, bd, ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12, isr_tm, i2c_int, srstflag;
  output tf1_gate, riti0_gate, iex7_gate, iex2_gate, int_vect_8b, int_vect_93,
         int_vect_9b, int_vect_a3, ext_sfr_sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341;

  INVX4 U2 ( .A(sfraddr[3]), .Y(n60) );
  NAND32X1 U3 ( .B(sfraddr[3]), .C(n94), .A(n42), .Y(n112) );
  NOR5XL U4 ( .A(n29), .B(n43), .C(n61), .D(n76), .E(sfraddr[3]), .Y(n48) );
  INVX2 U5 ( .A(n65), .Y(n77) );
  NAND21XL U6 ( .B(n85), .A(n49), .Y(n165) );
  NAND2X1 U7 ( .A(sfrdatai[4]), .B(n319), .Y(n5) );
  INVX1 U8 ( .A(n122), .Y(n313) );
  OR2X1 U9 ( .A(n71), .B(n60), .Y(n26) );
  NAND21X1 U10 ( .B(n92), .A(n91), .Y(n156) );
  INVXL U11 ( .A(n80), .Y(n91) );
  NAND21X1 U12 ( .B(n89), .A(n77), .Y(n190) );
  NAND21X1 U13 ( .B(sfraddr[4]), .A(n62), .Y(n94) );
  INVX3 U14 ( .A(sfraddr[2]), .Y(n59) );
  INVX2 U15 ( .A(n134), .Y(n233) );
  NOR5X1 U16 ( .A(n54), .B(n34), .C(n300), .D(n301), .E(n302), .Y(n88) );
  INVX1 U17 ( .A(n90), .Y(n73) );
  INVX1 U18 ( .A(n72), .Y(n75) );
  AND3X1 U19 ( .A(n1), .B(n2), .C(n3), .Y(n223) );
  NAND2X1 U20 ( .A(sfrdatai[2]), .B(n319), .Y(n2) );
  NAND32X1 U21 ( .B(n35), .C(n92), .A(n70), .Y(n134) );
  NOR43XL U22 ( .B(n151), .C(n150), .D(n149), .A(n148), .Y(n185) );
  NAND31X1 U23 ( .C(n183), .A(n182), .B(n181), .Y(n184) );
  NAND6XL U24 ( .A(n132), .B(n131), .C(n130), .D(n129), .E(n128), .F(n127), 
        .Y(sfrdatao[0]) );
  NAND42X1 U25 ( .C(n299), .D(n298), .A(n297), .B(n296), .Y(sfrdatao[6]) );
  NAND42X1 U26 ( .C(n338), .D(n337), .A(n336), .B(n335), .Y(sfrdatao[7]) );
  NAND6XL U27 ( .A(n264), .B(n263), .C(n262), .D(n261), .E(n260), .F(n259), 
        .Y(sfrdatao[4]) );
  NAND6XL U28 ( .A(n88), .B(n169), .C(n171), .D(n107), .E(n164), .F(n170), .Y(
        n101) );
  NAND6XL U29 ( .A(n69), .B(n140), .C(n122), .D(n121), .E(n141), .F(n120), .Y(
        n103) );
  INVX1 U30 ( .A(n114), .Y(n341) );
  INVX1 U31 ( .A(sfraddr[5]), .Y(n62) );
  NAND32X1 U32 ( .B(n94), .C(n60), .A(n43), .Y(n81) );
  NAND21X1 U33 ( .B(n56), .A(n75), .Y(n192) );
  NAND32X1 U34 ( .B(n112), .C(n23), .A(n56), .Y(n194) );
  NAND32XL U35 ( .B(sfraddr[1]), .C(sfraddr[0]), .A(n59), .Y(n37) );
  INVX1 U36 ( .A(n209), .Y(n7) );
  AOI221XL U37 ( .A(i2cadr_o[2]), .B(n331), .C(it1), .D(n41), .E(n215), .Y(
        n221) );
  INVX1 U38 ( .A(n25), .Y(n53) );
  NOR31XL U39 ( .C(n86), .A(n56), .B(n26), .Y(n30) );
  NAND42XL U40 ( .C(n318), .D(n317), .A(n316), .B(n315), .Y(n337) );
  NAND42X1 U41 ( .C(n289), .D(n288), .A(n287), .B(n286), .Y(n298) );
  NAND2X1 U42 ( .A(i2ccon_o[2]), .B(n323), .Y(n1) );
  NAND2X1 U43 ( .A(i2cdat_o[2]), .B(n321), .Y(n3) );
  INVX3 U44 ( .A(n96), .Y(n86) );
  NAND2XL U45 ( .A(n82), .B(n97), .Y(n146) );
  INVXL U46 ( .A(n67), .Y(n55) );
  AND2X2 U47 ( .A(n82), .B(n83), .Y(n54) );
  NAND32XL U48 ( .B(n29), .C(n21), .A(n61), .Y(n105) );
  NAND21XL U49 ( .B(sfraddr[6]), .A(n52), .Y(n191) );
  AND3X2 U50 ( .A(n82), .B(n27), .C(n56), .Y(n31) );
  INVX2 U51 ( .A(sfraddr[0]), .Y(n56) );
  NAND2X1 U52 ( .A(i2ccon_o[4]), .B(n323), .Y(n4) );
  NAND21X1 U53 ( .B(n61), .A(sfraddr[5]), .Y(n65) );
  NAND21XL U54 ( .B(n112), .A(n83), .Y(n120) );
  INVXL U55 ( .A(n153), .Y(n321) );
  NOR2X1 U56 ( .A(n112), .B(n92), .Y(n32) );
  NAND32XL U57 ( .B(n58), .C(n56), .A(n59), .Y(n93) );
  NAND4X1 U58 ( .A(n163), .B(n162), .C(n161), .D(n11), .Y(n8) );
  NOR31X1 U59 ( .C(n185), .A(n8), .B(n184), .Y(n209) );
  INVX1 U60 ( .A(n160), .Y(n11) );
  AO222XL U61 ( .A(ien1[5]), .B(n39), .C(dpl[5]), .D(n32), .E(dph[5]), .F(n314), .Y(n269) );
  NAND2X1 U62 ( .A(i2cdat_o[4]), .B(n321), .Y(n6) );
  AND3X2 U63 ( .A(n4), .B(n5), .C(n6), .Y(n254) );
  INVXL U64 ( .A(n154), .Y(n323) );
  INVX3 U65 ( .A(n152), .Y(n319) );
  INVXL U66 ( .A(n170), .Y(n266) );
  INVXL U67 ( .A(n171), .Y(n330) );
  INVXL U68 ( .A(n164), .Y(n334) );
  INVXL U69 ( .A(n39), .Y(n140) );
  NAND21X2 U70 ( .B(n43), .A(n73), .Y(n98) );
  NAND21XL U71 ( .B(n80), .A(n97), .Y(n169) );
  BUFX1 U72 ( .A(n311), .Y(n28) );
  INVXL U73 ( .A(n121), .Y(n283) );
  INVXL U74 ( .A(n141), .Y(n305) );
  NAND32XL U75 ( .B(sfraddr[6]), .C(n60), .A(n77), .Y(n80) );
  NAND32XL U76 ( .B(n43), .C(n93), .A(n51), .Y(n147) );
  NAND2XL U77 ( .A(n63), .B(n51), .Y(n40) );
  NAND32XL U78 ( .B(n35), .C(n93), .A(n70), .Y(n186) );
  INVXL U79 ( .A(n195), .Y(n309) );
  INVXL U80 ( .A(n196), .Y(n304) );
  INVXL U81 ( .A(n107), .Y(n333) );
  NOR2XL U82 ( .A(n71), .B(n60), .Y(n51) );
  NAND3XL U83 ( .A(n51), .B(n86), .C(n56), .Y(n154) );
  NAND32XL U84 ( .B(n92), .C(n42), .A(n51), .Y(n153) );
  NAND32XL U85 ( .B(n92), .C(n90), .A(n42), .Y(n155) );
  NAND32XL U86 ( .B(sfraddr[1]), .C(n57), .A(n59), .Y(n85) );
  INVX1 U87 ( .A(n68), .Y(n271) );
  NAND31XL U88 ( .C(sfraddr[0]), .A(sfraddr[1]), .B(n59), .Y(n92) );
  NAND43X1 U89 ( .B(n211), .C(n210), .D(n7), .A(n208), .Y(sfrdatao[1]) );
  NAND21XL U90 ( .B(sfraddr[0]), .A(n75), .Y(n176) );
  NAND21X1 U91 ( .B(n341), .A(n115), .Y(n339) );
  NAND21XL U92 ( .B(sfraddr[5]), .A(sfraddr[4]), .Y(n71) );
  OA21XL U93 ( .B(t1_tr1), .C(t0_tr1), .A(n41), .Y(n290) );
  AOI221XL U94 ( .A(tl1[7]), .B(n334), .C(tl0[7]), .D(n333), .E(n332), .Y(n335) );
  AOI22XL U95 ( .A(i2ccon_o[6]), .B(n323), .C(s0rell[6]), .D(n322), .Y(n293)
         );
  NOR42X2 U96 ( .C(n329), .D(n328), .A(n9), .B(n10), .Y(n336) );
  AO222XL U97 ( .A(i2csta_o[7]), .B(n30), .C(acc[7]), .D(n325), .E(s0relh[7]), 
        .F(n324), .Y(n9) );
  AO22XL U98 ( .A(md0[7]), .B(n327), .C(t2con[7]), .D(n326), .Y(n10) );
  NAND6X1 U99 ( .A(n248), .B(n247), .C(n246), .D(n245), .E(n244), .F(n243), 
        .Y(sfrdatao[3]) );
  AOI21BXL U100 ( .C(n25), .B(s0buf[1]), .A(n133), .Y(n136) );
  AOI21BXL U101 ( .C(n140), .B(ien1[1]), .A(n139), .Y(n143) );
  AND2XL U102 ( .A(tl0[1]), .B(n333), .Y(n168) );
  NAND2XL U103 ( .A(n41), .B(ie0), .Y(n150) );
  NAND21XL U104 ( .B(n141), .A(sp[1]), .Y(n142) );
  AND2XL U105 ( .A(f1), .B(n55), .Y(n137) );
  AND2XL U106 ( .A(acc[1]), .B(n325), .Y(n159) );
  AND2XL U107 ( .A(ip0[1]), .B(n283), .Y(n144) );
  AND2XL U108 ( .A(dph[1]), .B(n314), .Y(n145) );
  INVX1 U109 ( .A(n98), .Y(n82) );
  INVX1 U110 ( .A(n146), .Y(n327) );
  INVX1 U111 ( .A(n169), .Y(n265) );
  NAND21XL U112 ( .B(n36), .A(n79), .Y(n170) );
  INVX1 U113 ( .A(n120), .Y(n314) );
  INVX1 U114 ( .A(n147), .Y(n331) );
  INVX3 U115 ( .A(n165), .Y(n301) );
  INVX1 U116 ( .A(n40), .Y(n52) );
  INVX1 U117 ( .A(sfraddr[1]), .Y(n58) );
  INVX1 U118 ( .A(n191), .Y(n310) );
  INVX1 U119 ( .A(n105), .Y(n325) );
  INVX1 U120 ( .A(n186), .Y(n272) );
  NOR21XL U121 ( .B(n63), .A(n80), .Y(n39) );
  NAND3X1 U122 ( .A(n51), .B(n97), .C(n43), .Y(n25) );
  INVX1 U123 ( .A(sfraddr[6]), .Y(n42) );
  NAND21XL U124 ( .B(n112), .A(n97), .Y(n141) );
  OR2XL U125 ( .A(n112), .B(n76), .Y(n171) );
  NAND32XL U126 ( .B(n90), .C(n85), .A(n42), .Y(n121) );
  AND2XL U127 ( .A(n63), .B(n49), .Y(n41) );
  INVX1 U128 ( .A(n85), .Y(n97) );
  INVX1 U129 ( .A(n93), .Y(n83) );
  INVX1 U130 ( .A(n64), .Y(n115) );
  INVXL U131 ( .A(n192), .Y(n50) );
  INVX1 U132 ( .A(sfraddr[6]), .Y(n43) );
  NAND31X1 U133 ( .C(n59), .A(n49), .B(n58), .Y(n72) );
  INVX1 U134 ( .A(n66), .Y(n70) );
  NAND21X1 U135 ( .B(sfraddr[6]), .A(n60), .Y(n66) );
  INVX1 U136 ( .A(n31), .Y(n197) );
  INVX1 U137 ( .A(n155), .Y(n322) );
  INVXL U138 ( .A(n156), .Y(n324) );
  INVX1 U139 ( .A(n92), .Y(n74) );
  NAND42XL U140 ( .C(n37), .D(n29), .A(n61), .B(n70), .Y(n122) );
  NAND32XL U141 ( .B(n81), .C(n23), .A(n56), .Y(n196) );
  NAND32XL U142 ( .B(n56), .C(n98), .A(n27), .Y(n195) );
  INVX1 U143 ( .A(n95), .Y(n326) );
  NAND43X1 U144 ( .B(n36), .C(n37), .D(n60), .A(sfraddr[6]), .Y(n95) );
  INVX1 U145 ( .A(n37), .Y(n63) );
  INVX1 U146 ( .A(n176), .Y(n307) );
  NAND32XL U147 ( .B(n26), .C(n92), .A(n43), .Y(n68) );
  INVX3 U148 ( .A(n84), .Y(n300) );
  INVX1 U149 ( .A(sfraddr[4]), .Y(n61) );
  INVX1 U150 ( .A(n339), .Y(n306) );
  NAND42X1 U151 ( .C(n145), .D(n144), .A(n143), .B(n142), .Y(n210) );
  NAND42X1 U152 ( .C(n138), .D(n137), .A(n136), .B(n135), .Y(n211) );
  NOR21XL U153 ( .B(n207), .A(n206), .Y(n208) );
  AND2XL U154 ( .A(bd), .B(sfraddr[6]), .Y(n320) );
  AOI221XL U155 ( .A(tl0[6]), .B(n333), .C(t1_tmod[2]), .D(n301), .E(n295), 
        .Y(n296) );
  AO222XL U156 ( .A(ien1[4]), .B(n39), .C(dpl[4]), .D(n32), .E(dph[4]), .F(
        n314), .Y(n255) );
  AO222XL U157 ( .A(wdt_tm), .B(n330), .C(i2cadr_o[6]), .D(n331), .E(tl1[6]), 
        .F(n334), .Y(n295) );
  AO222X1 U158 ( .A(iex5), .B(n266), .C(ip1[4]), .D(n265), .E(pmw), .F(n330), 
        .Y(n249) );
  AO222X1 U159 ( .A(iex6), .B(n266), .C(ip1[5]), .D(n265), .E(isr_tm), .F(n330), .Y(n267) );
  AO222XL U160 ( .A(md0[2]), .B(n327), .C(i2csta_o[2]), .D(n30), .E(t2con[2]), 
        .F(n326), .Y(n215) );
  AO222XL U161 ( .A(md0[3]), .B(n327), .C(i2csta_o[3]), .D(n30), .E(t2con[3]), 
        .F(n326), .Y(n234) );
  AOI221XL U162 ( .A(ien2[5]), .B(n271), .C(f0), .D(n55), .E(n270), .Y(n278)
         );
  AOI221XL U163 ( .A(p2[5]), .B(n313), .C(sp[5]), .D(n305), .E(n269), .Y(n279)
         );
  AOI221XL U164 ( .A(tl1[5]), .B(n334), .C(tl0[5]), .D(n333), .E(n267), .Y(
        n282) );
  AOI222XL U165 ( .A(s0relh[0]), .B(n324), .C(s0rell[0]), .D(n322), .E(acc[0]), 
        .F(n325), .Y(n131) );
  AND4X1 U166 ( .A(n126), .B(n125), .C(n124), .D(n123), .Y(n127) );
  AND4X1 U167 ( .A(n294), .B(n293), .C(n292), .D(n291), .Y(n297) );
  AOI22XL U168 ( .A(md0[6]), .B(n327), .C(t2con[6]), .D(n326), .Y(n291) );
  AOI222XL U169 ( .A(i2csta_o[6]), .B(n30), .C(acc[6]), .D(n325), .E(s0relh[6]), .F(n324), .Y(n292) );
  AOI22X1 U170 ( .A(i2ccon_o[7]), .B(n323), .C(s0rell[7]), .D(n322), .Y(n328)
         );
  AOI221XL U171 ( .A(ien2[4]), .B(n271), .C(rs[1]), .D(n55), .E(n256), .Y(n260) );
  AOI221XL U172 ( .A(p2[4]), .B(n313), .C(sp[4]), .D(n305), .E(n255), .Y(n261)
         );
  AOI221XL U173 ( .A(tl1[4]), .B(n334), .C(tl0[4]), .D(n333), .E(n249), .Y(
        n264) );
  AOI222XL U174 ( .A(s0relh[2]), .B(n324), .C(s0rell[2]), .D(n322), .E(acc[2]), 
        .F(n325), .Y(n222) );
  AOI222XL U175 ( .A(s0relh[3]), .B(n324), .C(s0rell[3]), .D(n322), .E(acc[3]), 
        .F(n325), .Y(n241) );
  AOI221XL U176 ( .A(i2cadr_o[3]), .B(n331), .C(ie1), .D(n41), .E(n234), .Y(
        n240) );
  AOI22XL U177 ( .A(i2cadr_o[4]), .B(n331), .C(t0_tr0), .D(n41), .Y(n251) );
  AOI222XL U178 ( .A(s0relh[4]), .B(n324), .C(s0rell[4]), .D(n322), .E(acc[4]), 
        .F(n325), .Y(n253) );
  AOI222XL U179 ( .A(t2con[4]), .B(n326), .C(i2csta_o[4]), .D(n30), .E(md0[4]), 
        .F(n327), .Y(n252) );
  AOI222XL U180 ( .A(dpc[2]), .B(n272), .C(port0ff[2]), .D(n306), .E(port0[2]), 
        .F(n341), .Y(n229) );
  AOI221XL U181 ( .A(dps[2]), .B(n233), .C(ov), .D(n55), .E(n214), .Y(n225) );
  AOI222XL U182 ( .A(dpc[3]), .B(n272), .C(port0ff[3]), .D(n306), .E(port0[3]), 
        .F(n341), .Y(n248) );
  AOI221XL U183 ( .A(sp[3]), .B(n305), .C(ip0[3]), .D(n283), .E(n231), .Y(n245) );
  AND4X1 U184 ( .A(n119), .B(n118), .C(n117), .D(n116), .Y(n128) );
  NOR42XL U185 ( .C(n258), .D(n257), .A(n12), .B(n13), .Y(n259) );
  AO222XL U186 ( .A(th1[4]), .B(n50), .C(md5[4]), .D(n31), .E(b[4]), .F(n303), 
        .Y(n12) );
  AO22XL U187 ( .A(s0con[4]), .B(n310), .C(wdtrel[4]), .D(n311), .Y(n13) );
  AND4X1 U188 ( .A(n276), .B(n275), .C(n274), .D(n273), .Y(n277) );
  AOI221X1 U189 ( .A(arcon[6]), .B(n309), .C(ckcon[6]), .D(n304), .E(n284), 
        .Y(n287) );
  AO222XL U190 ( .A(port0ff[6]), .B(n306), .C(th0[6]), .D(n307), .E(port0[6]), 
        .F(n341), .Y(n284) );
  AOI221X1 U191 ( .A(port0[7]), .B(n341), .C(arcon[7]), .D(n309), .E(n308), 
        .Y(n316) );
  AOI221XL U192 ( .A(p2[6]), .B(n313), .C(sp[6]), .D(n305), .E(n285), .Y(n286)
         );
  AOI221XL U193 ( .A(dph[7]), .B(n314), .C(p2[7]), .D(n313), .E(n312), .Y(n315) );
  AO222XL U194 ( .A(wdtrel[7]), .B(n28), .C(s0con[7]), .D(n310), .E(dpl[7]), 
        .F(n32), .Y(n312) );
  AOI222XL U195 ( .A(port0[4]), .B(n341), .C(th0[4]), .D(n307), .E(port0ff[4]), 
        .F(n306), .Y(n258) );
  AOI222XL U196 ( .A(port0[5]), .B(n341), .C(th0[5]), .D(n307), .E(port0ff[5]), 
        .F(n306), .Y(n276) );
  AOI222XL U197 ( .A(dpc[0]), .B(n272), .C(port0ff[0]), .D(n306), .E(port0[0]), 
        .F(n341), .Y(n119) );
  AOI222XL U198 ( .A(p2sel), .B(n330), .C(ip1[3]), .D(n265), .E(iex4), .F(n266), .Y(n238) );
  AOI222XL U199 ( .A(idle), .B(n330), .C(ip1[0]), .D(n265), .E(iex7), .F(n266), 
        .Y(n111) );
  AOI222XL U200 ( .A(gf0), .B(n330), .C(ip1[2]), .D(n265), .E(iex3), .F(n266), 
        .Y(n219) );
  AOI222XL U201 ( .A(t0_tmod[3]), .B(n301), .C(tl1[3]), .D(n334), .E(tl0[3]), 
        .F(n333), .Y(n237) );
  AOI222XL U202 ( .A(t0_tmod[0]), .B(n301), .C(tl1[0]), .D(n334), .E(tl0[0]), 
        .F(n333), .Y(n110) );
  AOI222XL U203 ( .A(t0_tmod[2]), .B(n301), .C(tl1[2]), .D(n334), .E(tl0[2]), 
        .F(n333), .Y(n218) );
  AOI221XL U204 ( .A(dps[3]), .B(n233), .C(rs[0]), .D(n55), .E(n232), .Y(n244)
         );
  AOI221XL U205 ( .A(sp[2]), .B(n305), .C(ip0[2]), .D(n283), .E(n213), .Y(n226) );
  AO222XL U206 ( .A(dph[2]), .B(n314), .C(ien1[2]), .D(n39), .E(p2[2]), .F(
        n313), .Y(n213) );
  AOI221XL U207 ( .A(i2cadr_o[0]), .B(n331), .C(it0), .D(n41), .E(n106), .Y(
        n130) );
  AO222XL U208 ( .A(md0[0]), .B(n327), .C(i2csta_o[0]), .D(n30), .E(t2con[0]), 
        .F(n326), .Y(n106) );
  AND4X1 U209 ( .A(n180), .B(n179), .C(n178), .D(n14), .Y(n181) );
  AOI22XL U210 ( .A(md4[1]), .B(n302), .C(md3[1]), .D(n300), .Y(n14) );
  NAND31X1 U211 ( .C(n159), .A(n158), .B(n157), .Y(n160) );
  NAND21XL U212 ( .B(n155), .A(s0rell[1]), .Y(n158) );
  NAND21XL U213 ( .B(n156), .A(s0relh[1]), .Y(n157) );
  AND2X1 U214 ( .A(p2[1]), .B(n313), .Y(n139) );
  AO222XL U215 ( .A(dph[3]), .B(n314), .C(ien1[3]), .D(n39), .E(p2[3]), .F(
        n313), .Y(n231) );
  AO222XL U216 ( .A(n41), .B(tf1_gate), .C(i2cadr_o[7]), .D(n331), .E(smod), 
        .F(n330), .Y(n332) );
  NOR32XL U217 ( .B(n189), .C(n188), .A(n187), .Y(n207) );
  AND2XL U218 ( .A(port0[1]), .B(n341), .Y(n187) );
  NAND21XL U219 ( .B(n186), .A(dpc[1]), .Y(n188) );
  NAND21XL U220 ( .B(n339), .A(port0ff[1]), .Y(n189) );
  NAND8XL U221 ( .A(n205), .B(n204), .C(n203), .D(n202), .E(n201), .F(n200), 
        .G(n199), .H(n198), .Y(n206) );
  NAND21XL U222 ( .B(n191), .A(s0con[1]), .Y(n204) );
  NAND2XL U223 ( .A(n303), .B(b[1]), .Y(n205) );
  NAND21XL U224 ( .B(n134), .A(dps[1]), .Y(n135) );
  NAND21XL U225 ( .B(n153), .A(i2cdat_o[1]), .Y(n162) );
  NAND21XL U226 ( .B(n146), .A(md0[1]), .Y(n151) );
  NAND21XL U227 ( .B(n147), .A(i2cadr_o[1]), .Y(n149) );
  AND3X1 U228 ( .A(n174), .B(n173), .C(n172), .Y(n182) );
  NAND21XL U229 ( .B(n169), .A(ip1[1]), .Y(n174) );
  NAND21XL U230 ( .B(n197), .A(md5[1]), .Y(n198) );
  NAND21XL U231 ( .B(n154), .A(i2ccon_o[1]), .Y(n161) );
  AND2XL U232 ( .A(ien2[1]), .B(n271), .Y(n133) );
  AOI222XL U233 ( .A(dph[0]), .B(n314), .C(dpl[0]), .D(n32), .E(ien1[0]), .F(
        n39), .Y(n126) );
  AOI222XL U234 ( .A(ip0[0]), .B(n283), .C(p2[0]), .D(n313), .E(sp[0]), .F(
        n305), .Y(n125) );
  AND2XL U235 ( .A(ien0[1]), .B(n38), .Y(n138) );
  NAND31X1 U236 ( .C(n168), .A(n167), .B(n166), .Y(n183) );
  NAND21XL U237 ( .B(n164), .A(tl1[1]), .Y(n167) );
  AOI22XL U238 ( .A(dps[0]), .B(n233), .C(p), .D(n55), .Y(n123) );
  INVXL U239 ( .A(n32), .Y(n193) );
  OR2X1 U240 ( .A(t1_tf1), .B(t0_tf1), .Y(tf1_gate) );
  BUFX3 U241 ( .A(iex7), .Y(iex7_gate) );
  BUFX3 U242 ( .A(iex8), .Y(int_vect_8b) );
  BUFX3 U243 ( .A(iex2), .Y(iex2_gate) );
  BUFX3 U244 ( .A(iex9), .Y(int_vect_93) );
  OR2X1 U245 ( .A(s0con[1]), .B(s0con[0]), .Y(riti0_gate) );
  AO22XL U246 ( .A(i2csta_o[1]), .B(n30), .C(t2con[1]), .D(n326), .Y(n148) );
  BUFX3 U247 ( .A(iex11), .Y(int_vect_a3) );
  BUFX3 U248 ( .A(iex10), .Y(int_vect_9b) );
  INVX1 U249 ( .A(n194), .Y(n311) );
  NAND32X1 U250 ( .B(n113), .C(n42), .A(n60), .Y(n21) );
  NAND32X1 U251 ( .B(n113), .C(n42), .A(n60), .Y(n89) );
  BUFXL U252 ( .A(n311), .Y(n22) );
  NAND21X1 U253 ( .B(n58), .A(sfraddr[2]), .Y(n23) );
  INVXL U254 ( .A(sfraddr[5]), .Y(n24) );
  INVX1 U255 ( .A(n21), .Y(n79) );
  NAND21X1 U256 ( .B(n35), .A(n79), .Y(n67) );
  INVX1 U257 ( .A(sfraddr[0]), .Y(n57) );
  NOR5X2 U258 ( .A(n50), .B(n48), .C(n311), .D(n32), .E(n303), .Y(n78) );
  AO222X1 U259 ( .A(s0buf[4]), .B(n53), .C(ip0[4]), .D(n283), .E(ien0[4]), .F(
        n38), .Y(n256) );
  AO222X1 U260 ( .A(s0buf[5]), .B(n53), .C(ip0[5]), .D(n283), .E(ien0[5]), .F(
        n38), .Y(n270) );
  AO222XL U261 ( .A(ien0[3]), .B(n38), .C(s0buf[3]), .D(n53), .E(ien2[3]), .F(
        n271), .Y(n232) );
  INVX1 U262 ( .A(n23), .Y(n27) );
  BUFXL U263 ( .A(n71), .Y(n35) );
  BUFX3 U264 ( .A(n24), .Y(n29) );
  NAND32X1 U265 ( .B(n42), .C(n59), .A(n58), .Y(n96) );
  AOI22XL U266 ( .A(s0con[0]), .B(n310), .C(wdtrel[0]), .D(n311), .Y(n116) );
  AOI221XL U267 ( .A(wdtrel[2]), .B(n22), .C(dpl[2]), .D(n32), .E(n212), .Y(
        n227) );
  AOI221XL U268 ( .A(wdtrel[3]), .B(n22), .C(dpl[3]), .D(n32), .E(n230), .Y(
        n246) );
  AOI22XL U269 ( .A(s0con[5]), .B(n310), .C(wdtrel[5]), .D(n311), .Y(n273) );
  AO222X1 U270 ( .A(dpl[6]), .B(n32), .C(wdtrel[6]), .D(n28), .E(dph[6]), .F(
        n314), .Y(n285) );
  NAND32X2 U271 ( .B(n90), .C(n56), .A(n86), .Y(n87) );
  NAND32X1 U272 ( .B(sfraddr[1]), .C(sfraddr[0]), .A(n59), .Y(n113) );
  NAND21X1 U273 ( .B(n195), .A(arcon[1]), .Y(n200) );
  AND2XL U274 ( .A(n82), .B(n83), .Y(n33) );
  INVX1 U275 ( .A(n34), .Y(n177) );
  NAND6X1 U276 ( .A(n280), .B(n281), .C(n282), .D(n279), .E(n278), .F(n277), 
        .Y(sfrdatao[5]) );
  AOI222XL U277 ( .A(ckcon[5]), .B(n304), .C(dpc[5]), .D(n272), .E(arcon[5]), 
        .F(n309), .Y(n275) );
  AOI222XL U278 ( .A(ckcon[4]), .B(n304), .C(dpc[4]), .D(n272), .E(arcon[4]), 
        .F(n309), .Y(n257) );
  AOI222XL U279 ( .A(md5[3]), .B(n31), .C(arcon[3]), .D(n309), .E(ckcon[3]), 
        .F(n304), .Y(n247) );
  AOI222XL U280 ( .A(md5[2]), .B(n31), .C(arcon[2]), .D(n309), .E(ckcon[2]), 
        .F(n304), .Y(n228) );
  AOI222XL U281 ( .A(md5[0]), .B(n31), .C(arcon[0]), .D(n309), .E(ckcon[0]), 
        .F(n304), .Y(n118) );
  AO222XL U282 ( .A(th0[7]), .B(n307), .C(md2[7]), .D(n33), .E(port0ff[7]), 
        .F(n306), .Y(n308) );
  NAND21X1 U283 ( .B(n177), .A(md1[1]), .Y(n178) );
  AND4XL U284 ( .A(n111), .B(n110), .C(n109), .D(n108), .Y(n129) );
  AND4XL U285 ( .A(n238), .B(n237), .C(n236), .D(n235), .Y(n239) );
  AND4XL U286 ( .A(n219), .B(n218), .C(n217), .D(n216), .Y(n220) );
  NAND21X1 U287 ( .B(n112), .A(n63), .Y(n64) );
  INVX3 U288 ( .A(n190), .Y(n303) );
  NOR21X2 U289 ( .B(n74), .A(n98), .Y(n34) );
  INVXL U290 ( .A(n81), .Y(n49) );
  NAND21X1 U291 ( .B(n171), .A(stop), .Y(n172) );
  NAND21X1 U292 ( .B(n193), .A(dpl[1]), .Y(n202) );
  NAND21X1 U293 ( .B(n194), .A(wdtrel[1]), .Y(n201) );
  NAND21X1 U294 ( .B(n92), .A(n49), .Y(n107) );
  NAND21X1 U295 ( .B(n93), .A(n49), .Y(n164) );
  NAND21X1 U296 ( .B(n196), .A(ckcon[1]), .Y(n199) );
  NAND21X1 U297 ( .B(n170), .A(iex2), .Y(n173) );
  BUFXL U298 ( .A(n94), .Y(n36) );
  AND3X2 U299 ( .A(n63), .B(n73), .C(n43), .Y(n38) );
  AOI221XL U300 ( .A(md1[4]), .B(n34), .C(md2[4]), .D(n33), .E(n250), .Y(n263)
         );
  AOI22XL U301 ( .A(md2[0]), .B(n33), .C(th0[0]), .D(n307), .Y(n108) );
  AOI221XL U302 ( .A(md1[5]), .B(n34), .C(md2[5]), .D(n33), .E(n268), .Y(n281)
         );
  INVXL U303 ( .A(n33), .Y(n175) );
  AOI22XL U304 ( .A(md2[2]), .B(n33), .C(th0[2]), .D(n307), .Y(n216) );
  AO2222XL U305 ( .A(s0buf[7]), .B(n53), .C(sp[7]), .D(n305), .E(c), .F(n55), 
        .G(ien0[7]), .H(n38), .Y(n317) );
  AO2222XL U306 ( .A(s0buf[6]), .B(n53), .C(ip0wdts), .D(n283), .E(ac), .F(n55), .G(ien0[6]), .H(n38), .Y(n288) );
  AO222X1 U307 ( .A(ien0[2]), .B(n38), .C(s0buf[2]), .D(n53), .E(ien2[2]), .F(
        n271), .Y(n214) );
  AOI222XL U308 ( .A(ien2[0]), .B(n271), .C(s0buf[0]), .D(n53), .E(ien0[0]), 
        .F(n38), .Y(n124) );
  NOR5X1 U309 ( .A(n233), .B(n55), .C(n271), .D(n53), .E(n38), .Y(n69) );
  NOR4X1 U310 ( .A(n44), .B(n45), .C(n46), .D(n47), .Y(n280) );
  AO222X1 U311 ( .A(i2ccon_o[5]), .B(n323), .C(sfrdatai[5]), .D(n319), .E(
        i2cdat_o[5]), .F(n321), .Y(n44) );
  AO222X1 U312 ( .A(s0relh[5]), .B(n324), .C(s0rell[5]), .D(n322), .E(acc[5]), 
        .F(n325), .Y(n45) );
  AO222XL U313 ( .A(t2con[5]), .B(n326), .C(i2csta_o[5]), .D(n30), .E(md0[5]), 
        .F(n327), .Y(n46) );
  AO22XL U314 ( .A(i2cadr_o[5]), .B(n331), .C(t0_tf0), .D(n41), .Y(n47) );
  NAND32X2 U315 ( .B(n62), .C(n60), .A(n61), .Y(n90) );
  AOI22XL U316 ( .A(md2[3]), .B(n33), .C(th0[3]), .D(n307), .Y(n235) );
  AO2222XL U317 ( .A(md3[6]), .B(n300), .C(md4[6]), .D(n302), .E(md2[6]), .F(
        n33), .G(md1[6]), .H(n34), .Y(n299) );
  AO2222XL U318 ( .A(md4[7]), .B(n302), .C(t1_tmod[3]), .D(n301), .E(md1[7]), 
        .F(n34), .G(md3[7]), .H(n300), .Y(n338) );
  AOI222XL U319 ( .A(md1[0]), .B(n34), .C(md4[0]), .D(n302), .E(md3[0]), .F(
        n300), .Y(n109) );
  AOI222XL U320 ( .A(md1[3]), .B(n34), .C(md4[3]), .D(n302), .E(md3[3]), .F(
        n300), .Y(n236) );
  AO222XL U321 ( .A(md4[5]), .B(n302), .C(t1_tmod[1]), .D(n301), .E(md3[5]), 
        .F(n300), .Y(n268) );
  AO222XL U322 ( .A(md4[4]), .B(n302), .C(t1_tmod[0]), .D(n301), .E(md3[4]), 
        .F(n300), .Y(n250) );
  AOI222XL U323 ( .A(md1[2]), .B(n34), .C(md4[2]), .D(n302), .E(md3[2]), .F(
        n300), .Y(n217) );
  AND4X1 U324 ( .A(n242), .B(n241), .C(n240), .D(n239), .Y(n243) );
  INVX3 U325 ( .A(n87), .Y(n302) );
  NAND21XL U326 ( .B(n192), .A(th1[1]), .Y(n203) );
  AO2222XL U327 ( .A(md5[7]), .B(n31), .C(ckcon[7]), .D(n304), .E(th1[7]), .F(
        n50), .G(b[7]), .H(n303), .Y(n318) );
  AO2222XL U328 ( .A(b[6]), .B(n303), .C(md5[6]), .D(n31), .E(s0con[6]), .F(
        n310), .G(th1[6]), .H(n50), .Y(n289) );
  AOI222XL U329 ( .A(th1[5]), .B(n50), .C(md5[5]), .D(n31), .E(b[5]), .F(n303), 
        .Y(n274) );
  AO222XL U330 ( .A(th1[3]), .B(n50), .C(b[3]), .D(n303), .E(s0con[3]), .F(
        n310), .Y(n230) );
  AO222XL U331 ( .A(th1[2]), .B(n50), .C(b[2]), .D(n303), .E(s0con[2]), .F(
        n310), .Y(n212) );
  AOI222XL U332 ( .A(th1[0]), .B(n50), .C(srstflag), .D(n48), .E(b[0]), .F(
        n303), .Y(n117) );
  NAND21X1 U333 ( .B(n176), .A(th0[1]), .Y(n179) );
  NAND21X1 U334 ( .B(n175), .A(md2[1]), .Y(n180) );
  NAND21XL U335 ( .B(n165), .A(t0_tmod[1]), .Y(n166) );
  AOI221XL U336 ( .A(i2cdat_o[6]), .B(n321), .C(sfrdatai[6]), .D(n319), .E(
        n290), .Y(n294) );
  AOI222XL U337 ( .A(i2cdat_o[7]), .B(n321), .C(n52), .D(n320), .E(sfrdatai[7]), .F(n319), .Y(n329) );
  AOI222XL U338 ( .A(i2ccon_o[0]), .B(n323), .C(sfrdatai[0]), .D(n319), .E(
        i2cdat_o[0]), .F(n321), .Y(n132) );
  AOI222XL U339 ( .A(i2ccon_o[3]), .B(n323), .C(sfrdatai[3]), .D(n319), .E(
        i2cdat_o[3]), .F(n321), .Y(n242) );
  NAND6X1 U340 ( .A(n78), .B(n176), .C(n195), .D(n197), .E(n196), .F(n186), 
        .Y(n102) );
  NAND32X2 U341 ( .B(n96), .C(n90), .A(n56), .Y(n84) );
  NAND21X2 U342 ( .B(n115), .A(n104), .Y(n152) );
  NAND43X1 U343 ( .B(n103), .C(n101), .D(n102), .A(n100), .Y(n340) );
  INVX2 U344 ( .A(n340), .Y(n104) );
  NOR6XL U345 ( .A(n99), .B(n331), .C(n41), .D(n326), .E(n30), .F(n327), .Y(
        n100) );
  NAND6XL U346 ( .A(n153), .B(n40), .C(n154), .D(n105), .E(n155), .F(n156), 
        .Y(n99) );
  NAND21X2 U347 ( .B(n57), .A(n27), .Y(n76) );
  NAND32XL U348 ( .B(n341), .C(n340), .A(n339), .Y(ext_sfr_sel) );
  NAND21XL U349 ( .B(n152), .A(sfrdatai[1]), .Y(n163) );
  NAND32XL U350 ( .B(n37), .C(n112), .A(rmwinstr), .Y(n114) );
  AND4X1 U351 ( .A(n254), .B(n253), .C(n252), .D(n251), .Y(n262) );
  NAND6X2 U352 ( .A(n229), .B(n228), .C(n227), .D(n226), .E(n225), .F(n224), 
        .Y(sfrdatao[2]) );
  AND4X1 U353 ( .A(n223), .B(n222), .C(n221), .D(n220), .Y(n224) );
endmodule


module syncneg_a0 ( clk, reset, rsttowdt, rsttosrst, rst, int0, int1, port0i, 
        rxd0i, sdai, int0ff, int1ff, port0ff, t0ff, t1ff, rxd0ff, sdaiff, 
        rsttowdtff, rsttosrstff, rstff, resetff, test_si, test_se );
  input [7:0] port0i;
  output [7:0] port0ff;
  input clk, reset, rsttowdt, rsttosrst, rst, int0, int1, rxd0i, sdai, test_si,
         test_se;
  output int0ff, int1ff, t0ff, t1ff, rxd0ff, sdaiff, rsttowdtff, rsttosrstff,
         rstff, resetff;
  wire   reset_ff1, int0_ff1, int1_ff1, rxd0_ff1, sdai_ff1;
  wire   [7:0] p0_ff1;

  SDFFQX1 reset_ff2_reg ( .D(reset_ff1), .SIN(reset_ff1), .SMC(test_se), .C(
        clk), .Q(resetff) );
  SDFFQX1 rsttosrst_ff1_reg ( .D(rsttosrst), .SIN(rstff), .SMC(test_se), .C(
        clk), .Q(rsttosrstff) );
  SDFFQX1 rsttowdt_ff1_reg ( .D(rsttowdt), .SIN(rsttosrstff), .SMC(test_se), 
        .C(clk), .Q(rsttowdtff) );
  SDFFQX1 int0_ff2_reg ( .D(int0_ff1), .SIN(int0_ff1), .SMC(test_se), .C(clk), 
        .Q(int0ff) );
  SDFFQX1 int1_ff2_reg ( .D(int1_ff1), .SIN(int1_ff1), .SMC(test_se), .C(clk), 
        .Q(int1ff) );
  SDFFQX1 rxd0_ff2_reg ( .D(rxd0_ff1), .SIN(rxd0_ff1), .SMC(test_se), .C(clk), 
        .Q(rxd0ff) );
  SDFFQX1 sdai_ff2_reg ( .D(sdai_ff1), .SIN(sdai_ff1), .SMC(test_se), .C(clk), 
        .Q(sdaiff) );
  SDFFQX1 p0_ff2_reg_3_ ( .D(p0_ff1[3]), .SIN(port0ff[2]), .SMC(test_se), .C(
        clk), .Q(port0ff[3]) );
  SDFFQX1 p0_ff2_reg_2_ ( .D(p0_ff1[2]), .SIN(port0ff[1]), .SMC(test_se), .C(
        clk), .Q(port0ff[2]) );
  SDFFQX1 p0_ff2_reg_1_ ( .D(p0_ff1[1]), .SIN(port0ff[0]), .SMC(test_se), .C(
        clk), .Q(port0ff[1]) );
  SDFFQX1 p0_ff2_reg_7_ ( .D(p0_ff1[7]), .SIN(port0ff[6]), .SMC(test_se), .C(
        clk), .Q(port0ff[7]) );
  SDFFQX1 p0_ff2_reg_5_ ( .D(p0_ff1[5]), .SIN(port0ff[4]), .SMC(test_se), .C(
        clk), .Q(port0ff[5]) );
  SDFFQX1 p0_ff2_reg_4_ ( .D(p0_ff1[4]), .SIN(port0ff[3]), .SMC(test_se), .C(
        clk), .Q(port0ff[4]) );
  SDFFQX1 p0_ff2_reg_0_ ( .D(p0_ff1[0]), .SIN(p0_ff1[7]), .SMC(test_se), .C(
        clk), .Q(port0ff[0]) );
  SDFFQX1 p0_ff2_reg_6_ ( .D(p0_ff1[6]), .SIN(port0ff[5]), .SMC(test_se), .C(
        clk), .Q(port0ff[6]) );
  SDFFQX1 rst_ff1_reg ( .D(rst), .SIN(resetff), .SMC(test_se), .C(clk), .Q(
        rstff) );
  SDFFQX1 int0_ff1_reg ( .D(int0), .SIN(test_si), .SMC(test_se), .C(clk), .Q(
        int0_ff1) );
  SDFFQX1 int1_ff1_reg ( .D(int1), .SIN(int0ff), .SMC(test_se), .C(clk), .Q(
        int1_ff1) );
  SDFFQX1 p0_ff1_reg_6_ ( .D(port0i[6]), .SIN(p0_ff1[5]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[6]) );
  SDFFQX1 p0_ff1_reg_5_ ( .D(port0i[5]), .SIN(p0_ff1[4]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[5]) );
  SDFFQX1 p0_ff1_reg_4_ ( .D(port0i[4]), .SIN(p0_ff1[3]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[4]) );
  SDFFQX1 p0_ff1_reg_2_ ( .D(port0i[2]), .SIN(p0_ff1[1]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[2]) );
  SDFFQX1 p0_ff1_reg_1_ ( .D(port0i[1]), .SIN(p0_ff1[0]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[1]) );
  SDFFQX1 p0_ff1_reg_0_ ( .D(port0i[0]), .SIN(int1ff), .SMC(test_se), .C(clk), 
        .Q(p0_ff1[0]) );
  SDFFQX1 rxd0_ff1_reg ( .D(rxd0i), .SIN(rsttowdtff), .SMC(test_se), .C(clk), 
        .Q(rxd0_ff1) );
  SDFFQX1 p0_ff1_reg_7_ ( .D(port0i[7]), .SIN(p0_ff1[6]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[7]) );
  SDFFQX1 p0_ff1_reg_3_ ( .D(port0i[3]), .SIN(p0_ff1[2]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[3]) );
  SDFFQX1 sdai_ff1_reg ( .D(sdai), .SIN(rxd0ff), .SMC(test_se), .C(clk), .Q(
        sdai_ff1) );
  SDFFQX1 reset_ff1_reg ( .D(reset), .SIN(port0ff[7]), .SMC(test_se), .C(clk), 
        .Q(reset_ff1) );
  INVX1 U5 ( .A(1'b1), .Y(t1ff) );
  INVX1 U7 ( .A(1'b1), .Y(t0ff) );
endmodule


module mcu51_cpu_a0 ( clkcpu, rst, mempsack, memack, memdatai, memaddr, 
        mempsrd, mempswr, memrd, memwr, memaddr_comb, mempsrd_comb, 
        mempswr_comb, memrd_comb, memwr_comb, cpu_hold, cpu_resume, irq, 
        intvect, intcall, retiinstr, newinstr, rmwinstr, waitstaten, ramdatai, 
        sfrdatai, ramsfraddr, ramdatao, ramoe, ramwe, sfroe, sfrwe, sfroe_r, 
        sfrwe_r, sfroe_comb_s, sfrwe_comb_s, pc_o, pc_ini, cs_run, instr, 
        codefetch_s, sfrack, ramsfraddr_comb, ramdatao_comb, ramoe_comb, 
        ramwe_comb, ckcon, pmw, p2sel, gf0, stop, idle, acc, b, rs, c, ac, ov, 
        p, f0, f1, dph, dpl, dps, dpc, p2, sp, test_si, test_so, test_se );
  input [7:0] memdatai;
  output [15:0] memaddr;
  output [15:0] memaddr_comb;
  input [4:0] intvect;
  input [7:0] ramdatai;
  input [7:0] sfrdatai;
  output [7:0] ramsfraddr;
  output [7:0] ramdatao;
  output [15:0] pc_o;
  input [15:0] pc_ini;
  output [7:0] instr;
  output [7:0] ramsfraddr_comb;
  output [7:0] ramdatao_comb;
  output [7:0] ckcon;
  output [7:0] acc;
  output [7:0] b;
  output [1:0] rs;
  output [7:0] dph;
  output [7:0] dpl;
  output [3:0] dps;
  output [5:0] dpc;
  output [7:0] p2;
  output [7:0] sp;
  input clkcpu, rst, mempsack, memack, cpu_hold, cpu_resume, irq, sfrack,
         test_si, test_se;
  output mempsrd, mempswr, memrd, memwr, mempsrd_comb, mempswr_comb,
         memrd_comb, memwr_comb, intcall, retiinstr, newinstr, rmwinstr,
         waitstaten, ramoe, ramwe, sfroe, sfrwe, sfroe_r, sfrwe_r,
         sfroe_comb_s, sfrwe_comb_s, cs_run, codefetch_s, ramoe_comb,
         ramwe_comb, pmw, p2sel, gf0, stop, idle, c, ac, ov, p, f0, f1,
         test_so;
  wire   N343, N344, N345, n2482, n2481, finishmul, finishdiv, N370, N371,
         N372, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489,
         N490, N491, N492, N493, N494, N495, d_hold, idle_r, cpu_resume_fff,
         stop_r, ramsfrwe, N512, N515, N520, pdmode, interrupt, N582, N583,
         N584, N585, N589, N590, phase0_ff, newinstrlock, N670, N671, N672,
         N673, N674, N675, N676, N677, N679, N680, N681, N682, N683, N684,
         N685, N689, N690, accactv, N10562, N10563, N10564, N10565, N10566,
         N10567, N10568, N10569, N10570, N10571, N10572, N10573, N10574,
         N10575, N10576, N10577, N10578, N10581, N10582, N10583, N10584,
         N10585, N10586, N10587, N10588, N10589, N11478, N11479, N11480,
         N11481, N11482, N11483, N11484, N11486, N11487, N11488, N11489,
         N11491, N11498, N11499, N11500, N11501, N11502, N11503, N11504,
         N11505, N11524, N11525, N11543, N11544, N11555, N11584, N12469,
         N12470, N12472, N12477, N12478, N12479, N12480, N12481, N12482,
         N12483, N12484, N12485, N12486, N12487, N12488, N12489, N12490,
         N12491, N12492, N12493, N12494, N12495, N12496, N12497, N12498,
         N12499, N12500, N12501, N12502, N12503, N12504, N12505, N12506,
         N12507, N12508, N12509, N12510, N12511, N12512, N12513, N12514,
         N12515, N12516, N12517, N12518, N12519, N12520, N12521, N12522,
         N12523, N12524, N12525, N12526, N12527, N12528, N12529, N12530,
         N12531, N12532, N12533, N12534, N12535, N12536, N12537, N12538,
         N12539, N12540, N12541, N12542, N12543, N12544, N12545, N12546,
         N12547, N12548, N12549, N12550, N12551, N12552, N12553, N12554,
         N12555, N12556, N12557, N12558, N12559, N12560, N12561, N12562,
         N12563, N12564, N12566, N12567, N12568, N12569, N12570, N12571,
         N12572, N12573, N12575, N12576, N12577, N12578, N12579, N12580,
         N12581, N12582, N12584, N12585, N12586, N12587, N12588, N12589,
         N12590, N12591, N12593, N12594, N12595, N12596, N12597, N12598,
         N12599, N12600, N12602, N12603, N12604, N12605, N12606, N12607,
         N12608, N12609, N12611, N12612, N12613, N12614, N12615, N12616,
         N12617, N12618, N12620, N12621, N12622, N12623, N12624, N12625,
         N12626, N12627, N12629, N12630, N12631, N12632, N12633, N12634,
         N12635, N12636, N12637, N12644, N12651, N12658, N12665, N12672,
         N12679, N12686, N12690, N12691, N12692, N12693, N12694, N12695,
         N12697, N12698, N12699, N12700, N12701, N12702, N12703, N12704,
         N12705, N12706, N12709, N12710, N12711, N12714, N12715, N12716,
         N12717, N12718, N12719, N12720, N12721, N12722, N12723, N12724,
         N12725, N12726, N12727, N12728, N12729, N12730, N12770, N12771,
         N12772, N12773, N12801, N12802, N12803, N12804, N12805, N12806,
         N12807, N12808, N12824, N12825, N12826, N12827, N12828, N12829,
         N12830, N12831, N12841, N12842, N12843, N12844, N12845, N12846,
         N12847, N12848, N12849, N12850, N12851, N12852, N12853, N12854,
         N12855, N12856, N12905, israccess, N12912, waitcnt_1_, waitcnt_0_,
         N12965, N12966, N12967, N12968, N12969, N12970, N12971, N12972,
         N12974, N12975, N12976, N12977, N13014, N13023, N13032, N13041,
         N13050, N13059, N13068, N13077, N13086, N13095, N13104, N13113,
         N13122, N13131, N13140, N13149, N13158, N13167, N13176, N13185,
         N13194, N13203, N13212, N13221, N13230, N13239, N13248, N13257,
         N13266, N13275, N13284, N13293, multemp1_0_, N13324, N13325, N13326,
         N13327, N13328, N13329, N13330, N13331, N13332, N13336, N13337,
         N13338, N13339, N13340, N13341, N13342, N13343, N13345, N13346,
         N13347, N13348, N13349, N13350, N13351, N13352, N13353, N13366,
         N13367, N13368, N13369, N13370, N13371, N13372, N13373,
         cpu_resume_ff1, N13379, N13380, net12400, net12406, net12411,
         net12416, net12421, net12426, net12431, net12436, net12441, net12446,
         net12451, net12456, net12461, net12466, net12471, net12476, net12481,
         net12486, net12491, net12496, net12501, net12506, net12511, net12516,
         net12521, net12526, net12531, net12536, net12541, net12546, net12551,
         net12556, net12561, net12566, net12571, net12576, net12581, net12586,
         net12591, net12596, net12601, net12606, net12611, net12616, net12621,
         net12626, net12631, net12636, net12641, net12646, net12651, net12656,
         net12661, net12666, net12671, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, N14351, N14350, N14349, N14348, N14347, N14346, N14345,
         N14344, N14343, N14342, N14341, N14340, N14339, N14338, N14337,
         N14336, n2475, n2474, n2479, n2478, n2477, n184, n185, n186, n187,
         n188, n189, n2480, n2476, n1968, n1969, n1973, multemp1_8_,
         multemp1_7_, multemp1_6_, multemp1_5_, multemp1_4_, multemp1_3_,
         multemp1_2_, multemp1_1_, n106, n125, n217, n460, n461, n466, n469,
         n470, n471, n472, n474, n476, n477, n478, n483, n484, n485, n486,
         n487, n495, n496, n511, n512, n513, n514, n515, n516, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n601,
         n602, n606, n607, n608, n609, n610, n618, n620, n621, n645, n650,
         n655, n660, n670, n671, n678, n684, n690, n691, n692, n696, n697,
         n698, n699, n704, n712, n717, n722, n727, n732, n737, n742, n743,
         n744, n745, n749, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n786, n787, n788, n789, n790, n791, n792,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n897, n900, n901, n902, n909, n910,
         n911, n912, n915, n916, n917, n918, n919, n920, n921, n922, n925,
         n926, n927, n930, n931, n932, n935, n936, n937, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1005, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1382, n1386, n1387, n1388,
         n1390, n1391, n1393, n1394, n1395, n1396, n1400, n1401, n1402, n1403,
         n1412, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1435, n1437, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1478, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1507, n1508, n1509, n1517, n1520, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1548, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1640, n1643, n1655, n1657, n1669, n1679, n1680, n1681, n1682,
         n1683, n1684, n1686, n1687, n1690, n1691, n1692, n1693, n1694, n1695,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1725, n1726, n1727,
         n1728, n1729, n1730, n1732, n1733, n1734, n1735, n1737, n1738, n1739,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1753, n1754, n1755, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1768, n1769, n1770, n1771, n1773, n1774, n1775, n1776,
         n1777, n1780, n1781, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1876, n1877, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1970, n1971,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2073, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2141, n2142, n2143, n2148, n1, n2, n3, n10, n11, n12, n13, n14, n15,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n29, n31, n33,
         n35, n36, n38, n40, n42, n44, n45, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n62, n64, n65, n66, n67, n68, n69, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n122, n123, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n190, n191,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n462,
         n463, n464, n465, n467, n468, n473, n475, n479, n480, n481, n482,
         n488, n489, n490, n491, n492, n493, n494, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n517,
         n518, n597, n598, n599, n600, n603, n604, n605, n611, n612, n613,
         n614, n615, n616, n617, n619, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n646, n647, n648, n649, n651,
         n652, n653, n654, n656, n657, n658, n659, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n672, n673, n674, n675, n676, n677,
         n679, n680, n681, n682, n683, n685, n686, n687, n688, n689, n693,
         n694, n695, n700, n701, n702, n703, n705, n706, n707, n708, n709,
         n710, n711, n713, n714, n715, n716, n718, n719, n720, n721, n723,
         n724, n725, n726, n728, n729, n730, n731, n733, n734, n735, n736,
         n738, n739, n740, n741, n746, n747, n748, n750, n785, n793, n794,
         n795, n796, n797, n798, n799, n818, n833, n834, n835, n836, n837,
         n838, n866, n867, n868, n869, n870, n871, n881, n896, n898, n899,
         n903, n904, n905, n906, n907, n908, n913, n914, n923, n924, n928,
         n929, n933, n934, n938, n939, n1004, n1006, n1024, n1150, n1240,
         n1346, n1380, n1381, n1383, n1384, n1385, n1389, n1392, n1397, n1398,
         n1399, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1413,
         n1414, n1415, n1416, n1433, n1434, n1436, n1438, n1447, n1448, n1449,
         n1450, n1451, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1479, n1480, n1506, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1518, n1519, n1521, n1544, n1545, n1546, n1547, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1641, n1642, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1656,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1685, n1688, n1689, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1724, n1731, n1736, n1740, n1751, n1752,
         n1756, n1757, n1767, n1772, n1778, n1779, n1782, n1783, n1872, n1873,
         n1874, n1875, n1900, n1901, n1902, n1903, n1947, n1948, n1949, n1950,
         n1972, n1974, n1975, n1976, n2010, n2011, n2012, n2013, n2072, n2074,
         n2075, n2086, n2087, n2136, n2137, n2138, n2139, n2140, n2144, n2145,
         n2146, n2147, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, SYNOPSYS_UNCONNECTED_1;
  wire   [2:0] state;
  wire   [5:0] phase;
  wire   [15:0] alu_out;
  wire   [15:0] pc_i;
  wire   [7:0] temp;
  wire   [18:0] dec_accop;
  wire   [7:0] dec_cop;
  wire   [3:2] adder_out;
  wire   [9:1] multemp2;
  wire   [7:0] temp2_comb;
  wire   [7:0] dph_current;
  wire   [7:0] dpl_current;
  wire   [15:0] dptr_inc;
  wire   [63:0] dpl_reg;
  wire   [63:0] dph_reg;
  wire   [47:0] dpc_tab;
  wire   [255:0] rn_reg;
  wire   [7:0] multempreg;
  wire   [6:0] divtempreg;
  wire   [3:2] add_1_root_add_5140_2_carry;

  FAD1X1 add_1_root_add_5140_2_U1_2 ( .A(N11524), .B(N11543), .CI(
        add_1_root_add_5140_2_carry[2]), .CO(add_1_root_add_5140_2_carry[3]), 
        .SO(adder_out[2]) );
  FAD1X1 add_1_root_add_5140_2_U1_3 ( .A(N11525), .B(N11544), .CI(
        add_1_root_add_5140_2_carry[3]), .CO(N11555), .SO(adder_out[3]) );
  MAJ3X1 U2647 ( .A(n1463), .B(n1464), .C(n1465), .Y(n1426) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 clk_gate_finishmul_reg ( .CLK(clkcpu), 
        .EN(N370), .ENCLK(net12400), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 clk_gate_instr_reg ( .CLK(clkcpu), .EN(
        N685), .ENCLK(net12406), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 clk_gate_bitno_reg ( .CLK(clkcpu), .EN(
        N11491), .ENCLK(net12411), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 clk_gate_dph_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N12556), .ENCLK(net12416), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 clk_gate_dph_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N12547), .ENCLK(net12421), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 clk_gate_dph_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N12538), .ENCLK(net12426), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 clk_gate_dph_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N12529), .ENCLK(net12431), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 clk_gate_dph_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N12520), .ENCLK(net12436), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 clk_gate_dph_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N12511), .ENCLK(net12441), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 clk_gate_dph_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N12502), .ENCLK(net12446), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 clk_gate_dph_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N12493), .ENCLK(net12451), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 clk_gate_dpc_tab_reg_7_ ( .CLK(clkcpu), 
        .EN(N12686), .ENCLK(net12456), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 clk_gate_dpc_tab_reg_6_ ( .CLK(clkcpu), 
        .EN(N12679), .ENCLK(net12461), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 clk_gate_dpc_tab_reg_5_ ( .CLK(clkcpu), 
        .EN(N12672), .ENCLK(net12466), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 clk_gate_dpc_tab_reg_4_ ( .CLK(clkcpu), 
        .EN(N12665), .ENCLK(net12471), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 clk_gate_dpc_tab_reg_3_ ( .CLK(clkcpu), 
        .EN(N12658), .ENCLK(net12476), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 clk_gate_dpc_tab_reg_2_ ( .CLK(clkcpu), 
        .EN(N12651), .ENCLK(net12481), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 clk_gate_dpc_tab_reg_1_ ( .CLK(clkcpu), 
        .EN(N12644), .ENCLK(net12486), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 clk_gate_dpc_tab_reg_0_ ( .CLK(clkcpu), 
        .EN(N12637), .ENCLK(net12491), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 clk_gate_temp_reg ( .CLK(clkcpu), .EN(
        N12722), .ENCLK(net12496), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 clk_gate_waitcnt_reg ( .CLK(clkcpu), 
        .EN(N12977), .ENCLK(net12501), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 clk_gate_rn_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N13293), .ENCLK(net12506), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 clk_gate_rn_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N13284), .ENCLK(net12511), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 clk_gate_rn_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N13275), .ENCLK(net12516), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 clk_gate_rn_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N13266), .ENCLK(net12521), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 clk_gate_rn_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N13257), .ENCLK(net12526), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 clk_gate_rn_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N13248), .ENCLK(net12531), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 clk_gate_rn_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N13239), .ENCLK(net12536), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 clk_gate_rn_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N13230), .ENCLK(net12541), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 clk_gate_rn_reg_reg_8_ ( .CLK(clkcpu), 
        .EN(N13221), .ENCLK(net12546), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 clk_gate_rn_reg_reg_9_ ( .CLK(clkcpu), 
        .EN(N13212), .ENCLK(net12551), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 clk_gate_rn_reg_reg_10_ ( .CLK(clkcpu), 
        .EN(N13203), .ENCLK(net12556), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 clk_gate_rn_reg_reg_11_ ( .CLK(clkcpu), 
        .EN(N13194), .ENCLK(net12561), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 clk_gate_rn_reg_reg_12_ ( .CLK(clkcpu), 
        .EN(N13185), .ENCLK(net12566), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 clk_gate_rn_reg_reg_13_ ( .CLK(clkcpu), 
        .EN(N13176), .ENCLK(net12571), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 clk_gate_rn_reg_reg_14_ ( .CLK(clkcpu), 
        .EN(N13167), .ENCLK(net12576), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 clk_gate_rn_reg_reg_15_ ( .CLK(clkcpu), 
        .EN(N13158), .ENCLK(net12581), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 clk_gate_rn_reg_reg_16_ ( .CLK(clkcpu), 
        .EN(N13149), .ENCLK(net12586), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 clk_gate_rn_reg_reg_17_ ( .CLK(clkcpu), 
        .EN(N13140), .ENCLK(net12591), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 clk_gate_rn_reg_reg_18_ ( .CLK(clkcpu), 
        .EN(N13131), .ENCLK(net12596), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 clk_gate_rn_reg_reg_19_ ( .CLK(clkcpu), 
        .EN(N13122), .ENCLK(net12601), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 clk_gate_rn_reg_reg_20_ ( .CLK(clkcpu), 
        .EN(N13113), .ENCLK(net12606), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 clk_gate_rn_reg_reg_21_ ( .CLK(clkcpu), 
        .EN(N13104), .ENCLK(net12611), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 clk_gate_rn_reg_reg_22_ ( .CLK(clkcpu), 
        .EN(N13095), .ENCLK(net12616), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 clk_gate_rn_reg_reg_23_ ( .CLK(clkcpu), 
        .EN(N13086), .ENCLK(net12621), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 clk_gate_rn_reg_reg_24_ ( .CLK(clkcpu), 
        .EN(N13077), .ENCLK(net12626), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 clk_gate_rn_reg_reg_25_ ( .CLK(clkcpu), 
        .EN(N13068), .ENCLK(net12631), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 clk_gate_rn_reg_reg_26_ ( .CLK(clkcpu), 
        .EN(N13059), .ENCLK(net12636), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 clk_gate_rn_reg_reg_27_ ( .CLK(clkcpu), 
        .EN(N13050), .ENCLK(net12641), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 clk_gate_rn_reg_reg_28_ ( .CLK(clkcpu), 
        .EN(N13041), .ENCLK(net12646), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 clk_gate_rn_reg_reg_29_ ( .CLK(clkcpu), 
        .EN(N13032), .ENCLK(net12651), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 clk_gate_rn_reg_reg_30_ ( .CLK(clkcpu), 
        .EN(N13023), .ENCLK(net12656), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 clk_gate_rn_reg_reg_31_ ( .CLK(clkcpu), 
        .EN(N13014), .ENCLK(net12661), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 clk_gate_multempreg_reg ( .CLK(clkcpu), 
        .EN(N13324), .ENCLK(net12666), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 clk_gate_divtempreg_reg ( .CLK(clkcpu), 
        .EN(N13366), .ENCLK(net12671), .TE(test_se) );
  mcu51_cpu_a0_DW01_add_0 add_5586 ( .A({n2148, n2148, n2148, n2148, n2148, 
        n2148, n2148, n2148, N12831, N12830, N12829, N12828, N12827, N12826, 
        N12825, N12824}), .B({N12856, N12855, N12854, N12853, N12852, N12851, 
        N12850, N12849, N12848, N12847, N12846, N12845, N12844, N12843, N12842, 
        N12841}), .CI(1'b0), .SUM(alu_out), .CO() );
  mcu51_cpu_a0_DW01_sub_0 sub_5969 ( .A({1'b0, n189, n188, n187, n186, n185, 
        n184, n2135, acc[6]}), .B({1'b0, b}), .CI(1'b0), .DIFF({N13353, N13352, 
        N13351, N13350, N13349, N13348, N13347, N13346, N13345}), .CO() );
  mcu51_cpu_a0_DW01_sub_1 sub_5950 ( .A({1'b0, divtempreg, n2481}), .B({1'b0, 
        b}), .CI(1'b0), .DIFF({N13343, SYNOPSYS_UNCONNECTED_1, N13342, N13341, 
        N13340, N13339, N13338, N13337, N13336}), .CO() );
  mcu51_cpu_a0_DW01_inc_0 add_5525 ( .A({n106, n2250, n125, N12773, N12772, 
        N12771, N12770, n217}), .SUM({N12808, N12807, N12806, N12805, N12804, 
        N12803, N12802, N12801}) );
  mcu51_cpu_a0_DW01_inc_1 add_5286 ( .A({dph_current, dpl_current[7], n2143, 
        dpl_current[5], n2142, n2141, dpl_current[2:0]}), .SUM(dptr_inc) );
  mcu51_cpu_a0_DW01_inc_2 r715 ( .A({pc_o[15:7], memaddr[6:5], pc_o[4:0]}), 
        .SUM(pc_i) );
  mcu51_cpu_a0_DW01_add_8 add_5901_aco ( .A({1'b0, multempreg}), .B({1'b0, 
        N14343, N14342, N14341, N14340, N14339, N14338, N14337, N14336}), .CI(
        1'b0), .SUM({multemp1_8_, multemp1_7_, multemp1_6_, multemp1_5_, 
        multemp1_4_, multemp1_3_, multemp1_2_, multemp1_1_, multemp1_0_}), 
        .CO() );
  mcu51_cpu_a0_DW01_add_7 add_5907_aco ( .A({1'b0, multemp1_8_, multemp1_7_, 
        multemp1_6_, multemp1_5_, multemp1_4_, multemp1_3_, multemp1_2_, 
        multemp1_1_}), .B({1'b0, N14351, N14350, N14349, N14348, N14347, 
        N14346, N14345, N14344}), .CI(1'b0), .SUM(multemp2), .CO() );
  SDFFQX1 pc_reg_0_ ( .D(N480), .SIN(p), .SMC(test_se), .C(net12400), .Q(
        pc_o[0]) );
  SDFFQX1 pc_reg_1_ ( .D(N481), .SIN(pc_o[0]), .SMC(test_se), .C(net12400), 
        .Q(memaddr[1]) );
  SDFFQX1 pc_reg_2_ ( .D(N482), .SIN(pc_o[1]), .SMC(test_se), .C(net12400), 
        .Q(memaddr[2]) );
  SDFFQX1 pc_reg_3_ ( .D(N483), .SIN(memaddr[2]), .SMC(test_se), .C(net12400), 
        .Q(memaddr[3]) );
  SDFFQX1 pc_reg_4_ ( .D(N484), .SIN(pc_o[3]), .SMC(test_se), .C(net12400), 
        .Q(memaddr[4]) );
  SDFFQX1 pc_reg_5_ ( .D(N485), .SIN(memaddr[4]), .SMC(test_se), .C(net12400), 
        .Q(memaddr[5]) );
  SDFFQX1 pc_reg_6_ ( .D(N486), .SIN(pc_o[5]), .SMC(test_se), .C(net12400), 
        .Q(pc_o[6]) );
  SDFFQX1 pc_reg_7_ ( .D(N487), .SIN(pc_o[6]), .SMC(test_se), .C(net12400), 
        .Q(pc_o[7]) );
  SDFFQX1 pc_reg_8_ ( .D(N488), .SIN(pc_o[7]), .SMC(test_se), .C(net12400), 
        .Q(memaddr[8]) );
  SDFFQX1 pc_reg_9_ ( .D(N489), .SIN(pc_o[8]), .SMC(test_se), .C(net12400), 
        .Q(memaddr[9]) );
  SDFFQX1 pc_reg_10_ ( .D(N490), .SIN(pc_o[9]), .SMC(test_se), .C(net12400), 
        .Q(pc_o[10]) );
  SDFFQX1 pc_reg_11_ ( .D(N491), .SIN(memaddr[10]), .SMC(test_se), .C(net12400), .Q(memaddr[11]) );
  SDFFQX1 pc_reg_12_ ( .D(N492), .SIN(pc_o[11]), .SMC(test_se), .C(net12400), 
        .Q(memaddr[12]) );
  SDFFQX1 pc_reg_13_ ( .D(N493), .SIN(pc_o[12]), .SMC(test_se), .C(net12400), 
        .Q(pc_o[13]) );
  SDFFQX1 pc_reg_14_ ( .D(N494), .SIN(pc_o[13]), .SMC(test_se), .C(net12400), 
        .Q(pc_o[14]) );
  SDFFQX1 pc_reg_15_ ( .D(N495), .SIN(pc_o[14]), .SMC(test_se), .C(net12400), 
        .Q(pc_o[15]) );
  SDFFQX1 cpu_resume_ff1_reg ( .D(N13379), .SIN(ckcon[7]), .SMC(test_se), .C(
        clkcpu), .Q(cpu_resume_ff1) );
  SDFFQX1 newinstrlock_reg ( .D(n1878), .SIN(multempreg[7]), .SMC(test_se), 
        .C(net12400), .Q(newinstrlock) );
  SDFFQX1 phase0_ff_reg ( .D(N689), .SIN(pdmode), .SMC(test_se), .C(net12400), 
        .Q(phase0_ff) );
  SDFFQX1 finishdiv_reg ( .D(N372), .SIN(f1), .SMC(test_se), .C(net12400), .Q(
        finishdiv) );
  SDFFQX1 finishmul_reg ( .D(N371), .SIN(finishdiv), .SMC(test_se), .C(
        net12400), .Q(finishmul) );
  SDFFQX1 multempreg_reg_7_ ( .D(N13332), .SIN(multempreg[6]), .SMC(test_se), 
        .C(net12666), .Q(multempreg[7]) );
  SDFFQX1 multempreg_reg_6_ ( .D(N13331), .SIN(multempreg[5]), .SMC(test_se), 
        .C(net12666), .Q(multempreg[6]) );
  SDFFQX1 multempreg_reg_5_ ( .D(N13330), .SIN(multempreg[4]), .SMC(test_se), 
        .C(net12666), .Q(multempreg[5]) );
  SDFFQX1 multempreg_reg_4_ ( .D(N13329), .SIN(multempreg[3]), .SMC(test_se), 
        .C(net12666), .Q(multempreg[4]) );
  SDFFQX1 multempreg_reg_3_ ( .D(N13328), .SIN(multempreg[2]), .SMC(test_se), 
        .C(net12666), .Q(multempreg[3]) );
  SDFFQX1 multempreg_reg_2_ ( .D(N13327), .SIN(multempreg[1]), .SMC(test_se), 
        .C(net12666), .Q(multempreg[2]) );
  SDFFQX1 pdmode_reg ( .D(n1973), .SIN(pc_o[15]), .SMC(test_se), .C(net12400), 
        .Q(pdmode) );
  SDFFQX1 d_hold_reg ( .D(cpu_hold), .SIN(cpu_resume_fff), .SMC(test_se), .C(
        clkcpu), .Q(d_hold) );
  SDFFQX1 cpu_resume_fff_reg ( .D(N13380), .SIN(cpu_resume_ff1), .SMC(test_se), 
        .C(clkcpu), .Q(cpu_resume_fff) );
  SDFFQX1 idle_r_reg ( .D(N512), .SIN(gf0), .SMC(test_se), .C(net12400), .Q(
        idle_r) );
  SDFFQX1 stop_r_reg ( .D(N515), .SIN(state[2]), .SMC(test_se), .C(net12400), 
        .Q(stop_r) );
  SDFFQX1 israccess_reg ( .D(N12912), .SIN(interrupt), .SMC(test_se), .C(
        net12400), .Q(israccess) );
  SDFFQX1 state_reg_1_ ( .D(N589), .SIN(state[0]), .SMC(test_se), .C(net12400), 
        .Q(state[1]) );
  SDFFQX1 phase_reg_5_ ( .D(N684), .SIN(phase[4]), .SMC(test_se), .C(net12400), 
        .Q(phase[5]) );
  SDFFQX1 state_reg_2_ ( .D(N590), .SIN(state[1]), .SMC(test_se), .C(net12400), 
        .Q(state[2]) );
  SDFFQX1 state_reg_0_ ( .D(n1724), .SIN(sp[7]), .SMC(test_se), .C(net12400), 
        .Q(state[0]) );
  SDFFQX1 ramoe_r_reg ( .D(N11486), .SIN(ramdatao[7]), .SMC(test_se), .C(
        net12400), .Q(ramoe) );
  SDFFQX1 phase_reg_4_ ( .D(N683), .SIN(phase[3]), .SMC(test_se), .C(net12400), 
        .Q(phase[4]) );
  SDFFQX1 dec_cop_reg_0_ ( .D(N10582), .SIN(dec_accop[18]), .SMC(test_se), .C(
        net12400), .Q(dec_cop[0]) );
  SDFFQX1 phase_reg_3_ ( .D(N682), .SIN(phase[2]), .SMC(test_se), .C(net12400), 
        .Q(phase[3]) );
  SDFFQX1 f0_reg ( .D(n1882), .SIN(dps[3]), .SMC(test_se), .C(net12400), .Q(f0) );
  SDFFQX1 f1_reg ( .D(n1883), .SIN(f0), .SMC(test_se), .C(net12400), .Q(f1) );
  SDFFQX1 ov_reg_reg ( .D(N12711), .SIN(newinstrlock), .SMC(test_se), .C(
        net12400), .Q(ov) );
  SDFFQX1 p2_reg_reg_7_ ( .D(N12492), .SIN(p2[6]), .SMC(test_se), .C(net12400), 
        .Q(p2[7]) );
  SDFFQX1 p2_reg_reg_5_ ( .D(N12490), .SIN(p2[4]), .SMC(test_se), .C(net12400), 
        .Q(p2[5]) );
  SDFFQX1 p2_reg_reg_4_ ( .D(N12489), .SIN(p2[3]), .SMC(test_se), .C(net12400), 
        .Q(p2[4]) );
  SDFFQX1 p2_reg_reg_6_ ( .D(N12491), .SIN(p2[5]), .SMC(test_se), .C(net12400), 
        .Q(p2[6]) );
  SDFFQX1 stop_s_reg ( .D(n1880), .SIN(stop_r), .SMC(test_se), .C(net12400), 
        .Q(stop) );
  SDFFQX1 p2_reg_reg_1_ ( .D(N12486), .SIN(p2[0]), .SMC(test_se), .C(net12400), 
        .Q(p2[1]) );
  SDFFQX1 p_reg ( .D(N12905), .SIN(p2sel), .SMC(test_se), .C(net12400), .Q(p)
         );
  SDFFQX1 rn_reg_reg_7__2_ ( .D(n243), .SIN(rn_reg[193]), .SMC(test_se), .C(
        net12541), .Q(rn_reg[194]) );
  SDFFQX1 rn_reg_reg_7__6_ ( .D(n1778), .SIN(rn_reg[197]), .SMC(test_se), .C(
        net12541), .Q(rn_reg[198]) );
  SDFFQX1 rn_reg_reg_23__6_ ( .D(n230), .SIN(rn_reg[69]), .SMC(test_se), .C(
        net12621), .Q(rn_reg[70]) );
  SDFFQX1 rn_reg_reg_23__2_ ( .D(n243), .SIN(rn_reg[65]), .SMC(test_se), .C(
        net12621), .Q(rn_reg[66]) );
  SDFFQX1 dpc_tab_reg_3__2_ ( .D(n243), .SIN(dpc_tab[19]), .SMC(test_se), .C(
        net12476), .Q(dpc_tab[20]) );
  SDFFQX1 dpc_tab_reg_7__2_ ( .D(n243), .SIN(dpc_tab[43]), .SMC(test_se), .C(
        net12456), .Q(dpc_tab[44]) );
  SDFFQX1 rn_reg_reg_31__6_ ( .D(n230), .SIN(rn_reg[5]), .SMC(test_se), .C(
        net12661), .Q(rn_reg[6]) );
  SDFFQX1 rn_reg_reg_31__2_ ( .D(n243), .SIN(rn_reg[1]), .SMC(test_se), .C(
        net12661), .Q(rn_reg[2]) );
  SDFFQX1 rn_reg_reg_15__6_ ( .D(n230), .SIN(rn_reg[133]), .SMC(test_se), .C(
        net12581), .Q(rn_reg[134]) );
  SDFFQX1 rn_reg_reg_15__2_ ( .D(n243), .SIN(rn_reg[129]), .SMC(test_se), .C(
        net12581), .Q(rn_reg[130]) );
  SDFFQX1 rn_reg_reg_5__2_ ( .D(n241), .SIN(rn_reg[209]), .SMC(test_se), .C(
        net12531), .Q(rn_reg[210]) );
  SDFFQX1 rn_reg_reg_5__6_ ( .D(n229), .SIN(rn_reg[213]), .SMC(test_se), .C(
        net12531), .Q(rn_reg[214]) );
  SDFFQX1 rn_reg_reg_21__6_ ( .D(n229), .SIN(rn_reg[85]), .SMC(test_se), .C(
        net12611), .Q(rn_reg[86]) );
  SDFFQX1 rn_reg_reg_21__2_ ( .D(n241), .SIN(rn_reg[81]), .SMC(test_se), .C(
        net12611), .Q(rn_reg[82]) );
  SDFFQX1 rn_reg_reg_29__6_ ( .D(n229), .SIN(rn_reg[21]), .SMC(test_se), .C(
        net12651), .Q(rn_reg[22]) );
  SDFFQX1 rn_reg_reg_29__2_ ( .D(n241), .SIN(rn_reg[17]), .SMC(test_se), .C(
        net12651), .Q(rn_reg[18]) );
  SDFFQX1 rn_reg_reg_13__6_ ( .D(n229), .SIN(rn_reg[149]), .SMC(test_se), .C(
        net12571), .Q(rn_reg[150]) );
  SDFFQX1 rn_reg_reg_13__2_ ( .D(n241), .SIN(rn_reg[145]), .SMC(test_se), .C(
        net12571), .Q(rn_reg[146]) );
  SDFFQX1 rn_reg_reg_6__2_ ( .D(n240), .SIN(rn_reg[201]), .SMC(test_se), .C(
        net12536), .Q(rn_reg[202]) );
  SDFFQX1 rn_reg_reg_6__6_ ( .D(n228), .SIN(rn_reg[205]), .SMC(test_se), .C(
        net12536), .Q(rn_reg[206]) );
  SDFFQX1 rn_reg_reg_22__6_ ( .D(n228), .SIN(rn_reg[77]), .SMC(test_se), .C(
        net12616), .Q(rn_reg[78]) );
  SDFFQX1 rn_reg_reg_22__2_ ( .D(n240), .SIN(rn_reg[73]), .SMC(test_se), .C(
        net12616), .Q(rn_reg[74]) );
  SDFFQX1 dpc_tab_reg_2__2_ ( .D(n240), .SIN(dpc_tab[13]), .SMC(test_se), .C(
        net12481), .Q(dpc_tab[14]) );
  SDFFQX1 dpc_tab_reg_6__2_ ( .D(n240), .SIN(dpc_tab[37]), .SMC(test_se), .C(
        net12461), .Q(dpc_tab[38]) );
  SDFFQX1 rn_reg_reg_30__6_ ( .D(n228), .SIN(rn_reg[13]), .SMC(test_se), .C(
        net12656), .Q(rn_reg[14]) );
  SDFFQX1 rn_reg_reg_30__2_ ( .D(n240), .SIN(rn_reg[9]), .SMC(test_se), .C(
        net12656), .Q(rn_reg[10]) );
  SDFFQX1 rn_reg_reg_14__6_ ( .D(n228), .SIN(rn_reg[141]), .SMC(test_se), .C(
        net12576), .Q(rn_reg[142]) );
  SDFFQX1 rn_reg_reg_14__2_ ( .D(n240), .SIN(rn_reg[137]), .SMC(test_se), .C(
        net12576), .Q(rn_reg[138]) );
  SDFFQX1 rn_reg_reg_23__5_ ( .D(n233), .SIN(rn_reg[68]), .SMC(test_se), .C(
        net12621), .Q(rn_reg[69]) );
  SDFFQX1 dpc_tab_reg_3__3_ ( .D(N12690), .SIN(dpc_tab[20]), .SMC(test_se), 
        .C(net12476), .Q(dpc_tab[21]) );
  SDFFQX1 dpc_tab_reg_3__1_ ( .D(n247), .SIN(dpc_tab[18]), .SMC(test_se), .C(
        net12476), .Q(dpc_tab[19]) );
  SDFFQX1 dpc_tab_reg_7__3_ ( .D(N12690), .SIN(dpc_tab[44]), .SMC(test_se), 
        .C(net12456), .Q(dpc_tab[45]) );
  SDFFQX1 dpc_tab_reg_7__1_ ( .D(n247), .SIN(dpc_tab[42]), .SMC(test_se), .C(
        net12456), .Q(dpc_tab[43]) );
  SDFFQX1 rn_reg_reg_31__5_ ( .D(n233), .SIN(rn_reg[4]), .SMC(test_se), .C(
        net12661), .Q(rn_reg[5]) );
  SDFFQX1 rn_reg_reg_21__5_ ( .D(n232), .SIN(rn_reg[84]), .SMC(test_se), .C(
        net12611), .Q(rn_reg[85]) );
  SDFFQX1 rn_reg_reg_29__5_ ( .D(n232), .SIN(rn_reg[20]), .SMC(test_se), .C(
        net12651), .Q(rn_reg[21]) );
  SDFFQX1 rn_reg_reg_22__5_ ( .D(n231), .SIN(rn_reg[76]), .SMC(test_se), .C(
        net12616), .Q(rn_reg[77]) );
  SDFFQX1 dpc_tab_reg_2__3_ ( .D(n238), .SIN(dpc_tab[14]), .SMC(test_se), .C(
        net12481), .Q(dpc_tab[15]) );
  SDFFQX1 dpc_tab_reg_2__1_ ( .D(n244), .SIN(dpc_tab[12]), .SMC(test_se), .C(
        net12481), .Q(dpc_tab[13]) );
  SDFFQX1 dpc_tab_reg_6__3_ ( .D(n238), .SIN(dpc_tab[38]), .SMC(test_se), .C(
        net12461), .Q(dpc_tab[39]) );
  SDFFQX1 dpc_tab_reg_6__1_ ( .D(n244), .SIN(dpc_tab[36]), .SMC(test_se), .C(
        net12461), .Q(dpc_tab[37]) );
  SDFFQX1 rn_reg_reg_30__5_ ( .D(n231), .SIN(rn_reg[12]), .SMC(test_se), .C(
        net12656), .Q(rn_reg[13]) );
  SDFFQX1 rn_reg_reg_27__6_ ( .D(n230), .SIN(rn_reg[37]), .SMC(test_se), .C(
        net12641), .Q(rn_reg[38]) );
  SDFFQX1 rn_reg_reg_27__2_ ( .D(n243), .SIN(rn_reg[33]), .SMC(test_se), .C(
        net12641), .Q(rn_reg[34]) );
  SDFFQX1 rn_reg_reg_11__6_ ( .D(n230), .SIN(rn_reg[165]), .SMC(test_se), .C(
        net12561), .Q(rn_reg[166]) );
  SDFFQX1 rn_reg_reg_11__2_ ( .D(n243), .SIN(rn_reg[161]), .SMC(test_se), .C(
        net12561), .Q(rn_reg[162]) );
  SDFFQX1 rn_reg_reg_0__2_ ( .D(n243), .SIN(rn_reg[249]), .SMC(test_se), .C(
        net12506), .Q(rn_reg[250]) );
  SDFFQX1 rn_reg_reg_0__6_ ( .D(n230), .SIN(rn_reg[253]), .SMC(test_se), .C(
        net12506), .Q(rn_reg[254]) );
  SDFFQX1 rn_reg_reg_16__6_ ( .D(n230), .SIN(rn_reg[125]), .SMC(test_se), .C(
        net12586), .Q(rn_reg[126]) );
  SDFFQX1 rn_reg_reg_16__2_ ( .D(n242), .SIN(rn_reg[121]), .SMC(test_se), .C(
        net12586), .Q(rn_reg[122]) );
  SDFFQX1 dpc_tab_reg_0__2_ ( .D(n242), .SIN(dpc_tab[1]), .SMC(test_se), .C(
        net12491), .Q(dpc_tab[2]) );
  SDFFQX1 dpc_tab_reg_4__2_ ( .D(n242), .SIN(dpc_tab[25]), .SMC(test_se), .C(
        net12471), .Q(dpc_tab[26]) );
  SDFFQX1 rn_reg_reg_1__2_ ( .D(n242), .SIN(rn_reg[241]), .SMC(test_se), .C(
        net12511), .Q(rn_reg[242]) );
  SDFFQX1 rn_reg_reg_1__6_ ( .D(n229), .SIN(rn_reg[245]), .SMC(test_se), .C(
        net12511), .Q(rn_reg[246]) );
  SDFFQX1 rn_reg_reg_17__6_ ( .D(n229), .SIN(rn_reg[117]), .SMC(test_se), .C(
        net12591), .Q(rn_reg[118]) );
  SDFFQX1 rn_reg_reg_17__2_ ( .D(n241), .SIN(rn_reg[113]), .SMC(test_se), .C(
        net12591), .Q(rn_reg[114]) );
  SDFFQX1 dpc_tab_reg_1__2_ ( .D(n241), .SIN(dpc_tab[7]), .SMC(test_se), .C(
        net12486), .Q(dpc_tab[8]) );
  SDFFQX1 dpc_tab_reg_5__2_ ( .D(n241), .SIN(dpc_tab[31]), .SMC(test_se), .C(
        net12466), .Q(dpc_tab[32]) );
  SDFFQX1 rn_reg_reg_25__2_ ( .D(n241), .SIN(rn_reg[49]), .SMC(test_se), .C(
        net12631), .Q(rn_reg[50]) );
  SDFFQX1 rn_reg_reg_9__6_ ( .D(n229), .SIN(rn_reg[181]), .SMC(test_se), .C(
        net12551), .Q(rn_reg[182]) );
  SDFFQX1 rn_reg_reg_9__2_ ( .D(n241), .SIN(rn_reg[177]), .SMC(test_se), .C(
        net12551), .Q(rn_reg[178]) );
  SDFFQX1 rn_reg_reg_2__2_ ( .D(n241), .SIN(rn_reg[233]), .SMC(test_se), .C(
        net12516), .Q(rn_reg[234]) );
  SDFFQX1 rn_reg_reg_2__6_ ( .D(n228), .SIN(rn_reg[237]), .SMC(test_se), .C(
        net12516), .Q(rn_reg[238]) );
  SDFFQX1 rn_reg_reg_18__6_ ( .D(n228), .SIN(rn_reg[109]), .SMC(test_se), .C(
        net12596), .Q(rn_reg[110]) );
  SDFFQX1 rn_reg_reg_18__2_ ( .D(n240), .SIN(rn_reg[105]), .SMC(test_se), .C(
        net12596), .Q(rn_reg[106]) );
  SDFFQX1 rn_reg_reg_26__6_ ( .D(n228), .SIN(rn_reg[45]), .SMC(test_se), .C(
        net12636), .Q(rn_reg[46]) );
  SDFFQX1 rn_reg_reg_26__2_ ( .D(n240), .SIN(rn_reg[41]), .SMC(test_se), .C(
        net12636), .Q(rn_reg[42]) );
  SDFFQX1 rn_reg_reg_10__6_ ( .D(n228), .SIN(rn_reg[173]), .SMC(test_se), .C(
        net12556), .Q(rn_reg[174]) );
  SDFFQX1 rn_reg_reg_10__2_ ( .D(n240), .SIN(rn_reg[169]), .SMC(test_se), .C(
        net12556), .Q(rn_reg[170]) );
  SDFFQX1 rn_reg_reg_27__5_ ( .D(n233), .SIN(rn_reg[36]), .SMC(test_se), .C(
        net12641), .Q(rn_reg[37]) );
  SDFFQX1 rn_reg_reg_0__5_ ( .D(n233), .SIN(rn_reg[252]), .SMC(test_se), .C(
        net12506), .Q(rn_reg[253]) );
  SDFFQX1 rn_reg_reg_16__5_ ( .D(n233), .SIN(rn_reg[124]), .SMC(test_se), .C(
        net12586), .Q(rn_reg[125]) );
  SDFFQX1 dpc_tab_reg_0__3_ ( .D(n239), .SIN(dpc_tab[2]), .SMC(test_se), .C(
        net12491), .Q(dpc_tab[3]) );
  SDFFQX1 dpc_tab_reg_0__1_ ( .D(n246), .SIN(dpc_tab[0]), .SMC(test_se), .C(
        net12491), .Q(dpc_tab[1]) );
  SDFFQX1 dpc_tab_reg_4__3_ ( .D(n239), .SIN(dpc_tab[26]), .SMC(test_se), .C(
        net12471), .Q(dpc_tab[27]) );
  SDFFQX1 dpc_tab_reg_4__1_ ( .D(n246), .SIN(dpc_tab[24]), .SMC(test_se), .C(
        net12471), .Q(dpc_tab[25]) );
  SDFFQX1 rn_reg_reg_1__5_ ( .D(n232), .SIN(rn_reg[244]), .SMC(test_se), .C(
        net12511), .Q(rn_reg[245]) );
  SDFFQX1 rn_reg_reg_17__5_ ( .D(n232), .SIN(rn_reg[116]), .SMC(test_se), .C(
        net12591), .Q(rn_reg[117]) );
  SDFFQX1 rn_reg_reg_17__0_ ( .D(n249), .SIN(rn_reg[127]), .SMC(test_se), .C(
        net12591), .Q(rn_reg[112]) );
  SDFFQX1 dpc_tab_reg_1__3_ ( .D(N12690), .SIN(dpc_tab[8]), .SMC(test_se), .C(
        net12486), .Q(dpc_tab[9]) );
  SDFFQX1 dpc_tab_reg_1__1_ ( .D(n245), .SIN(dpc_tab[6]), .SMC(test_se), .C(
        net12486), .Q(dpc_tab[7]) );
  SDFFQX1 dpc_tab_reg_5__3_ ( .D(N12690), .SIN(dpc_tab[32]), .SMC(test_se), 
        .C(net12466), .Q(dpc_tab[33]) );
  SDFFQX1 dpc_tab_reg_5__1_ ( .D(n245), .SIN(dpc_tab[30]), .SMC(test_se), .C(
        net12466), .Q(dpc_tab[31]) );
  SDFFQX1 rn_reg_reg_25__6_ ( .D(n228), .SIN(rn_reg[53]), .SMC(test_se), .C(
        net12631), .Q(rn_reg[54]) );
  SDFFQX1 rn_reg_reg_25__5_ ( .D(n232), .SIN(rn_reg[52]), .SMC(test_se), .C(
        net12631), .Q(rn_reg[53]) );
  SDFFQX1 rn_reg_reg_9__5_ ( .D(n232), .SIN(rn_reg[180]), .SMC(test_se), .C(
        net12551), .Q(rn_reg[181]) );
  SDFFQX1 rn_reg_reg_18__5_ ( .D(n231), .SIN(rn_reg[108]), .SMC(test_se), .C(
        net12596), .Q(rn_reg[109]) );
  SDFFQX1 rn_reg_reg_26__5_ ( .D(n231), .SIN(rn_reg[44]), .SMC(test_se), .C(
        net12636), .Q(rn_reg[45]) );
  SDFFQX1 rn_reg_reg_3__2_ ( .D(n1872), .SIN(rn_reg[225]), .SMC(test_se), .C(
        net12521), .Q(rn_reg[226]) );
  SDFFQX1 rn_reg_reg_3__6_ ( .D(n1778), .SIN(rn_reg[229]), .SMC(test_se), .C(
        net12521), .Q(rn_reg[230]) );
  SDFFQX1 rn_reg_reg_19__6_ ( .D(n1778), .SIN(rn_reg[101]), .SMC(test_se), .C(
        net12601), .Q(rn_reg[102]) );
  SDFFQX1 rn_reg_reg_19__2_ ( .D(n243), .SIN(rn_reg[97]), .SMC(test_se), .C(
        net12601), .Q(rn_reg[98]) );
  SDFFQX1 rn_reg_reg_3__5_ ( .D(n1779), .SIN(rn_reg[228]), .SMC(test_se), .C(
        net12521), .Q(rn_reg[229]) );
  SDFFQX1 rn_reg_reg_19__5_ ( .D(n1779), .SIN(rn_reg[100]), .SMC(test_se), .C(
        net12601), .Q(rn_reg[101]) );
  SDFFQX1 rn_reg_reg_24__6_ ( .D(n230), .SIN(rn_reg[61]), .SMC(test_se), .C(
        net12626), .Q(rn_reg[62]) );
  SDFFQX1 rn_reg_reg_24__2_ ( .D(n242), .SIN(rn_reg[57]), .SMC(test_se), .C(
        net12626), .Q(rn_reg[58]) );
  SDFFQX1 rn_reg_reg_8__6_ ( .D(n229), .SIN(rn_reg[189]), .SMC(test_se), .C(
        net12546), .Q(rn_reg[190]) );
  SDFFQX1 rn_reg_reg_8__2_ ( .D(n242), .SIN(rn_reg[185]), .SMC(test_se), .C(
        net12546), .Q(rn_reg[186]) );
  SDFFQX1 rn_reg_reg_28__6_ ( .D(n229), .SIN(rn_reg[29]), .SMC(test_se), .C(
        net12646), .Q(rn_reg[30]) );
  SDFFQX1 rn_reg_reg_28__2_ ( .D(n242), .SIN(rn_reg[25]), .SMC(test_se), .C(
        net12646), .Q(rn_reg[26]) );
  SDFFQX1 rn_reg_reg_12__6_ ( .D(n229), .SIN(rn_reg[157]), .SMC(test_se), .C(
        net12566), .Q(rn_reg[158]) );
  SDFFQX1 rn_reg_reg_12__2_ ( .D(n242), .SIN(rn_reg[153]), .SMC(test_se), .C(
        net12566), .Q(rn_reg[154]) );
  SDFFQX1 rn_reg_reg_28__5_ ( .D(n232), .SIN(rn_reg[28]), .SMC(test_se), .C(
        net12646), .Q(rn_reg[29]) );
  SDFFQX1 rn_reg_reg_4__2_ ( .D(n242), .SIN(rn_reg[217]), .SMC(test_se), .C(
        net12526), .Q(rn_reg[218]) );
  SDFFQX1 rn_reg_reg_4__6_ ( .D(n230), .SIN(rn_reg[221]), .SMC(test_se), .C(
        net12526), .Q(rn_reg[222]) );
  SDFFQX1 rn_reg_reg_20__6_ ( .D(n230), .SIN(rn_reg[93]), .SMC(test_se), .C(
        net12606), .Q(rn_reg[94]) );
  SDFFQX1 rn_reg_reg_20__2_ ( .D(n242), .SIN(rn_reg[89]), .SMC(test_se), .C(
        net12606), .Q(rn_reg[90]) );
  SDFFQX1 rn_reg_reg_20__5_ ( .D(n233), .SIN(rn_reg[92]), .SMC(test_se), .C(
        net12606), .Q(rn_reg[93]) );
  SDFFQX1 dec_cop_reg_5_ ( .D(N10587), .SIN(dec_cop[4]), .SMC(test_se), .C(
        net12400), .Q(dec_cop[5]) );
  SDFFQX1 dpl_reg_reg_3__3_ ( .D(N12596), .SIN(dpl_reg[26]), .SMC(test_se), 
        .C(net12436), .Q(dpl_reg[27]) );
  SDFFQX1 dph_reg_reg_3__1_ ( .D(N12522), .SIN(dph_reg[24]), .SMC(test_se), 
        .C(net12436), .Q(dph_reg[25]) );
  SDFFQX1 dpl_reg_reg_7__3_ ( .D(N12632), .SIN(dpl_reg[58]), .SMC(test_se), 
        .C(net12416), .Q(dpl_reg[59]) );
  SDFFQX1 dph_reg_reg_3__7_ ( .D(N12528), .SIN(dph_reg[30]), .SMC(test_se), 
        .C(net12436), .Q(dph_reg[31]) );
  SDFFQX1 dph_reg_reg_7__7_ ( .D(N12564), .SIN(dph_reg[62]), .SMC(test_se), 
        .C(net12416), .Q(dph_reg[63]) );
  SDFFQX1 dph_reg_reg_7__1_ ( .D(N12558), .SIN(dph_reg[56]), .SMC(test_se), 
        .C(net12416), .Q(dph_reg[57]) );
  SDFFQX1 dpl_reg_reg_2__3_ ( .D(N12587), .SIN(dpl_reg[18]), .SMC(test_se), 
        .C(net12441), .Q(dpl_reg[19]) );
  SDFFQX1 dpl_reg_reg_1__3_ ( .D(N12578), .SIN(dpl_reg[10]), .SMC(test_se), 
        .C(net12446), .Q(dpl_reg[11]) );
  SDFFQX1 dpl_reg_reg_5__3_ ( .D(N12614), .SIN(dpl_reg[42]), .SMC(test_se), 
        .C(net12426), .Q(dpl_reg[43]) );
  SDFFQX1 dph_reg_reg_2__1_ ( .D(N12513), .SIN(dph_reg[16]), .SMC(test_se), 
        .C(net12441), .Q(dph_reg[17]) );
  SDFFQX1 dpl_reg_reg_6__3_ ( .D(N12623), .SIN(dpl_reg[50]), .SMC(test_se), 
        .C(net12421), .Q(dpl_reg[51]) );
  SDFFQX1 dph_reg_reg_1__7_ ( .D(N12510), .SIN(dph_reg[14]), .SMC(test_se), 
        .C(net12446), .Q(dph_reg[15]) );
  SDFFQX1 dph_reg_reg_1__1_ ( .D(N12504), .SIN(dph_reg[8]), .SMC(test_se), .C(
        net12446), .Q(dph_reg[9]) );
  SDFFQX1 dph_reg_reg_5__7_ ( .D(N12546), .SIN(dph_reg[46]), .SMC(test_se), 
        .C(net12426), .Q(dph_reg[47]) );
  SDFFQX1 dph_reg_reg_5__1_ ( .D(N12540), .SIN(dph_reg[40]), .SMC(test_se), 
        .C(net12426), .Q(dph_reg[41]) );
  SDFFQX1 dph_reg_reg_2__7_ ( .D(N12519), .SIN(dph_reg[22]), .SMC(test_se), 
        .C(net12441), .Q(dph_reg[23]) );
  SDFFQX1 dph_reg_reg_6__7_ ( .D(N12555), .SIN(dph_reg[54]), .SMC(test_se), 
        .C(net12421), .Q(dph_reg[55]) );
  SDFFQX1 dph_reg_reg_6__1_ ( .D(N12549), .SIN(dph_reg[48]), .SMC(test_se), 
        .C(net12421), .Q(dph_reg[49]) );
  SDFFQX1 dpl_reg_reg_0__3_ ( .D(N12569), .SIN(dpl_reg[2]), .SMC(test_se), .C(
        net12451), .Q(dpl_reg[3]) );
  SDFFQX1 dpl_reg_reg_4__3_ ( .D(N12605), .SIN(dpl_reg[34]), .SMC(test_se), 
        .C(net12431), .Q(dpl_reg[35]) );
  SDFFQX1 dph_reg_reg_0__7_ ( .D(N12501), .SIN(dph_reg[6]), .SMC(test_se), .C(
        net12451), .Q(dph_reg[7]) );
  SDFFQX1 dph_reg_reg_0__1_ ( .D(N12495), .SIN(dph_reg[0]), .SMC(test_se), .C(
        net12451), .Q(dph_reg[1]) );
  SDFFQX1 dph_reg_reg_4__7_ ( .D(N12537), .SIN(dph_reg[38]), .SMC(test_se), 
        .C(net12431), .Q(dph_reg[39]) );
  SDFFQX1 dph_reg_reg_4__1_ ( .D(N12531), .SIN(dph_reg[32]), .SMC(test_se), 
        .C(net12431), .Q(dph_reg[33]) );
  SDFFQX1 gf0_reg ( .D(n1881), .SIN(finishmul), .SMC(test_se), .C(net12400), 
        .Q(gf0) );
  SDFFQX1 dec_cop_reg_7_ ( .D(N10589), .SIN(dec_cop[6]), .SMC(test_se), .C(
        net12400), .Q(dec_cop[7]) );
  SDFFQX1 ckcon_r_reg_7_ ( .D(N12972), .SIN(ckcon[6]), .SMC(test_se), .C(
        net12400), .Q(ckcon[7]) );
  SDFFQX1 ckcon_r_reg_3_ ( .D(N12968), .SIN(ckcon[2]), .SMC(test_se), .C(
        net12400), .Q(ckcon[3]) );
  SDFFQX1 p2sel_s_reg ( .D(N520), .SIN(p2[7]), .SMC(test_se), .C(net12400), 
        .Q(p2sel) );
  SDFFQX1 p2_reg_reg_3_ ( .D(N12488), .SIN(p2[2]), .SMC(test_se), .C(net12400), 
        .Q(p2[3]) );
  SDFFQX1 dec_cop_reg_6_ ( .D(N10588), .SIN(dec_cop[5]), .SMC(test_se), .C(
        net12400), .Q(dec_cop[6]) );
  SDFFQX1 idle_s_reg ( .D(n1879), .SIN(idle_r), .SMC(test_se), .C(net12400), 
        .Q(idle) );
  SDFFQX1 bitno_reg_2_ ( .D(n1740), .SIN(N344), .SMC(test_se), .C(net12411), 
        .Q(N345) );
  SDFFQX1 p2_reg_reg_0_ ( .D(N12485), .SIN(ov), .SMC(test_se), .C(net12400), 
        .Q(p2[0]) );
  SDFFQX1 dpc_tab_reg_3__5_ ( .D(n1779), .SIN(dpc_tab[22]), .SMC(test_se), .C(
        net12476), .Q(dpc_tab[23]) );
  SDFFQX1 dpc_tab_reg_3__4_ ( .D(N12691), .SIN(dpc_tab[21]), .SMC(test_se), 
        .C(net12476), .Q(dpc_tab[22]) );
  SDFFQX1 dpc_tab_reg_7__5_ ( .D(N12692), .SIN(dpc_tab[46]), .SMC(test_se), 
        .C(net12456), .Q(dpc_tab[47]) );
  SDFFQX1 dpc_tab_reg_2__5_ ( .D(n1779), .SIN(dpc_tab[16]), .SMC(test_se), .C(
        net12481), .Q(dpc_tab[17]) );
  SDFFQX1 dpc_tab_reg_2__4_ ( .D(N12691), .SIN(dpc_tab[15]), .SMC(test_se), 
        .C(net12481), .Q(dpc_tab[16]) );
  SDFFQX1 dpc_tab_reg_6__5_ ( .D(N12692), .SIN(dpc_tab[40]), .SMC(test_se), 
        .C(net12461), .Q(dpc_tab[41]) );
  SDFFQX1 rn_reg_reg_7__7_ ( .D(n225), .SIN(rn_reg[198]), .SMC(test_se), .C(
        net12541), .Q(rn_reg[199]) );
  SDFFQX1 rn_reg_reg_23__7_ ( .D(n225), .SIN(rn_reg[70]), .SMC(test_se), .C(
        net12621), .Q(rn_reg[71]) );
  SDFFQX1 dpc_tab_reg_3__0_ ( .D(n1874), .SIN(dpc_tab[17]), .SMC(test_se), .C(
        net12476), .Q(dpc_tab[18]) );
  SDFFQX1 dpc_tab_reg_7__4_ ( .D(N12691), .SIN(dpc_tab[45]), .SMC(test_se), 
        .C(net12456), .Q(dpc_tab[46]) );
  SDFFQX1 dpc_tab_reg_7__0_ ( .D(n251), .SIN(dpc_tab[41]), .SMC(test_se), .C(
        net12456), .Q(dpc_tab[42]) );
  SDFFQX1 rn_reg_reg_31__7_ ( .D(n225), .SIN(rn_reg[6]), .SMC(test_se), .C(
        net12661), .Q(rn_reg[7]) );
  SDFFQX1 rn_reg_reg_15__7_ ( .D(n225), .SIN(rn_reg[134]), .SMC(test_se), .C(
        net12581), .Q(rn_reg[135]) );
  SDFFQX1 rn_reg_reg_5__7_ ( .D(n226), .SIN(rn_reg[214]), .SMC(test_se), .C(
        net12531), .Q(rn_reg[215]) );
  SDFFQX1 rn_reg_reg_21__7_ ( .D(n226), .SIN(rn_reg[86]), .SMC(test_se), .C(
        net12611), .Q(rn_reg[87]) );
  SDFFQX1 rn_reg_reg_29__7_ ( .D(n227), .SIN(rn_reg[22]), .SMC(test_se), .C(
        net12651), .Q(rn_reg[23]) );
  SDFFQX1 rn_reg_reg_13__7_ ( .D(n227), .SIN(rn_reg[150]), .SMC(test_se), .C(
        net12571), .Q(rn_reg[151]) );
  SDFFQX1 rn_reg_reg_6__7_ ( .D(n227), .SIN(rn_reg[206]), .SMC(test_se), .C(
        net12536), .Q(rn_reg[207]) );
  SDFFQX1 rn_reg_reg_22__7_ ( .D(n227), .SIN(rn_reg[78]), .SMC(test_se), .C(
        net12616), .Q(rn_reg[79]) );
  SDFFQX1 dpc_tab_reg_2__0_ ( .D(n251), .SIN(dpc_tab[11]), .SMC(test_se), .C(
        net12481), .Q(dpc_tab[12]) );
  SDFFQX1 dpc_tab_reg_6__4_ ( .D(N12691), .SIN(dpc_tab[39]), .SMC(test_se), 
        .C(net12461), .Q(dpc_tab[40]) );
  SDFFQX1 dpc_tab_reg_6__0_ ( .D(n251), .SIN(dpc_tab[35]), .SMC(test_se), .C(
        net12461), .Q(dpc_tab[36]) );
  SDFFQX1 rn_reg_reg_30__7_ ( .D(n227), .SIN(rn_reg[14]), .SMC(test_se), .C(
        net12656), .Q(rn_reg[15]) );
  SDFFQX1 rn_reg_reg_14__7_ ( .D(n1772), .SIN(rn_reg[142]), .SMC(test_se), .C(
        net12576), .Q(rn_reg[143]) );
  SDFFQX1 rn_reg_reg_7__3_ ( .D(n1783), .SIN(rn_reg[194]), .SMC(test_se), .C(
        net12541), .Q(rn_reg[195]) );
  SDFFQX1 rn_reg_reg_7__1_ ( .D(n247), .SIN(rn_reg[192]), .SMC(test_se), .C(
        net12541), .Q(rn_reg[193]) );
  SDFFQX1 rn_reg_reg_7__0_ ( .D(n251), .SIN(rn_reg[207]), .SMC(test_se), .C(
        net12541), .Q(rn_reg[192]) );
  SDFFQX1 rn_reg_reg_7__4_ ( .D(n1782), .SIN(rn_reg[195]), .SMC(test_se), .C(
        net12541), .Q(rn_reg[196]) );
  SDFFQX1 rn_reg_reg_7__5_ ( .D(n1779), .SIN(rn_reg[196]), .SMC(test_se), .C(
        net12541), .Q(rn_reg[197]) );
  SDFFQX1 rn_reg_reg_23__4_ ( .D(n236), .SIN(rn_reg[67]), .SMC(test_se), .C(
        net12621), .Q(rn_reg[68]) );
  SDFFQX1 rn_reg_reg_23__3_ ( .D(n1783), .SIN(rn_reg[66]), .SMC(test_se), .C(
        net12621), .Q(rn_reg[67]) );
  SDFFQX1 rn_reg_reg_23__1_ ( .D(n247), .SIN(rn_reg[64]), .SMC(test_se), .C(
        net12621), .Q(rn_reg[65]) );
  SDFFQX1 rn_reg_reg_23__0_ ( .D(n250), .SIN(rn_reg[79]), .SMC(test_se), .C(
        net12621), .Q(rn_reg[64]) );
  SDFFQX1 rn_reg_reg_31__4_ ( .D(n236), .SIN(rn_reg[3]), .SMC(test_se), .C(
        net12661), .Q(rn_reg[4]) );
  SDFFQX1 rn_reg_reg_31__3_ ( .D(n1783), .SIN(rn_reg[2]), .SMC(test_se), .C(
        net12661), .Q(rn_reg[3]) );
  SDFFQX1 rn_reg_reg_31__1_ ( .D(n247), .SIN(rn_reg[0]), .SMC(test_se), .C(
        net12661), .Q(rn_reg[1]) );
  SDFFQX1 rn_reg_reg_31__0_ ( .D(n250), .SIN(rn_reg[15]), .SMC(test_se), .C(
        net12661), .Q(rn_reg[0]) );
  SDFFQX1 rn_reg_reg_15__5_ ( .D(n233), .SIN(rn_reg[132]), .SMC(test_se), .C(
        net12581), .Q(rn_reg[133]) );
  SDFFQX1 rn_reg_reg_15__4_ ( .D(n236), .SIN(rn_reg[131]), .SMC(test_se), .C(
        net12581), .Q(rn_reg[132]) );
  SDFFQX1 rn_reg_reg_15__3_ ( .D(n1783), .SIN(rn_reg[130]), .SMC(test_se), .C(
        net12581), .Q(rn_reg[131]) );
  SDFFQX1 rn_reg_reg_15__1_ ( .D(n247), .SIN(rn_reg[128]), .SMC(test_se), .C(
        net12581), .Q(rn_reg[129]) );
  SDFFQX1 rn_reg_reg_15__0_ ( .D(n250), .SIN(rn_reg[143]), .SMC(test_se), .C(
        net12581), .Q(rn_reg[128]) );
  SDFFQX1 rn_reg_reg_5__3_ ( .D(n239), .SIN(rn_reg[210]), .SMC(test_se), .C(
        net12531), .Q(rn_reg[211]) );
  SDFFQX1 rn_reg_reg_5__1_ ( .D(n245), .SIN(rn_reg[208]), .SMC(test_se), .C(
        net12531), .Q(rn_reg[209]) );
  SDFFQX1 rn_reg_reg_5__0_ ( .D(n249), .SIN(rn_reg[223]), .SMC(test_se), .C(
        net12531), .Q(rn_reg[208]) );
  SDFFQX1 rn_reg_reg_5__4_ ( .D(n235), .SIN(rn_reg[211]), .SMC(test_se), .C(
        net12531), .Q(rn_reg[212]) );
  SDFFQX1 rn_reg_reg_5__5_ ( .D(n232), .SIN(rn_reg[212]), .SMC(test_se), .C(
        net12531), .Q(rn_reg[213]) );
  SDFFQX1 rn_reg_reg_21__4_ ( .D(n235), .SIN(rn_reg[83]), .SMC(test_se), .C(
        net12611), .Q(rn_reg[84]) );
  SDFFQX1 rn_reg_reg_21__1_ ( .D(n245), .SIN(rn_reg[80]), .SMC(test_se), .C(
        net12611), .Q(rn_reg[81]) );
  SDFFQX1 rn_reg_reg_21__0_ ( .D(n249), .SIN(rn_reg[95]), .SMC(test_se), .C(
        net12611), .Q(rn_reg[80]) );
  SDFFQX1 rn_reg_reg_29__4_ ( .D(n235), .SIN(rn_reg[19]), .SMC(test_se), .C(
        net12651), .Q(rn_reg[20]) );
  SDFFQX1 rn_reg_reg_29__1_ ( .D(n245), .SIN(rn_reg[16]), .SMC(test_se), .C(
        net12651), .Q(rn_reg[17]) );
  SDFFQX1 rn_reg_reg_29__0_ ( .D(n249), .SIN(rn_reg[31]), .SMC(test_se), .C(
        net12651), .Q(rn_reg[16]) );
  SDFFQX1 rn_reg_reg_13__5_ ( .D(n231), .SIN(rn_reg[148]), .SMC(test_se), .C(
        net12571), .Q(rn_reg[149]) );
  SDFFQX1 rn_reg_reg_13__4_ ( .D(n234), .SIN(rn_reg[147]), .SMC(test_se), .C(
        net12571), .Q(rn_reg[148]) );
  SDFFQX1 rn_reg_reg_13__3_ ( .D(n239), .SIN(rn_reg[146]), .SMC(test_se), .C(
        net12571), .Q(rn_reg[147]) );
  SDFFQX1 rn_reg_reg_13__1_ ( .D(n245), .SIN(rn_reg[144]), .SMC(test_se), .C(
        net12571), .Q(rn_reg[145]) );
  SDFFQX1 rn_reg_reg_13__0_ ( .D(n248), .SIN(rn_reg[159]), .SMC(test_se), .C(
        net12571), .Q(rn_reg[144]) );
  SDFFQX1 rn_reg_reg_6__3_ ( .D(n238), .SIN(rn_reg[202]), .SMC(test_se), .C(
        net12536), .Q(rn_reg[203]) );
  SDFFQX1 rn_reg_reg_6__1_ ( .D(n244), .SIN(rn_reg[200]), .SMC(test_se), .C(
        net12536), .Q(rn_reg[201]) );
  SDFFQX1 rn_reg_reg_6__0_ ( .D(n248), .SIN(rn_reg[215]), .SMC(test_se), .C(
        net12536), .Q(rn_reg[200]) );
  SDFFQX1 rn_reg_reg_6__4_ ( .D(n234), .SIN(rn_reg[203]), .SMC(test_se), .C(
        net12536), .Q(rn_reg[204]) );
  SDFFQX1 rn_reg_reg_6__5_ ( .D(n231), .SIN(rn_reg[204]), .SMC(test_se), .C(
        net12536), .Q(rn_reg[205]) );
  SDFFQX1 rn_reg_reg_22__4_ ( .D(n234), .SIN(rn_reg[75]), .SMC(test_se), .C(
        net12616), .Q(rn_reg[76]) );
  SDFFQX1 rn_reg_reg_22__3_ ( .D(n238), .SIN(rn_reg[74]), .SMC(test_se), .C(
        net12616), .Q(rn_reg[75]) );
  SDFFQX1 rn_reg_reg_22__1_ ( .D(n244), .SIN(rn_reg[72]), .SMC(test_se), .C(
        net12616), .Q(rn_reg[73]) );
  SDFFQX1 rn_reg_reg_22__0_ ( .D(n248), .SIN(rn_reg[87]), .SMC(test_se), .C(
        net12616), .Q(rn_reg[72]) );
  SDFFQX1 rn_reg_reg_30__4_ ( .D(n234), .SIN(rn_reg[11]), .SMC(test_se), .C(
        net12656), .Q(rn_reg[12]) );
  SDFFQX1 rn_reg_reg_30__3_ ( .D(n238), .SIN(rn_reg[10]), .SMC(test_se), .C(
        net12656), .Q(rn_reg[11]) );
  SDFFQX1 rn_reg_reg_30__1_ ( .D(n244), .SIN(rn_reg[8]), .SMC(test_se), .C(
        net12656), .Q(rn_reg[9]) );
  SDFFQX1 rn_reg_reg_30__0_ ( .D(n248), .SIN(rn_reg[23]), .SMC(test_se), .C(
        net12656), .Q(rn_reg[8]) );
  SDFFQX1 rn_reg_reg_14__5_ ( .D(n231), .SIN(rn_reg[140]), .SMC(test_se), .C(
        net12576), .Q(rn_reg[141]) );
  SDFFQX1 rn_reg_reg_14__4_ ( .D(n234), .SIN(rn_reg[139]), .SMC(test_se), .C(
        net12576), .Q(rn_reg[140]) );
  SDFFQX1 rn_reg_reg_14__3_ ( .D(n238), .SIN(rn_reg[138]), .SMC(test_se), .C(
        net12576), .Q(rn_reg[139]) );
  SDFFQX1 rn_reg_reg_14__1_ ( .D(n244), .SIN(rn_reg[136]), .SMC(test_se), .C(
        net12576), .Q(rn_reg[137]) );
  SDFFQX1 rn_reg_reg_14__0_ ( .D(n248), .SIN(rn_reg[151]), .SMC(test_se), .C(
        net12576), .Q(rn_reg[136]) );
  SDFFQX1 rn_reg_reg_21__3_ ( .D(n237), .SIN(rn_reg[82]), .SMC(test_se), .C(
        net12611), .Q(rn_reg[83]) );
  SDFFQX1 rn_reg_reg_29__3_ ( .D(n237), .SIN(rn_reg[18]), .SMC(test_se), .C(
        net12651), .Q(rn_reg[19]) );
  SDFFQX1 dpc_tab_reg_0__5_ ( .D(n1779), .SIN(dpc_tab[4]), .SMC(test_se), .C(
        net12491), .Q(dpc_tab[5]) );
  SDFFQX1 dpc_tab_reg_0__4_ ( .D(n1782), .SIN(dpc_tab[3]), .SMC(test_se), .C(
        net12491), .Q(dpc_tab[4]) );
  SDFFQX1 dpc_tab_reg_4__5_ ( .D(N12692), .SIN(dpc_tab[28]), .SMC(test_se), 
        .C(net12471), .Q(dpc_tab[29]) );
  SDFFQX1 dpc_tab_reg_1__5_ ( .D(n1779), .SIN(dpc_tab[10]), .SMC(test_se), .C(
        net12486), .Q(dpc_tab[11]) );
  SDFFQX1 rn_reg_reg_27__7_ ( .D(n225), .SIN(rn_reg[38]), .SMC(test_se), .C(
        net12641), .Q(rn_reg[39]) );
  SDFFQX1 rn_reg_reg_11__7_ ( .D(n225), .SIN(rn_reg[166]), .SMC(test_se), .C(
        net12561), .Q(rn_reg[167]) );
  SDFFQX1 rn_reg_reg_0__7_ ( .D(n225), .SIN(rn_reg[254]), .SMC(test_se), .C(
        net12506), .Q(rn_reg[255]) );
  SDFFQX1 rn_reg_reg_16__7_ ( .D(n226), .SIN(rn_reg[126]), .SMC(test_se), .C(
        net12586), .Q(rn_reg[127]) );
  SDFFQX1 dpc_tab_reg_0__0_ ( .D(n251), .SIN(divtempreg[6]), .SMC(test_se), 
        .C(net12491), .Q(dpc_tab[0]) );
  SDFFQX1 dpc_tab_reg_4__4_ ( .D(n1782), .SIN(dpc_tab[27]), .SMC(test_se), .C(
        net12471), .Q(dpc_tab[28]) );
  SDFFQX1 dpc_tab_reg_4__0_ ( .D(n251), .SIN(dpc_tab[23]), .SMC(test_se), .C(
        net12471), .Q(dpc_tab[24]) );
  SDFFQX1 rn_reg_reg_1__7_ ( .D(n226), .SIN(rn_reg[246]), .SMC(test_se), .C(
        net12511), .Q(rn_reg[247]) );
  SDFFQX1 rn_reg_reg_17__7_ ( .D(n226), .SIN(rn_reg[118]), .SMC(test_se), .C(
        net12591), .Q(rn_reg[119]) );
  SDFFQX1 dpc_tab_reg_1__4_ ( .D(n1782), .SIN(dpc_tab[9]), .SMC(test_se), .C(
        net12486), .Q(dpc_tab[10]) );
  SDFFQX1 dpc_tab_reg_1__0_ ( .D(n251), .SIN(dpc_tab[5]), .SMC(test_se), .C(
        net12486), .Q(dpc_tab[6]) );
  SDFFQX1 dpc_tab_reg_5__5_ ( .D(N12692), .SIN(dpc_tab[34]), .SMC(test_se), 
        .C(net12466), .Q(dpc_tab[35]) );
  SDFFQX1 dpc_tab_reg_5__4_ ( .D(n1782), .SIN(dpc_tab[33]), .SMC(test_se), .C(
        net12466), .Q(dpc_tab[34]) );
  SDFFQX1 dpc_tab_reg_5__0_ ( .D(n251), .SIN(dpc_tab[29]), .SMC(test_se), .C(
        net12466), .Q(dpc_tab[30]) );
  SDFFQX1 rn_reg_reg_25__7_ ( .D(n227), .SIN(rn_reg[54]), .SMC(test_se), .C(
        net12631), .Q(rn_reg[55]) );
  SDFFQX1 rn_reg_reg_9__7_ ( .D(n227), .SIN(rn_reg[182]), .SMC(test_se), .C(
        net12551), .Q(rn_reg[183]) );
  SDFFQX1 rn_reg_reg_2__7_ ( .D(n227), .SIN(rn_reg[238]), .SMC(test_se), .C(
        net12516), .Q(rn_reg[239]) );
  SDFFQX1 rn_reg_reg_18__7_ ( .D(n227), .SIN(rn_reg[110]), .SMC(test_se), .C(
        net12596), .Q(rn_reg[111]) );
  SDFFQX1 rn_reg_reg_26__7_ ( .D(n227), .SIN(rn_reg[46]), .SMC(test_se), .C(
        net12636), .Q(rn_reg[47]) );
  SDFFQX1 rn_reg_reg_10__7_ ( .D(n1772), .SIN(rn_reg[174]), .SMC(test_se), .C(
        net12556), .Q(rn_reg[175]) );
  SDFFQX1 rn_reg_reg_27__4_ ( .D(n236), .SIN(rn_reg[35]), .SMC(test_se), .C(
        net12641), .Q(rn_reg[36]) );
  SDFFQX1 rn_reg_reg_27__1_ ( .D(n247), .SIN(rn_reg[32]), .SMC(test_se), .C(
        net12641), .Q(rn_reg[33]) );
  SDFFQX1 rn_reg_reg_27__0_ ( .D(n250), .SIN(rn_reg[47]), .SMC(test_se), .C(
        net12641), .Q(rn_reg[32]) );
  SDFFQX1 rn_reg_reg_11__5_ ( .D(n233), .SIN(rn_reg[164]), .SMC(test_se), .C(
        net12561), .Q(rn_reg[165]) );
  SDFFQX1 rn_reg_reg_11__4_ ( .D(n236), .SIN(rn_reg[163]), .SMC(test_se), .C(
        net12561), .Q(rn_reg[164]) );
  SDFFQX1 rn_reg_reg_11__3_ ( .D(n1783), .SIN(rn_reg[162]), .SMC(test_se), .C(
        net12561), .Q(rn_reg[163]) );
  SDFFQX1 rn_reg_reg_11__1_ ( .D(n247), .SIN(rn_reg[160]), .SMC(test_se), .C(
        net12561), .Q(rn_reg[161]) );
  SDFFQX1 rn_reg_reg_11__0_ ( .D(n250), .SIN(rn_reg[175]), .SMC(test_se), .C(
        net12561), .Q(rn_reg[160]) );
  SDFFQX1 rn_reg_reg_0__3_ ( .D(n1783), .SIN(rn_reg[250]), .SMC(test_se), .C(
        net12506), .Q(rn_reg[251]) );
  SDFFQX1 rn_reg_reg_0__1_ ( .D(n247), .SIN(rn_reg[248]), .SMC(test_se), .C(
        net12506), .Q(rn_reg[249]) );
  SDFFQX1 rn_reg_reg_0__0_ ( .D(n250), .SIN(rmwinstr), .SMC(test_se), .C(
        net12506), .Q(rn_reg[248]) );
  SDFFQX1 rn_reg_reg_0__4_ ( .D(n236), .SIN(rn_reg[251]), .SMC(test_se), .C(
        net12506), .Q(rn_reg[252]) );
  SDFFQX1 rn_reg_reg_16__4_ ( .D(n236), .SIN(rn_reg[123]), .SMC(test_se), .C(
        net12586), .Q(rn_reg[124]) );
  SDFFQX1 rn_reg_reg_16__1_ ( .D(n246), .SIN(rn_reg[120]), .SMC(test_se), .C(
        net12586), .Q(rn_reg[121]) );
  SDFFQX1 rn_reg_reg_16__0_ ( .D(n250), .SIN(rn_reg[135]), .SMC(test_se), .C(
        net12586), .Q(rn_reg[120]) );
  SDFFQX1 rn_reg_reg_1__3_ ( .D(n239), .SIN(rn_reg[242]), .SMC(test_se), .C(
        net12511), .Q(rn_reg[243]) );
  SDFFQX1 rn_reg_reg_1__1_ ( .D(n246), .SIN(rn_reg[240]), .SMC(test_se), .C(
        net12511), .Q(rn_reg[241]) );
  SDFFQX1 rn_reg_reg_1__0_ ( .D(n249), .SIN(rn_reg[255]), .SMC(test_se), .C(
        net12511), .Q(rn_reg[240]) );
  SDFFQX1 rn_reg_reg_1__4_ ( .D(n235), .SIN(rn_reg[243]), .SMC(test_se), .C(
        net12511), .Q(rn_reg[244]) );
  SDFFQX1 rn_reg_reg_17__4_ ( .D(n235), .SIN(rn_reg[115]), .SMC(test_se), .C(
        net12591), .Q(rn_reg[116]) );
  SDFFQX1 rn_reg_reg_17__1_ ( .D(n245), .SIN(rn_reg[112]), .SMC(test_se), .C(
        net12591), .Q(rn_reg[113]) );
  SDFFQX1 rn_reg_reg_25__4_ ( .D(n235), .SIN(rn_reg[51]), .SMC(test_se), .C(
        net12631), .Q(rn_reg[52]) );
  SDFFQX1 rn_reg_reg_25__1_ ( .D(n245), .SIN(rn_reg[48]), .SMC(test_se), .C(
        net12631), .Q(rn_reg[49]) );
  SDFFQX1 rn_reg_reg_25__0_ ( .D(n249), .SIN(rn_reg[63]), .SMC(test_se), .C(
        net12631), .Q(rn_reg[48]) );
  SDFFQX1 rn_reg_reg_9__4_ ( .D(n235), .SIN(rn_reg[179]), .SMC(test_se), .C(
        net12551), .Q(rn_reg[180]) );
  SDFFQX1 rn_reg_reg_9__3_ ( .D(n239), .SIN(rn_reg[178]), .SMC(test_se), .C(
        net12551), .Q(rn_reg[179]) );
  SDFFQX1 rn_reg_reg_9__1_ ( .D(n245), .SIN(rn_reg[176]), .SMC(test_se), .C(
        net12551), .Q(rn_reg[177]) );
  SDFFQX1 rn_reg_reg_9__0_ ( .D(n249), .SIN(rn_reg[191]), .SMC(test_se), .C(
        net12551), .Q(rn_reg[176]) );
  SDFFQX1 rn_reg_reg_2__3_ ( .D(n239), .SIN(rn_reg[234]), .SMC(test_se), .C(
        net12516), .Q(rn_reg[235]) );
  SDFFQX1 rn_reg_reg_2__1_ ( .D(n245), .SIN(rn_reg[232]), .SMC(test_se), .C(
        net12516), .Q(rn_reg[233]) );
  SDFFQX1 rn_reg_reg_2__0_ ( .D(n248), .SIN(rn_reg[247]), .SMC(test_se), .C(
        net12516), .Q(rn_reg[232]) );
  SDFFQX1 rn_reg_reg_2__4_ ( .D(n234), .SIN(rn_reg[235]), .SMC(test_se), .C(
        net12516), .Q(rn_reg[236]) );
  SDFFQX1 rn_reg_reg_2__5_ ( .D(n231), .SIN(rn_reg[236]), .SMC(test_se), .C(
        net12516), .Q(rn_reg[237]) );
  SDFFQX1 rn_reg_reg_18__4_ ( .D(n234), .SIN(rn_reg[107]), .SMC(test_se), .C(
        net12596), .Q(rn_reg[108]) );
  SDFFQX1 rn_reg_reg_18__1_ ( .D(n244), .SIN(rn_reg[104]), .SMC(test_se), .C(
        net12596), .Q(rn_reg[105]) );
  SDFFQX1 rn_reg_reg_18__0_ ( .D(n248), .SIN(rn_reg[119]), .SMC(test_se), .C(
        net12596), .Q(rn_reg[104]) );
  SDFFQX1 rn_reg_reg_26__4_ ( .D(n234), .SIN(rn_reg[43]), .SMC(test_se), .C(
        net12636), .Q(rn_reg[44]) );
  SDFFQX1 rn_reg_reg_26__1_ ( .D(n244), .SIN(rn_reg[40]), .SMC(test_se), .C(
        net12636), .Q(rn_reg[41]) );
  SDFFQX1 rn_reg_reg_26__0_ ( .D(n248), .SIN(rn_reg[55]), .SMC(test_se), .C(
        net12636), .Q(rn_reg[40]) );
  SDFFQX1 rn_reg_reg_10__5_ ( .D(n231), .SIN(rn_reg[172]), .SMC(test_se), .C(
        net12556), .Q(rn_reg[173]) );
  SDFFQX1 rn_reg_reg_10__4_ ( .D(n234), .SIN(rn_reg[171]), .SMC(test_se), .C(
        net12556), .Q(rn_reg[172]) );
  SDFFQX1 rn_reg_reg_10__3_ ( .D(n238), .SIN(rn_reg[170]), .SMC(test_se), .C(
        net12556), .Q(rn_reg[171]) );
  SDFFQX1 rn_reg_reg_10__1_ ( .D(n244), .SIN(rn_reg[168]), .SMC(test_se), .C(
        net12556), .Q(rn_reg[169]) );
  SDFFQX1 rn_reg_reg_10__0_ ( .D(n248), .SIN(rn_reg[183]), .SMC(test_se), .C(
        net12556), .Q(rn_reg[168]) );
  SDFFQX1 rn_reg_reg_27__3_ ( .D(n238), .SIN(rn_reg[34]), .SMC(test_se), .C(
        net12641), .Q(rn_reg[35]) );
  SDFFQX1 rn_reg_reg_16__3_ ( .D(n238), .SIN(rn_reg[122]), .SMC(test_se), .C(
        net12586), .Q(rn_reg[123]) );
  SDFFQX1 rn_reg_reg_17__3_ ( .D(n237), .SIN(rn_reg[114]), .SMC(test_se), .C(
        net12591), .Q(rn_reg[115]) );
  SDFFQX1 rn_reg_reg_25__3_ ( .D(n237), .SIN(rn_reg[50]), .SMC(test_se), .C(
        net12631), .Q(rn_reg[51]) );
  SDFFQX1 rn_reg_reg_18__3_ ( .D(n237), .SIN(rn_reg[106]), .SMC(test_se), .C(
        net12596), .Q(rn_reg[107]) );
  SDFFQX1 rn_reg_reg_26__3_ ( .D(n237), .SIN(rn_reg[42]), .SMC(test_se), .C(
        net12636), .Q(rn_reg[43]) );
  SDFFQX1 rn_reg_reg_3__7_ ( .D(n225), .SIN(rn_reg[230]), .SMC(test_se), .C(
        net12521), .Q(rn_reg[231]) );
  SDFFQX1 rn_reg_reg_19__7_ ( .D(n225), .SIN(rn_reg[102]), .SMC(test_se), .C(
        net12601), .Q(rn_reg[103]) );
  SDFFQX1 rn_reg_reg_3__3_ ( .D(n1783), .SIN(rn_reg[226]), .SMC(test_se), .C(
        net12521), .Q(rn_reg[227]) );
  SDFFQX1 rn_reg_reg_3__1_ ( .D(n1873), .SIN(rn_reg[224]), .SMC(test_se), .C(
        net12521), .Q(rn_reg[225]) );
  SDFFQX1 rn_reg_reg_3__0_ ( .D(n251), .SIN(rn_reg[239]), .SMC(test_se), .C(
        net12521), .Q(rn_reg[224]) );
  SDFFQX1 rn_reg_reg_3__4_ ( .D(n1782), .SIN(rn_reg[227]), .SMC(test_se), .C(
        net12521), .Q(rn_reg[228]) );
  SDFFQX1 rn_reg_reg_19__4_ ( .D(n1782), .SIN(rn_reg[99]), .SMC(test_se), .C(
        net12601), .Q(rn_reg[100]) );
  SDFFQX1 rn_reg_reg_19__1_ ( .D(n247), .SIN(rn_reg[96]), .SMC(test_se), .C(
        net12601), .Q(rn_reg[97]) );
  SDFFQX1 rn_reg_reg_19__0_ ( .D(n251), .SIN(rn_reg[111]), .SMC(test_se), .C(
        net12601), .Q(rn_reg[96]) );
  SDFFQX1 rn_reg_reg_19__3_ ( .D(n238), .SIN(rn_reg[98]), .SMC(test_se), .C(
        net12601), .Q(rn_reg[99]) );
  SDFFQX1 rn_reg_reg_24__7_ ( .D(n226), .SIN(rn_reg[62]), .SMC(test_se), .C(
        net12626), .Q(rn_reg[63]) );
  SDFFQX1 rn_reg_reg_8__7_ ( .D(n226), .SIN(rn_reg[190]), .SMC(test_se), .C(
        net12546), .Q(rn_reg[191]) );
  SDFFQX1 rn_reg_reg_24__5_ ( .D(n233), .SIN(rn_reg[60]), .SMC(test_se), .C(
        net12626), .Q(rn_reg[61]) );
  SDFFQX1 rn_reg_reg_24__1_ ( .D(n246), .SIN(rn_reg[56]), .SMC(test_se), .C(
        net12626), .Q(rn_reg[57]) );
  SDFFQX1 rn_reg_reg_24__0_ ( .D(n250), .SIN(rn_reg[71]), .SMC(test_se), .C(
        net12626), .Q(rn_reg[56]) );
  SDFFQX1 rn_reg_reg_8__5_ ( .D(n232), .SIN(rn_reg[188]), .SMC(test_se), .C(
        net12546), .Q(rn_reg[189]) );
  SDFFQX1 rn_reg_reg_8__1_ ( .D(n246), .SIN(rn_reg[184]), .SMC(test_se), .C(
        net12546), .Q(rn_reg[185]) );
  SDFFQX1 rn_reg_reg_8__0_ ( .D(n249), .SIN(rn_reg[199]), .SMC(test_se), .C(
        net12546), .Q(rn_reg[184]) );
  SDFFQX1 rn_reg_reg_28__7_ ( .D(n226), .SIN(rn_reg[30]), .SMC(test_se), .C(
        net12646), .Q(rn_reg[31]) );
  SDFFQX1 rn_reg_reg_12__7_ ( .D(n226), .SIN(rn_reg[158]), .SMC(test_se), .C(
        net12566), .Q(rn_reg[159]) );
  SDFFQX1 rn_reg_reg_28__4_ ( .D(n235), .SIN(rn_reg[27]), .SMC(test_se), .C(
        net12646), .Q(rn_reg[28]) );
  SDFFQX1 rn_reg_reg_28__1_ ( .D(n246), .SIN(rn_reg[24]), .SMC(test_se), .C(
        net12646), .Q(rn_reg[25]) );
  SDFFQX1 rn_reg_reg_28__0_ ( .D(n249), .SIN(rn_reg[39]), .SMC(test_se), .C(
        net12646), .Q(rn_reg[24]) );
  SDFFQX1 rn_reg_reg_12__5_ ( .D(n232), .SIN(rn_reg[156]), .SMC(test_se), .C(
        net12566), .Q(rn_reg[157]) );
  SDFFQX1 rn_reg_reg_12__1_ ( .D(n246), .SIN(rn_reg[152]), .SMC(test_se), .C(
        net12566), .Q(rn_reg[153]) );
  SDFFQX1 rn_reg_reg_12__0_ ( .D(n249), .SIN(rn_reg[167]), .SMC(test_se), .C(
        net12566), .Q(rn_reg[152]) );
  SDFFQX1 rn_reg_reg_4__7_ ( .D(n225), .SIN(rn_reg[222]), .SMC(test_se), .C(
        net12526), .Q(rn_reg[223]) );
  SDFFQX1 rn_reg_reg_20__7_ ( .D(n226), .SIN(rn_reg[94]), .SMC(test_se), .C(
        net12606), .Q(rn_reg[95]) );
  SDFFQX1 rn_reg_reg_4__3_ ( .D(n239), .SIN(rn_reg[218]), .SMC(test_se), .C(
        net12526), .Q(rn_reg[219]) );
  SDFFQX1 rn_reg_reg_4__1_ ( .D(n246), .SIN(rn_reg[216]), .SMC(test_se), .C(
        net12526), .Q(rn_reg[217]) );
  SDFFQX1 rn_reg_reg_4__0_ ( .D(n250), .SIN(rn_reg[231]), .SMC(test_se), .C(
        net12526), .Q(rn_reg[216]) );
  SDFFQX1 rn_reg_reg_4__4_ ( .D(n236), .SIN(rn_reg[219]), .SMC(test_se), .C(
        net12526), .Q(rn_reg[220]) );
  SDFFQX1 rn_reg_reg_4__5_ ( .D(n233), .SIN(rn_reg[220]), .SMC(test_se), .C(
        net12526), .Q(rn_reg[221]) );
  SDFFQX1 rn_reg_reg_20__4_ ( .D(n236), .SIN(rn_reg[91]), .SMC(test_se), .C(
        net12606), .Q(rn_reg[92]) );
  SDFFQX1 rn_reg_reg_20__1_ ( .D(n246), .SIN(rn_reg[88]), .SMC(test_se), .C(
        net12606), .Q(rn_reg[89]) );
  SDFFQX1 rn_reg_reg_20__0_ ( .D(n250), .SIN(rn_reg[103]), .SMC(test_se), .C(
        net12606), .Q(rn_reg[88]) );
  SDFFQX1 sp_reg_reg_7_ ( .D(N12704), .SIN(sp[6]), .SMC(test_se), .C(net12400), 
        .Q(sp[7]) );
  SDFFQX1 dph_reg_reg_3__6_ ( .D(N12527), .SIN(dph_reg[29]), .SMC(test_se), 
        .C(net12436), .Q(dph_reg[30]) );
  SDFFQX1 dph_reg_reg_3__3_ ( .D(N12524), .SIN(dph_reg[26]), .SMC(test_se), 
        .C(net12436), .Q(dph_reg[27]) );
  SDFFQX1 dph_reg_reg_3__2_ ( .D(N12523), .SIN(dph_reg[25]), .SMC(test_se), 
        .C(net12436), .Q(dph_reg[26]) );
  SDFFQX1 dpl_reg_reg_3__5_ ( .D(N12598), .SIN(dpl_reg[28]), .SMC(test_se), 
        .C(net12436), .Q(dpl_reg[29]) );
  SDFFQX1 dpl_reg_reg_3__2_ ( .D(N12595), .SIN(dpl_reg[25]), .SMC(test_se), 
        .C(net12436), .Q(dpl_reg[26]) );
  SDFFQX1 dph_reg_reg_7__6_ ( .D(N12563), .SIN(dph_reg[61]), .SMC(test_se), 
        .C(net12416), .Q(dph_reg[62]) );
  SDFFQX1 dph_reg_reg_7__5_ ( .D(N12562), .SIN(dph_reg[60]), .SMC(test_se), 
        .C(net12416), .Q(dph_reg[61]) );
  SDFFQX1 dph_reg_reg_7__2_ ( .D(N12559), .SIN(dph_reg[57]), .SMC(test_se), 
        .C(net12416), .Q(dph_reg[58]) );
  SDFFQX1 dpl_reg_reg_7__5_ ( .D(N12634), .SIN(dpl_reg[60]), .SMC(test_se), 
        .C(net12416), .Q(dpl_reg[61]) );
  SDFFQX1 dpl_reg_reg_7__4_ ( .D(N12633), .SIN(dpl_reg[59]), .SMC(test_se), 
        .C(net12416), .Q(dpl_reg[60]) );
  SDFFQX1 dpl_reg_reg_7__2_ ( .D(N12631), .SIN(dpl_reg[57]), .SMC(test_se), 
        .C(net12416), .Q(dpl_reg[58]) );
  SDFFQX1 dph_reg_reg_7__0_ ( .D(N12557), .SIN(dph_reg[55]), .SMC(test_se), 
        .C(net12416), .Q(dph_reg[56]) );
  SDFFQX1 dph_reg_reg_3__0_ ( .D(N12521), .SIN(dph_reg[23]), .SMC(test_se), 
        .C(net12436), .Q(dph_reg[24]) );
  SDFFQX1 dpl_reg_reg_3__7_ ( .D(N12600), .SIN(dpl_reg[30]), .SMC(test_se), 
        .C(net12436), .Q(dpl_reg[31]) );
  SDFFQX1 dpl_reg_reg_3__6_ ( .D(N12599), .SIN(dpl_reg[29]), .SMC(test_se), 
        .C(net12436), .Q(dpl_reg[30]) );
  SDFFQX1 dpl_reg_reg_3__1_ ( .D(N12594), .SIN(dpl_reg[24]), .SMC(test_se), 
        .C(net12436), .Q(dpl_reg[25]) );
  SDFFQX1 dpl_reg_reg_3__0_ ( .D(N12593), .SIN(dpl_reg[23]), .SMC(test_se), 
        .C(net12436), .Q(dpl_reg[24]) );
  SDFFQX1 dph_reg_reg_7__3_ ( .D(N12560), .SIN(dph_reg[58]), .SMC(test_se), 
        .C(net12416), .Q(dph_reg[59]) );
  SDFFQX1 dpl_reg_reg_7__7_ ( .D(N12636), .SIN(dpl_reg[62]), .SMC(test_se), 
        .C(net12416), .Q(dpl_reg[63]) );
  SDFFQX1 dpl_reg_reg_7__6_ ( .D(N12635), .SIN(dpl_reg[61]), .SMC(test_se), 
        .C(net12416), .Q(dpl_reg[62]) );
  SDFFQX1 dpl_reg_reg_7__1_ ( .D(N12630), .SIN(dpl_reg[56]), .SMC(test_se), 
        .C(net12416), .Q(dpl_reg[57]) );
  SDFFQX1 dpl_reg_reg_7__0_ ( .D(N12629), .SIN(dpl_reg[55]), .SMC(test_se), 
        .C(net12416), .Q(dpl_reg[56]) );
  SDFFQX1 dph_reg_reg_1__6_ ( .D(N12509), .SIN(dph_reg[13]), .SMC(test_se), 
        .C(net12446), .Q(dph_reg[14]) );
  SDFFQX1 dph_reg_reg_1__5_ ( .D(N12508), .SIN(dph_reg[12]), .SMC(test_se), 
        .C(net12446), .Q(dph_reg[13]) );
  SDFFQX1 dph_reg_reg_1__2_ ( .D(N12505), .SIN(dph_reg[9]), .SMC(test_se), .C(
        net12446), .Q(dph_reg[10]) );
  SDFFQX1 dpl_reg_reg_1__5_ ( .D(N12580), .SIN(dpl_reg[12]), .SMC(test_se), 
        .C(net12446), .Q(dpl_reg[13]) );
  SDFFQX1 dpl_reg_reg_1__4_ ( .D(N12579), .SIN(dpl_reg[11]), .SMC(test_se), 
        .C(net12446), .Q(dpl_reg[12]) );
  SDFFQX1 dpl_reg_reg_1__2_ ( .D(N12577), .SIN(dpl_reg[9]), .SMC(test_se), .C(
        net12446), .Q(dpl_reg[10]) );
  SDFFQX1 dph_reg_reg_5__6_ ( .D(N12545), .SIN(dph_reg[45]), .SMC(test_se), 
        .C(net12426), .Q(dph_reg[46]) );
  SDFFQX1 dph_reg_reg_5__5_ ( .D(N12544), .SIN(dph_reg[44]), .SMC(test_se), 
        .C(net12426), .Q(dph_reg[45]) );
  SDFFQX1 dph_reg_reg_5__4_ ( .D(N12543), .SIN(dph_reg[43]), .SMC(test_se), 
        .C(net12426), .Q(dph_reg[44]) );
  SDFFQX1 dph_reg_reg_5__2_ ( .D(N12541), .SIN(dph_reg[41]), .SMC(test_se), 
        .C(net12426), .Q(dph_reg[42]) );
  SDFFQX1 dpl_reg_reg_5__5_ ( .D(N12616), .SIN(dpl_reg[44]), .SMC(test_se), 
        .C(net12426), .Q(dpl_reg[45]) );
  SDFFQX1 dpl_reg_reg_5__4_ ( .D(N12615), .SIN(dpl_reg[43]), .SMC(test_se), 
        .C(net12426), .Q(dpl_reg[44]) );
  SDFFQX1 dpl_reg_reg_5__2_ ( .D(N12613), .SIN(dpl_reg[41]), .SMC(test_se), 
        .C(net12426), .Q(dpl_reg[42]) );
  SDFFQX1 dph_reg_reg_5__0_ ( .D(N12539), .SIN(dph_reg[39]), .SMC(test_se), 
        .C(net12426), .Q(dph_reg[40]) );
  SDFFQX1 dph_reg_reg_1__0_ ( .D(N12503), .SIN(dph_reg[7]), .SMC(test_se), .C(
        net12446), .Q(dph_reg[8]) );
  SDFFQX1 dph_reg_reg_2__6_ ( .D(N12518), .SIN(dph_reg[21]), .SMC(test_se), 
        .C(net12441), .Q(dph_reg[22]) );
  SDFFQX1 dph_reg_reg_2__3_ ( .D(N12515), .SIN(dph_reg[18]), .SMC(test_se), 
        .C(net12441), .Q(dph_reg[19]) );
  SDFFQX1 dph_reg_reg_2__2_ ( .D(N12514), .SIN(dph_reg[17]), .SMC(test_se), 
        .C(net12441), .Q(dph_reg[18]) );
  SDFFQX1 dpl_reg_reg_2__5_ ( .D(N12589), .SIN(dpl_reg[20]), .SMC(test_se), 
        .C(net12441), .Q(dpl_reg[21]) );
  SDFFQX1 dpl_reg_reg_2__2_ ( .D(N12586), .SIN(dpl_reg[17]), .SMC(test_se), 
        .C(net12441), .Q(dpl_reg[18]) );
  SDFFQX1 dph_reg_reg_6__6_ ( .D(N12554), .SIN(dph_reg[53]), .SMC(test_se), 
        .C(net12421), .Q(dph_reg[54]) );
  SDFFQX1 dph_reg_reg_6__2_ ( .D(N12550), .SIN(dph_reg[49]), .SMC(test_se), 
        .C(net12421), .Q(dph_reg[50]) );
  SDFFQX1 dpl_reg_reg_6__5_ ( .D(N12625), .SIN(dpl_reg[52]), .SMC(test_se), 
        .C(net12421), .Q(dpl_reg[53]) );
  SDFFQX1 dpl_reg_reg_6__2_ ( .D(N12622), .SIN(dpl_reg[49]), .SMC(test_se), 
        .C(net12421), .Q(dpl_reg[50]) );
  SDFFQX1 dph_reg_reg_6__0_ ( .D(N12548), .SIN(dph_reg[47]), .SMC(test_se), 
        .C(net12421), .Q(dph_reg[48]) );
  SDFFQX1 dph_reg_reg_2__0_ ( .D(N12512), .SIN(dph_reg[15]), .SMC(test_se), 
        .C(net12441), .Q(dph_reg[16]) );
  SDFFQX1 dph_reg_reg_1__3_ ( .D(N12506), .SIN(dph_reg[10]), .SMC(test_se), 
        .C(net12446), .Q(dph_reg[11]) );
  SDFFQX1 dpl_reg_reg_1__7_ ( .D(N12582), .SIN(dpl_reg[14]), .SMC(test_se), 
        .C(net12446), .Q(dpl_reg[15]) );
  SDFFQX1 dpl_reg_reg_1__6_ ( .D(N12581), .SIN(dpl_reg[13]), .SMC(test_se), 
        .C(net12446), .Q(dpl_reg[14]) );
  SDFFQX1 dpl_reg_reg_1__1_ ( .D(N12576), .SIN(dpl_reg[8]), .SMC(test_se), .C(
        net12446), .Q(dpl_reg[9]) );
  SDFFQX1 dpl_reg_reg_1__0_ ( .D(N12575), .SIN(dpl_reg[7]), .SMC(test_se), .C(
        net12446), .Q(dpl_reg[8]) );
  SDFFQX1 dph_reg_reg_5__3_ ( .D(N12542), .SIN(dph_reg[42]), .SMC(test_se), 
        .C(net12426), .Q(dph_reg[43]) );
  SDFFQX1 dpl_reg_reg_5__7_ ( .D(N12618), .SIN(dpl_reg[46]), .SMC(test_se), 
        .C(net12426), .Q(dpl_reg[47]) );
  SDFFQX1 dpl_reg_reg_5__6_ ( .D(N12617), .SIN(dpl_reg[45]), .SMC(test_se), 
        .C(net12426), .Q(dpl_reg[46]) );
  SDFFQX1 dpl_reg_reg_5__1_ ( .D(N12612), .SIN(dpl_reg[40]), .SMC(test_se), 
        .C(net12426), .Q(dpl_reg[41]) );
  SDFFQX1 dpl_reg_reg_5__0_ ( .D(N12611), .SIN(dpl_reg[39]), .SMC(test_se), 
        .C(net12426), .Q(dpl_reg[40]) );
  SDFFQX1 dpl_reg_reg_2__7_ ( .D(N12591), .SIN(dpl_reg[22]), .SMC(test_se), 
        .C(net12441), .Q(dpl_reg[23]) );
  SDFFQX1 dpl_reg_reg_2__6_ ( .D(N12590), .SIN(dpl_reg[21]), .SMC(test_se), 
        .C(net12441), .Q(dpl_reg[22]) );
  SDFFQX1 dpl_reg_reg_2__1_ ( .D(N12585), .SIN(dpl_reg[16]), .SMC(test_se), 
        .C(net12441), .Q(dpl_reg[17]) );
  SDFFQX1 dpl_reg_reg_2__0_ ( .D(N12584), .SIN(dpl_reg[15]), .SMC(test_se), 
        .C(net12441), .Q(dpl_reg[16]) );
  SDFFQX1 dph_reg_reg_6__3_ ( .D(N12551), .SIN(dph_reg[50]), .SMC(test_se), 
        .C(net12421), .Q(dph_reg[51]) );
  SDFFQX1 dpl_reg_reg_6__7_ ( .D(N12627), .SIN(dpl_reg[54]), .SMC(test_se), 
        .C(net12421), .Q(dpl_reg[55]) );
  SDFFQX1 dpl_reg_reg_6__6_ ( .D(N12626), .SIN(dpl_reg[53]), .SMC(test_se), 
        .C(net12421), .Q(dpl_reg[54]) );
  SDFFQX1 dpl_reg_reg_6__1_ ( .D(N12621), .SIN(dpl_reg[48]), .SMC(test_se), 
        .C(net12421), .Q(dpl_reg[49]) );
  SDFFQX1 dpl_reg_reg_6__0_ ( .D(N12620), .SIN(dpl_reg[47]), .SMC(test_se), 
        .C(net12421), .Q(dpl_reg[48]) );
  SDFFQX1 dph_reg_reg_0__6_ ( .D(N12500), .SIN(dph_reg[5]), .SMC(test_se), .C(
        net12451), .Q(dph_reg[6]) );
  SDFFQX1 dph_reg_reg_0__5_ ( .D(N12499), .SIN(dph_reg[4]), .SMC(test_se), .C(
        net12451), .Q(dph_reg[5]) );
  SDFFQX1 dph_reg_reg_0__2_ ( .D(N12496), .SIN(dph_reg[1]), .SMC(test_se), .C(
        net12451), .Q(dph_reg[2]) );
  SDFFQX1 dpl_reg_reg_0__5_ ( .D(N12571), .SIN(dpl_reg[4]), .SMC(test_se), .C(
        net12451), .Q(dpl_reg[5]) );
  SDFFQX1 dpl_reg_reg_0__4_ ( .D(N12570), .SIN(dpl_reg[3]), .SMC(test_se), .C(
        net12451), .Q(dpl_reg[4]) );
  SDFFQX1 dpl_reg_reg_0__2_ ( .D(N12568), .SIN(dpl_reg[1]), .SMC(test_se), .C(
        net12451), .Q(dpl_reg[2]) );
  SDFFQX1 dph_reg_reg_4__6_ ( .D(N12536), .SIN(dph_reg[37]), .SMC(test_se), 
        .C(net12431), .Q(dph_reg[38]) );
  SDFFQX1 dph_reg_reg_4__5_ ( .D(N12535), .SIN(dph_reg[36]), .SMC(test_se), 
        .C(net12431), .Q(dph_reg[37]) );
  SDFFQX1 dph_reg_reg_4__4_ ( .D(N12534), .SIN(dph_reg[35]), .SMC(test_se), 
        .C(net12431), .Q(dph_reg[36]) );
  SDFFQX1 dph_reg_reg_4__2_ ( .D(N12532), .SIN(dph_reg[33]), .SMC(test_se), 
        .C(net12431), .Q(dph_reg[34]) );
  SDFFQX1 dpl_reg_reg_4__5_ ( .D(N12607), .SIN(dpl_reg[36]), .SMC(test_se), 
        .C(net12431), .Q(dpl_reg[37]) );
  SDFFQX1 dpl_reg_reg_4__4_ ( .D(N12606), .SIN(dpl_reg[35]), .SMC(test_se), 
        .C(net12431), .Q(dpl_reg[36]) );
  SDFFQX1 dpl_reg_reg_4__2_ ( .D(N12604), .SIN(dpl_reg[33]), .SMC(test_se), 
        .C(net12431), .Q(dpl_reg[34]) );
  SDFFQX1 dph_reg_reg_4__0_ ( .D(N12530), .SIN(dph_reg[31]), .SMC(test_se), 
        .C(net12431), .Q(dph_reg[32]) );
  SDFFQX1 dph_reg_reg_0__0_ ( .D(N12494), .SIN(dpc_tab[47]), .SMC(test_se), 
        .C(net12451), .Q(dph_reg[0]) );
  SDFFQX1 dph_reg_reg_0__3_ ( .D(N12497), .SIN(dph_reg[2]), .SMC(test_se), .C(
        net12451), .Q(dph_reg[3]) );
  SDFFQX1 dpl_reg_reg_0__7_ ( .D(N12573), .SIN(dpl_reg[6]), .SMC(test_se), .C(
        net12451), .Q(dpl_reg[7]) );
  SDFFQX1 dpl_reg_reg_0__6_ ( .D(N12572), .SIN(dpl_reg[5]), .SMC(test_se), .C(
        net12451), .Q(dpl_reg[6]) );
  SDFFQX1 dpl_reg_reg_0__1_ ( .D(N12567), .SIN(dpl_reg[0]), .SMC(test_se), .C(
        net12451), .Q(dpl_reg[1]) );
  SDFFQX1 dpl_reg_reg_0__0_ ( .D(N12566), .SIN(dph_reg[63]), .SMC(test_se), 
        .C(net12451), .Q(dpl_reg[0]) );
  SDFFQX1 dph_reg_reg_4__3_ ( .D(N12533), .SIN(dph_reg[34]), .SMC(test_se), 
        .C(net12431), .Q(dph_reg[35]) );
  SDFFQX1 dpl_reg_reg_4__7_ ( .D(N12609), .SIN(dpl_reg[38]), .SMC(test_se), 
        .C(net12431), .Q(dpl_reg[39]) );
  SDFFQX1 dpl_reg_reg_4__6_ ( .D(N12608), .SIN(dpl_reg[37]), .SMC(test_se), 
        .C(net12431), .Q(dpl_reg[38]) );
  SDFFQX1 dpl_reg_reg_4__1_ ( .D(N12603), .SIN(dpl_reg[32]), .SMC(test_se), 
        .C(net12431), .Q(dpl_reg[33]) );
  SDFFQX1 dpl_reg_reg_4__0_ ( .D(N12602), .SIN(dpl_reg[31]), .SMC(test_se), 
        .C(net12431), .Q(dpl_reg[32]) );
  SDFFQX1 sp_reg_reg_5_ ( .D(N12702), .SIN(sp[4]), .SMC(test_se), .C(net12400), 
        .Q(sp[5]) );
  SDFFQX1 sp_reg_reg_6_ ( .D(N12703), .SIN(sp[5]), .SMC(test_se), .C(net12400), 
        .Q(sp[6]) );
  SDFFQX1 dec_cop_reg_4_ ( .D(N10586), .SIN(dec_cop[3]), .SMC(test_se), .C(
        net12400), .Q(dec_cop[4]) );
  SDFFQX1 dec_cop_reg_2_ ( .D(N10584), .SIN(dec_cop[1]), .SMC(test_se), .C(
        net12400), .Q(dec_cop[2]) );
  SDFFQX1 dec_cop_reg_1_ ( .D(N10583), .SIN(dec_cop[0]), .SMC(test_se), .C(
        net12400), .Q(dec_cop[1]) );
  SDFFQX1 dec_cop_reg_3_ ( .D(N10585), .SIN(dec_cop[2]), .SMC(test_se), .C(
        net12400), .Q(dec_cop[3]) );
  SDFFQX1 pmw_reg_reg ( .D(n1756), .SIN(phase[5]), .SMC(test_se), .C(net12400), 
        .Q(pmw) );
  SDFFQX1 temp_reg_3_ ( .D(N12717), .SIN(temp[2]), .SMC(test_se), .C(net12496), 
        .Q(temp[3]) );
  SDFFQX1 temp_reg_7_ ( .D(N12721), .SIN(temp[6]), .SMC(test_se), .C(net12496), 
        .Q(temp[7]) );
  SDFFQX1 temp_reg_6_ ( .D(N12720), .SIN(temp[5]), .SMC(test_se), .C(net12496), 
        .Q(temp[6]) );
  SDFFQX1 temp_reg_0_ ( .D(N12714), .SIN(temp2_comb[7]), .SMC(test_se), .C(
        net12496), .Q(temp[0]) );
  SDFFQX1 temp2_reg_7_ ( .D(N12730), .SIN(temp2_comb[6]), .SMC(test_se), .C(
        net12400), .Q(temp2_comb[7]) );
  SDFFQX1 temp_reg_4_ ( .D(N12718), .SIN(temp[3]), .SMC(test_se), .C(net12496), 
        .Q(temp[4]) );
  SDFFQX1 temp_reg_5_ ( .D(N12719), .SIN(temp[4]), .SMC(test_se), .C(net12496), 
        .Q(temp[5]) );
  SDFFQX1 p2_reg_reg_2_ ( .D(N12487), .SIN(p2[1]), .SMC(test_se), .C(net12400), 
        .Q(p2[2]) );
  SDFFQX1 bitno_reg_1_ ( .D(n1751), .SIN(N343), .SMC(test_se), .C(net12411), 
        .Q(N344) );
  SDFFQX1 temp_reg_1_ ( .D(N12715), .SIN(temp[0]), .SMC(test_se), .C(net12496), 
        .Q(temp[1]) );
  SDFFQX1 ramdatao_r_reg_6_ ( .D(N11504), .SIN(ramdatao[5]), .SMC(test_se), 
        .C(net12400), .Q(ramdatao[6]) );
  SDFFQX1 temp_reg_2_ ( .D(N12716), .SIN(temp[1]), .SMC(test_se), .C(net12496), 
        .Q(temp[2]) );
  SDFFQX1 ramdatao_r_reg_7_ ( .D(N11505), .SIN(ramdatao[6]), .SMC(test_se), 
        .C(net12400), .Q(ramdatao[7]) );
  SDFFQX1 rmwinstr_reg ( .D(N690), .SIN(ramwe), .SMC(test_se), .C(net12400), 
        .Q(rmwinstr) );
  SDFFQX1 rn_reg_reg_24__4_ ( .D(n236), .SIN(rn_reg[59]), .SMC(test_se), .C(
        net12626), .Q(rn_reg[60]) );
  SDFFQX1 rn_reg_reg_8__4_ ( .D(n235), .SIN(rn_reg[187]), .SMC(test_se), .C(
        net12546), .Q(rn_reg[188]) );
  SDFFQX1 rn_reg_reg_8__3_ ( .D(n239), .SIN(rn_reg[186]), .SMC(test_se), .C(
        net12546), .Q(rn_reg[187]) );
  SDFFQX1 rn_reg_reg_24__3_ ( .D(n237), .SIN(rn_reg[58]), .SMC(test_se), .C(
        net12626), .Q(rn_reg[59]) );
  SDFFQX1 rn_reg_reg_12__4_ ( .D(n235), .SIN(rn_reg[155]), .SMC(test_se), .C(
        net12566), .Q(rn_reg[156]) );
  SDFFQX1 rn_reg_reg_12__3_ ( .D(n239), .SIN(rn_reg[154]), .SMC(test_se), .C(
        net12566), .Q(rn_reg[155]) );
  SDFFQX1 rn_reg_reg_28__3_ ( .D(n237), .SIN(rn_reg[26]), .SMC(test_se), .C(
        net12646), .Q(rn_reg[27]) );
  SDFFQX1 rn_reg_reg_20__3_ ( .D(n237), .SIN(rn_reg[90]), .SMC(test_se), .C(
        net12606), .Q(rn_reg[91]) );
  SDFFQX1 dph_reg_reg_3__5_ ( .D(N12526), .SIN(dph_reg[28]), .SMC(test_se), 
        .C(net12436), .Q(dph_reg[29]) );
  SDFFQX1 dph_reg_reg_3__4_ ( .D(N12525), .SIN(dph_reg[27]), .SMC(test_se), 
        .C(net12436), .Q(dph_reg[28]) );
  SDFFQX1 dpl_reg_reg_3__4_ ( .D(N12597), .SIN(dpl_reg[27]), .SMC(test_se), 
        .C(net12436), .Q(dpl_reg[28]) );
  SDFFQX1 dph_reg_reg_7__4_ ( .D(N12561), .SIN(dph_reg[59]), .SMC(test_se), 
        .C(net12416), .Q(dph_reg[60]) );
  SDFFQX1 dph_reg_reg_1__4_ ( .D(N12507), .SIN(dph_reg[11]), .SMC(test_se), 
        .C(net12446), .Q(dph_reg[12]) );
  SDFFQX1 dph_reg_reg_2__5_ ( .D(N12517), .SIN(dph_reg[20]), .SMC(test_se), 
        .C(net12441), .Q(dph_reg[21]) );
  SDFFQX1 dph_reg_reg_2__4_ ( .D(N12516), .SIN(dph_reg[19]), .SMC(test_se), 
        .C(net12441), .Q(dph_reg[20]) );
  SDFFQX1 dpl_reg_reg_2__4_ ( .D(N12588), .SIN(dpl_reg[19]), .SMC(test_se), 
        .C(net12441), .Q(dpl_reg[20]) );
  SDFFQX1 dph_reg_reg_6__5_ ( .D(N12553), .SIN(dph_reg[52]), .SMC(test_se), 
        .C(net12421), .Q(dph_reg[53]) );
  SDFFQX1 dph_reg_reg_6__4_ ( .D(N12552), .SIN(dph_reg[51]), .SMC(test_se), 
        .C(net12421), .Q(dph_reg[52]) );
  SDFFQX1 dpl_reg_reg_6__4_ ( .D(N12624), .SIN(dpl_reg[51]), .SMC(test_se), 
        .C(net12421), .Q(dpl_reg[52]) );
  SDFFQX1 sp_reg_reg_4_ ( .D(N12701), .SIN(sp[3]), .SMC(test_se), .C(net12400), 
        .Q(sp[4]) );
  SDFFQX1 dph_reg_reg_0__4_ ( .D(N12498), .SIN(dph_reg[3]), .SMC(test_se), .C(
        net12451), .Q(dph_reg[4]) );
  SDFFQX1 sp_reg_reg_3_ ( .D(N12700), .SIN(sp[2]), .SMC(test_se), .C(net12400), 
        .Q(sp[3]) );
  SDFFQX1 sp_reg_reg_2_ ( .D(N12699), .SIN(sp[1]), .SMC(test_se), .C(net12400), 
        .Q(sp[2]) );
  SDFFQX1 multempreg_reg_0_ ( .D(N13325), .SIN(memwr), .SMC(test_se), .C(
        net12666), .Q(multempreg[0]) );
  SDFFQX1 multempreg_reg_1_ ( .D(N13326), .SIN(multempreg[0]), .SMC(test_se), 
        .C(net12666), .Q(multempreg[1]) );
  SDFFQX1 dec_accop_reg_17_ ( .D(n1757), .SIN(dec_accop[16]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[17]) );
  SDFFQX1 phase_reg_2_ ( .D(N681), .SIN(n259), .SMC(test_se), .C(net12400), 
        .Q(phase[2]) );
  SDFFQX1 bitno_reg_0_ ( .D(n1752), .SIN(b[7]), .SMC(test_se), .C(net12411), 
        .Q(N343) );
  SDFFQX1 ramdatao_r_reg_5_ ( .D(N11503), .SIN(ramdatao[4]), .SMC(test_se), 
        .C(net12400), .Q(ramdatao[5]) );
  SDFFQX1 sp_reg_reg_0_ ( .D(N12697), .SIN(sfrwe_r), .SMC(test_se), .C(
        net12400), .Q(sp[0]) );
  SDFFQX1 dec_accop_reg_11_ ( .D(N10574), .SIN(dec_accop[10]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[11]) );
  SDFFQX1 sp_reg_reg_1_ ( .D(N12698), .SIN(sp[0]), .SMC(test_se), .C(net12400), 
        .Q(sp[1]) );
  SDFFQX1 dec_accop_reg_12_ ( .D(N10575), .SIN(dec_accop[11]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[12]) );
  SDFFQX1 ramwe_r_reg ( .D(N11487), .SIN(ramsfrwe), .SMC(test_se), .C(net12400), .Q(ramwe) );
  SDFFQX1 sfroe_r_reg ( .D(N11488), .SIN(rs[1]), .SMC(test_se), .C(net12400), 
        .Q(sfroe_r) );
  SDFFQX1 sfrwe_r_reg ( .D(N11489), .SIN(sfroe_r), .SMC(test_se), .C(net12400), 
        .Q(sfrwe_r) );
  SDFFQX1 mempsrd_r_reg ( .D(N582), .SIN(israccess), .SMC(test_se), .C(
        net12400), .Q(mempsrd) );
  SDFFQX1 dps_reg_reg_0_ ( .D(N12693), .SIN(dpl_reg[63]), .SMC(test_se), .C(
        net12400), .Q(dps[0]) );
  SDFFQX1 dps_reg_reg_1_ ( .D(N12694), .SIN(dps[0]), .SMC(test_se), .C(
        net12400), .Q(dps[1]) );
  SDFFQX1 temp2_reg_5_ ( .D(N12728), .SIN(temp2_comb[4]), .SMC(test_se), .C(
        net12400), .Q(temp2_comb[5]) );
  SDFFQX1 temp2_reg_6_ ( .D(N12729), .SIN(temp2_comb[5]), .SMC(test_se), .C(
        net12400), .Q(temp2_comb[6]) );
  SDFFQX1 ramdatao_r_reg_0_ ( .D(N11498), .SIN(pmw), .SMC(test_se), .C(
        net12400), .Q(ramdatao[0]) );
  SDFFQX1 dps_reg_reg_2_ ( .D(N12695), .SIN(dps[1]), .SMC(test_se), .C(
        net12400), .Q(n2482) );
  SDFFQX1 dec_accop_reg_14_ ( .D(N10577), .SIN(dec_accop[13]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[14]) );
  SDFFQX1 dec_accop_reg_2_ ( .D(N10565), .SIN(dec_accop[1]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[2]) );
  SDFFQX1 dec_accop_reg_3_ ( .D(N10566), .SIN(dec_accop[2]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[3]) );
  SDFFQX1 dec_accop_reg_4_ ( .D(N10567), .SIN(dec_accop[3]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[4]) );
  SDFFQX1 dec_accop_reg_1_ ( .D(N10564), .SIN(dec_accop[0]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[1]) );
  SDFFQX1 dec_accop_reg_15_ ( .D(N10578), .SIN(dec_accop[14]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[15]) );
  SDFFQX1 dec_accop_reg_13_ ( .D(N10576), .SIN(dec_accop[12]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[13]) );
  SDFFQX1 rs_reg_reg_1_ ( .D(N12710), .SIN(rs[0]), .SMC(test_se), .C(net12400), 
        .Q(rs[1]) );
  SDFFQX1 rs_reg_reg_0_ ( .D(N12709), .SIN(rn_reg[7]), .SMC(test_se), .C(
        net12400), .Q(rs[0]) );
  SDFFQX1 ckcon_r_reg_2_ ( .D(N12967), .SIN(ckcon[1]), .SMC(test_se), .C(
        net12400), .Q(ckcon[2]) );
  SDFFQX1 interrupt_reg ( .D(n2193), .SIN(instr[7]), .SMC(test_se), .C(
        net12406), .Q(interrupt) );
  SDFFQX1 dps_reg_reg_3_ ( .D(n1884), .SIN(dps[2]), .SMC(test_se), .C(net12400), .Q(dps[3]) );
  SDFFQX1 memrd_s_reg ( .D(N584), .SIN(mempswr), .SMC(test_se), .C(net12400), 
        .Q(memrd) );
  SDFFQX1 memwr_s_reg ( .D(N585), .SIN(memrd), .SMC(test_se), .C(net12400), 
        .Q(memwr) );
  SDFFQX1 ckcon_r_reg_6_ ( .D(N12971), .SIN(ckcon[5]), .SMC(test_se), .C(
        net12400), .Q(ckcon[6]) );
  SDFFQX1 temp2_reg_4_ ( .D(N12727), .SIN(temp2_comb[3]), .SMC(test_se), .C(
        net12400), .Q(temp2_comb[4]) );
  SDFFQX1 ramdatao_r_reg_4_ ( .D(N11502), .SIN(ramdatao[3]), .SMC(test_se), 
        .C(net12400), .Q(ramdatao[4]) );
  SDFFQX1 phase_reg_0_ ( .D(N679), .SIN(phase0_ff), .SMC(test_se), .C(net12400), .Q(phase[0]) );
  SDFFQX1 ramdatao_r_reg_3_ ( .D(N11501), .SIN(ramdatao[2]), .SMC(test_se), 
        .C(net12400), .Q(ramdatao[3]) );
  SDFFQX1 acc_reg_reg_4_ ( .D(n1902), .SIN(n126), .SMC(test_se), .C(net12400), 
        .Q(acc[4]) );
  SDFFQX1 mempswr_s_reg ( .D(N583), .SIN(mempsrd), .SMC(test_se), .C(net12400), 
        .Q(mempswr) );
  SDFFQX1 ramdatao_r_reg_1_ ( .D(N11499), .SIN(ramdatao[0]), .SMC(test_se), 
        .C(net12400), .Q(ramdatao[1]) );
  SDFFQX1 ramdatao_r_reg_2_ ( .D(N11500), .SIN(ramdatao[1]), .SMC(test_se), 
        .C(net12400), .Q(ramdatao[2]) );
  SDFFQX1 phase_reg_1_ ( .D(N680), .SIN(n254), .SMC(test_se), .C(net12400), 
        .Q(phase[1]) );
  SDFFQX1 instr_reg_4_ ( .D(N674), .SIN(instr[3]), .SMC(test_se), .C(net12406), 
        .Q(n2477) );
  SDFFQX1 dec_accop_reg_0_ ( .D(N10563), .SIN(d_hold), .SMC(test_se), .C(
        net12400), .Q(dec_accop[0]) );
  SDFFQX1 ckcon_r_reg_0_ ( .D(N12965), .SIN(c), .SMC(test_se), .C(net12400), 
        .Q(ckcon[0]) );
  SDFFQX1 ckcon_r_reg_4_ ( .D(N12969), .SIN(ckcon[3]), .SMC(test_se), .C(
        net12400), .Q(ckcon[4]) );
  SDFFQX1 ckcon_r_reg_5_ ( .D(N12970), .SIN(ckcon[4]), .SMC(test_se), .C(
        net12400), .Q(ckcon[5]) );
  SDFFQX1 ckcon_r_reg_1_ ( .D(N12966), .SIN(ckcon[0]), .SMC(test_se), .C(
        net12400), .Q(ckcon[1]) );
  SDFFQX1 waitcnt_reg_2_ ( .D(N12976), .SIN(waitcnt_1_), .SMC(test_se), .C(
        net12501), .Q(test_so) );
  SDFFQX1 waitcnt_reg_1_ ( .D(N12975), .SIN(waitcnt_0_), .SMC(test_se), .C(
        net12501), .Q(waitcnt_1_) );
  SDFFQX1 waitcnt_reg_0_ ( .D(N12974), .SIN(temp[7]), .SMC(test_se), .C(
        net12501), .Q(waitcnt_0_) );
  SDFFQX1 instr_reg_2_ ( .D(N672), .SIN(instr[1]), .SMC(test_se), .C(net12406), 
        .Q(instr[2]) );
  SDFFQX1 temp2_reg_3_ ( .D(N12726), .SIN(temp2_comb[2]), .SMC(test_se), .C(
        net12400), .Q(temp2_comb[3]) );
  SDFFQX1 temp2_reg_2_ ( .D(N12725), .SIN(temp2_comb[1]), .SMC(test_se), .C(
        net12400), .Q(temp2_comb[2]) );
  SDFFQX1 ramsfraddr_s_reg_5_ ( .D(N11483), .SIN(ramsfraddr[4]), .SMC(test_se), 
        .C(net12400), .Q(ramsfraddr[5]) );
  SDFFQX1 acc_reg_reg_5_ ( .D(n1901), .SIN(acc[4]), .SMC(test_se), .C(net12400), .Q(acc[5]) );
  SDFFQX1 instr_reg_1_ ( .D(N671), .SIN(instr[0]), .SMC(test_se), .C(net12406), 
        .Q(n2479) );
  SDFFQX1 instr_reg_7_ ( .D(N677), .SIN(instr[6]), .SMC(test_se), .C(net12406), 
        .Q(n2474) );
  SDFFQX1 instr_reg_0_ ( .D(N670), .SIN(idle), .SMC(test_se), .C(net12406), 
        .Q(n2480) );
  SDFFQX1 instr_reg_3_ ( .D(N673), .SIN(instr[2]), .SMC(test_se), .C(net12406), 
        .Q(n2478) );
  SDFFQX1 acc_reg_reg_6_ ( .D(n1900), .SIN(acc[5]), .SMC(test_se), .C(net12400), .Q(acc[6]) );
  SDFFQX1 accactv_reg ( .D(N10562), .SIN(acc[7]), .SMC(test_se), .C(net12400), 
        .Q(accactv) );
  SDFFQX1 ramsfrwe_reg ( .D(n1731), .SIN(ramsfraddr[7]), .SMC(test_se), .C(
        net12400), .Q(ramsfrwe) );
  SDFFQX1 divtempreg_reg_6_ ( .D(N13373), .SIN(divtempreg[5]), .SMC(test_se), 
        .C(net12671), .Q(divtempreg[6]) );
  SDFFQX1 temp2_reg_1_ ( .D(N12724), .SIN(temp2_comb[0]), .SMC(test_se), .C(
        net12400), .Q(temp2_comb[1]) );
  SDFFQX1 ramsfraddr_s_reg_1_ ( .D(N11479), .SIN(ramsfraddr[0]), .SMC(test_se), 
        .C(net12400), .Q(ramsfraddr[1]) );
  SDFFQX1 ramsfraddr_s_reg_4_ ( .D(N11482), .SIN(ramsfraddr[3]), .SMC(test_se), 
        .C(net12400), .Q(ramsfraddr[4]) );
  SDFFQX1 ramsfraddr_s_reg_7_ ( .D(n1736), .SIN(ramsfraddr[6]), .SMC(test_se), 
        .C(net12400), .Q(ramsfraddr[7]) );
  SDFFQX1 ramsfraddr_s_reg_0_ ( .D(N11478), .SIN(ramoe), .SMC(test_se), .C(
        net12400), .Q(ramsfraddr[0]) );
  SDFFQX1 ramsfraddr_s_reg_6_ ( .D(N11484), .SIN(ramsfraddr[5]), .SMC(test_se), 
        .C(net12400), .Q(ramsfraddr[6]) );
  SDFFQX1 ramsfraddr_s_reg_2_ ( .D(N11480), .SIN(ramsfraddr[1]), .SMC(test_se), 
        .C(net12400), .Q(ramsfraddr[2]) );
  SDFFQX1 ramsfraddr_s_reg_3_ ( .D(N11481), .SIN(ramsfraddr[2]), .SMC(test_se), 
        .C(net12400), .Q(ramsfraddr[3]) );
  SDFFQX1 b_reg_reg_7_ ( .D(N12484), .SIN(b[6]), .SMC(test_se), .C(net12400), 
        .Q(b[7]) );
  SDFFQX1 instr_reg_6_ ( .D(N676), .SIN(n2476), .SMC(test_se), .C(net12406), 
        .Q(n2475) );
  SDFFQX1 instr_reg_5_ ( .D(N675), .SIN(instr[4]), .SMC(test_se), .C(net12406), 
        .Q(n2476) );
  SDFFQX1 ac_reg_reg ( .D(N12706), .SIN(test_si), .SMC(test_se), .C(net12400), 
        .Q(ac) );
  SDFFQX1 divtempreg_reg_5_ ( .D(N13372), .SIN(divtempreg[4]), .SMC(test_se), 
        .C(net12671), .Q(divtempreg[5]) );
  SDFFQX1 temp2_reg_0_ ( .D(N12723), .SIN(stop), .SMC(test_se), .C(net12400), 
        .Q(temp2_comb[0]) );
  SDFFQX1 acc_reg_reg_0_ ( .D(N12469), .SIN(ac), .SMC(test_se), .C(net12400), 
        .Q(acc[0]) );
  SDFFQX1 acc_reg_reg_3_ ( .D(N12472), .SIN(acc[2]), .SMC(test_se), .C(
        net12400), .Q(acc[3]) );
  SDFFQX1 b_reg_reg_6_ ( .D(N12483), .SIN(b[5]), .SMC(test_se), .C(net12400), 
        .Q(b[6]) );
  SDFFQX1 dec_accop_reg_16_ ( .D(n1767), .SIN(dec_accop[15]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[16]) );
  SDFFQX1 divtempreg_reg_4_ ( .D(N13371), .SIN(divtempreg[3]), .SMC(test_se), 
        .C(net12671), .Q(divtempreg[4]) );
  SDFFQX1 divtempreg_reg_3_ ( .D(N13370), .SIN(divtempreg[2]), .SMC(test_se), 
        .C(net12671), .Q(divtempreg[3]) );
  SDFFQX1 dec_accop_reg_7_ ( .D(N10570), .SIN(dec_accop[6]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[7]) );
  SDFFQX1 dec_accop_reg_6_ ( .D(N10569), .SIN(dec_accop[5]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[6]) );
  SDFFQX1 dec_accop_reg_18_ ( .D(N10581), .SIN(dec_accop[17]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[18]) );
  SDFFQX1 dec_accop_reg_5_ ( .D(N10568), .SIN(dec_accop[4]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[5]) );
  SDFFQX1 acc_reg_reg_1_ ( .D(N12470), .SIN(n69), .SMC(test_se), .C(net12400), 
        .Q(acc[1]) );
  SDFFQX1 c_reg_reg ( .D(N12705), .SIN(N345), .SMC(test_se), .C(net12400), .Q(
        c) );
  SDFFQX1 acc_reg_reg_2_ ( .D(n1947), .SIN(acc[1]), .SMC(test_se), .C(net12400), .Q(acc[2]) );
  SDFFQX1 b_reg_reg_5_ ( .D(N12482), .SIN(b[4]), .SMC(test_se), .C(net12400), 
        .Q(b[5]) );
  SDFFQX1 dec_accop_reg_8_ ( .D(N10571), .SIN(dec_accop[7]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[8]) );
  SDFFQX1 divtempreg_reg_2_ ( .D(N13369), .SIN(divtempreg[1]), .SMC(test_se), 
        .C(net12671), .Q(divtempreg[2]) );
  SDFFQX1 dec_accop_reg_10_ ( .D(N10573), .SIN(dec_accop[9]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[10]) );
  SDFFQX1 dec_accop_reg_9_ ( .D(N10572), .SIN(dec_accop[8]), .SMC(test_se), 
        .C(net12400), .Q(dec_accop[9]) );
  SDFFQX1 b_reg_reg_3_ ( .D(N12480), .SIN(b[2]), .SMC(test_se), .C(net12400), 
        .Q(b[3]) );
  SDFFQX1 b_reg_reg_4_ ( .D(N12481), .SIN(b[3]), .SMC(test_se), .C(net12400), 
        .Q(b[4]) );
  SDFFQX1 divtempreg_reg_1_ ( .D(N13368), .SIN(divtempreg[0]), .SMC(test_se), 
        .C(net12671), .Q(divtempreg[1]) );
  SDFFQX1 divtempreg_reg_0_ ( .D(N13367), .SIN(dec_cop[7]), .SMC(test_se), .C(
        net12671), .Q(divtempreg[0]) );
  SDFFQX1 b_reg_reg_2_ ( .D(N12479), .SIN(b[1]), .SMC(test_se), .C(net12400), 
        .Q(b[2]) );
  SDFFQX1 b_reg_reg_1_ ( .D(N12478), .SIN(b[0]), .SMC(test_se), .C(net12400), 
        .Q(b[1]) );
  SDFFQX1 b_reg_reg_0_ ( .D(N12477), .SIN(n151), .SMC(test_se), .C(net12400), 
        .Q(b[0]) );
  SDFFQX1 acc_reg_reg_7_ ( .D(n1875), .SIN(acc[6]), .SMC(test_se), .C(net12400), .Q(n2481) );
  MUX4X1 U2268 ( .D0(temp[4]), .D1(temp[5]), .D2(temp[6]), .D3(temp[7]), .S0(
        N343), .S1(N344), .Y(n1968) );
  MUX4X1 U2267 ( .D0(temp[0]), .D1(temp[1]), .D2(temp[2]), .D3(temp[3]), .S0(
        N343), .S1(N344), .Y(n1969) );
  MUX2X1 U2266 ( .D0(n1969), .D1(n1968), .S(N345), .Y(N11584) );
  NAND21XL U9 ( .B(n449), .A(n2075), .Y(n632) );
  INVXL U10 ( .A(n449), .Y(n260) );
  INVX3 U11 ( .A(n449), .Y(n262) );
  NAND4X2 U12 ( .A(n279), .B(n159), .C(n277), .D(n276), .Y(n449) );
  AND2X4 U13 ( .A(n923), .B(waitstaten), .Y(n155) );
  NAND2X2 U14 ( .A(n707), .B(n709), .Y(n923) );
  MUX2X2 U15 ( .D0(pc_o[1]), .D1(n1557), .S(n155), .Y(memaddr_comb[1]) );
  OAI222X1 U16 ( .A(n946), .B(n353), .C(n354), .D(n715), .E(n355), .F(n1639), 
        .Y(n433) );
  INVX3 U17 ( .A(sfrdatai[2]), .Y(n1639) );
  OAI222X1 U18 ( .A(n936), .B(n353), .C(n2468), .D(n354), .E(n355), .F(n1648), 
        .Y(n455) );
  MUX2IX1 U19 ( .D0(n359), .D1(n358), .S(N345), .Y(n360) );
  NAND21X1 U20 ( .B(n1407), .A(n380), .Y(n397) );
  MUX2X1 U21 ( .D0(n432), .D1(n1666), .S(n2075), .Y(n1675) );
  OAI22X1 U22 ( .A(n355), .B(n1646), .C(n354), .D(n735), .Y(n506) );
  NAND32X1 U23 ( .B(n362), .C(n366), .A(n361), .Y(n456) );
  NAND21X1 U24 ( .B(n1643), .A(n360), .Y(n361) );
  OR2X1 U25 ( .A(n355), .B(n1647), .Y(n162) );
  GEN2XL U26 ( .D(n419), .E(n2138), .C(n1392), .B(n181), .A(n417), .Y(n422) );
  INVX2 U27 ( .A(n363), .Y(n1406) );
  NAND32X1 U28 ( .B(N345), .C(n256), .A(n456), .Y(n363) );
  INVX1 U29 ( .A(n708), .Y(n709) );
  INVX1 U30 ( .A(sfrdatai[4]), .Y(n1648) );
  INVX1 U31 ( .A(sfrdatai[6]), .Y(n1646) );
  NAND31X1 U32 ( .C(n398), .A(n397), .B(n396), .Y(n405) );
  MUX2IX1 U33 ( .D0(stop), .D1(n1675), .S(n1661), .Y(n654) );
  MUX2X1 U34 ( .D0(pc_o[2]), .D1(n1579), .S(n155), .Y(memaddr_comb[2]) );
  MUX2X2 U35 ( .D0(pc_o[0]), .D1(n1571), .S(n155), .Y(memaddr_comb[0]) );
  NOR2X1 U36 ( .A(n1110), .B(n2482), .Y(n1) );
  NOR2X1 U37 ( .A(n1107), .B(n2482), .Y(n2) );
  OAI222XL U38 ( .A(n730), .B(n1868), .C(n2247), .D(n1794), .E(n1945), .F(
        n2199), .Y(n3) );
  MUX2X1 U39 ( .D0(n405), .D1(n1664), .S(n2075), .Y(n10) );
  OA22X1 U40 ( .A(n1501), .B(n156), .C(n440), .D(n439), .Y(n11) );
  NAND2X1 U41 ( .A(n2242), .B(n882), .Y(n12) );
  OR4X1 U42 ( .A(n2263), .B(ramsfraddr[5]), .C(ramsfraddr[6]), .D(
        ramsfraddr[7]), .Y(n13) );
  AND4X1 U43 ( .A(phase[1]), .B(n1744), .C(n51), .D(n102), .Y(n14) );
  INVXL U44 ( .A(pc_o[15]), .Y(n15) );
  INVXL U45 ( .A(n15), .Y(memaddr[15]) );
  INVXL U46 ( .A(n516), .Y(n17) );
  INVXL U47 ( .A(n17), .Y(n18) );
  INVXL U48 ( .A(n207), .Y(n19) );
  INVXL U49 ( .A(n19), .Y(n20) );
  INVXL U50 ( .A(n1556), .Y(n21) );
  INVXL U51 ( .A(n1556), .Y(n22) );
  INVXL U52 ( .A(n1554), .Y(n23) );
  INVXL U53 ( .A(n1554), .Y(n24) );
  INVXL U54 ( .A(instr[2]), .Y(n25) );
  INVXL U55 ( .A(instr[2]), .Y(n26) );
  INVXL U56 ( .A(memaddr[12]), .Y(n27) );
  INVXL U57 ( .A(n27), .Y(pc_o[12]) );
  INVXL U58 ( .A(memaddr[5]), .Y(n29) );
  INVXL U59 ( .A(n29), .Y(pc_o[5]) );
  INVXL U60 ( .A(pc_o[13]), .Y(n31) );
  INVXL U61 ( .A(n31), .Y(memaddr[13]) );
  INVXL U62 ( .A(pc_o[0]), .Y(n33) );
  INVXL U63 ( .A(n33), .Y(memaddr[0]) );
  INVXL U64 ( .A(pc_o[6]), .Y(n35) );
  INVXL U65 ( .A(memaddr[3]), .Y(n36) );
  INVXL U66 ( .A(n36), .Y(pc_o[3]) );
  INVXL U67 ( .A(pc_o[14]), .Y(n38) );
  INVXL U68 ( .A(n38), .Y(memaddr[14]) );
  INVXL U69 ( .A(pc_o[7]), .Y(n40) );
  INVXL U70 ( .A(n40), .Y(memaddr[7]) );
  INVXL U71 ( .A(pc_o[10]), .Y(n42) );
  INVXL U72 ( .A(n42), .Y(memaddr[10]) );
  INVX1 U73 ( .A(instr[0]), .Y(n44) );
  INVX1 U74 ( .A(n50), .Y(n45) );
  INVX1 U75 ( .A(n102), .Y(instr[1]) );
  BUFX3 U76 ( .A(n2475), .Y(instr[6]) );
  BUFX3 U77 ( .A(n1130), .Y(n48) );
  BUFX3 U78 ( .A(n206), .Y(n49) );
  BUFX3 U79 ( .A(n2231), .Y(n50) );
  INVX1 U80 ( .A(instr[3]), .Y(n51) );
  BUFX3 U81 ( .A(n1136), .Y(n52) );
  BUFX3 U82 ( .A(n205), .Y(n53) );
  INVX1 U83 ( .A(n2388), .Y(n54) );
  INVX1 U84 ( .A(n62), .Y(n55) );
  INVX1 U85 ( .A(instr[7]), .Y(n56) );
  BUFX3 U86 ( .A(n1132), .Y(n57) );
  NAND2X1 U87 ( .A(n2027), .B(n2032), .Y(n1809) );
  INVX1 U88 ( .A(n1809), .Y(n58) );
  INVX1 U89 ( .A(n1809), .Y(n59) );
  INVX1 U90 ( .A(n69), .Y(n60) );
  INVX1 U91 ( .A(n127), .Y(dps[2]) );
  BUFX3 U92 ( .A(n1146), .Y(n62) );
  BUFX3 U93 ( .A(n2480), .Y(instr[0]) );
  BUFX3 U94 ( .A(n1117), .Y(n64) );
  NAND2X1 U95 ( .A(n2030), .B(n2031), .Y(n1810) );
  INVX1 U96 ( .A(n1810), .Y(n65) );
  INVX1 U97 ( .A(n1810), .Y(n66) );
  INVX1 U98 ( .A(n1974), .Y(n67) );
  NAND2X1 U99 ( .A(phase[2]), .B(n1976), .Y(n68) );
  BUFX3 U100 ( .A(acc[0]), .Y(n69) );
  BUFX3 U101 ( .A(n2478), .Y(instr[3]) );
  BUFX3 U102 ( .A(n1138), .Y(n71) );
  AOI21X1 U103 ( .B(n196), .C(n122), .A(n221), .Y(n1129) );
  INVX1 U104 ( .A(n1129), .Y(n72) );
  INVX1 U105 ( .A(n1129), .Y(n73) );
  AOI21X1 U106 ( .B(n195), .C(n146), .A(n216), .Y(n1131) );
  INVX1 U107 ( .A(n1131), .Y(n74) );
  INVX1 U108 ( .A(n1131), .Y(n75) );
  NAND2X1 U109 ( .A(n1239), .B(n123), .Y(n76) );
  NAND2X1 U110 ( .A(n2028), .B(n2045), .Y(n1819) );
  INVX1 U111 ( .A(n1819), .Y(n77) );
  INVX1 U112 ( .A(n1819), .Y(n78) );
  NAND2X1 U113 ( .A(n2030), .B(n2029), .Y(n1811) );
  INVX1 U114 ( .A(n1811), .Y(n79) );
  INVX1 U115 ( .A(n1811), .Y(n80) );
  NAND2X1 U116 ( .A(n2046), .B(n2032), .Y(n1826) );
  INVX1 U117 ( .A(n1826), .Y(n81) );
  INVX1 U118 ( .A(n1826), .Y(n82) );
  INVX1 U119 ( .A(n2418), .Y(pc_o[11]) );
  BUFX3 U120 ( .A(n2474), .Y(instr[7]) );
  INVX1 U121 ( .A(n2302), .Y(n85) );
  NOR3XL U122 ( .A(n1344), .B(n1101), .C(n1345), .Y(n1158) );
  INVX1 U123 ( .A(n2297), .Y(n86) );
  NOR3XL U124 ( .A(n2391), .B(n2298), .C(n2393), .Y(n1163) );
  BUFX3 U125 ( .A(n155), .Y(n87) );
  INVX1 U126 ( .A(n1365), .Y(n88) );
  AOI21X1 U127 ( .B(n195), .C(n1447), .A(n221), .Y(n1127) );
  INVX1 U128 ( .A(n1127), .Y(n89) );
  INVX1 U129 ( .A(n1127), .Y(n90) );
  AOI21X1 U130 ( .B(n196), .C(n1448), .A(n221), .Y(n1125) );
  INVX1 U131 ( .A(n1125), .Y(n91) );
  INVX1 U132 ( .A(n1125), .Y(n92) );
  INVX1 U133 ( .A(n2234), .Y(n93) );
  BUFX3 U134 ( .A(n1134), .Y(n94) );
  NAND2X1 U135 ( .A(n2029), .B(n2045), .Y(n1821) );
  INVX1 U136 ( .A(n1821), .Y(n95) );
  INVX1 U137 ( .A(n1821), .Y(n96) );
  NAND2X1 U138 ( .A(n2027), .B(n2028), .Y(n1808) );
  INVX1 U139 ( .A(n1808), .Y(n97) );
  INVX1 U140 ( .A(n1808), .Y(n98) );
  NAND2X1 U141 ( .A(n2046), .B(n2031), .Y(n1823) );
  INVX1 U142 ( .A(n1823), .Y(n99) );
  INVX1 U143 ( .A(n1823), .Y(n100) );
  BUFX3 U144 ( .A(n913), .Y(n101) );
  BUFX3 U145 ( .A(n2417), .Y(n102) );
  INVX1 U146 ( .A(n2299), .Y(n103) );
  NOR3XL U147 ( .A(n1344), .B(n2393), .C(n1345), .Y(n1157) );
  INVX1 U148 ( .A(n2296), .Y(n104) );
  NOR3XL U149 ( .A(n1101), .B(n2298), .C(n2391), .Y(n1164) );
  INVX1 U150 ( .A(n2477), .Y(n105) );
  INVX1 U151 ( .A(n612), .Y(acc[7]) );
  AOI21X1 U152 ( .B(n196), .C(n104), .A(n221), .Y(n1115) );
  INVX1 U153 ( .A(n1115), .Y(n108) );
  INVX1 U154 ( .A(n1115), .Y(n109) );
  AOI21X1 U155 ( .B(n195), .C(n86), .A(n220), .Y(n1123) );
  INVX1 U156 ( .A(n1123), .Y(n110) );
  INVX1 U157 ( .A(n1123), .Y(n111) );
  NAND2X1 U158 ( .A(n2030), .B(n2032), .Y(n1813) );
  INVX1 U159 ( .A(n1813), .Y(n112) );
  INVX1 U160 ( .A(n1813), .Y(n113) );
  NAND2X1 U161 ( .A(n1239), .B(n147), .Y(n114) );
  NAND2X1 U162 ( .A(n2045), .B(n2031), .Y(n1820) );
  INVX1 U163 ( .A(n1820), .Y(n115) );
  INVX1 U164 ( .A(n1820), .Y(n116) );
  NAND2X1 U165 ( .A(n2027), .B(n2029), .Y(n1807) );
  INVX1 U166 ( .A(n1807), .Y(n117) );
  INVX1 U167 ( .A(n1807), .Y(n118) );
  NAND2X1 U168 ( .A(n2046), .B(n2028), .Y(n1825) );
  INVX1 U169 ( .A(n1825), .Y(n119) );
  INVX1 U170 ( .A(n1825), .Y(n120) );
  INVX1 U171 ( .A(n2423), .Y(pc_o[9]) );
  INVX1 U172 ( .A(n2301), .Y(n122) );
  NOR3XL U173 ( .A(n2391), .B(n1101), .C(n1345), .Y(n1160) );
  INVX1 U174 ( .A(n2295), .Y(n123) );
  NOR3XL U175 ( .A(n2393), .B(n2298), .C(n1344), .Y(n1161) );
  BUFX3 U176 ( .A(n2477), .Y(instr[4]) );
  INVX1 U177 ( .A(n2446), .Y(n126) );
  BUFX3 U178 ( .A(n2293), .Y(n127) );
  INVX1 U179 ( .A(acc[1]), .Y(n128) );
  AOI21X1 U180 ( .B(n195), .C(n103), .A(n221), .Y(n1135) );
  INVX1 U181 ( .A(n1135), .Y(n129) );
  INVX1 U182 ( .A(n1135), .Y(n130) );
  AOI21X1 U183 ( .B(n196), .C(n85), .A(n221), .Y(n1133) );
  INVX1 U184 ( .A(n1133), .Y(n131) );
  INVX1 U185 ( .A(n1133), .Y(n132) );
  BUFX3 U186 ( .A(n1124), .Y(n133) );
  BUFX3 U187 ( .A(n1844), .Y(n134) );
  NAND2X1 U188 ( .A(n2030), .B(n2028), .Y(n1812) );
  INVX1 U189 ( .A(n1812), .Y(n135) );
  INVX1 U190 ( .A(n1812), .Y(n136) );
  NAND2X1 U191 ( .A(n2027), .B(n2031), .Y(n1827) );
  INVX1 U192 ( .A(n1827), .Y(n137) );
  INVX1 U193 ( .A(n1827), .Y(n138) );
  NAND2X1 U194 ( .A(n2032), .B(n2045), .Y(n1822) );
  INVX1 U195 ( .A(n1822), .Y(n139) );
  INVX1 U196 ( .A(n1822), .Y(n140) );
  NAND2X1 U197 ( .A(n2046), .B(n2029), .Y(n1824) );
  INVX1 U198 ( .A(n1824), .Y(n141) );
  INVX1 U199 ( .A(n1824), .Y(n142) );
  INVX1 U200 ( .A(n2437), .Y(pc_o[1]) );
  INVX1 U201 ( .A(n2422), .Y(pc_o[8]) );
  INVX1 U202 ( .A(n2317), .Y(n145) );
  AOI211X1 U203 ( .C(n2412), .D(n2406), .A(n253), .B(n911), .Y(n909) );
  INVX1 U204 ( .A(n2300), .Y(n146) );
  NOR3XL U205 ( .A(n2393), .B(n2391), .C(n1345), .Y(n1159) );
  INVX1 U206 ( .A(n2294), .Y(n147) );
  NOR3XL U207 ( .A(n1101), .B(n2298), .C(n1344), .Y(n1162) );
  INVX1 U208 ( .A(n680), .Y(n148) );
  INVX1 U209 ( .A(accactv), .Y(n149) );
  INVX1 U210 ( .A(n149), .Y(n150) );
  INVX1 U211 ( .A(n149), .Y(n151) );
  INVX1 U212 ( .A(n2476), .Y(n152) );
  INVX1 U213 ( .A(n152), .Y(n153) );
  INVX1 U214 ( .A(n152), .Y(instr[5]) );
  INVX1 U215 ( .A(sfrdatai[7]), .Y(n1638) );
  AOI211XL U216 ( .C(n1406), .D(n357), .A(n422), .B(n421), .Y(n424) );
  NAND3X1 U217 ( .A(n160), .B(n161), .C(n162), .Y(n482) );
  MUX2XL U218 ( .D0(pc_o[4]), .D1(n1585), .S(n155), .Y(memaddr_comb[4]) );
  NAND2X1 U219 ( .A(n1699), .B(n654), .Y(n1703) );
  MUX2X1 U220 ( .D0(memaddr[6]), .D1(n1634), .S(n155), .Y(memaddr_comb[6]) );
  NOR2X2 U221 ( .A(n165), .B(n157), .Y(n156) );
  INVX1 U222 ( .A(n386), .Y(n157) );
  OAI22X1 U223 ( .A(n1644), .B(n355), .C(n2470), .D(n354), .Y(n364) );
  XOR3X1 U224 ( .A(n2149), .B(n156), .C(n439), .Y(n423) );
  INVX1 U225 ( .A(n281), .Y(n159) );
  AND2X1 U226 ( .A(sfrwe_r), .B(n262), .Y(sfrwe) );
  INVXL U227 ( .A(n449), .Y(n261) );
  INVXL U228 ( .A(n449), .Y(waitstaten) );
  INVXL U229 ( .A(n416), .Y(n419) );
  NAND21XL U230 ( .B(n386), .A(n165), .Y(n387) );
  NAND21XL U231 ( .B(n507), .A(n372), .Y(n373) );
  AND2XL U232 ( .A(n156), .B(n1501), .Y(n440) );
  INVXL U233 ( .A(n614), .Y(n611) );
  OAI222XL U234 ( .A(n1346), .B(n1639), .C(n1240), .D(n715), .E(n946), .F(n438), .Y(n1380) );
  OAI31XL U235 ( .A(n1472), .B(n253), .C(n2384), .D(n679), .Y(n2318) );
  XNOR3X1 U236 ( .A(n897), .B(n900), .C(n158), .Y(n1667) );
  XNOR2XL U237 ( .A(n1666), .B(n1665), .Y(n158) );
  AND2XL U238 ( .A(n213), .B(n1666), .Y(N12470) );
  MUX2IX1 U239 ( .D0(n1452), .D1(n2138), .S(n375), .Y(n370) );
  AOI31XL U240 ( .A(n1399), .B(n480), .C(n420), .D(n419), .Y(n421) );
  NAND3XL U241 ( .A(n279), .B(memack), .C(n278), .Y(n1480) );
  OR4X1 U242 ( .A(n283), .B(n282), .C(n270), .D(n281), .Y(N12977) );
  NOR3XL U243 ( .A(n2248), .B(dpc[1]), .C(n1182), .Y(n1138) );
  NAND32X1 U244 ( .B(n428), .C(n427), .A(n426), .Y(n432) );
  MUX2XL U245 ( .D0(pc_o[3]), .D1(n1593), .S(n155), .Y(memaddr_comb[3]) );
  OAI222XL U246 ( .A(n1799), .B(n1798), .C(ramdatao[7]), .D(n1802), .E(n1801), 
        .F(n1800), .Y(n917) );
  AOI222XL U247 ( .A(n1148), .B(temp[1]), .C(n1149), .D(dpl_current[1]), .E(
        dptr_inc[1]), .F(n1972), .Y(n737) );
  AOI222XL U248 ( .A(n1148), .B(temp[0]), .C(n1149), .D(dpl_current[0]), .E(
        dptr_inc[0]), .F(n1972), .Y(n742) );
  AOI222XL U249 ( .A(n1148), .B(temp[3]), .C(n1149), .D(n2141), .E(dptr_inc[3]), .F(n1972), .Y(n727) );
  AOI222XL U250 ( .A(n1148), .B(temp[2]), .C(n1149), .D(dpl_current[2]), .E(
        dptr_inc[2]), .F(n1972), .Y(n732) );
  OAI222XL U251 ( .A(n1924), .B(n1923), .C(ramdatao[3]), .D(n1802), .E(n1926), 
        .F(n1925), .Y(n941) );
  AOI22AXL U252 ( .A(sp[0]), .B(n1844), .D(n1844), .C(ramdatao[0]), .Y(n1994)
         );
  AOI222XL U253 ( .A(n1148), .B(temp[6]), .C(n1149), .D(n2143), .E(dptr_inc[6]), .F(n1972), .Y(n712) );
  AOI222XL U254 ( .A(n1148), .B(temp[4]), .C(n1149), .D(n2142), .E(dptr_inc[4]), .F(n1972), .Y(n722) );
  AOI222XL U255 ( .A(n1148), .B(temp[5]), .C(n1149), .D(dpl_current[5]), .E(
        dptr_inc[5]), .F(n1972), .Y(n717) );
  OAI222XL U256 ( .A(n1846), .B(n1845), .C(ramdatao[6]), .D(n1802), .E(n1848), 
        .F(n1847), .Y(n926) );
  AOI22AXL U257 ( .A(sp[5]), .B(n134), .D(n1844), .C(ramdatao[5]), .Y(n1871)
         );
  OAI31XL U258 ( .A(n642), .B(n620), .C(n1518), .D(mempsrd), .Y(n596) );
  AOI22AXL U259 ( .A(sp[7]), .B(n134), .D(n134), .C(ramdatao[7]), .Y(n1840) );
  AOI22AXL U260 ( .A(sp[6]), .B(n134), .D(n134), .C(ramdatao[6]), .Y(n1842) );
  AOI222XL U261 ( .A(n1148), .B(temp[7]), .C(n1149), .D(dpl_current[7]), .E(
        dptr_inc[7]), .F(n1972), .Y(n704) );
  OAI222XL U262 ( .A(n590), .B(n2275), .C(n253), .D(n169), .E(n1773), .F(n257), 
        .Y(n667) );
  NOR3XL U263 ( .A(n2440), .B(ramsfraddr[2]), .C(n2444), .Y(n865) );
  OR2X1 U264 ( .A(n931), .B(n353), .Y(n160) );
  OR2X1 U265 ( .A(n2467), .B(n354), .Y(n161) );
  INVX1 U266 ( .A(n218), .Y(n210) );
  INVX1 U267 ( .A(n218), .Y(n209) );
  INVX1 U268 ( .A(n218), .Y(n211) );
  INVX1 U269 ( .A(n216), .Y(n212) );
  INVX1 U270 ( .A(n216), .Y(n213) );
  INVX1 U271 ( .A(n216), .Y(n214) );
  INVX1 U272 ( .A(n216), .Y(n215) );
  INVX1 U273 ( .A(n224), .Y(n218) );
  INVX1 U274 ( .A(n223), .Y(n219) );
  INVX1 U275 ( .A(n222), .Y(n220) );
  INVX1 U276 ( .A(n224), .Y(n216) );
  INVX1 U277 ( .A(n222), .Y(n221) );
  INVX1 U278 ( .A(n1671), .Y(n224) );
  INVX1 U279 ( .A(n1671), .Y(n223) );
  INVX1 U280 ( .A(n1671), .Y(n222) );
  NAND21X1 U281 ( .B(n262), .A(n264), .Y(N370) );
  NOR2X1 U282 ( .A(n285), .B(n2378), .Y(n1693) );
  INVX1 U283 ( .A(n2350), .Y(n1976) );
  INVX1 U284 ( .A(n481), .Y(n1392) );
  INVX1 U285 ( .A(n2341), .Y(n805) );
  INVX1 U286 ( .A(n388), .Y(n404) );
  INVX1 U287 ( .A(n1542), .Y(n390) );
  INVX1 U288 ( .A(n608), .Y(n2352) );
  INVX1 U289 ( .A(n2311), .Y(n391) );
  INVX1 U290 ( .A(n934), .Y(n392) );
  INVX1 U291 ( .A(n965), .Y(n2345) );
  NAND21X1 U292 ( .B(n270), .A(n260), .Y(n1671) );
  INVX1 U293 ( .A(n2205), .Y(n240) );
  INVX1 U294 ( .A(n2206), .Y(n244) );
  INVX1 U295 ( .A(n2207), .Y(n248) );
  INVX1 U296 ( .A(n2204), .Y(n238) );
  INVX1 U297 ( .A(n2206), .Y(n245) );
  INVX1 U298 ( .A(n2207), .Y(n249) );
  INVX1 U299 ( .A(n2203), .Y(n235) );
  INVX1 U300 ( .A(n2202), .Y(n232) );
  INVX1 U301 ( .A(n2206), .Y(n246) );
  INVX1 U302 ( .A(n2204), .Y(n239) );
  INVX1 U303 ( .A(n2207), .Y(n250) );
  INVX1 U304 ( .A(n2203), .Y(n236) );
  INVX1 U305 ( .A(n2202), .Y(n233) );
  INVX1 U306 ( .A(n2206), .Y(n247) );
  INVX1 U307 ( .A(n2200), .Y(n227) );
  INVX1 U308 ( .A(n2205), .Y(n241) );
  INVX1 U309 ( .A(n2201), .Y(n229) );
  INVX1 U310 ( .A(n2200), .Y(n226) );
  INVX1 U311 ( .A(n2205), .Y(n242) );
  INVX1 U312 ( .A(n2207), .Y(n251) );
  INVX1 U313 ( .A(n2201), .Y(n230) );
  INVX1 U314 ( .A(n2205), .Y(n243) );
  AO21X1 U315 ( .B(n215), .C(n86), .A(n272), .Y(N12547) );
  NOR21XL U316 ( .B(n223), .A(n806), .Y(N10572) );
  AND2X1 U317 ( .A(n213), .B(n1549), .Y(N11482) );
  AND2X1 U318 ( .A(n213), .B(n1553), .Y(N11484) );
  INVX1 U319 ( .A(n1552), .Y(n1736) );
  NAND21X1 U320 ( .B(n1551), .A(n211), .Y(n1552) );
  INVX1 U321 ( .A(n2194), .Y(n1752) );
  INVX1 U322 ( .A(n2196), .Y(n1751) );
  INVX1 U323 ( .A(n2198), .Y(n1740) );
  NOR2X1 U324 ( .A(n2378), .B(n2057), .Y(N10583) );
  INVX1 U325 ( .A(n1541), .Y(n2086) );
  INVX1 U326 ( .A(n2338), .Y(n2074) );
  INVX1 U327 ( .A(n271), .Y(n264) );
  INVX1 U328 ( .A(n273), .Y(n265) );
  INVX1 U329 ( .A(rst), .Y(n267) );
  INVX1 U330 ( .A(rst), .Y(n266) );
  INVX1 U331 ( .A(n270), .Y(n268) );
  INVX1 U332 ( .A(n923), .Y(n1555) );
  INVX1 U333 ( .A(n364), .Y(n372) );
  NAND21X1 U334 ( .B(n1392), .A(n373), .Y(n374) );
  INVX1 U335 ( .A(n700), .Y(n740) );
  NAND21X1 U336 ( .B(n799), .A(n166), .Y(n700) );
  INVX1 U337 ( .A(n793), .Y(n1949) );
  NAND21X1 U338 ( .B(n913), .A(n1436), .Y(n793) );
  INVX1 U339 ( .A(n1651), .Y(n1551) );
  OAI22X1 U340 ( .A(n1501), .B(n11), .C(n1381), .D(n1380), .Y(n1533) );
  AND2X1 U341 ( .A(n11), .B(n1501), .Y(n1381) );
  INVX1 U342 ( .A(n1659), .Y(n676) );
  INVX1 U343 ( .A(n1696), .Y(n1661) );
  INVX1 U344 ( .A(n1867), .Y(n648) );
  NAND32X1 U345 ( .B(n389), .C(n331), .A(n2359), .Y(n1686) );
  NAND2X1 U346 ( .A(n1640), .B(n2004), .Y(n1796) );
  NOR2X1 U347 ( .A(n2337), .B(n2394), .Y(n2031) );
  NAND21X1 U348 ( .B(n2410), .A(n2147), .Y(n2350) );
  NAND2X1 U349 ( .A(n2004), .B(n2339), .Y(n1795) );
  INVX1 U350 ( .A(n2005), .Y(n2312) );
  INVX1 U351 ( .A(n775), .Y(n2378) );
  AO21X1 U352 ( .B(n611), .C(n2138), .A(n1392), .Y(n617) );
  INVX1 U353 ( .A(n1016), .Y(n2185) );
  INVX1 U354 ( .A(n1568), .Y(n2178) );
  OR4X1 U355 ( .A(n334), .B(n349), .C(n1150), .D(n163), .Y(n1542) );
  AOI21X1 U356 ( .B(n1652), .C(n2186), .A(n257), .Y(n163) );
  NAND21X1 U357 ( .B(n2342), .A(n2161), .Y(n2341) );
  NAND43X1 U358 ( .B(n366), .C(n1392), .D(n2349), .A(n2339), .Y(n1411) );
  AO21X1 U359 ( .B(n929), .C(n365), .A(n368), .Y(n481) );
  NAND21X1 U360 ( .B(n1640), .A(n347), .Y(n349) );
  INVX1 U361 ( .A(n2339), .Y(n1640) );
  INVX1 U362 ( .A(n346), .Y(n366) );
  INVX1 U363 ( .A(n1026), .Y(n928) );
  INVX1 U364 ( .A(n1668), .Y(n1724) );
  INVX1 U365 ( .A(n1380), .Y(n441) );
  NOR2X1 U366 ( .A(n2195), .B(n602), .Y(N673) );
  NOR2X1 U367 ( .A(n725), .B(n602), .Y(N674) );
  INVXL U368 ( .A(n506), .Y(n517) );
  INVX1 U369 ( .A(n1669), .Y(n383) );
  INVX1 U370 ( .A(n1797), .Y(n2321) );
  NAND21X1 U371 ( .B(n2145), .A(n1543), .Y(n388) );
  INVX1 U372 ( .A(n953), .Y(n2145) );
  NOR2X1 U373 ( .A(n2357), .B(n2430), .Y(n608) );
  INVX1 U374 ( .A(n1501), .Y(n2149) );
  INVX1 U375 ( .A(n2318), .Y(n1974) );
  INVX1 U376 ( .A(n766), .Y(n2188) );
  INVX1 U377 ( .A(n1691), .Y(n2346) );
  INVX1 U378 ( .A(n964), .Y(n2375) );
  INVX1 U379 ( .A(n2001), .Y(n2342) );
  INVX1 U380 ( .A(n778), .Y(n289) );
  NAND21X1 U381 ( .B(n332), .A(n331), .Y(n1541) );
  AND2X1 U382 ( .A(n801), .B(n2345), .Y(n806) );
  INVX1 U383 ( .A(n507), .Y(n2138) );
  INVX1 U384 ( .A(n2359), .Y(n2159) );
  NOR3XL U385 ( .A(n2174), .B(n1976), .C(n749), .Y(n164) );
  INVX1 U386 ( .A(n1750), .Y(n2405) );
  NAND21X1 U387 ( .B(n2159), .A(n389), .Y(n934) );
  NAND21X1 U388 ( .B(n2184), .A(n953), .Y(n2311) );
  NOR2X1 U389 ( .A(n2188), .B(n2404), .Y(n965) );
  INVX1 U390 ( .A(n749), .Y(n2348) );
  INVX1 U391 ( .A(n1472), .Y(n1975) );
  INVX1 U392 ( .A(n1543), .Y(n2146) );
  INVX1 U393 ( .A(n1024), .Y(n1947) );
  NAND21X1 U394 ( .B(n1006), .A(n209), .Y(n1024) );
  INVX1 U395 ( .A(n1414), .Y(n1902) );
  NAND21X1 U396 ( .B(n1413), .A(n209), .Y(n1414) );
  NAND21X1 U397 ( .B(n2075), .A(n260), .Y(n633) );
  INVX1 U398 ( .A(n669), .Y(n2354) );
  INVX1 U399 ( .A(n2204), .Y(n237) );
  NAND21X1 U400 ( .B(n2197), .A(n211), .Y(n2196) );
  NAND21X1 U401 ( .B(n1516), .A(n210), .Y(n2194) );
  NAND21X1 U402 ( .B(n2199), .A(n211), .Y(n2198) );
  INVX1 U403 ( .A(n1438), .Y(n1239) );
  NAND21X1 U404 ( .B(n1436), .A(n210), .Y(n1438) );
  NAND2X1 U405 ( .A(n1239), .B(n86), .Y(n1124) );
  INVX1 U406 ( .A(n2203), .Y(n234) );
  INVX1 U407 ( .A(n2201), .Y(n228) );
  INVX1 U408 ( .A(n1471), .Y(n1028) );
  NAND21X1 U409 ( .B(n2428), .A(n210), .Y(n1471) );
  INVX1 U410 ( .A(n2202), .Y(n231) );
  INVX1 U411 ( .A(n2200), .Y(n225) );
  NAND21X1 U412 ( .B(n221), .A(n2071), .Y(n2057) );
  AO21X1 U413 ( .B(n222), .C(n103), .A(n270), .Y(N12493) );
  AO21X1 U414 ( .B(n222), .C(n85), .A(n272), .Y(N12502) );
  AO21X1 U415 ( .B(n222), .C(n146), .A(n272), .Y(N12511) );
  AO21X1 U416 ( .B(n222), .C(n122), .A(n273), .Y(N12520) );
  AO21X1 U417 ( .B(n215), .C(n1447), .A(n272), .Y(N12529) );
  AO21X1 U418 ( .B(n223), .C(n1448), .A(n272), .Y(N12538) );
  AO21X1 U419 ( .B(n215), .C(n104), .A(n273), .Y(N12556) );
  AND3X1 U420 ( .A(n212), .B(n1781), .C(n1633), .Y(N10577) );
  AND2X1 U421 ( .A(n1731), .B(n1651), .Y(N11489) );
  AND2X1 U422 ( .A(n213), .B(n1572), .Y(N11481) );
  AND2X1 U423 ( .A(n1867), .B(n214), .Y(N11483) );
  AND2X1 U424 ( .A(n1620), .B(n1633), .Y(N10568) );
  NOR21XL U425 ( .B(n212), .A(n2394), .Y(N12709) );
  NOR21XL U426 ( .B(n212), .A(n2309), .Y(N12710) );
  INVX1 U427 ( .A(n1670), .Y(n1731) );
  NOR2X1 U428 ( .A(n2060), .B(n2067), .Y(N10570) );
  INVX1 U429 ( .A(n460), .Y(n1553) );
  INVX1 U430 ( .A(n461), .Y(n1549) );
  INVX1 U431 ( .A(n1240), .Y(n2150) );
  INVX1 U432 ( .A(n1346), .Y(n2151) );
  INVX1 U433 ( .A(n939), .Y(n2154) );
  NAND4X1 U434 ( .A(n2216), .B(n2215), .C(n2214), .D(n2213), .Y(n1042) );
  NAND21X1 U435 ( .B(n2340), .A(n2161), .Y(n2338) );
  NAND4X1 U436 ( .A(n2220), .B(n2219), .C(n2218), .D(n2217), .Y(n1043) );
  INVX1 U437 ( .A(n967), .Y(n2323) );
  INVX1 U438 ( .A(n947), .Y(n2314) );
  INVX1 U439 ( .A(n915), .Y(n2344) );
  INVX1 U440 ( .A(n1163), .Y(n2297) );
  INVX1 U441 ( .A(n274), .Y(n270) );
  OAI21X1 U442 ( .B(n2404), .C(n2346), .A(n2341), .Y(n2084) );
  INVX1 U443 ( .A(n275), .Y(n273) );
  NOR2X1 U444 ( .A(n2428), .B(n269), .Y(n485) );
  INVX1 U445 ( .A(n275), .Y(n271) );
  INVX1 U446 ( .A(n275), .Y(n272) );
  OAI22X1 U447 ( .A(n355), .B(n1638), .C(n2466), .D(n354), .Y(n614) );
  OAI22X1 U448 ( .A(n355), .B(n1641), .C(n2469), .D(n354), .Y(n416) );
  OAI222XL U449 ( .A(n1346), .B(n1641), .C(n2469), .D(n1240), .E(n952), .F(
        n438), .Y(n439) );
  INVX1 U450 ( .A(sfrdatai[1]), .Y(n1641) );
  OA222X1 U451 ( .A(n2470), .B(n1240), .C(n1346), .D(n1644), .E(n959), .F(n438), .Y(n165) );
  NAND21X1 U452 ( .B(n2318), .A(n707), .Y(n913) );
  INVX1 U453 ( .A(n701), .Y(n739) );
  NAND21X1 U454 ( .B(n796), .A(n166), .Y(n701) );
  AND2X1 U455 ( .A(n743), .B(n2236), .Y(n166) );
  OAI22X1 U456 ( .A(n895), .B(n1794), .C(n1793), .D(n2209), .Y(n1651) );
  INVX1 U457 ( .A(memdatai[7]), .Y(n2209) );
  NAND2X1 U458 ( .A(n743), .B(n744), .Y(n167) );
  OAI21X1 U459 ( .B(n1444), .C(n1445), .A(n1446), .Y(n1402) );
  NAND21X1 U460 ( .B(n1678), .A(cs_run), .Y(n1659) );
  OAI21BBX1 U461 ( .A(n1533), .B(n1534), .C(n1535), .Y(n1502) );
  OAI21X1 U462 ( .B(n1534), .C(n1533), .A(n2149), .Y(n1535) );
  AOI22AXL U463 ( .A(n1502), .B(n1503), .D(n1504), .C(n2149), .Y(n1444) );
  NOR2X1 U464 ( .A(n1503), .B(n1502), .Y(n1504) );
  AOI22X1 U465 ( .A(n2146), .B(n1137), .C(n1393), .D(n2320), .Y(n1390) );
  XNOR2XL U466 ( .A(n1394), .B(n1395), .Y(n1393) );
  XNOR2XL U467 ( .A(n2149), .B(n1396), .Y(n1395) );
  AOI22X1 U468 ( .A(n2149), .B(n1400), .C(n1401), .D(n1402), .Y(n1394) );
  INVX1 U469 ( .A(n1377), .Y(n2449) );
  OR2X1 U470 ( .A(n1401), .B(n1402), .Y(n1400) );
  OAI222XL U471 ( .A(n1868), .B(n2208), .C(n1793), .D(n2195), .E(n1794), .F(
        n637), .Y(n1572) );
  INVX1 U472 ( .A(n888), .Y(n637) );
  OAI221X1 U473 ( .A(n885), .B(n1794), .C(n1793), .D(n730), .E(n1868), .Y(
        n1867) );
  NAND5XL U474 ( .A(n460), .B(n461), .C(sfrwe_comb_s), .D(n651), .E(n649), .Y(
        n1696) );
  INVX1 U475 ( .A(n1572), .Y(n651) );
  INVX1 U476 ( .A(n643), .Y(sfrwe_comb_s) );
  AND4X1 U477 ( .A(n1550), .B(n174), .C(n3), .D(n648), .Y(n649) );
  INVX1 U478 ( .A(memdatai[2]), .Y(n2199) );
  INVX1 U479 ( .A(memdatai[3]), .Y(n2195) );
  INVX1 U480 ( .A(memdatai[1]), .Y(n2197) );
  OA22X1 U481 ( .A(n1793), .B(n2208), .C(n889), .D(n1794), .Y(n460) );
  AOI22BXL U482 ( .B(n1793), .A(memdatai[4]), .D(n1794), .C(n893), .Y(n461) );
  INVX1 U483 ( .A(memdatai[0]), .Y(n1516) );
  NOR21XL U484 ( .B(n1949), .A(n691), .Y(n670) );
  NAND32X1 U485 ( .B(n692), .C(n799), .A(n798), .Y(n896) );
  XNOR2XL U486 ( .A(n888), .B(n893), .Y(n894) );
  INVX1 U487 ( .A(n795), .Y(n798) );
  NAND32X1 U488 ( .B(n2175), .C(n794), .A(n1949), .Y(n795) );
  INVX1 U489 ( .A(n691), .Y(n794) );
  NAND2X1 U490 ( .A(n2018), .B(n1802), .Y(n1814) );
  NAND2X1 U491 ( .A(n1802), .B(n2309), .Y(n1832) );
  INVX1 U492 ( .A(n797), .Y(n1948) );
  NAND32X1 U493 ( .B(n692), .C(n796), .A(n798), .Y(n797) );
  INVX1 U494 ( .A(n796), .Y(n799) );
  INVX1 U495 ( .A(n752), .Y(n2430) );
  INVX1 U496 ( .A(n1432), .Y(n2262) );
  INVX1 U497 ( .A(n895), .Y(n2242) );
  NOR2X1 U498 ( .A(n883), .B(n884), .Y(n882) );
  OR2X1 U499 ( .A(n2175), .B(n1948), .Y(n168) );
  INVX1 U500 ( .A(n1364), .Y(n2327) );
  INVX1 U501 ( .A(n1362), .Y(n2303) );
  NAND21X1 U502 ( .B(n255), .A(n175), .Y(n2359) );
  OAI211X1 U503 ( .C(n2008), .D(n253), .A(n2185), .B(n2313), .Y(n2005) );
  AOI21X1 U504 ( .B(n2161), .C(n1737), .A(n1976), .Y(n2008) );
  XNOR2XL U505 ( .A(n583), .B(n586), .Y(n1608) );
  INVX1 U506 ( .A(n753), .Y(n2404) );
  INVX1 U507 ( .A(n2047), .Y(n2394) );
  INVX1 U508 ( .A(n2018), .Y(n2309) );
  INVX1 U509 ( .A(n2351), .Y(n2147) );
  INVX1 U510 ( .A(n959), .Y(n634) );
  NOR3XL U511 ( .A(n2007), .B(n2002), .C(n2005), .Y(n2004) );
  INVX1 U512 ( .A(n1866), .Y(n2276) );
  INVX1 U513 ( .A(n1802), .Y(n406) );
  NOR2X1 U514 ( .A(n2394), .B(n2039), .Y(n2029) );
  NOR2X1 U515 ( .A(n2337), .B(n2047), .Y(n2028) );
  INVX1 U516 ( .A(n313), .Y(n331) );
  NAND21X1 U517 ( .B(n256), .A(n312), .Y(n313) );
  INVX1 U518 ( .A(n311), .Y(n389) );
  NAND21X1 U519 ( .B(n252), .A(n175), .Y(n311) );
  INVX1 U520 ( .A(n484), .Y(n2427) );
  INVX1 U521 ( .A(n1027), .Y(n2428) );
  INVX1 U522 ( .A(n890), .Y(n2258) );
  INVX1 U523 ( .A(n1459), .Y(n2181) );
  INVX1 U524 ( .A(n1687), .Y(n2184) );
  NAND32X1 U525 ( .B(n310), .C(n2404), .A(n2189), .Y(n953) );
  INVX1 U526 ( .A(intcall), .Y(n310) );
  NAND21X1 U527 ( .B(n252), .A(n312), .Y(n1543) );
  NOR21XL U528 ( .B(n1710), .A(n1711), .Y(n1374) );
  NOR2X1 U529 ( .A(n2358), .B(n2388), .Y(n1737) );
  INVX1 U530 ( .A(n1044), .Y(n2306) );
  NOR2X1 U531 ( .A(n2402), .B(n2379), .Y(n775) );
  INVX1 U532 ( .A(n2373), .Y(n2161) );
  XNOR2XL U533 ( .A(n1534), .B(n1501), .Y(n1548) );
  NOR2X1 U534 ( .A(n2350), .B(n255), .Y(n1016) );
  NOR2X1 U535 ( .A(n1056), .B(n1073), .Y(n1568) );
  INVX1 U536 ( .A(n258), .Y(n256) );
  NOR2X1 U537 ( .A(n2047), .B(n2039), .Y(n2032) );
  INVX1 U538 ( .A(n774), .Y(n2189) );
  INVX1 U539 ( .A(n505), .Y(n619) );
  INVX1 U540 ( .A(memdatai[4]), .Y(n725) );
  INVX1 U541 ( .A(memdatai[5]), .Y(n730) );
  ENOX1 U542 ( .A(n470), .B(n1379), .C(n2075), .D(n1901), .Y(N11503) );
  INVX1 U543 ( .A(n1742), .Y(n2410) );
  INVX1 U544 ( .A(n1843), .Y(n2277) );
  INVX1 U545 ( .A(n2039), .Y(n2337) );
  INVX1 U546 ( .A(n1682), .Y(n2402) );
  NAND21X1 U547 ( .B(n1678), .A(n209), .Y(n1668) );
  AO21X1 U548 ( .B(n1701), .C(n1659), .A(n273), .Y(n1660) );
  NAND2X1 U549 ( .A(n2322), .B(n2007), .Y(n1797) );
  INVX1 U550 ( .A(n1748), .Y(n2377) );
  OAI21X1 U551 ( .B(n601), .C(n2194), .A(n474), .Y(N670) );
  OAI21X1 U552 ( .B(n601), .C(n2198), .A(n474), .Y(N672) );
  OAI31XL U553 ( .A(n730), .B(n601), .C(n220), .D(n474), .Y(N675) );
  OAI31XL U554 ( .A(n601), .B(n2209), .C(n219), .D(n474), .Y(N677) );
  INVX1 U555 ( .A(n2002), .Y(n2322) );
  NOR2X1 U556 ( .A(n1789), .B(n1693), .Y(n1768) );
  ENOX1 U557 ( .A(n471), .B(n1379), .C(n2075), .D(n1902), .Y(N11502) );
  INVX1 U558 ( .A(n1498), .Y(n2180) );
  INVX1 U559 ( .A(n780), .Y(n2382) );
  NAND21X1 U560 ( .B(n255), .A(n318), .Y(n2339) );
  NAND21X1 U561 ( .B(n2351), .A(n2161), .Y(n346) );
  OAI211X1 U562 ( .C(n2050), .D(n2404), .A(n315), .B(n314), .Y(n2349) );
  INVX1 U563 ( .A(n1693), .Y(n315) );
  INVX1 U564 ( .A(n1692), .Y(n314) );
  OR2X1 U565 ( .A(n350), .B(n349), .Y(n353) );
  NOR2X1 U566 ( .A(n2413), .B(n2358), .Y(n1026) );
  NAND32X1 U567 ( .B(n2379), .C(n2384), .A(n1026), .Y(n929) );
  NAND32X1 U568 ( .B(n2379), .C(n2389), .A(n1026), .Y(n365) );
  INVX1 U569 ( .A(n339), .Y(n1655) );
  NAND32X1 U570 ( .B(n338), .C(n366), .A(n369), .Y(n339) );
  INVX1 U571 ( .A(n365), .Y(n338) );
  NAND2X1 U572 ( .A(n353), .B(n355), .Y(n354) );
  NAND21X1 U573 ( .B(n255), .A(n2349), .Y(n347) );
  NAND32X1 U574 ( .B(n1452), .C(n2349), .A(n2339), .Y(n368) );
  NOR2X1 U575 ( .A(n2347), .B(n2385), .Y(n1691) );
  OR3XL U576 ( .A(n2320), .B(n332), .C(n1686), .Y(n334) );
  NAND21X1 U577 ( .B(n2351), .A(n775), .Y(n340) );
  INVX1 U578 ( .A(n1004), .Y(n2075) );
  NOR2X1 U579 ( .A(n2406), .B(n774), .Y(n1692) );
  NOR2X1 U580 ( .A(n2340), .B(n2379), .Y(n1669) );
  NOR2X1 U581 ( .A(n2343), .B(n2386), .Y(n2001) );
  NOR2X1 U582 ( .A(n1972), .B(n1148), .Y(n1149) );
  INVX1 U583 ( .A(n1452), .Y(n2140) );
  INVX1 U584 ( .A(n758), .Y(n2347) );
  INVX1 U585 ( .A(n2372), .Y(n809) );
  OR2X1 U586 ( .A(n601), .B(n593), .Y(n602) );
  INVX1 U587 ( .A(n367), .Y(n2139) );
  AND3X1 U588 ( .A(n768), .B(n769), .C(n770), .Y(n762) );
  NOR32XL U589 ( .B(n169), .C(n786), .A(n787), .Y(n768) );
  NOR4XL U590 ( .A(n318), .B(n782), .C(n2174), .D(n783), .Y(n769) );
  NOR4XL U591 ( .A(n771), .B(n772), .C(n2349), .D(n592), .Y(n770) );
  AND2X1 U592 ( .A(n213), .B(n1662), .Y(N11501) );
  INVX1 U593 ( .A(n1151), .Y(n2426) );
  INVX1 U594 ( .A(n474), .Y(n2193) );
  INVX1 U595 ( .A(n764), .Y(n2340) );
  INVX1 U596 ( .A(n910), .Y(n2384) );
  AND2X1 U597 ( .A(n929), .B(n933), .Y(n1657) );
  INVX1 U598 ( .A(n591), .Y(n2186) );
  INVX1 U599 ( .A(n482), .Y(n492) );
  NOR2X1 U600 ( .A(n2208), .B(n602), .Y(N676) );
  GEN2XL U601 ( .D(n337), .E(n336), .C(n2361), .B(n335), .A(n334), .Y(n1407)
         );
  AND2X1 U602 ( .A(n2160), .B(n2186), .Y(n337) );
  AND2X1 U603 ( .A(n333), .B(n1652), .Y(n336) );
  INVX1 U604 ( .A(n2349), .Y(n333) );
  AO21X1 U605 ( .B(n933), .C(n369), .A(n368), .Y(n507) );
  INVX1 U606 ( .A(n1476), .Y(n1413) );
  OAI22X1 U607 ( .A(n253), .B(n308), .C(n257), .D(n307), .Y(n1501) );
  INVX1 U608 ( .A(n306), .Y(n308) );
  AND2X1 U609 ( .A(n587), .B(n2188), .Y(n307) );
  OR2X1 U610 ( .A(n2152), .B(n382), .Y(n1346) );
  NAND21X1 U611 ( .B(n2152), .A(n382), .Y(n1240) );
  NOR2X1 U612 ( .A(n2416), .B(n2347), .Y(n766) );
  NAND21X1 U613 ( .B(n1687), .A(n404), .Y(n332) );
  NOR2X1 U614 ( .A(n2346), .B(n2412), .Y(n778) );
  NOR2X1 U615 ( .A(n2376), .B(n2407), .Y(n964) );
  OAI211X1 U616 ( .C(n256), .D(n385), .A(n384), .B(n2149), .Y(n386) );
  AND2X1 U617 ( .A(n589), .B(n383), .Y(n385) );
  NOR2X1 U618 ( .A(n2130), .B(n1742), .Y(n1750) );
  INVX1 U619 ( .A(n2325), .Y(n628) );
  INVX1 U620 ( .A(n909), .Y(n679) );
  INVX1 U621 ( .A(n438), .Y(n2152) );
  AOI21X1 U622 ( .B(n2066), .C(n753), .A(n964), .Y(n801) );
  INVX1 U623 ( .A(n258), .Y(n257) );
  INVX1 U624 ( .A(n342), .Y(n1384) );
  NAND32X1 U625 ( .B(n2349), .C(n350), .A(n2339), .Y(n342) );
  AOI21AX1 U626 ( .B(n1691), .C(n1781), .A(n296), .Y(n169) );
  INVX1 U627 ( .A(n592), .Y(n1652) );
  INVX1 U628 ( .A(n1449), .Y(n1436) );
  INVX1 U629 ( .A(n1561), .Y(n429) );
  NAND2X1 U630 ( .A(n2406), .B(n1694), .Y(n2130) );
  INVX1 U631 ( .A(n784), .Y(n2174) );
  INVX1 U632 ( .A(n1681), .Y(n2376) );
  INVX1 U633 ( .A(n1336), .Y(n2357) );
  NAND21X1 U634 ( .B(n1743), .A(n628), .Y(n939) );
  NAND21X1 U635 ( .B(n2379), .A(n2157), .Y(n1472) );
  NAND21X1 U636 ( .B(n2384), .A(n2156), .Y(n669) );
  XNOR2XL U637 ( .A(n170), .B(n171), .Y(n897) );
  XNOR2XL U638 ( .A(n1474), .B(n1473), .Y(n170) );
  XNOR2XL U639 ( .A(n1476), .B(n1475), .Y(n171) );
  INVX1 U640 ( .A(n909), .Y(n2317) );
  INVX1 U641 ( .A(n335), .Y(n1150) );
  OAI221X1 U642 ( .A(n2409), .B(n2346), .C(n2413), .D(n2376), .E(n589), .Y(
        n782) );
  INVX1 U643 ( .A(n318), .Y(n2160) );
  NAND3X1 U644 ( .A(n1026), .B(n2377), .C(n910), .Y(n590) );
  NOR2X1 U645 ( .A(n2358), .B(n2386), .Y(n777) );
  NOR3XL U646 ( .A(n2411), .B(n285), .C(n2377), .Y(n803) );
  NAND2X1 U647 ( .A(n2059), .B(n774), .Y(n2063) );
  INVX1 U648 ( .A(n2320), .Y(n1410) );
  AND2X1 U649 ( .A(n223), .B(n1667), .Y(N12905) );
  XNOR2XL U650 ( .A(n901), .B(n902), .Y(n900) );
  ENOX1 U651 ( .A(n472), .B(n1379), .C(n2075), .D(n1947), .Y(N11500) );
  INVX1 U652 ( .A(n384), .Y(n2158) );
  NAND3X1 U653 ( .A(n2413), .B(n2430), .C(n2406), .Y(n2108) );
  INVX1 U654 ( .A(n902), .Y(n1006) );
  INVX1 U655 ( .A(n810), .Y(n2374) );
  NOR2X1 U656 ( .A(n2059), .B(n2407), .Y(n749) );
  NOR2X1 U657 ( .A(n2384), .B(n2358), .Y(n2071) );
  INVX1 U658 ( .A(n1781), .Y(n2401) );
  AND2X1 U659 ( .A(n213), .B(n10), .Y(N11498) );
  INVX1 U660 ( .A(n744), .Y(n2236) );
  INVX1 U661 ( .A(n1664), .Y(n1665) );
  INVX1 U662 ( .A(n2050), .Y(n2187) );
  INVX1 U663 ( .A(n1433), .Y(n1875) );
  NAND21X1 U664 ( .B(n1473), .A(n209), .Y(n1433) );
  INVX1 U665 ( .A(n1416), .Y(n1900) );
  NAND21X1 U666 ( .B(n1474), .A(n209), .Y(n1416) );
  INVX1 U667 ( .A(n1415), .Y(n1901) );
  NAND21X1 U668 ( .B(n1475), .A(n209), .Y(n1415) );
  NOR3XL U669 ( .A(n2351), .B(n256), .C(n2409), .Y(n698) );
  NOR2X1 U670 ( .A(n2175), .B(n698), .Y(n788) );
  INVX1 U671 ( .A(n692), .Y(n2176) );
  AND2X1 U672 ( .A(n212), .B(n1664), .Y(N12469) );
  AND2X1 U673 ( .A(n213), .B(n901), .Y(N12472) );
  INVX1 U674 ( .A(n818), .Y(n833) );
  NAND21X1 U675 ( .B(n2176), .A(n691), .Y(n818) );
  NOR2X1 U676 ( .A(n1022), .B(n1972), .Y(n1247) );
  INVX1 U677 ( .A(n2204), .Y(n1783) );
  INVX1 U678 ( .A(n2205), .Y(n1872) );
  INVX1 U679 ( .A(n1248), .Y(n2425) );
  NOR21XL U680 ( .B(n1356), .A(n1355), .Y(n1359) );
  NAND21X1 U681 ( .B(n1573), .A(n209), .Y(n1670) );
  NAND21X1 U682 ( .B(n1434), .A(n210), .Y(n1350) );
  NAND21X1 U683 ( .B(n216), .A(n1742), .Y(n2067) );
  NAND2X1 U684 ( .A(n1239), .B(n147), .Y(n1126) );
  NAND2X1 U685 ( .A(n1239), .B(n85), .Y(n1134) );
  NAND2X1 U686 ( .A(n1239), .B(n123), .Y(n1128) );
  NAND2X1 U687 ( .A(n1239), .B(n146), .Y(n1132) );
  NAND2X1 U688 ( .A(n1239), .B(n103), .Y(n1136) );
  NAND2X1 U689 ( .A(n1239), .B(n122), .Y(n1130) );
  NAND2X1 U690 ( .A(n1239), .B(n104), .Y(n1117) );
  OAI32X1 U691 ( .A(n2411), .B(n2376), .C(n220), .D(n2065), .E(n2067), .Y(
        N10571) );
  INVX1 U692 ( .A(n2202), .Y(n1779) );
  OAI21X1 U693 ( .B(n1450), .C(n861), .A(n267), .Y(N13122) );
  OAI21X1 U694 ( .B(n2439), .C(n861), .A(n266), .Y(N13131) );
  OAI21X1 U695 ( .B(n851), .C(n861), .A(n266), .Y(N13149) );
  OAI21X1 U696 ( .B(n1450), .C(n852), .A(n265), .Y(N13266) );
  OAI21X1 U697 ( .B(n2439), .C(n852), .A(n265), .Y(N13275) );
  OAI21X1 U698 ( .B(n851), .C(n852), .A(n265), .Y(N13293) );
  OAI21X1 U699 ( .B(n1111), .C(n1113), .A(n274), .Y(N12637) );
  INVX1 U700 ( .A(n2203), .Y(n1782) );
  INVX1 U701 ( .A(n2200), .Y(n1772) );
  INVX1 U702 ( .A(n2206), .Y(n1873) );
  INVX1 U703 ( .A(n2201), .Y(n1778) );
  INVX1 U704 ( .A(n2207), .Y(n1874) );
  NAND2X1 U705 ( .A(n264), .B(n2204), .Y(N12690) );
  NAND2X1 U706 ( .A(n264), .B(n2202), .Y(N12692) );
  NAND2X1 U707 ( .A(n264), .B(n2203), .Y(N12691) );
  NOR2X1 U708 ( .A(n848), .B(n2220), .Y(N13325) );
  NOR2X1 U709 ( .A(n848), .B(n2219), .Y(N13326) );
  NOR2X1 U710 ( .A(n848), .B(n2218), .Y(N13327) );
  NOR2X1 U711 ( .A(n848), .B(n2217), .Y(N13328) );
  NOR2X1 U712 ( .A(n848), .B(n2216), .Y(N13329) );
  NOR2X1 U713 ( .A(n848), .B(n2215), .Y(N13330) );
  NOR2X1 U714 ( .A(n848), .B(n2214), .Y(N13331) );
  NOR2X1 U715 ( .A(n848), .B(n2213), .Y(N13332) );
  NOR21XL U716 ( .B(n1756), .A(n495), .Y(N583) );
  NOR21XL U717 ( .B(n215), .A(n2062), .Y(N10574) );
  AOI21BX1 U718 ( .C(n1694), .B(n2063), .A(n2064), .Y(n2062) );
  NAND21X1 U719 ( .B(n219), .A(n1004), .Y(n1379) );
  NAND21X1 U720 ( .B(n220), .A(n2177), .Y(n1091) );
  NAND32X1 U721 ( .B(n216), .C(n1519), .A(n1544), .Y(n594) );
  AO21X1 U722 ( .B(n215), .C(n1628), .A(n273), .Y(N12699) );
  INVX1 U723 ( .A(n1088), .Y(n1628) );
  AO21X1 U724 ( .B(n215), .C(n1631), .A(n273), .Y(N12698) );
  INVX1 U725 ( .A(n1089), .Y(n1631) );
  AO21X1 U726 ( .B(n222), .C(n1632), .A(n273), .Y(N12697) );
  INVX1 U727 ( .A(n1090), .Y(n1632) );
  NOR31X1 U728 ( .C(n212), .A(n2412), .B(n2060), .Y(N10576) );
  AND3X1 U729 ( .A(n212), .B(n1630), .C(n1629), .Y(N10575) );
  INVX1 U730 ( .A(n1694), .Y(n1630) );
  AND3X1 U731 ( .A(n211), .B(n753), .C(n1653), .Y(N10589) );
  NOR32XL U732 ( .B(n212), .C(n1629), .A(n2406), .Y(N10573) );
  AND2X1 U733 ( .A(n1620), .B(n1653), .Y(N10564) );
  AND2X1 U734 ( .A(n1619), .B(n214), .Y(N584) );
  AND2X1 U735 ( .A(n2058), .B(n214), .Y(N10578) );
  AND2X1 U736 ( .A(n213), .B(n1550), .Y(N11478) );
  AND2X1 U737 ( .A(n213), .B(n3), .Y(N11480) );
  AND2X1 U738 ( .A(n223), .B(n174), .Y(N11479) );
  NOR21XL U739 ( .B(n222), .A(n1087), .Y(N12700) );
  NOR21XL U740 ( .B(n223), .A(n1086), .Y(N12701) );
  NOR21XL U741 ( .B(n223), .A(n1084), .Y(N12703) );
  NOR21XL U742 ( .B(n223), .A(n1085), .Y(N12702) );
  NOR21XL U743 ( .B(n223), .A(n1013), .Y(N10585) );
  NOR21XL U744 ( .B(n223), .A(n1083), .Y(N12704) );
  NOR3XL U745 ( .A(n2055), .B(n2343), .C(n2373), .Y(N10581) );
  NOR3XL U746 ( .A(n2055), .B(n2343), .C(n2378), .Y(N10565) );
  NOR3XL U747 ( .A(n2057), .B(n2379), .C(n2411), .Y(N10563) );
  INVX1 U748 ( .A(n1547), .Y(n1620) );
  NAND21X1 U749 ( .B(n2409), .A(n210), .Y(n1547) );
  AOI31X1 U750 ( .A(n588), .B(n587), .C(n1652), .D(n1671), .Y(N690) );
  NOR32XL U751 ( .B(n589), .C(n590), .A(n591), .Y(n588) );
  NOR2X1 U752 ( .A(n2373), .B(n2057), .Y(N10582) );
  NOR2X1 U753 ( .A(n846), .B(n841), .Y(N13368) );
  NOR2X1 U754 ( .A(n844), .B(n841), .Y(N13370) );
  NOR2X1 U755 ( .A(n845), .B(n841), .Y(N13369) );
  NOR2X1 U756 ( .A(n843), .B(n841), .Y(N13371) );
  NOR2X1 U757 ( .A(n842), .B(n841), .Y(N13372) );
  NOR2X1 U758 ( .A(n840), .B(n841), .Y(N13373) );
  NOR2X1 U759 ( .A(n252), .B(n595), .Y(N680) );
  NOR2X1 U760 ( .A(n255), .B(n595), .Y(N681) );
  NAND3X1 U761 ( .A(n593), .B(n264), .C(n594), .Y(N685) );
  INVX1 U762 ( .A(N13353), .Y(n2190) );
  INVX1 U763 ( .A(n618), .Y(n663) );
  OAI22X1 U764 ( .A(n936), .B(n2323), .C(n725), .D(n918), .Y(n935) );
  INVX1 U765 ( .A(n1515), .Y(n1544) );
  INVX1 U766 ( .A(n1519), .Y(n2010) );
  NAND2X1 U767 ( .A(n1509), .B(n2338), .Y(n1386) );
  INVX1 U768 ( .A(n1144), .Y(n2231) );
  INVX1 U769 ( .A(n1146), .Y(n2232) );
  AOI21X1 U770 ( .B(n2370), .C(n2232), .A(n1182), .Y(n1169) );
  AOI21X1 U771 ( .B(n1204), .C(n2232), .A(n1182), .Y(n1192) );
  INVX1 U772 ( .A(n1509), .Y(n2153) );
  INVX1 U773 ( .A(n1182), .Y(n2233) );
  AOI221XL U774 ( .A(n2287), .B(n2231), .C(n2292), .D(n1138), .E(n1182), .Y(
        n1271) );
  INVX1 U775 ( .A(multemp2[9]), .Y(n2213) );
  INVX1 U776 ( .A(multemp2[8]), .Y(n2214) );
  INVX1 U777 ( .A(n1138), .Y(n2235) );
  OAI21X1 U778 ( .B(n1181), .C(n1144), .A(n1169), .Y(n1180) );
  INVX1 U779 ( .A(n938), .Y(n2155) );
  INVX1 U780 ( .A(multemp2[7]), .Y(n2215) );
  INVX1 U781 ( .A(multemp2[6]), .Y(n2216) );
  OAI21X1 U782 ( .B(n1142), .C(n62), .A(n1312), .Y(n1321) );
  NOR2X1 U783 ( .A(n1138), .B(n2231), .Y(n1221) );
  INVX1 U784 ( .A(multemp2[5]), .Y(n2217) );
  INVX1 U785 ( .A(multemp2[4]), .Y(n2218) );
  INVX1 U786 ( .A(n1189), .Y(n452) );
  INVX1 U787 ( .A(n1267), .Y(n2291) );
  NAND31X1 U788 ( .C(n1020), .A(n590), .B(n1021), .Y(n1019) );
  INVX1 U789 ( .A(multemp2[3]), .Y(n2219) );
  OAI21X1 U790 ( .B(n2353), .C(n257), .A(n1008), .Y(n985) );
  INVX1 U791 ( .A(n1211), .Y(n2419) );
  INVX1 U792 ( .A(n993), .Y(n2281) );
  INVX1 U793 ( .A(n1269), .Y(n2292) );
  INVX1 U794 ( .A(multemp2[2]), .Y(n2220) );
  NOR2X1 U795 ( .A(n2345), .B(n255), .Y(n915) );
  INVX1 U796 ( .A(n921), .Y(n2282) );
  NOR2X1 U797 ( .A(n2375), .B(n252), .Y(n967) );
  NAND2X1 U798 ( .A(n960), .B(n2319), .Y(n947) );
  INVX1 U799 ( .A(n495), .Y(n1596) );
  INVX1 U800 ( .A(n2295), .Y(n1447) );
  INVX1 U801 ( .A(n1161), .Y(n2295) );
  INVX1 U802 ( .A(n1159), .Y(n2300) );
  INVX1 U803 ( .A(n1157), .Y(n2299) );
  INVX1 U804 ( .A(n2294), .Y(n1448) );
  INVX1 U805 ( .A(n1162), .Y(n2294) );
  INVX1 U806 ( .A(n1158), .Y(n2302) );
  INVX1 U807 ( .A(n1160), .Y(n2301) );
  INVX1 U808 ( .A(n1164), .Y(n2296) );
  AOI21BBXL U809 ( .B(n1669), .C(n2158), .A(n2413), .Y(n2064) );
  INVX1 U810 ( .A(rst), .Y(n274) );
  INVX1 U811 ( .A(n2061), .Y(n1629) );
  NOR21XL U812 ( .B(n2065), .A(n972), .Y(n2061) );
  NOR2X1 U813 ( .A(n2066), .B(n766), .Y(n2065) );
  INVX1 U814 ( .A(n1204), .Y(n2421) );
  NOR21XL U815 ( .B(n2068), .A(n2063), .Y(n2060) );
  NAND2X1 U816 ( .A(n264), .B(n2424), .Y(n878) );
  INVX1 U817 ( .A(n275), .Y(n269) );
  INVX1 U818 ( .A(rst), .Y(n275) );
  INVX1 U819 ( .A(n2059), .Y(n1633) );
  MUX2X1 U820 ( .D0(memwr), .D1(n644), .S(n261), .Y(memwr_comb) );
  AND2X1 U821 ( .A(n496), .B(n1596), .Y(n647) );
  NAND21X1 U822 ( .B(mempsack), .A(n280), .Y(n276) );
  NAND21X1 U823 ( .B(memack), .A(n278), .Y(n277) );
  OA2222XL U824 ( .A(n1541), .B(n425), .C(n1542), .D(n2260), .E(n424), .F(
        n1407), .G(n1410), .H(n423), .Y(n426) );
  INVX1 U825 ( .A(pc_i[9]), .Y(n425) );
  NOR21XL U826 ( .B(n2156), .A(n345), .Y(n362) );
  NOR21X1 U827 ( .B(n1406), .A(n2273), .Y(n378) );
  NAND21X1 U828 ( .B(n596), .A(n1703), .Y(n708) );
  NOR21XL U829 ( .B(pc_i[8]), .A(n1541), .Y(n398) );
  NAND21X1 U830 ( .B(n372), .A(n371), .Y(n377) );
  NAND31X1 U831 ( .C(n418), .A(n370), .B(n454), .Y(n371) );
  INVX1 U832 ( .A(sfrdatai[5]), .Y(n1647) );
  INVX1 U833 ( .A(sfrdatai[3]), .Y(n1649) );
  INVX1 U834 ( .A(sfrdatai[0]), .Y(n1644) );
  MUX2X1 U835 ( .D0(n507), .D1(n2140), .S(n181), .Y(n420) );
  OAI211X1 U836 ( .C(n628), .D(n1516), .A(n402), .B(n401), .Y(n1664) );
  OA222X1 U837 ( .A(n1509), .B(n2261), .C(n959), .D(n939), .E(n2470), .F(n429), 
        .Y(n401) );
  OA22XL U838 ( .A(n703), .B(n627), .C(n1644), .D(n938), .Y(n402) );
  OAI211X1 U839 ( .C(n628), .D(n2197), .A(n431), .B(n430), .Y(n1666) );
  OA222X1 U840 ( .A(n1509), .B(n2260), .C(n952), .D(n939), .E(n2469), .F(n429), 
        .Y(n430) );
  OA22XL U841 ( .A(n2433), .B(n627), .C(n1641), .D(n938), .Y(n431) );
  NOR2XL U842 ( .A(n1555), .B(n870), .Y(n172) );
  NOR2XL U843 ( .A(n1555), .B(n881), .Y(n173) );
  OAI22X1 U844 ( .A(n2259), .B(n1974), .C(n2264), .D(n2318), .Y(N12827) );
  OAI22X1 U845 ( .A(n909), .B(n36), .C(n727), .D(n679), .Y(N12844) );
  OAI22X1 U846 ( .A(n909), .B(n2371), .C(n722), .D(n2317), .Y(N12845) );
  ENOX1 U847 ( .A(n2265), .B(n2318), .C(n829), .D(n2318), .Y(N12828) );
  OAI22X1 U848 ( .A(n437), .B(n1974), .C(n2270), .D(n67), .Y(N12826) );
  OAI22X1 U849 ( .A(n909), .B(n2420), .C(n732), .D(n2317), .Y(N12843) );
  OAI22X1 U850 ( .A(n909), .B(n29), .C(n717), .D(n679), .Y(N12846) );
  ENOX1 U851 ( .A(n2266), .B(n2318), .C(n830), .D(n2318), .Y(N12829) );
  MUX2X1 U852 ( .D0(n826), .D1(temp[1]), .S(n1974), .Y(N12825) );
  OAI22X1 U853 ( .A(n909), .B(n2437), .C(n737), .D(n679), .Y(N12842) );
  NAND21X1 U854 ( .B(n686), .A(n685), .Y(n707) );
  OAI221X1 U855 ( .A(n2166), .B(n2345), .C(n784), .D(n2275), .E(n683), .Y(n685) );
  AND3X1 U856 ( .A(n812), .B(n1472), .C(n682), .Y(n686) );
  GEN2XL U857 ( .D(n1472), .E(n928), .C(n2388), .B(n800), .A(n2361), .Y(n683)
         );
  AND4X1 U858 ( .A(n788), .B(n1949), .C(n697), .D(n2176), .Y(n743) );
  OAI22X1 U859 ( .A(n909), .B(n35), .C(n712), .D(n2317), .Y(N12847) );
  OAI22X1 U860 ( .A(n2252), .B(n1974), .C(n2267), .D(n2318), .Y(N12830) );
  OA22X1 U861 ( .A(n807), .B(n681), .C(n811), .D(n928), .Y(n682) );
  AND3X1 U862 ( .A(n806), .B(n800), .C(n2341), .Y(n681) );
  AOI222XL U863 ( .A(n819), .B(n820), .C(n2237), .D(n821), .E(n807), .F(n822), 
        .Y(n811) );
  AND2X1 U864 ( .A(n823), .B(n824), .Y(n807) );
  INVX1 U865 ( .A(N13343), .Y(n2191) );
  NOR4XL U866 ( .A(n825), .B(n826), .C(n827), .D(n828), .Y(n824) );
  OAI22X1 U867 ( .A(n2317), .B(n671), .C(n145), .D(n2418), .Y(N12852) );
  OAI22X1 U868 ( .A(n679), .B(n660), .C(n145), .D(n27), .Y(N12853) );
  OAI22X1 U869 ( .A(n2317), .B(n655), .C(n145), .D(n31), .Y(N12854) );
  OAI22X1 U870 ( .A(n145), .B(n2422), .C(n699), .D(n679), .Y(N12849) );
  OAI22X1 U871 ( .A(n145), .B(n2423), .C(n684), .D(n2317), .Y(N12850) );
  OAI22X1 U872 ( .A(n909), .B(n40), .C(n704), .D(n679), .Y(N12848) );
  AO21X1 U873 ( .B(n832), .C(n2318), .A(n2148), .Y(N12831) );
  OAI22X1 U874 ( .A(n145), .B(n42), .C(n678), .D(n679), .Y(N12851) );
  OAI22X1 U875 ( .A(n679), .B(n650), .C(n145), .D(n38), .Y(N12855) );
  OAI21BBX1 U876 ( .A(n2209), .B(n1945), .C(n1794), .Y(n1793) );
  AOI22X1 U877 ( .A(N11555), .B(n1466), .C(n1467), .D(n2333), .Y(n1464) );
  NAND2X1 U878 ( .A(n1468), .B(n2336), .Y(n1466) );
  INVX1 U879 ( .A(N11555), .Y(n2399) );
  XNOR2XL U880 ( .A(n1426), .B(n1423), .Y(n1461) );
  OAI22X1 U881 ( .A(n1423), .B(n1424), .C(n1425), .D(n1426), .Y(n1040) );
  AND2X1 U882 ( .A(n1424), .B(n1423), .Y(n1425) );
  OAI222XL U883 ( .A(n466), .B(n633), .C(n1473), .D(n632), .E(n2257), .F(n262), 
        .Y(ramdatao_comb[7]) );
  NOR2X1 U884 ( .A(n2450), .B(n1725), .Y(n1377) );
  AND4X1 U885 ( .A(n2162), .B(n2168), .C(n1518), .D(n1705), .Y(n672) );
  OAI21X1 U886 ( .B(n1611), .C(n1612), .A(n1613), .Y(n583) );
  OAI21BBX1 U887 ( .A(n1612), .B(n1611), .C(n1614), .Y(n1613) );
  OAI21X1 U888 ( .B(n1377), .C(n2433), .A(n2438), .Y(n586) );
  OAI21X1 U889 ( .B(n1422), .C(n1040), .A(n1082), .Y(n1081) );
  INVX1 U890 ( .A(n1702), .Y(n1678) );
  INVX1 U891 ( .A(n825), .Y(n2261) );
  XNOR2XL U892 ( .A(n1490), .B(n1463), .Y(n1489) );
  AOI21X1 U893 ( .B(n2333), .C(n1467), .A(n1496), .Y(n1490) );
  AOI21X1 U894 ( .B(n2336), .C(n1468), .A(n2399), .Y(n1496) );
  OAI21X1 U895 ( .B(n583), .C(n584), .A(n586), .Y(n585) );
  NOR4XL U896 ( .A(n829), .B(n830), .C(n831), .D(n832), .Y(n823) );
  AOI32XL U897 ( .A(n1705), .B(n2164), .C(codefetch_s), .D(n708), .E(n1521), 
        .Y(n657) );
  NAND2X1 U898 ( .A(n1422), .B(n1040), .Y(n1082) );
  INVX1 U899 ( .A(n1378), .Y(n2451) );
  INVX1 U900 ( .A(n1610), .Y(n2450) );
  NAND31X1 U901 ( .C(n1755), .A(n2209), .B(n1945), .Y(n1868) );
  NAND21X1 U902 ( .B(n1551), .A(n667), .Y(n643) );
  MUX2X1 U903 ( .D0(ramsfraddr[0]), .D1(n1550), .S(n261), .Y(
        ramsfraddr_comb[0]) );
  MUX2X1 U904 ( .D0(ramsfraddr[1]), .D1(n174), .S(n261), .Y(ramsfraddr_comb[1]) );
  MUX2X1 U905 ( .D0(ramsfraddr[2]), .D1(n3), .S(n261), .Y(ramsfraddr_comb[2])
         );
  XNOR2XL U906 ( .A(n2399), .B(n1468), .Y(n1528) );
  OAI222XL U907 ( .A(n1945), .B(n1516), .C(n1794), .D(n892), .E(n1868), .F(
        n2195), .Y(n1550) );
  OAI21X1 U908 ( .B(n1080), .C(n1081), .A(n1082), .Y(n1041) );
  INVX1 U909 ( .A(n884), .Y(n2247) );
  OAI222XL U910 ( .A(n725), .B(n1868), .C(n2258), .D(n1794), .E(n1945), .F(
        n2197), .Y(n174) );
  NAND2X1 U911 ( .A(n2458), .B(n2459), .Y(n1495) );
  INVX1 U912 ( .A(n820), .Y(n2237) );
  AO222X1 U913 ( .A(n1176), .B(n2146), .C(n830), .D(n479), .E(n1482), .F(n2320), .Y(n500) );
  INVX1 U914 ( .A(n624), .Y(n479) );
  XNOR2XL U915 ( .A(n1444), .B(n1500), .Y(n1482) );
  OAI222XL U916 ( .A(n469), .B(n633), .C(n1474), .D(n632), .E(n2255), .F(
        waitstaten), .Y(ramdatao_comb[6]) );
  OAI222XL U917 ( .A(n470), .B(n633), .C(n1475), .D(n632), .E(n2256), .F(
        waitstaten), .Y(ramdatao_comb[5]) );
  AOI22X1 U918 ( .A(n1441), .B(n2320), .C(n2146), .D(n1165), .Y(n1439) );
  XOR2X1 U919 ( .A(n1402), .B(n1443), .Y(n1441) );
  XNOR2XL U920 ( .A(n1401), .B(n2149), .Y(n1443) );
  AOI222XL U921 ( .A(n2150), .B(ramdatai[3]), .C(n2151), .D(sfrdatai[3]), .E(
        n2152), .F(n1950), .Y(n1534) );
  INVX1 U922 ( .A(memdatai[6]), .Y(n2208) );
  INVX1 U923 ( .A(n501), .Y(n470) );
  NAND41X1 U924 ( .D(n500), .A(n499), .B(n498), .C(n497), .Y(n501) );
  OA222X1 U925 ( .A(n29), .B(n953), .C(n934), .D(n493), .E(n2359), .F(n2315), 
        .Y(n498) );
  OA222X1 U926 ( .A(n2467), .B(n2338), .C(n1541), .D(n494), .E(n31), .F(n2311), 
        .Y(n497) );
  INVX1 U927 ( .A(n936), .Y(n2136) );
  NAND31X1 U928 ( .C(n1729), .A(n1718), .B(n1717), .Y(n1711) );
  AO222X1 U929 ( .A(n326), .B(n325), .C(n324), .D(n323), .E(n406), .F(n2169), 
        .Y(n936) );
  AND4X1 U930 ( .A(n1910), .B(n1911), .C(n1908), .D(n1909), .Y(n325) );
  AND4X1 U931 ( .A(n1918), .B(n1919), .C(n1916), .D(n1917), .Y(n323) );
  AND4X1 U932 ( .A(n1906), .B(n1907), .C(n1904), .D(n1905), .Y(n326) );
  NAND41X1 U933 ( .D(n13), .A(n2033), .B(n2034), .C(n2035), .Y(n1802) );
  XNOR2XL U934 ( .A(n2432), .B(n2394), .Y(n2033) );
  XNOR2XL U935 ( .A(n2447), .B(n2309), .Y(n2034) );
  NOR3XL U936 ( .A(n2036), .B(n2037), .C(n2038), .Y(n2035) );
  MUX2BXL U937 ( .D0(n695), .D1(n694), .S(codefetch_s), .Y(n796) );
  NAND21X1 U938 ( .B(n693), .A(n689), .Y(n695) );
  AND2X1 U939 ( .A(n1515), .B(n2164), .Y(n694) );
  OAI221X1 U940 ( .A(n2275), .B(n688), .C(n2166), .D(n164), .E(n745), .Y(n689)
         );
  OAI221X1 U941 ( .A(n2432), .B(n1795), .C(n2322), .D(n2394), .E(n1922), .Y(
        n888) );
  OA222X1 U942 ( .A(n2264), .B(n1796), .C(n1087), .D(n2312), .E(n941), .F(
        n1797), .Y(n1922) );
  OAI211X1 U943 ( .C(n1573), .D(n12), .A(irq), .B(n182), .Y(n1515) );
  OAI221X1 U944 ( .A(n2447), .B(n1795), .C(n2322), .D(n2309), .E(n1899), .Y(
        n893) );
  OA222X1 U945 ( .A(n2265), .B(n1796), .C(n1086), .D(n2312), .E(n936), .F(
        n1797), .Y(n1899) );
  OAI211X1 U946 ( .C(n149), .D(n2308), .A(n1713), .B(n1712), .Y(n1715) );
  NOR2X1 U947 ( .A(n2172), .B(n2436), .Y(n752) );
  NOR3XL U948 ( .A(n1374), .B(n1373), .C(n2303), .Y(n1459) );
  XNOR2XL U949 ( .A(n2440), .B(n2360), .Y(n2038) );
  OAI222XL U950 ( .A(n471), .B(n633), .C(n1413), .D(n632), .E(n2169), .F(
        waitstaten), .Y(ramdatao_comb[4]) );
  NOR2X1 U951 ( .A(n2430), .B(n2408), .Y(n1781) );
  NOR2X1 U952 ( .A(n1429), .B(n2182), .Y(n1364) );
  NOR2X1 U953 ( .A(n1037), .B(n1370), .Y(n1432) );
  NOR2X1 U954 ( .A(n1715), .B(n149), .Y(n1369) );
  NOR2X1 U955 ( .A(n1035), .B(n1038), .Y(n1362) );
  NAND3X1 U956 ( .A(n2440), .B(n2443), .C(n2444), .Y(n851) );
  INVX1 U957 ( .A(n1365), .Y(n2305) );
  INVX1 U958 ( .A(n1430), .Y(n2182) );
  AOI33X1 U959 ( .A(n885), .B(n2258), .C(n886), .D(n887), .E(n888), .F(n889), 
        .Y(n883) );
  OAI21X1 U960 ( .B(n885), .C(n890), .A(n891), .Y(n887) );
  NOR3XL U961 ( .A(n894), .B(n889), .C(n892), .Y(n886) );
  NAND4X1 U962 ( .A(n892), .B(n885), .C(n890), .D(n893), .Y(n891) );
  INVX1 U963 ( .A(n2040), .Y(n2360) );
  INVX1 U964 ( .A(n468), .Y(n471) );
  NAND41X1 U965 ( .D(n467), .A(n465), .B(n464), .C(n463), .Y(n468) );
  OA222X1 U966 ( .A(n2371), .B(n953), .C(n934), .D(n450), .E(n2359), .F(n2332), 
        .Y(n465) );
  OA222X1 U967 ( .A(n2468), .B(n2338), .C(n624), .D(n453), .E(n1543), .F(n452), 
        .Y(n464) );
  GEN2XL U968 ( .D(n2249), .E(n1842), .C(n2276), .B(n1843), .A(n1840), .Y(
        n1841) );
  INVX1 U969 ( .A(n1839), .Y(n2249) );
  NOR21XL U970 ( .B(n1712), .A(n1713), .Y(n1370) );
  OA2222XL U971 ( .A(n1795), .B(n2173), .C(n2271), .D(n1796), .E(n1083), .F(
        n2312), .G(n1797), .H(n917), .Y(n895) );
  INVX1 U972 ( .A(n931), .Y(n2087) );
  AO222X1 U973 ( .A(n295), .B(n294), .C(n293), .D(n292), .E(n406), .F(n2414), 
        .Y(n959) );
  AND4X1 U974 ( .A(n2021), .B(n2022), .C(n2019), .D(n2020), .Y(n294) );
  AND4X1 U975 ( .A(n2043), .B(n2044), .C(n2041), .D(n2042), .Y(n292) );
  AND4X1 U976 ( .A(n2016), .B(n2017), .C(n2014), .D(n2015), .Y(n295) );
  AO222X1 U977 ( .A(n410), .B(n409), .C(n408), .D(n407), .E(n406), .F(n2415), 
        .Y(n952) );
  AND4X1 U978 ( .A(n1983), .B(n1984), .C(n1981), .D(n1982), .Y(n409) );
  AND4X1 U979 ( .A(n1991), .B(n1992), .C(n1989), .D(n1990), .Y(n407) );
  AND4X1 U980 ( .A(n1979), .B(n1980), .C(n1977), .D(n1978), .Y(n410) );
  AO222X1 U981 ( .A(n322), .B(n321), .C(n320), .D(n319), .E(n406), .F(n2316), 
        .Y(n946) );
  AND4X1 U982 ( .A(n1957), .B(n1958), .C(n1955), .D(n1956), .Y(n321) );
  AND4X1 U983 ( .A(n1965), .B(n1966), .C(n1963), .D(n1964), .Y(n319) );
  AND4X1 U984 ( .A(n1953), .B(n1954), .C(n1951), .D(n1952), .Y(n322) );
  OA2222XL U985 ( .A(n2445), .B(n1795), .C(n2266), .D(n1796), .E(n931), .F(
        n1797), .G(n1085), .H(n2312), .Y(n885) );
  NAND21X1 U986 ( .B(n853), .A(n1234), .Y(n1844) );
  NAND21X1 U987 ( .B(n2358), .A(n1014), .Y(n2351) );
  AOI21X1 U988 ( .B(n697), .C(n2006), .A(n1837), .Y(n1866) );
  AO21X1 U989 ( .B(n280), .C(n1479), .A(n1477), .Y(n281) );
  NOR21XL U990 ( .B(n1944), .A(N12772), .Y(n1921) );
  NOR21XL U991 ( .B(n1970), .A(N12771), .Y(n1944) );
  NOR2X1 U992 ( .A(n2172), .B(n2407), .Y(n753) );
  OAI221X1 U993 ( .A(n2440), .B(n1795), .C(n2322), .D(n102), .E(n1971), .Y(
        n890) );
  OA222X1 U994 ( .A(n2269), .B(n1796), .C(n1089), .D(n2312), .E(n952), .F(
        n1797), .Y(n1971) );
  AND2X1 U995 ( .A(n1766), .B(n1791), .Y(n175) );
  AND3X1 U996 ( .A(n2445), .B(n1352), .C(n2441), .Y(n1114) );
  AOI22X1 U997 ( .A(n2395), .B(n1027), .C(n2435), .D(n2428), .Y(n2047) );
  OAI221X1 U998 ( .A(n2443), .B(n1795), .C(n2322), .D(n26), .E(n1946), .Y(n884) );
  OA222X1 U999 ( .A(n2270), .B(n1796), .C(n1088), .D(n2312), .E(n946), .F(
        n1797), .Y(n1946) );
  MUX2AXL U1000 ( .D0(n2435), .D1(n1662), .S(n262), .Y(ramdatao_comb[3]) );
  OAI22X1 U1001 ( .A(n909), .B(n33), .C(n742), .D(n2317), .Y(N12841) );
  AOI22X1 U1002 ( .A(n2310), .B(n1027), .C(n2169), .D(n2428), .Y(n2018) );
  AOI222XL U1003 ( .A(n1866), .B(n1870), .C(n1920), .D(N12773), .E(N12805), 
        .F(n1837), .Y(n1086) );
  OAI21X1 U1004 ( .B(n1921), .C(n2276), .A(n1843), .Y(n1920) );
  AOI222XL U1005 ( .A(n1866), .B(n1970), .C(n1993), .D(N12770), .E(N12802), 
        .F(n1837), .Y(n1089) );
  OAI21X1 U1006 ( .B(n1994), .C(n2276), .A(n1843), .Y(n1993) );
  AOI222XL U1007 ( .A(n1866), .B(n1921), .C(n1943), .D(N12772), .E(N12804), 
        .F(n1837), .Y(n1087) );
  OAI21X1 U1008 ( .B(n1944), .C(n2276), .A(n1843), .Y(n1943) );
  AOI211X1 U1009 ( .C(N12808), .D(n1837), .A(n2243), .B(n1838), .Y(n1083) );
  NOR4XL U1010 ( .A(n2276), .B(n1839), .C(n2250), .D(n106), .Y(n1838) );
  INVX1 U1011 ( .A(n1841), .Y(n2243) );
  AND2X1 U1012 ( .A(n1114), .B(n859), .Y(n1234) );
  NOR2X1 U1013 ( .A(n26), .B(n2048), .Y(n2039) );
  XNOR2XL U1014 ( .A(n2443), .B(n2039), .Y(n2037) );
  NAND3X1 U1015 ( .A(n1114), .B(n862), .C(n864), .Y(n484) );
  NOR4XL U1016 ( .A(n2168), .B(n255), .C(n774), .D(n2404), .Y(n1687) );
  NAND2X1 U1017 ( .A(n979), .B(n1791), .Y(n774) );
  NAND3X1 U1018 ( .A(n2313), .B(n68), .C(n2006), .Y(n1843) );
  NAND3X1 U1019 ( .A(n1375), .B(n2445), .C(n862), .Y(n1027) );
  INVX1 U1020 ( .A(n1994), .Y(n217) );
  OAI222XL U1021 ( .A(n1410), .B(n1409), .C(n1408), .D(n1407), .E(n1199), .F(
        n1543), .Y(n1537) );
  AOI211XL U1022 ( .C(n1406), .D(n351), .A(n1405), .B(n1404), .Y(n1408) );
  XOR2X1 U1023 ( .A(n1533), .B(n1548), .Y(n1409) );
  GEN2XL U1024 ( .D(n1397), .E(n2138), .C(n1392), .B(n1389), .A(n1385), .Y(
        n1405) );
  INVX1 U1025 ( .A(n1738), .Y(n2407) );
  INVX1 U1026 ( .A(n808), .Y(n2358) );
  INVX1 U1027 ( .A(n309), .Y(n312) );
  NAND32X1 U1028 ( .B(n2170), .C(n2409), .A(n2147), .Y(n309) );
  INVX1 U1029 ( .A(n1467), .Y(n2336) );
  INVX1 U1030 ( .A(n765), .Y(n2411) );
  NOR2X1 U1031 ( .A(n2387), .B(n2360), .Y(n2027) );
  INVX1 U1032 ( .A(n1690), .Y(n2409) );
  AOI22AXL U1033 ( .A(N11584), .B(n1058), .D(N11584), .C(n1059), .Y(n1057) );
  INVX1 U1034 ( .A(n776), .Y(n2386) );
  MUX2AXL U1035 ( .D0(n1536), .D1(n901), .S(n2075), .Y(n1662) );
  NOR4XL U1036 ( .A(n1537), .B(n1538), .C(n1539), .D(n1540), .Y(n1536) );
  OAI22X1 U1037 ( .A(n2359), .B(n2400), .C(n953), .D(n36), .Y(n1540) );
  ENOX1 U1038 ( .A(n2311), .B(n2418), .C(n392), .D(pc_i[3]), .Y(n1539) );
  INVX1 U1039 ( .A(n1344), .Y(n2391) );
  INVX1 U1040 ( .A(n1345), .Y(n2298) );
  ENOX1 U1041 ( .A(n466), .B(n1379), .C(n2075), .D(n1875), .Y(N11505) );
  NOR2X1 U1042 ( .A(n217), .B(N12770), .Y(n1970) );
  NAND4X1 U1043 ( .A(n1074), .B(n1037), .C(n1067), .D(n1075), .Y(n1059) );
  INVX1 U1044 ( .A(n831), .Y(n2252) );
  INVX1 U1045 ( .A(n1468), .Y(n2333) );
  INVX1 U1046 ( .A(n1716), .Y(n2307) );
  INVX1 U1047 ( .A(n1837), .Y(n2313) );
  NOR32XL U1048 ( .B(n849), .C(n1716), .A(n1715), .Y(n1044) );
  NOR21XL U1049 ( .B(n1717), .A(n1718), .Y(n1073) );
  NAND21X1 U1050 ( .B(n2170), .A(n1684), .Y(n2373) );
  NOR21XL U1051 ( .B(n1921), .A(N12773), .Y(n1870) );
  OA2222XL U1052 ( .A(n2312), .B(n1084), .C(n926), .D(n1797), .E(n1795), .F(
        n2441), .G(n2267), .H(n1796), .Y(n889) );
  NAND32XL U1053 ( .B(n256), .C(n2167), .A(n456), .Y(n505) );
  NOR2X1 U1054 ( .A(n2168), .B(n252), .Y(intcall) );
  AOI222XL U1055 ( .A(n2277), .B(n125), .C(N12806), .D(n1837), .E(n1866), .F(
        n1869), .Y(n1085) );
  OAI21X1 U1056 ( .B(n1870), .C(n1871), .A(n1839), .Y(n1869) );
  AOI222XL U1057 ( .A(n1866), .B(n1944), .C(n1967), .D(N12771), .E(N12803), 
        .F(n1837), .Y(n1088) );
  OAI21X1 U1058 ( .B(n1970), .C(n2276), .A(n1843), .Y(n1967) );
  AOI222XL U1059 ( .A(n1866), .B(n1994), .C(n2277), .D(n217), .E(N12801), .F(
        n1837), .Y(n1090) );
  AOI222XL U1060 ( .A(n2277), .B(n2250), .C(N12807), .D(n1837), .E(n1865), .F(
        n1866), .Y(n1084) );
  XNOR2XL U1061 ( .A(n2250), .B(n1839), .Y(n1865) );
  NOR2X1 U1062 ( .A(n2411), .B(n2172), .Y(n1742) );
  OA222X1 U1063 ( .A(n612), .B(n297), .C(n1498), .D(n2459), .E(n2458), .F(
        n2306), .Y(n298) );
  INVX1 U1064 ( .A(n1073), .Y(n297) );
  XNOR2XL U1065 ( .A(n1376), .B(n2369), .Y(n1424) );
  XNOR2XL U1066 ( .A(n1376), .B(n2334), .Y(n1465) );
  NOR2X1 U1067 ( .A(n2431), .B(n2408), .Y(n1684) );
  INVX1 U1068 ( .A(n1871), .Y(n125) );
  AND3X1 U1069 ( .A(n1717), .B(n1718), .C(n1729), .Y(n1056) );
  NOR2X1 U1070 ( .A(n2436), .B(n2408), .Y(n1682) );
  OAI222XL U1071 ( .A(n472), .B(n633), .C(n1006), .D(n632), .E(n2316), .F(
        waitstaten), .Y(ramdatao_comb[2]) );
  INVX1 U1072 ( .A(n1372), .Y(n411) );
  NAND2X1 U1073 ( .A(n1870), .B(n1871), .Y(n1839) );
  INVX1 U1074 ( .A(n259), .Y(n255) );
  INVX1 U1075 ( .A(n2361), .Y(n259) );
  INVX1 U1076 ( .A(n254), .Y(n252) );
  INVX1 U1077 ( .A(n819), .Y(n2379) );
  INVX1 U1078 ( .A(ramdatai[4]), .Y(n2468) );
  INVX1 U1079 ( .A(ramdatai[5]), .Y(n2467) );
  OAI222XL U1080 ( .A(n2466), .B(n2338), .C(n624), .D(n623), .E(n622), .F(
        n1407), .Y(n625) );
  INVX1 U1081 ( .A(n832), .Y(n623) );
  AOI222XL U1082 ( .A(n619), .B(n351), .C(n617), .D(n616), .E(n615), .F(n614), 
        .Y(n622) );
  INVX1 U1083 ( .A(n2012), .Y(n616) );
  INVX1 U1084 ( .A(n1015), .Y(n2388) );
  INVX1 U1085 ( .A(ramdatai[7]), .Y(n2466) );
  INVX1 U1086 ( .A(n448), .Y(n472) );
  NAND43X1 U1087 ( .B(n447), .C(n446), .D(n445), .A(n444), .Y(n448) );
  OAI22X1 U1088 ( .A(n1543), .B(n1211), .C(n1542), .D(n437), .Y(n445) );
  AOI31X1 U1089 ( .A(n1399), .B(n509), .C(n434), .D(n436), .Y(n447) );
  NOR2X1 U1090 ( .A(n2040), .B(n2387), .Y(n2030) );
  INVX1 U1091 ( .A(ramdatai[0]), .Y(n2470) );
  INVX1 U1092 ( .A(ramdatai[1]), .Y(n2469) );
  INVX1 U1093 ( .A(ramdatai[6]), .Y(n735) );
  INVX1 U1094 ( .A(ramdatai[2]), .Y(n715) );
  INVX1 U1095 ( .A(n1047), .Y(n2179) );
  ENOX1 U1096 ( .A(n469), .B(n1379), .C(n2075), .D(n1900), .Y(N11504) );
  INVX1 U1097 ( .A(n1101), .Y(n2393) );
  NOR2X1 U1098 ( .A(n2454), .B(n149), .Y(n1710) );
  INVX1 U1099 ( .A(n2361), .Y(n258) );
  INVX1 U1100 ( .A(n1368), .Y(n2304) );
  INVX1 U1101 ( .A(n828), .Y(n2259) );
  INVX1 U1102 ( .A(n1777), .Y(n2431) );
  NOR32XL U1103 ( .B(n979), .C(n753), .A(n2417), .Y(n1789) );
  NOR21XL U1104 ( .B(n1234), .A(n857), .Y(n487) );
  AOI21X1 U1105 ( .B(n1430), .C(n1429), .A(n1055), .Y(n1498) );
  NOR21XL U1106 ( .B(n275), .A(n1700), .Y(N512) );
  AOI21BBXL U1107 ( .B(n1699), .C(n1698), .A(n1697), .Y(n1700) );
  NOR21XL U1108 ( .B(n10), .A(n1696), .Y(n1697) );
  OAI31XL U1109 ( .A(n252), .B(n2052), .C(n2171), .D(n1758), .Y(n2002) );
  NOR4XL U1110 ( .A(n775), .B(n2161), .C(n1690), .D(n2054), .Y(n2052) );
  MUX2AXL U1111 ( .D0(n2415), .D1(n1675), .S(n262), .Y(ramdatao_comb[1]) );
  MUX2AXL U1112 ( .D0(n2414), .D1(n10), .S(n262), .Y(ramdatao_comb[0]) );
  OR2X1 U1113 ( .A(n219), .B(n176), .Y(n474) );
  AOI21X1 U1114 ( .B(n1544), .C(n1622), .A(n596), .Y(n176) );
  GEN2XL U1115 ( .D(n436), .E(n2138), .C(n1392), .B(n191), .A(n435), .Y(n446)
         );
  AND2XL U1116 ( .A(n1406), .B(n356), .Y(n435) );
  GEN2XL U1117 ( .D(n619), .E(n356), .C(n598), .B(n597), .A(n518), .Y(n599) );
  INVX1 U1118 ( .A(n1407), .Y(n597) );
  OAI22X1 U1119 ( .A(n2338), .B(n735), .C(n624), .D(n2252), .Y(n518) );
  GEN2XL U1120 ( .D(n517), .E(n2138), .C(n1392), .B(n190), .A(n510), .Y(n598)
         );
  NOR2X1 U1121 ( .A(n2416), .B(n25), .Y(n764) );
  OA222X1 U1122 ( .A(n462), .B(n459), .C(n458), .D(n457), .E(n2273), .F(n505), 
        .Y(n463) );
  INVX1 U1123 ( .A(n1517), .Y(n458) );
  AND3X1 U1124 ( .A(n1520), .B(n183), .C(n454), .Y(n459) );
  OA22X1 U1125 ( .A(n1544), .B(n1622), .C(n1705), .D(n1521), .Y(n1546) );
  NAND32X1 U1126 ( .B(n1677), .C(n220), .A(n1678), .Y(n1704) );
  NAND2X1 U1127 ( .A(n2053), .B(n753), .Y(n780) );
  XNOR2XL U1128 ( .A(n177), .B(n1614), .Y(n1721) );
  XNOR2XL U1129 ( .A(n1612), .B(n1611), .Y(n177) );
  NOR2X1 U1130 ( .A(n2172), .B(n2170), .Y(n1748) );
  AOI222XL U1131 ( .A(n2150), .B(ramdatai[6]), .C(n2151), .D(sfrdatai[6]), .E(
        n2152), .F(n2072), .Y(n1401) );
  INVX1 U1132 ( .A(n926), .Y(n2072) );
  INVX1 U1133 ( .A(n2011), .Y(n496) );
  NAND2X1 U1134 ( .A(n2390), .B(n2392), .Y(n1111) );
  INVX1 U1135 ( .A(n596), .Y(codefetch_s) );
  AOI222XL U1136 ( .A(n2151), .B(sfrdatai[7]), .C(ramdatai[7]), .D(n2150), .E(
        n2013), .F(n2152), .Y(n1396) );
  INVX1 U1137 ( .A(n917), .Y(n2013) );
  NOR2X1 U1138 ( .A(n1109), .B(n2293), .Y(n204) );
  NAND2X1 U1139 ( .A(n1945), .B(n1755), .Y(n1794) );
  OAI31XL U1140 ( .A(n1678), .B(cs_run), .C(n1677), .D(n1696), .Y(n1698) );
  OAI32X1 U1141 ( .A(n1616), .B(n1603), .C(n1668), .D(n1602), .E(n220), .Y(
        N582) );
  INVX1 U1142 ( .A(n1600), .Y(n1616) );
  INVX1 U1143 ( .A(n1601), .Y(n1602) );
  OAI32X1 U1144 ( .A(n476), .B(n270), .C(n2192), .D(n477), .E(n2162), .Y(n1973) );
  INVX1 U1145 ( .A(n477), .Y(n2192) );
  OAI211X1 U1146 ( .C(n478), .D(codefetch_s), .A(n265), .B(n1622), .Y(n477) );
  OA21X1 U1147 ( .B(n1546), .C(n1545), .A(n596), .Y(n476) );
  INVX1 U1148 ( .A(n826), .Y(n2260) );
  OAI22X1 U1149 ( .A(n2164), .B(n1704), .C(n1660), .D(n1676), .Y(n1880) );
  NOR2X1 U1150 ( .A(n2377), .B(n2436), .Y(n2054) );
  AND2X1 U1151 ( .A(n1689), .B(n264), .Y(N515) );
  OAI22X1 U1152 ( .A(n1688), .B(n1696), .C(n1685), .D(n1698), .Y(n1689) );
  AND2X1 U1153 ( .A(n1676), .B(n2164), .Y(n1685) );
  INVXL U1154 ( .A(n1675), .Y(n1688) );
  INVX1 U1155 ( .A(ramdatai[3]), .Y(n720) );
  OAI32X1 U1156 ( .A(n2050), .B(n2404), .C(n256), .D(n2051), .E(n2324), .Y(
        n2007) );
  AOI21X1 U1157 ( .B(n1781), .C(n2048), .A(n764), .Y(n2051) );
  INVX1 U1158 ( .A(n2048), .Y(n2416) );
  AOI31X1 U1159 ( .A(n1558), .B(n1399), .C(n1398), .D(n1397), .Y(n1404) );
  EORX1 U1160 ( .A(n1903), .B(n2138), .C(n1903), .D(n2140), .Y(n1558) );
  NAND21X1 U1161 ( .B(n1544), .A(n1622), .Y(n601) );
  NAND2X1 U1162 ( .A(n317), .B(n911), .Y(n1452) );
  NAND21X1 U1163 ( .B(n2171), .A(n2161), .Y(n2372) );
  AO21X1 U1164 ( .B(n348), .C(n347), .A(n2173), .Y(n355) );
  INVX1 U1165 ( .A(n350), .Y(n348) );
  OR2X1 U1166 ( .A(n252), .B(n178), .Y(n438) );
  AOI21X1 U1167 ( .B(n765), .C(n2158), .A(n306), .Y(n178) );
  AO21X1 U1168 ( .B(n972), .C(n1690), .A(n809), .Y(n306) );
  OAI211X1 U1169 ( .C(n256), .D(n305), .A(n381), .B(n438), .Y(n2320) );
  OA22X1 U1170 ( .A(n2411), .B(n383), .C(n2409), .D(n2188), .Y(n305) );
  NAND3X1 U1171 ( .A(n1695), .B(n792), .C(n1026), .Y(n933) );
  OAI22X1 U1172 ( .A(n2373), .B(n285), .C(n383), .D(n2407), .Y(n318) );
  INVX1 U1173 ( .A(n1737), .Y(n285) );
  OAI221X1 U1174 ( .A(n257), .B(n1655), .C(n1657), .D(n2275), .E(n341), .Y(
        n350) );
  AND2X1 U1175 ( .A(n2139), .B(n2140), .Y(n341) );
  NAND5XL U1176 ( .A(n404), .B(n1410), .C(n1407), .D(n2359), .E(n403), .Y(
        n1004) );
  AND4X1 U1177 ( .A(n2311), .B(n1541), .C(n451), .D(n934), .Y(n403) );
  AOI21X1 U1178 ( .B(n1690), .C(n1691), .A(n805), .Y(n587) );
  OAI211X1 U1179 ( .C(n344), .D(n343), .A(n340), .B(n316), .Y(n592) );
  AND2X1 U1180 ( .A(n2117), .B(n317), .Y(n316) );
  AND2X1 U1181 ( .A(n1643), .B(n1655), .Y(n2117) );
  OAI211X1 U1182 ( .C(n2356), .D(n344), .A(n2186), .B(n340), .Y(n367) );
  OA222X1 U1183 ( .A(n492), .B(n491), .C(n490), .D(n489), .E(n488), .F(n505), 
        .Y(n499) );
  INVX1 U1184 ( .A(n1478), .Y(n490) );
  AND3X1 U1185 ( .A(n1481), .B(n183), .C(n480), .Y(n491) );
  OAI211X1 U1186 ( .C(n2412), .D(n2416), .A(n762), .B(n763), .Y(n618) );
  AOI221XL U1187 ( .A(n764), .B(n765), .C(n766), .D(n152), .E(n2187), .Y(n763)
         );
  NAND21X1 U1188 ( .B(n2056), .A(n1026), .Y(n369) );
  NOR3XL U1189 ( .A(n285), .B(n2170), .C(n2409), .Y(n591) );
  NOR2X1 U1190 ( .A(n2358), .B(n2408), .Y(n1336) );
  NOR2X1 U1191 ( .A(n26), .B(n2170), .Y(n758) );
  INVX1 U1192 ( .A(n2356), .Y(n2157) );
  NAND2X1 U1193 ( .A(n864), .B(n1234), .Y(n1151) );
  NOR2X1 U1194 ( .A(n2417), .B(n2387), .Y(n910) );
  NOR2X1 U1195 ( .A(n1023), .B(n2275), .Y(n1148) );
  INVX1 U1196 ( .A(n980), .Y(n2406) );
  INVX1 U1197 ( .A(n781), .Y(n2412) );
  INVX1 U1198 ( .A(n343), .Y(n2156) );
  NAND2X1 U1199 ( .A(n2048), .B(n979), .Y(n2050) );
  NOR2X1 U1200 ( .A(n1111), .B(n2293), .Y(n202) );
  NOR2X1 U1201 ( .A(n1110), .B(n2293), .Y(n198) );
  INVX1 U1202 ( .A(n982), .Y(n2413) );
  NOR2X1 U1203 ( .A(n1107), .B(n2293), .Y(n200) );
  INVX1 U1204 ( .A(n418), .Y(n1399) );
  NOR2X1 U1205 ( .A(n1111), .B(n2293), .Y(n201) );
  NOR2X1 U1206 ( .A(n1110), .B(n2293), .Y(n197) );
  NOR2X1 U1207 ( .A(n1111), .B(n127), .Y(n519) );
  NOR2X1 U1208 ( .A(n1110), .B(n127), .Y(n521) );
  NOR2X1 U1209 ( .A(n1109), .B(n2293), .Y(n203) );
  NOR2X1 U1210 ( .A(n1107), .B(n2293), .Y(n199) );
  NOR2X1 U1211 ( .A(n1109), .B(n2293), .Y(n520) );
  NOR2X1 U1212 ( .A(n1107), .B(n127), .Y(n522) );
  INVX1 U1213 ( .A(n254), .Y(n253) );
  INVX1 U1214 ( .A(n1842), .Y(n2250) );
  OAI22X1 U1215 ( .A(n593), .B(n1623), .C(n594), .D(codefetch_s), .Y(N679) );
  INVX1 U1216 ( .A(n1622), .Y(n1623) );
  INVX1 U1217 ( .A(n1683), .Y(n2343) );
  NOR3XL U1218 ( .A(n2196), .B(n596), .C(n601), .Y(N671) );
  INVX1 U1219 ( .A(n621), .Y(n688) );
  GEN2XL U1220 ( .D(n751), .E(n752), .C(n753), .B(n754), .A(n755), .Y(n621) );
  EORX1 U1221 ( .A(n756), .B(n2436), .C(n757), .D(n2436), .Y(n754) );
  OAI211X1 U1222 ( .C(n758), .D(n102), .A(n759), .B(n760), .Y(n756) );
  INVX1 U1223 ( .A(n1840), .Y(n106) );
  NOR2X1 U1224 ( .A(n60), .B(n2464), .Y(N14336) );
  AOI31X1 U1225 ( .A(n509), .B(n183), .C(n508), .D(n517), .Y(n510) );
  MUX2X1 U1226 ( .D0(n507), .D1(n2140), .S(n190), .Y(n508) );
  INVX1 U1227 ( .A(n880), .Y(n2424) );
  INVX1 U1228 ( .A(n1014), .Y(n2389) );
  INVX1 U1229 ( .A(n1791), .Y(n2385) );
  OA21X1 U1230 ( .B(n627), .C(n2332), .A(n1505), .Y(n475) );
  OA22X1 U1231 ( .A(n628), .B(n725), .C(n936), .D(n939), .Y(n473) );
  AOI22X1 U1232 ( .A(n829), .B(n1386), .C(ramdatai[4]), .D(n1387), .Y(n1505)
         );
  INVX1 U1233 ( .A(n504), .Y(n1475) );
  OA21X1 U1234 ( .B(n627), .C(n2315), .A(n1469), .Y(n503) );
  OA22X1 U1235 ( .A(n628), .B(n730), .C(n931), .D(n939), .Y(n502) );
  GEN2XL U1236 ( .D(n1749), .E(n1750), .C(n51), .B(n2372), .A(n2324), .Y(n1743) );
  AOI21X1 U1237 ( .B(n752), .C(n2170), .A(n775), .Y(n1749) );
  NAND31X1 U1238 ( .C(n1739), .A(n400), .B(n399), .Y(n1509) );
  OR2X1 U1239 ( .A(n2173), .B(n381), .Y(n382) );
  NAND21X1 U1240 ( .B(n2171), .A(n819), .Y(n384) );
  NAND2X1 U1241 ( .A(n1508), .B(n1507), .Y(n1561) );
  NAND21X1 U1242 ( .B(n384), .A(n1738), .Y(n296) );
  OAI22X1 U1243 ( .A(n253), .B(n291), .C(n257), .D(n290), .Y(n2325) );
  AND3X1 U1244 ( .A(n1730), .B(n1753), .C(n986), .Y(n291) );
  AND3X1 U1245 ( .A(n669), .B(n668), .C(n289), .Y(n290) );
  AOI32X1 U1246 ( .A(n1683), .B(n981), .C(n1015), .D(n1738), .E(n1754), .Y(
        n1753) );
  NAND32X1 U1247 ( .B(n1739), .C(n400), .A(n399), .Y(n627) );
  OAI31XL U1248 ( .A(n687), .B(n2324), .C(n2352), .D(n1102), .Y(n1449) );
  NOR42XL U1249 ( .C(n801), .D(n802), .A(n803), .B(n804), .Y(n784) );
  NOR2X1 U1250 ( .A(n591), .B(n805), .Y(n802) );
  INVX1 U1251 ( .A(n631), .Y(n1473) );
  OAI211XL U1252 ( .C(n1638), .D(n938), .A(n630), .B(n629), .Y(n631) );
  OA22X1 U1253 ( .A(n2209), .B(n628), .C(n917), .D(n939), .Y(n629) );
  OA21X1 U1254 ( .B(n627), .C(n746), .A(n1382), .Y(n630) );
  INVX1 U1255 ( .A(n680), .Y(n1972) );
  NAND32X1 U1256 ( .B(n2384), .C(n2356), .A(n822), .Y(n680) );
  NAND31X1 U1257 ( .C(n14), .A(n1743), .B(n628), .Y(n1739) );
  NAND32X1 U1258 ( .B(n2172), .C(n344), .A(n2157), .Y(n1643) );
  INVX1 U1259 ( .A(n871), .Y(n671) );
  INVX1 U1260 ( .A(n899), .Y(n660) );
  INVX1 U1261 ( .A(n904), .Y(n655) );
  NOR2X1 U1262 ( .A(n2377), .B(n2171), .Y(n1681) );
  NAND2X1 U1263 ( .A(n1777), .B(n56), .Y(n1694) );
  NOR2X1 U1264 ( .A(n2172), .B(n2387), .Y(n1695) );
  OAI211X1 U1265 ( .C(n2400), .D(n627), .A(n1559), .B(n1560), .Y(n901) );
  AOI222XL U1266 ( .A(memdatai[3]), .B(n2325), .C(n2154), .D(n1950), .E(
        ramdatai[3]), .F(n1561), .Y(n1560) );
  AOI22X1 U1267 ( .A(n2153), .B(n828), .C(sfrdatai[3]), .D(n2155), .Y(n1559)
         );
  NAND2X1 U1268 ( .A(n1690), .B(n2189), .Y(n589) );
  OAI21X1 U1269 ( .B(n2351), .C(n2409), .A(n1023), .Y(n783) );
  INVX1 U1270 ( .A(n344), .Y(n2144) );
  NOR2X1 U1271 ( .A(n2171), .B(n2170), .Y(n972) );
  AND2X1 U1272 ( .A(n2053), .B(n1738), .Y(n1999) );
  AOI32X1 U1273 ( .A(n1738), .B(n2170), .C(n1014), .D(n1683), .E(n2122), .Y(
        n2119) );
  OAI21X1 U1274 ( .B(n1695), .C(n2413), .A(n2410), .Y(n2122) );
  INVX1 U1275 ( .A(n822), .Y(n2380) );
  NOR3XL U1276 ( .A(n1067), .B(n2244), .C(n2241), .Y(n1064) );
  NOR2X1 U1277 ( .A(n2459), .B(n2464), .Y(N14344) );
  OR2X1 U1278 ( .A(n1754), .B(n1691), .Y(n2066) );
  INVX1 U1279 ( .A(n727), .Y(n719) );
  INVX1 U1280 ( .A(n732), .Y(n714) );
  INVX1 U1281 ( .A(n609), .Y(n2253) );
  NOR2X1 U1282 ( .A(n1684), .B(n1690), .Y(n1763) );
  INVX1 U1283 ( .A(n1075), .Y(n2244) );
  INVX1 U1284 ( .A(n1066), .Y(n2241) );
  OAI211X1 U1285 ( .C(n2434), .D(n627), .A(n1569), .B(n1570), .Y(n902) );
  AOI222XL U1286 ( .A(memdatai[2]), .B(n2325), .C(n2154), .D(n2137), .E(
        ramdatai[2]), .F(n1561), .Y(n1570) );
  INVX1 U1287 ( .A(n946), .Y(n2137) );
  NAND32X1 U1288 ( .B(n2173), .C(n2325), .A(n14), .Y(n938) );
  NAND32X1 U1289 ( .B(n152), .C(n928), .A(n2144), .Y(n1013) );
  NAND21X1 U1290 ( .B(n2275), .A(n787), .Y(n335) );
  NAND42X1 U1291 ( .C(n777), .D(n778), .A(n779), .B(n780), .Y(n771) );
  NAND2X1 U1292 ( .A(n766), .B(n781), .Y(n779) );
  OAI21X1 U1293 ( .B(n911), .C(n1694), .A(n1657), .Y(n787) );
  NAND21X1 U1294 ( .B(n978), .A(n2413), .Y(n981) );
  NAND3X1 U1295 ( .A(n979), .B(n2171), .C(n1015), .Y(n2059) );
  INVX1 U1296 ( .A(n906), .Y(n650) );
  AND3X1 U1297 ( .A(n2131), .B(n1013), .C(n2132), .Y(n786) );
  OAI21BBX1 U1298 ( .A(n1694), .B(n2128), .C(n2063), .Y(n2131) );
  AOI22X1 U1299 ( .A(n2157), .B(n2133), .C(n2066), .D(n2405), .Y(n2132) );
  OAI211X1 U1300 ( .C(n2379), .D(n2389), .A(n2134), .B(n2056), .Y(n2133) );
  AND2X1 U1301 ( .A(n979), .B(n776), .Y(n1770) );
  NAND2X1 U1302 ( .A(n2054), .B(n1015), .Y(n810) );
  OAI22X1 U1303 ( .A(n773), .B(n2343), .C(n774), .D(n2401), .Y(n772) );
  AOI22X1 U1304 ( .A(n2374), .B(n56), .C(n775), .D(n776), .Y(n773) );
  OAI211X1 U1305 ( .C(n2347), .D(n2092), .A(n2341), .B(n2375), .Y(n1020) );
  NAND2X1 U1306 ( .A(n753), .B(n2417), .Y(n2092) );
  INVX1 U1307 ( .A(n792), .Y(n2381) );
  OAI21X1 U1308 ( .B(n822), .C(n1748), .A(n1015), .Y(n2134) );
  AND2XL U1309 ( .A(n213), .B(n1675), .Y(N11499) );
  AOI211X1 U1310 ( .C(n910), .D(n25), .A(n2408), .B(n1770), .Y(n2097) );
  NAND3X1 U1311 ( .A(n1737), .B(n2379), .C(n765), .Y(n1021) );
  AOI31X1 U1312 ( .A(n2348), .B(n2186), .C(n2091), .D(n2166), .Y(n2090) );
  AOI31X1 U1313 ( .A(n808), .B(n2387), .C(n1742), .D(n1020), .Y(n2091) );
  NAND2X1 U1314 ( .A(n1015), .B(n26), .Y(n1785) );
  INVX1 U1315 ( .A(n667), .Y(n1573) );
  INVX1 U1316 ( .A(n605), .Y(n1474) );
  OAI211XL U1317 ( .C(n1646), .D(n938), .A(n604), .B(n603), .Y(n605) );
  OA22X1 U1318 ( .A(n2208), .B(n628), .C(n926), .D(n939), .Y(n603) );
  OA21X1 U1319 ( .B(n627), .C(n2283), .A(n1435), .Y(n604) );
  NOR2X1 U1320 ( .A(n1742), .B(n781), .Y(n2128) );
  INVX1 U1321 ( .A(n1792), .Y(n2383) );
  MUX2X1 U1322 ( .D0(n2448), .D1(n2268), .S(n1150), .Y(n375) );
  INVX1 U1323 ( .A(n646), .Y(n1619) );
  NAND32X1 U1324 ( .B(n253), .C(n668), .A(n2011), .Y(n646) );
  NAND31X1 U1325 ( .C(n256), .A(n764), .B(n2183), .Y(n399) );
  OAI31XL U1326 ( .A(n687), .B(n2324), .C(n2352), .D(n1102), .Y(n196) );
  OAI31XL U1327 ( .A(n687), .B(n2324), .C(n2352), .D(n1102), .Y(n195) );
  OAI211X1 U1328 ( .C(n789), .D(n257), .A(n790), .B(n2184), .Y(n744) );
  AOI21X1 U1329 ( .B(n608), .C(n792), .A(n2354), .Y(n789) );
  OR4X1 U1330 ( .A(n791), .B(n610), .C(n2401), .D(n2358), .Y(n790) );
  NAND21X1 U1331 ( .B(n2139), .A(n2273), .Y(n454) );
  NAND21X1 U1332 ( .B(n2139), .A(n488), .Y(n480) );
  INVX1 U1333 ( .A(n908), .Y(n645) );
  OAI222XL U1334 ( .A(n2369), .B(n2274), .C(n612), .D(n2272), .E(n2334), .F(
        n488), .Y(n816) );
  OAI221X1 U1335 ( .A(n2446), .B(n2272), .C(n2274), .D(n2458), .E(n2167), .Y(
        n814) );
  AOI31X1 U1336 ( .A(n2374), .B(n56), .C(n808), .D(n809), .Y(n800) );
  OAI22X1 U1337 ( .A(n2448), .B(n2273), .C(n488), .D(n2459), .Y(n815) );
  OAI21X1 U1338 ( .B(n44), .C(n2343), .A(n2416), .Y(n760) );
  AOI32X1 U1339 ( .A(n1682), .B(n2108), .C(n766), .D(n972), .E(n1780), .Y(
        n2104) );
  NAND2X1 U1340 ( .A(n2372), .B(n1025), .Y(n767) );
  OAI21X1 U1341 ( .B(n1975), .C(n1026), .A(n1015), .Y(n1025) );
  INVX1 U1342 ( .A(pc_i[1]), .Y(n415) );
  INVX1 U1343 ( .A(n2272), .Y(n351) );
  INVX1 U1344 ( .A(n2274), .Y(n356) );
  INVX1 U1345 ( .A(n488), .Y(n357) );
  NOR32XL U1346 ( .B(n697), .C(n2236), .A(n698), .Y(n691) );
  MUX2AXL U1347 ( .D0(n2447), .D1(n1549), .S(n261), .Y(ramsfraddr_comb[4]) );
  NOR3XL U1348 ( .A(n252), .B(n102), .C(n2352), .Y(n692) );
  INVX1 U1349 ( .A(n696), .Y(n2175) );
  AOI221XL U1350 ( .A(n989), .B(n830), .C(memdatai[5]), .D(n990), .E(n997), 
        .Y(n996) );
  OAI22X1 U1351 ( .A(n2278), .B(n2467), .C(n31), .D(n2281), .Y(n997) );
  AOI221XL U1352 ( .A(n989), .B(n829), .C(memdatai[4]), .D(n990), .E(n999), 
        .Y(n998) );
  OAI22X1 U1353 ( .A(n2278), .B(n2468), .C(n27), .D(n2281), .Y(n999) );
  MUX2AXL U1354 ( .D0(n2441), .D1(n1553), .S(n261), .Y(ramsfraddr_comb[6]) );
  NAND21X1 U1355 ( .B(n2435), .A(n210), .Y(n2204) );
  MUX2AXL U1356 ( .D0(n2445), .D1(n1867), .S(n261), .Y(ramsfraddr_comb[5]) );
  MUX2AXL U1357 ( .D0(n2432), .D1(n1572), .S(n261), .Y(ramsfraddr_comb[3]) );
  NAND21X1 U1358 ( .B(n2316), .A(n209), .Y(n2205) );
  NOR2X1 U1359 ( .A(n2318), .B(n2271), .Y(n2148) );
  NOR2X1 U1360 ( .A(n1023), .B(n255), .Y(n1022) );
  NAND2X1 U1361 ( .A(n865), .B(n1234), .Y(n1248) );
  INVX1 U1362 ( .A(n1677), .Y(n1701) );
  INVX1 U1363 ( .A(n1545), .Y(n1518) );
  OAI22XL U1364 ( .A(n270), .B(n1645), .C(n987), .D(n1644), .Y(N12714) );
  AOI221XL U1365 ( .A(n989), .B(n825), .C(n990), .D(memdatai[0]), .E(n1007), 
        .Y(n1645) );
  OAI22X1 U1366 ( .A(n2278), .B(n2470), .C(n2422), .D(n2281), .Y(n1007) );
  OAI22XL U1367 ( .A(n987), .B(n1638), .C(n988), .D(n271), .Y(N12721) );
  AOI221XL U1368 ( .A(n989), .B(n832), .C(memdatai[7]), .D(n990), .E(n991), 
        .Y(n988) );
  OAI22X1 U1369 ( .A(n2278), .B(n2466), .C(n15), .D(n2281), .Y(n991) );
  OAI22XL U1370 ( .A(n270), .B(n1642), .C(n987), .D(n1641), .Y(N12715) );
  AOI221XL U1371 ( .A(n989), .B(n826), .C(n990), .D(memdatai[1]), .E(n1005), 
        .Y(n1642) );
  OAI22X1 U1372 ( .A(n2278), .B(n2469), .C(n2423), .D(n2281), .Y(n1005) );
  INVX1 U1373 ( .A(n54), .Y(n687) );
  NAND3X1 U1374 ( .A(n849), .B(n2212), .C(n211), .Y(n848) );
  NAND21X1 U1375 ( .B(n2256), .A(n209), .Y(n2202) );
  NAND21X1 U1376 ( .B(n2169), .A(n210), .Y(n2203) );
  NAND21X1 U1377 ( .B(n2257), .A(n210), .Y(n2200) );
  NAND21X1 U1378 ( .B(n2415), .A(n210), .Y(n2206) );
  NAND21X1 U1379 ( .B(n2255), .A(n210), .Y(n2201) );
  NAND21X1 U1380 ( .B(n2414), .A(n209), .Y(n2207) );
  NAND21X1 U1381 ( .B(n219), .A(n1353), .Y(n1355) );
  NAND21X1 U1382 ( .B(n596), .A(n211), .Y(n593) );
  NOR3XL U1383 ( .A(n2212), .B(n2306), .C(n1355), .Y(n1360) );
  NOR3XL U1384 ( .A(n2211), .B(n1047), .C(n1355), .Y(n1361) );
  INVX1 U1385 ( .A(n1470), .Y(n1112) );
  NAND43X1 U1386 ( .B(n220), .C(n1451), .D(n1450), .A(n862), .Y(n1470) );
  INVX1 U1387 ( .A(n1114), .Y(n1451) );
  INVX1 U1388 ( .A(n865), .Y(n1450) );
  NAND2X1 U1389 ( .A(n858), .B(n859), .Y(n852) );
  NAND2X1 U1390 ( .A(n858), .B(n862), .Y(n861) );
  INVX1 U1391 ( .A(n1506), .Y(n858) );
  NAND21X1 U1392 ( .B(n13), .A(n211), .Y(n1506) );
  AND2X1 U1393 ( .A(n1673), .B(n1672), .Y(N12912) );
  OAI22X1 U1394 ( .A(n182), .B(n220), .C(n1670), .D(n12), .Y(n1673) );
  OAI22X1 U1395 ( .A(n645), .B(n111), .C(n1235), .D(n133), .Y(N12555) );
  OAI22X1 U1396 ( .A(n645), .B(n75), .C(n1235), .D(n57), .Y(N12519) );
  OAI22X1 U1397 ( .A(n645), .B(n92), .C(n1235), .D(n114), .Y(N12546) );
  OAI22X1 U1398 ( .A(n645), .B(n132), .C(n1235), .D(n94), .Y(N12510) );
  OAI22X1 U1399 ( .A(n645), .B(n90), .C(n1235), .D(n76), .Y(N12537) );
  OAI22X1 U1400 ( .A(n645), .B(n130), .C(n1235), .D(n52), .Y(N12501) );
  OAI22X1 U1401 ( .A(n645), .B(n109), .C(n1235), .D(n64), .Y(N12564) );
  OAI22X1 U1402 ( .A(n645), .B(n73), .C(n1235), .D(n48), .Y(N12528) );
  OAI22X1 U1403 ( .A(n742), .B(n110), .C(n1122), .D(n1124), .Y(N12620) );
  OAI22X1 U1404 ( .A(n737), .B(n110), .C(n1121), .D(n1124), .Y(N12621) );
  OAI22X1 U1405 ( .A(n712), .B(n110), .C(n1118), .D(n1124), .Y(N12626) );
  OAI22X1 U1406 ( .A(n704), .B(n110), .C(n1116), .D(n1124), .Y(N12627) );
  OAI22X1 U1407 ( .A(n684), .B(n111), .C(n1238), .D(n1124), .Y(N12549) );
  OAI22X1 U1408 ( .A(n671), .B(n111), .C(n1237), .D(n133), .Y(N12551) );
  OAI22X1 U1409 ( .A(n742), .B(n74), .C(n1122), .D(n1132), .Y(N12584) );
  OAI22X1 U1410 ( .A(n737), .B(n74), .C(n1121), .D(n1132), .Y(N12585) );
  OAI22X1 U1411 ( .A(n712), .B(n74), .C(n1118), .D(n1132), .Y(N12590) );
  OAI22X1 U1412 ( .A(n704), .B(n74), .C(n1116), .D(n1132), .Y(N12591) );
  OAI22X1 U1413 ( .A(n742), .B(n91), .C(n1122), .D(n1126), .Y(N12611) );
  OAI22X1 U1414 ( .A(n737), .B(n91), .C(n1121), .D(n114), .Y(N12612) );
  OAI22X1 U1415 ( .A(n712), .B(n91), .C(n1118), .D(n1126), .Y(N12617) );
  OAI22X1 U1416 ( .A(n704), .B(n91), .C(n1116), .D(n114), .Y(N12618) );
  OAI22X1 U1417 ( .A(n684), .B(n92), .C(n1238), .D(n1126), .Y(N12540) );
  OAI22X1 U1418 ( .A(n671), .B(n92), .C(n1237), .D(n1126), .Y(N12542) );
  OAI22X1 U1419 ( .A(n742), .B(n131), .C(n1122), .D(n1134), .Y(N12575) );
  OAI22X1 U1420 ( .A(n737), .B(n131), .C(n1121), .D(n1134), .Y(N12576) );
  OAI22X1 U1421 ( .A(n712), .B(n131), .C(n1118), .D(n1134), .Y(N12581) );
  OAI22X1 U1422 ( .A(n704), .B(n131), .C(n1116), .D(n1134), .Y(N12582) );
  OAI22X1 U1423 ( .A(n684), .B(n132), .C(n1238), .D(n1134), .Y(N12504) );
  OAI22X1 U1424 ( .A(n671), .B(n132), .C(n1237), .D(n94), .Y(N12506) );
  OAI22X1 U1425 ( .A(n742), .B(n89), .C(n1122), .D(n1128), .Y(N12602) );
  OAI22X1 U1426 ( .A(n737), .B(n89), .C(n1121), .D(n76), .Y(N12603) );
  OAI22X1 U1427 ( .A(n712), .B(n89), .C(n1118), .D(n1128), .Y(N12608) );
  OAI22X1 U1428 ( .A(n704), .B(n89), .C(n1116), .D(n76), .Y(N12609) );
  OAI22X1 U1429 ( .A(n684), .B(n90), .C(n1238), .D(n1128), .Y(N12531) );
  OAI22X1 U1430 ( .A(n671), .B(n90), .C(n1237), .D(n1128), .Y(N12533) );
  OAI22X1 U1431 ( .A(n742), .B(n129), .C(n1122), .D(n1136), .Y(N12566) );
  OAI22X1 U1432 ( .A(n737), .B(n129), .C(n1121), .D(n1136), .Y(N12567) );
  OAI22X1 U1433 ( .A(n712), .B(n129), .C(n1118), .D(n1136), .Y(N12572) );
  OAI22X1 U1434 ( .A(n704), .B(n129), .C(n1116), .D(n1136), .Y(N12573) );
  OAI22X1 U1435 ( .A(n684), .B(n130), .C(n1238), .D(n1136), .Y(N12495) );
  OAI22X1 U1436 ( .A(n671), .B(n130), .C(n1237), .D(n52), .Y(N12497) );
  OAI22X1 U1437 ( .A(n742), .B(n108), .C(n1122), .D(n1117), .Y(N12629) );
  OAI22X1 U1438 ( .A(n737), .B(n108), .C(n1121), .D(n1117), .Y(N12630) );
  OAI22X1 U1439 ( .A(n712), .B(n108), .C(n1118), .D(n1117), .Y(N12635) );
  OAI22X1 U1440 ( .A(n704), .B(n108), .C(n1116), .D(n1117), .Y(N12636) );
  OAI22X1 U1441 ( .A(n684), .B(n109), .C(n1238), .D(n1117), .Y(N12558) );
  OAI22X1 U1442 ( .A(n671), .B(n109), .C(n1237), .D(n64), .Y(N12560) );
  OAI22X1 U1443 ( .A(n742), .B(n72), .C(n1122), .D(n1130), .Y(N12593) );
  OAI22X1 U1444 ( .A(n737), .B(n72), .C(n1121), .D(n1130), .Y(N12594) );
  OAI22X1 U1445 ( .A(n712), .B(n72), .C(n1118), .D(n1130), .Y(N12599) );
  OAI22X1 U1446 ( .A(n704), .B(n72), .C(n1116), .D(n1130), .Y(N12600) );
  OAI22X1 U1447 ( .A(n699), .B(n75), .C(n2230), .D(n1132), .Y(N12512) );
  OAI22X1 U1448 ( .A(n699), .B(n111), .C(n2230), .D(n133), .Y(N12548) );
  OAI22X1 U1449 ( .A(n732), .B(n110), .C(n1120), .D(n1124), .Y(N12622) );
  OAI22X1 U1450 ( .A(n727), .B(n110), .C(n2223), .D(n1124), .Y(N12623) );
  OAI22X1 U1451 ( .A(n722), .B(n110), .C(n1119), .D(n1124), .Y(N12624) );
  OAI22X1 U1452 ( .A(n717), .B(n110), .C(n2222), .D(n1124), .Y(N12625) );
  OAI22X1 U1453 ( .A(n678), .B(n111), .C(n2228), .D(n133), .Y(N12550) );
  OAI22X1 U1454 ( .A(n660), .B(n111), .C(n2226), .D(n133), .Y(N12552) );
  OAI22X1 U1455 ( .A(n655), .B(n111), .C(n2224), .D(n133), .Y(N12553) );
  OAI22X1 U1456 ( .A(n650), .B(n111), .C(n1236), .D(n133), .Y(N12554) );
  OAI22X1 U1457 ( .A(n732), .B(n74), .C(n1120), .D(n1132), .Y(N12586) );
  OAI22X1 U1458 ( .A(n722), .B(n74), .C(n1119), .D(n1132), .Y(N12588) );
  OAI22X1 U1459 ( .A(n717), .B(n74), .C(n2222), .D(n1132), .Y(N12589) );
  OAI22X1 U1460 ( .A(n684), .B(n75), .C(n1238), .D(n57), .Y(N12513) );
  OAI22X1 U1461 ( .A(n678), .B(n75), .C(n2228), .D(n57), .Y(N12514) );
  OAI22X1 U1462 ( .A(n671), .B(n75), .C(n1237), .D(n57), .Y(N12515) );
  OAI22X1 U1463 ( .A(n660), .B(n75), .C(n2226), .D(n57), .Y(N12516) );
  OAI22X1 U1464 ( .A(n655), .B(n75), .C(n2224), .D(n57), .Y(N12517) );
  OAI22X1 U1465 ( .A(n650), .B(n75), .C(n1236), .D(n57), .Y(N12518) );
  OAI22X1 U1466 ( .A(n699), .B(n132), .C(n2230), .D(n94), .Y(N12503) );
  OAI22X1 U1467 ( .A(n699), .B(n92), .C(n2230), .D(n114), .Y(N12539) );
  OAI22X1 U1468 ( .A(n732), .B(n91), .C(n1120), .D(n1126), .Y(N12613) );
  OAI22X1 U1469 ( .A(n727), .B(n91), .C(n2223), .D(n114), .Y(N12614) );
  OAI22X1 U1470 ( .A(n722), .B(n91), .C(n1119), .D(n1126), .Y(N12615) );
  OAI22X1 U1471 ( .A(n717), .B(n91), .C(n2222), .D(n114), .Y(N12616) );
  OAI22X1 U1472 ( .A(n678), .B(n92), .C(n2228), .D(n1126), .Y(N12541) );
  OAI22X1 U1473 ( .A(n660), .B(n92), .C(n2226), .D(n1126), .Y(N12543) );
  OAI22X1 U1474 ( .A(n655), .B(n92), .C(n2224), .D(n114), .Y(N12544) );
  OAI22X1 U1475 ( .A(n650), .B(n92), .C(n1236), .D(n114), .Y(N12545) );
  OAI22X1 U1476 ( .A(n732), .B(n131), .C(n1120), .D(n1134), .Y(N12577) );
  OAI22X1 U1477 ( .A(n727), .B(n131), .C(n2223), .D(n1134), .Y(N12578) );
  OAI22X1 U1478 ( .A(n722), .B(n131), .C(n1119), .D(n1134), .Y(N12579) );
  OAI22X1 U1479 ( .A(n717), .B(n131), .C(n2222), .D(n1134), .Y(N12580) );
  OAI22X1 U1480 ( .A(n678), .B(n132), .C(n2228), .D(n94), .Y(N12505) );
  OAI22X1 U1481 ( .A(n660), .B(n132), .C(n2226), .D(n94), .Y(N12507) );
  OAI22X1 U1482 ( .A(n655), .B(n132), .C(n2224), .D(n94), .Y(N12508) );
  OAI22X1 U1483 ( .A(n650), .B(n132), .C(n1236), .D(n94), .Y(N12509) );
  OAI22X1 U1484 ( .A(n699), .B(n130), .C(n2230), .D(n52), .Y(N12494) );
  OAI22X1 U1485 ( .A(n699), .B(n90), .C(n2230), .D(n76), .Y(N12530) );
  OAI22X1 U1486 ( .A(n732), .B(n89), .C(n1120), .D(n1128), .Y(N12604) );
  OAI22X1 U1487 ( .A(n727), .B(n89), .C(n2223), .D(n76), .Y(N12605) );
  OAI22X1 U1488 ( .A(n722), .B(n89), .C(n1119), .D(n1128), .Y(N12606) );
  OAI22X1 U1489 ( .A(n717), .B(n89), .C(n2222), .D(n76), .Y(N12607) );
  OAI22X1 U1490 ( .A(n678), .B(n90), .C(n2228), .D(n1128), .Y(N12532) );
  OAI22X1 U1491 ( .A(n660), .B(n90), .C(n2226), .D(n1128), .Y(N12534) );
  OAI22X1 U1492 ( .A(n655), .B(n90), .C(n2224), .D(n76), .Y(N12535) );
  OAI22X1 U1493 ( .A(n650), .B(n90), .C(n1236), .D(n76), .Y(N12536) );
  OAI22X1 U1494 ( .A(n732), .B(n129), .C(n1120), .D(n1136), .Y(N12568) );
  OAI22X1 U1495 ( .A(n722), .B(n129), .C(n1119), .D(n1136), .Y(N12570) );
  OAI22X1 U1496 ( .A(n717), .B(n129), .C(n2222), .D(n1136), .Y(N12571) );
  OAI22X1 U1497 ( .A(n678), .B(n130), .C(n2228), .D(n52), .Y(N12496) );
  OAI22X1 U1498 ( .A(n660), .B(n130), .C(n2226), .D(n52), .Y(N12498) );
  OAI22X1 U1499 ( .A(n655), .B(n130), .C(n2224), .D(n52), .Y(N12499) );
  OAI22X1 U1500 ( .A(n650), .B(n130), .C(n1236), .D(n52), .Y(N12500) );
  OAI22X1 U1501 ( .A(n699), .B(n73), .C(n2230), .D(n1130), .Y(N12521) );
  OAI22X1 U1502 ( .A(n699), .B(n109), .C(n2230), .D(n64), .Y(N12557) );
  OAI22X1 U1503 ( .A(n732), .B(n108), .C(n1120), .D(n1117), .Y(N12631) );
  OAI22X1 U1504 ( .A(n727), .B(n108), .C(n2223), .D(n1117), .Y(N12632) );
  OAI22X1 U1505 ( .A(n722), .B(n108), .C(n1119), .D(n1117), .Y(N12633) );
  OAI22X1 U1506 ( .A(n717), .B(n108), .C(n2222), .D(n1117), .Y(N12634) );
  OAI22X1 U1507 ( .A(n678), .B(n109), .C(n2228), .D(n64), .Y(N12559) );
  OAI22X1 U1508 ( .A(n660), .B(n109), .C(n2226), .D(n64), .Y(N12561) );
  OAI22X1 U1509 ( .A(n655), .B(n109), .C(n2224), .D(n64), .Y(N12562) );
  OAI22X1 U1510 ( .A(n650), .B(n109), .C(n1236), .D(n64), .Y(N12563) );
  OAI22X1 U1511 ( .A(n732), .B(n72), .C(n1120), .D(n1130), .Y(N12595) );
  OAI22X1 U1512 ( .A(n722), .B(n72), .C(n1119), .D(n1130), .Y(N12597) );
  OAI22X1 U1513 ( .A(n717), .B(n72), .C(n2222), .D(n1130), .Y(N12598) );
  OAI22X1 U1514 ( .A(n684), .B(n73), .C(n1238), .D(n48), .Y(N12522) );
  OAI22X1 U1515 ( .A(n678), .B(n73), .C(n2228), .D(n48), .Y(N12523) );
  OAI22X1 U1516 ( .A(n671), .B(n73), .C(n1237), .D(n48), .Y(N12524) );
  OAI22X1 U1517 ( .A(n660), .B(n73), .C(n2226), .D(n48), .Y(N12525) );
  OAI22X1 U1518 ( .A(n655), .B(n73), .C(n2224), .D(n48), .Y(N12526) );
  OAI22X1 U1519 ( .A(n650), .B(n73), .C(n1236), .D(n48), .Y(N12527) );
  OAI22X1 U1520 ( .A(n727), .B(n74), .C(n2223), .D(n1132), .Y(N12587) );
  OAI22X1 U1521 ( .A(n727), .B(n129), .C(n2223), .D(n1136), .Y(N12569) );
  OAI22X1 U1522 ( .A(n727), .B(n72), .C(n2223), .D(n1130), .Y(N12596) );
  OAI22X1 U1523 ( .A(n955), .B(n221), .C(n918), .D(n2194), .Y(N12723) );
  NOR3XL U1524 ( .A(n956), .B(n957), .C(n958), .Y(n955) );
  OAI211X1 U1525 ( .C(n33), .D(n947), .A(n953), .B(n963), .Y(n956) );
  OAI22X1 U1526 ( .A(n2470), .B(n2344), .C(n959), .D(n2323), .Y(n958) );
  OAI22X1 U1527 ( .A(n948), .B(n216), .C(n918), .D(n2196), .Y(N12724) );
  NOR3XL U1528 ( .A(n949), .B(n950), .C(n951), .Y(n948) );
  OAI211X1 U1529 ( .C(n2437), .D(n947), .A(n953), .B(n954), .Y(n949) );
  OAI22X1 U1530 ( .A(n2469), .B(n2344), .C(n952), .D(n2323), .Y(n951) );
  OAI22X1 U1531 ( .A(n270), .B(n483), .C(n484), .D(n2204), .Y(n1884) );
  OAI22AX1 U1532 ( .D(n1650), .C(n219), .A(n1651), .B(n1670), .Y(N11487) );
  OAI21X1 U1533 ( .B(n857), .C(n861), .A(n267), .Y(N13086) );
  OAI21X1 U1534 ( .B(n856), .C(n861), .A(n267), .Y(N13095) );
  OAI21X1 U1535 ( .B(n855), .C(n861), .A(n267), .Y(N13104) );
  OAI21X1 U1536 ( .B(n854), .C(n861), .A(n267), .Y(N13113) );
  OAI21X1 U1537 ( .B(n853), .C(n861), .A(n266), .Y(N13140) );
  OAI21X1 U1538 ( .B(n857), .C(n852), .A(n266), .Y(N13230) );
  OAI21X1 U1539 ( .B(n856), .C(n852), .A(n265), .Y(N13239) );
  OAI21X1 U1540 ( .B(n852), .C(n855), .A(n266), .Y(N13248) );
  OAI21X1 U1541 ( .B(n852), .C(n854), .A(n265), .Y(N13257) );
  OAI21X1 U1542 ( .B(n853), .C(n852), .A(n265), .Y(N13284) );
  OAI21X1 U1543 ( .B(n857), .C(n863), .A(n268), .Y(N13014) );
  OAI21X1 U1544 ( .B(n856), .C(n863), .A(n268), .Y(N13023) );
  OAI21X1 U1545 ( .B(n855), .C(n863), .A(n267), .Y(N13032) );
  OAI21X1 U1546 ( .B(n854), .C(n863), .A(n268), .Y(N13041) );
  OAI21X1 U1547 ( .B(n1450), .C(n863), .A(n267), .Y(N13050) );
  OAI21X1 U1548 ( .B(n2439), .C(n863), .A(n267), .Y(N13059) );
  OAI21X1 U1549 ( .B(n853), .C(n863), .A(n267), .Y(N13068) );
  OAI21X1 U1550 ( .B(n851), .C(n863), .A(n267), .Y(N13077) );
  OAI21X1 U1551 ( .B(n857), .C(n860), .A(n266), .Y(N13158) );
  OAI21X1 U1552 ( .B(n856), .C(n860), .A(n266), .Y(N13167) );
  OAI21X1 U1553 ( .B(n855), .C(n860), .A(n266), .Y(N13176) );
  OAI21X1 U1554 ( .B(n854), .C(n860), .A(n265), .Y(N13185) );
  OAI21X1 U1555 ( .B(n1450), .C(n860), .A(n266), .Y(N13194) );
  OAI21X1 U1556 ( .B(n2439), .C(n860), .A(n265), .Y(N13203) );
  OAI21X1 U1557 ( .B(n853), .C(n860), .A(n266), .Y(N13212) );
  OAI21X1 U1558 ( .B(n851), .C(n860), .A(n265), .Y(N13221) );
  OAI21X1 U1559 ( .B(n1110), .C(n1113), .A(n268), .Y(N12644) );
  OAI21X1 U1560 ( .B(n1109), .C(n1113), .A(n268), .Y(N12651) );
  OAI21X1 U1561 ( .B(n1107), .C(n1113), .A(n268), .Y(N12658) );
  OAI21X1 U1562 ( .B(n1111), .C(n1108), .A(n268), .Y(N12665) );
  OAI21X1 U1563 ( .B(n1110), .C(n1108), .A(n268), .Y(N12672) );
  OAI21X1 U1564 ( .B(n1109), .C(n1108), .A(n268), .Y(N12679) );
  OAI21X1 U1565 ( .B(n1107), .C(n1108), .A(n268), .Y(N12686) );
  ENOX1 U1566 ( .A(n1027), .B(n2200), .C(n820), .D(n1028), .Y(N12705) );
  ENOX1 U1567 ( .A(n1027), .B(n2205), .C(n1028), .D(n1029), .Y(N12711) );
  NAND3X1 U1568 ( .A(n1030), .B(n1031), .C(n1032), .Y(n1029) );
  NAND4X1 U1569 ( .A(n2462), .B(n2461), .C(n1045), .D(n1046), .Y(n1030) );
  OAI21X1 U1570 ( .B(n1042), .C(n1043), .A(n1044), .Y(n1031) );
  NAND2X1 U1571 ( .A(n1112), .B(n127), .Y(n1113) );
  NAND32X1 U1572 ( .B(n220), .C(finishdiv), .A(n1511), .Y(n841) );
  INVX1 U1573 ( .A(n1510), .Y(n1511) );
  NAND32X1 U1574 ( .B(n1518), .C(n221), .A(n596), .Y(n595) );
  NOR21XL U1575 ( .B(n215), .A(n2069), .Y(N10569) );
  AOI211X1 U1576 ( .C(n1690), .D(n1754), .A(n809), .B(n805), .Y(n2069) );
  NAND21X1 U1577 ( .B(n219), .A(n54), .Y(n2055) );
  NAND21X1 U1578 ( .B(n219), .A(n1102), .Y(n1092) );
  AO21X1 U1579 ( .B(n215), .C(n284), .A(n272), .Y(N11491) );
  INVX1 U1580 ( .A(n1755), .Y(n284) );
  OR2X1 U1581 ( .A(n270), .B(n179), .Y(N13366) );
  AOI21X1 U1582 ( .B(n2211), .C(n1510), .A(n219), .Y(n179) );
  AND3X1 U1583 ( .A(n212), .B(n2011), .C(n1596), .Y(N585) );
  NOR32XL U1584 ( .B(n212), .C(n2157), .A(n2056), .Y(N10584) );
  AND3X1 U1585 ( .A(n1975), .B(n1014), .C(n214), .Y(N10586) );
  OAI22AX1 U1586 ( .D(dpc[3]), .C(n1091), .A(n1101), .B(n1092), .Y(N12693) );
  OAI22AX1 U1587 ( .D(dpc[4]), .C(n1091), .A(n2391), .B(n1092), .Y(N12694) );
  OAI22AX1 U1588 ( .D(dpc[5]), .C(n1091), .A(n2298), .B(n1092), .Y(N12695) );
  AND2X1 U1589 ( .A(n1767), .B(n620), .Y(N371) );
  AND2X1 U1590 ( .A(n1757), .B(n620), .Y(N372) );
  OAI21X1 U1591 ( .B(n983), .C(n219), .A(n274), .Y(N12722) );
  NOR3XL U1592 ( .A(n984), .B(n2319), .C(n985), .Y(n983) );
  OAI21X1 U1593 ( .B(n986), .C(n2324), .A(n953), .Y(n984) );
  AND2X1 U1594 ( .A(n1736), .B(n1627), .Y(N11488) );
  AND2X1 U1595 ( .A(n224), .B(n1674), .Y(N11486) );
  AOI22X1 U1596 ( .A(n1386), .B(n832), .C(ramdatai[7]), .D(n1387), .Y(n1382)
         );
  AOI22X1 U1597 ( .A(n831), .B(n1386), .C(ramdatai[6]), .D(n1387), .Y(n1435)
         );
  AOI22X1 U1598 ( .A(n830), .B(n1386), .C(ramdatai[5]), .D(n1387), .Y(n1469)
         );
  INVX1 U1599 ( .A(n1512), .Y(n1767) );
  NAND32X1 U1600 ( .B(n152), .C(n220), .A(n749), .Y(n1512) );
  NOR3XL U1601 ( .A(n2055), .B(n2377), .C(n2356), .Y(N10588) );
  NOR3XL U1602 ( .A(n2055), .B(n2356), .C(n2380), .Y(N10587) );
  INVX1 U1603 ( .A(n941), .Y(n1950) );
  INVX1 U1604 ( .A(n1514), .Y(n1756) );
  NAND21X1 U1605 ( .B(n2011), .A(n211), .Y(n1514) );
  NOR2X1 U1606 ( .A(n847), .B(n841), .Y(N13367) );
  NOR2X1 U1607 ( .A(n2275), .B(n595), .Y(N682) );
  NOR2X1 U1608 ( .A(n2166), .B(n595), .Y(N683) );
  NOR2X1 U1609 ( .A(n2165), .B(n595), .Y(N684) );
  NOR2X1 U1610 ( .A(n911), .B(n2067), .Y(N10567) );
  NAND2X1 U1611 ( .A(n264), .B(n875), .Y(n873) );
  AO21X1 U1612 ( .B(n1480), .C(n1479), .A(n1477), .Y(n875) );
  INVX1 U1613 ( .A(n620), .Y(n1672) );
  OAI211X1 U1614 ( .C(n2166), .D(n666), .A(n665), .B(n664), .Y(n1600) );
  INVX1 U1615 ( .A(n662), .Y(n666) );
  OA222X1 U1616 ( .A(n256), .B(n688), .C(n2275), .D(n164), .E(n253), .F(n663), 
        .Y(n664) );
  AND2X1 U1617 ( .A(n596), .B(n1672), .Y(n665) );
  NOR2X1 U1618 ( .A(n105), .B(n2185), .Y(retiinstr) );
  AOI21BBXL U1619 ( .B(cpu_resume), .C(irq), .A(n269), .Y(N13379) );
  NOR2X1 U1620 ( .A(n874), .B(n873), .Y(N12975) );
  XNOR2XL U1621 ( .A(n2329), .B(n2328), .Y(n874) );
  AND3X1 U1622 ( .A(mempsack), .B(n280), .C(n279), .Y(n282) );
  INVX1 U1623 ( .A(n1480), .Y(n283) );
  OAI22X1 U1624 ( .A(n2261), .B(n942), .C(n2268), .D(n2282), .Y(n957) );
  INVX1 U1625 ( .A(n829), .Y(n453) );
  AOI22X1 U1626 ( .A(n184), .B(N13353), .C(N13347), .D(n2190), .Y(n845) );
  AOI22X1 U1627 ( .A(n2135), .B(N13353), .C(N13346), .D(n2190), .Y(n846) );
  AOI22X1 U1628 ( .A(n185), .B(N13353), .C(N13348), .D(n2190), .Y(n844) );
  AOI22X1 U1629 ( .A(n186), .B(N13353), .C(N13349), .D(n2190), .Y(n843) );
  AOI22X1 U1630 ( .A(n188), .B(N13353), .C(N13351), .D(n2190), .Y(n840) );
  AOI22X1 U1631 ( .A(n187), .B(N13353), .C(N13350), .D(n2190), .Y(n842) );
  INVX1 U1632 ( .A(n690), .Y(n1434) );
  OAI22X1 U1633 ( .A(n1541), .B(n2285), .C(n2259), .D(n1542), .Y(n1538) );
  INVX1 U1634 ( .A(pc_i[11]), .Y(n2285) );
  INVX1 U1635 ( .A(n1352), .Y(n750) );
  NAND2X1 U1636 ( .A(n1521), .B(n1518), .Y(n1519) );
  NOR32XL U1637 ( .B(n1384), .C(n1950), .A(n2446), .Y(n1385) );
  OAI22X1 U1638 ( .A(n941), .B(n2323), .C(n2195), .D(n918), .Y(n940) );
  INVX1 U1639 ( .A(n827), .Y(n437) );
  OR2X1 U1640 ( .A(n2074), .B(n451), .Y(n624) );
  INVX1 U1641 ( .A(pc_i[13]), .Y(n494) );
  NAND32X1 U1642 ( .B(n1412), .C(n613), .A(n183), .Y(n615) );
  INVX1 U1643 ( .A(n1398), .Y(n613) );
  ENOX1 U1644 ( .A(n2140), .B(n2012), .C(n2012), .D(n2138), .Y(n1412) );
  OAI21X1 U1645 ( .B(n2074), .C(n1507), .A(n1508), .Y(n1387) );
  MUX2X1 U1646 ( .D0(n612), .D1(n2271), .S(n1150), .Y(n2012) );
  NAND21X1 U1647 ( .B(n2139), .A(n2272), .Y(n1398) );
  NAND3X1 U1648 ( .A(dpc[1]), .B(n2248), .C(n2233), .Y(n1146) );
  NAND3X1 U1649 ( .A(dpc[1]), .B(dpc[2]), .C(n2233), .Y(n1144) );
  NAND2X1 U1650 ( .A(n2177), .B(dpc[0]), .Y(n1182) );
  AOI221XL U1651 ( .A(n1147), .B(n2231), .C(n1302), .D(n1138), .E(n1182), .Y(
        n1312) );
  AOI221XL U1652 ( .A(n2288), .B(n2231), .C(n1281), .D(n1138), .E(n1182), .Y(
        n1290) );
  INVX1 U1653 ( .A(n1102), .Y(n2177) );
  NOR2X1 U1654 ( .A(n128), .B(n2442), .Y(N14351) );
  NOR2X1 U1655 ( .A(n2459), .B(n2465), .Y(N14346) );
  NOR2X1 U1656 ( .A(n128), .B(n2462), .Y(N14347) );
  NOR2X1 U1657 ( .A(n128), .B(n2461), .Y(N14348) );
  NOR2X1 U1658 ( .A(n128), .B(n2456), .Y(N14349) );
  NOR2X1 U1659 ( .A(n128), .B(n2457), .Y(N14350) );
  NOR2X1 U1660 ( .A(n2459), .B(n2463), .Y(N14345) );
  NAND21X1 U1661 ( .B(n2139), .A(n2274), .Y(n509) );
  OAI21X1 U1662 ( .B(n33), .C(n1146), .A(n2233), .Y(n1212) );
  INVX1 U1663 ( .A(n1903), .Y(n1389) );
  OAI211X1 U1664 ( .C(n1243), .D(n2235), .A(n2233), .B(n1255), .Y(n1245) );
  AOI21X1 U1665 ( .B(n2231), .C(n1256), .A(n1257), .Y(n1255) );
  AOI21X1 U1666 ( .B(n2291), .C(n31), .A(n1146), .Y(n1257) );
  OAI21X1 U1667 ( .B(n1203), .C(n1144), .A(n1192), .Y(n1202) );
  AOI22AXL U1668 ( .A(n1517), .B(n1452), .D(n1517), .C(n2138), .Y(n1520) );
  AOI22AXL U1669 ( .A(n1478), .B(n1452), .D(n1478), .C(n2138), .Y(n1481) );
  AOI211X1 U1670 ( .C(n1138), .D(n38), .A(n1245), .B(n1246), .Y(n1241) );
  AOI21X1 U1671 ( .B(n1144), .C(n62), .A(n38), .Y(n1246) );
  AOI211X1 U1672 ( .C(n1138), .D(n27), .A(n1270), .B(n2225), .Y(n1264) );
  OAI22X1 U1673 ( .A(n27), .B(n45), .C(n2291), .D(n62), .Y(n1270) );
  INVX1 U1674 ( .A(n1271), .Y(n2225) );
  NOR3XL U1675 ( .A(dpc[1]), .B(dpc[2]), .C(n1182), .Y(n1139) );
  OA21X1 U1676 ( .B(n1227), .C(n33), .A(n1228), .Y(n1122) );
  OAI21X1 U1677 ( .B(n55), .C(n93), .A(n33), .Y(n1228) );
  NOR21XL U1678 ( .B(n1221), .A(n1182), .Y(n1227) );
  MUX2X1 U1679 ( .D0(n507), .D1(n2140), .S(n191), .Y(n434) );
  NOR42XL U1680 ( .C(n1364), .D(n1071), .A(n2178), .B(n1055), .Y(n1039) );
  INVX1 U1681 ( .A(pc_i[4]), .Y(n450) );
  INVX1 U1682 ( .A(pc_i[5]), .Y(n493) );
  INVX1 U1683 ( .A(n1603), .Y(cs_run) );
  NOR2X1 U1684 ( .A(n36), .B(n1214), .Y(n1442) );
  OAI22X1 U1685 ( .A(n2260), .B(n942), .C(n2269), .D(n2282), .Y(n950) );
  OAI21X1 U1686 ( .B(n1301), .C(n62), .A(n1290), .Y(n1299) );
  XNOR2XL U1687 ( .A(n40), .B(n1403), .Y(n1137) );
  NOR2X1 U1688 ( .A(n1323), .B(n35), .Y(n1403) );
  XNOR2XL U1689 ( .A(n2371), .B(n1442), .Y(n1189) );
  XNOR2XL U1690 ( .A(n1214), .B(n36), .Y(n1199) );
  AND2X1 U1691 ( .A(n1145), .B(n40), .Y(n1142) );
  AND2X1 U1692 ( .A(n1168), .B(n35), .Y(n1143) );
  NAND2X1 U1693 ( .A(n1143), .B(n40), .Y(n1147) );
  NAND2X1 U1694 ( .A(n1203), .B(n33), .Y(n1204) );
  NAND2X1 U1695 ( .A(n1301), .B(n42), .Y(n1292) );
  NAND2X1 U1696 ( .A(n1142), .B(n2422), .Y(n1314) );
  AND2X1 U1697 ( .A(n1191), .B(n2371), .Y(n1181) );
  AND2X1 U1698 ( .A(n1203), .B(n36), .Y(n1191) );
  AND2X1 U1699 ( .A(n1181), .B(n29), .Y(n1168) );
  NAND2X1 U1700 ( .A(n1280), .B(n27), .Y(n1267) );
  NAND3X1 U1701 ( .A(n1039), .B(n1362), .C(n1363), .Y(n1356) );
  AOI221XL U1702 ( .A(n1044), .B(n2212), .C(n2179), .D(n2211), .E(n1037), .Y(
        n1363) );
  NAND3X1 U1703 ( .A(n27), .B(n31), .C(n1268), .Y(n1256) );
  INVX1 U1704 ( .A(n1303), .Y(n2288) );
  INVX1 U1705 ( .A(n1179), .Y(n2370) );
  XNOR2XL U1706 ( .A(n2420), .B(n2437), .Y(n1211) );
  NOR3XL U1707 ( .A(n42), .B(n2418), .C(n1281), .Y(n1269) );
  NOR2X1 U1708 ( .A(n985), .B(n961), .Y(n993) );
  NOR3XL U1709 ( .A(n27), .B(n31), .C(n2292), .Y(n1243) );
  INVX1 U1710 ( .A(n990), .Y(n2279) );
  AOI21X1 U1711 ( .B(n2164), .C(n2163), .A(n2010), .Y(n478) );
  NOR2X1 U1712 ( .A(n990), .B(n1016), .Y(n1008) );
  INVX1 U1713 ( .A(n989), .Y(n2280) );
  INVX1 U1714 ( .A(n994), .Y(n2278) );
  INVX1 U1715 ( .A(n1268), .Y(n2287) );
  INVX1 U1716 ( .A(dpc[2]), .Y(n2248) );
  NOR32XL U1717 ( .B(n960), .C(n961), .A(n962), .Y(n921) );
  NOR43XL U1718 ( .B(n960), .C(n962), .D(n961), .A(n919), .Y(n920) );
  AND3X1 U1719 ( .A(n942), .B(n966), .C(n953), .Y(n960) );
  AND3X1 U1720 ( .A(n918), .B(n2344), .C(n2323), .Y(n966) );
  NAND3X1 U1721 ( .A(n606), .B(n607), .C(n608), .Y(n495) );
  OAI21X1 U1722 ( .B(n105), .C(n2388), .A(n610), .Y(n606) );
  OAI22X1 U1723 ( .A(n2253), .B(n257), .C(n253), .D(n609), .Y(n607) );
  NAND2X1 U1724 ( .A(n698), .B(n105), .Y(n918) );
  AOI22X1 U1725 ( .A(n978), .B(n979), .C(n980), .D(n758), .Y(n977) );
  AOI22X1 U1726 ( .A(n978), .B(n2388), .C(n982), .D(n152), .Y(n975) );
  AOI21X1 U1727 ( .B(n758), .C(n776), .A(n972), .Y(n971) );
  INVX1 U1728 ( .A(n961), .Y(n2319) );
  INVX1 U1729 ( .A(n942), .Y(n2326) );
  INVX1 U1730 ( .A(n1010), .Y(n2353) );
  NOR2X1 U1731 ( .A(n696), .B(n105), .Y(n919) );
  OAI221X1 U1732 ( .A(n2404), .B(n911), .C(n2128), .D(n2068), .E(n2129), .Y(
        n2125) );
  OAI21X1 U1733 ( .B(n2071), .C(n1681), .A(n765), .Y(n2129) );
  NOR3XL U1734 ( .A(n2343), .B(n56), .C(n810), .Y(n2058) );
  AOI21X1 U1735 ( .B(n54), .C(n1683), .A(n2071), .Y(n2127) );
  NOR2X1 U1736 ( .A(n2187), .B(n2053), .Y(n2068) );
  NAND4X1 U1737 ( .A(n786), .B(n2059), .C(n2123), .D(n2124), .Y(n2083) );
  AOI222XL U1738 ( .A(n766), .B(n2405), .C(n1690), .D(n1754), .E(n972), .F(
        n2130), .Y(n2123) );
  NOR4XL U1739 ( .A(n2125), .B(n2126), .C(n2064), .D(n2058), .Y(n2124) );
  AOI21X1 U1740 ( .B(n2373), .C(n2378), .A(n2127), .Y(n2126) );
  NAND2X1 U1741 ( .A(n880), .B(n264), .Y(n879) );
  OAI22X1 U1742 ( .A(n2255), .B(n879), .C(n2398), .D(n878), .Y(N12971) );
  OAI22X1 U1743 ( .A(n2316), .B(n879), .C(n2330), .D(n878), .Y(N12967) );
  INVX1 U1744 ( .A(n1353), .Y(n2429) );
  INVX1 U1745 ( .A(n911), .Y(n1653) );
  INVX1 U1746 ( .A(n864), .Y(n2439) );
  MUX2AXL U1747 ( .D0(n2331), .D1(n647), .S(n260), .Y(mempswr_comb) );
  AND2X1 U1748 ( .A(n2011), .B(n1596), .Y(n644) );
  AND2X1 U1749 ( .A(n1627), .B(n1651), .Y(sfroe_comb_s) );
  NAND4X1 U1750 ( .A(n539), .B(n540), .C(n541), .D(n542), .Y(dpl[2]) );
  AOI22X1 U1751 ( .A(n198), .B(dpl_reg[42]), .C(n200), .D(dpl_reg[58]), .Y(
        n539) );
  NAND4X1 U1752 ( .A(n535), .B(n536), .C(n537), .D(n538), .Y(dpl[3]) );
  AOI22X1 U1753 ( .A(n521), .B(dpl_reg[43]), .C(n522), .D(dpl_reg[59]), .Y(
        n535) );
  INVX1 U1754 ( .A(n2273), .Y(n352) );
  OAI21AX1 U1755 ( .B(sfrwe_r), .C(sfroe_r), .A(sfrack), .Y(n279) );
  AO21X1 U1756 ( .B(n2159), .C(temp2_comb[1]), .A(n414), .Y(n428) );
  OAI22X1 U1757 ( .A(n934), .B(n415), .C(n2423), .D(n2311), .Y(n427) );
  NOR32XL U1758 ( .B(n653), .C(n2163), .A(n652), .Y(n1699) );
  AND2X1 U1759 ( .A(cpu_hold), .B(n620), .Y(n652) );
  MUX2IX1 U1760 ( .D0(idle), .D1(n10), .S(n1661), .Y(n653) );
  NOR32XL U1761 ( .B(n395), .C(n394), .A(n393), .Y(n396) );
  NAND2X1 U1762 ( .A(n388), .B(pc_o[0]), .Y(n394) );
  AO2222XL U1763 ( .A(n392), .B(pc_i[0]), .C(memaddr[8]), .D(n391), .E(n2159), 
        .F(temp2_comb[0]), .G(n390), .H(n825), .Y(n393) );
  NAND32XL U1764 ( .B(n1410), .C(n156), .A(n387), .Y(n395) );
  NAND4X1 U1765 ( .A(n531), .B(n532), .C(n533), .D(n534), .Y(dpl[4]) );
  NAND4X1 U1766 ( .A(n563), .B(n564), .C(n565), .D(n566), .Y(dph[4]) );
  AOI22X1 U1767 ( .A(n197), .B(dpl_reg[44]), .C(n199), .D(dpl_reg[60]), .Y(
        n531) );
  NAND4X1 U1768 ( .A(n527), .B(n528), .C(n529), .D(n530), .Y(dpl[5]) );
  NAND4X1 U1769 ( .A(n559), .B(n560), .C(n561), .D(n562), .Y(dph[5]) );
  AOI22X1 U1770 ( .A(n198), .B(dpl_reg[45]), .C(n200), .D(dpl_reg[61]), .Y(
        n527) );
  NOR32XL U1771 ( .B(n1384), .C(acc[1]), .A(n952), .Y(n417) );
  NOR32XL U1772 ( .B(n69), .C(n1384), .A(n959), .Y(n379) );
  NAND21X1 U1773 ( .B(n375), .A(n374), .Y(n376) );
  NAND4X1 U1774 ( .A(n523), .B(n524), .C(n525), .D(n526), .Y(dpl[6]) );
  NAND4X1 U1775 ( .A(n555), .B(n556), .C(n557), .D(n558), .Y(dph[6]) );
  NAND4X1 U1776 ( .A(n551), .B(n552), .C(n553), .D(n554), .Y(dph[7]) );
  AOI22X1 U1777 ( .A(n198), .B(dph_reg[47]), .C(n200), .D(dph_reg[63]), .Y(
        n551) );
  NAND4X1 U1778 ( .A(n571), .B(n572), .C(n573), .D(n574), .Y(dph[2]) );
  AOI22X1 U1779 ( .A(n521), .B(dph_reg[42]), .C(n522), .D(dph_reg[58]), .Y(
        n571) );
  NAND4X1 U1780 ( .A(n567), .B(n568), .C(n569), .D(n570), .Y(dph[3]) );
  AOI22X1 U1781 ( .A(n197), .B(dph_reg[43]), .C(n199), .D(dph_reg[59]), .Y(
        n567) );
  AOI22X1 U1782 ( .A(n53), .B(dph_reg[11]), .C(n49), .D(dph_reg[27]), .Y(n569)
         );
  NAND4X1 U1783 ( .A(n579), .B(n580), .C(n581), .D(n582), .Y(dph[0]) );
  NAND4X1 U1784 ( .A(n547), .B(n548), .C(n549), .D(n550), .Y(dpl[0]) );
  AOI22X1 U1785 ( .A(n197), .B(dph_reg[40]), .C(n199), .D(dph_reg[56]), .Y(
        n579) );
  NAND4X1 U1786 ( .A(n575), .B(n576), .C(n577), .D(n578), .Y(dph[1]) );
  AOI22X1 U1787 ( .A(n198), .B(dph_reg[41]), .C(n200), .D(dph_reg[57]), .Y(
        n575) );
  AOI22X1 U1788 ( .A(n202), .B(dph_reg[33]), .C(n204), .D(dph_reg[49]), .Y(
        n576) );
  NAND4X1 U1789 ( .A(n543), .B(n544), .C(n545), .D(n546), .Y(dpl[1]) );
  AOI22X1 U1790 ( .A(n197), .B(dpl_reg[41]), .C(n199), .D(dpl_reg[57]), .Y(
        n543) );
  MUX2XL U1791 ( .D0(pc_o[7]), .D1(n1574), .S(n155), .Y(memaddr_comb[7]) );
  MUX2XL U1792 ( .D0(pc_o[9]), .D1(n1576), .S(n87), .Y(memaddr_comb[9]) );
  MUX2X1 U1793 ( .D0(pc_o[11]), .D1(n1581), .S(n260), .Y(memaddr_comb[11]) );
  MUX2XL U1794 ( .D0(pc_o[8]), .D1(n1578), .S(n155), .Y(memaddr_comb[8]) );
  AO2222XL U1795 ( .A(alu_out[12]), .B(n101), .C(n899), .D(n196), .E(pc_i[12]), 
        .F(n168), .G(n670), .H(temp[4]), .Y(n903) );
  AO2222XL U1796 ( .A(alu_out[11]), .B(n101), .C(n871), .D(n195), .E(pc_i[11]), 
        .F(n168), .G(n670), .H(temp[3]), .Y(n898) );
  MUX2X1 U1797 ( .D0(pc_o[12]), .D1(n1580), .S(n260), .Y(memaddr_comb[12]) );
  MUX2BXL U1798 ( .D0(ramwe), .D1(n180), .S(n262), .Y(ramwe_comb) );
  AOI21X1 U1799 ( .B(n1551), .C(n667), .A(n1650), .Y(n180) );
  MUX2XL U1800 ( .D0(ramoe), .D1(n1674), .S(n262), .Y(ramoe_comb) );
  MUX2X1 U1801 ( .D0(pc_o[13]), .D1(n1575), .S(n260), .Y(memaddr_comb[13]) );
  MUX2XL U1802 ( .D0(memaddr[10]), .D1(n1577), .S(n87), .Y(memaddr_comb[10])
         );
  AO2222XL U1803 ( .A(alu_out[13]), .B(n101), .C(n904), .D(n195), .E(pc_i[13]), 
        .F(n168), .G(n670), .H(temp[5]), .Y(n905) );
  NAND32X1 U1804 ( .B(n302), .C(n301), .A(n300), .Y(n825) );
  AO22X1 U1805 ( .A(n1721), .B(n2181), .C(n1056), .D(c), .Y(n302) );
  OAI211X1 U1806 ( .C(n1708), .D(n703), .A(n299), .B(n298), .Y(n301) );
  OA222X1 U1807 ( .A(n2335), .B(n411), .C(n1047), .D(N13353), .E(n1430), .F(
        n2414), .Y(n300) );
  MUX2X1 U1808 ( .D0(memrd), .D1(n1619), .S(n261), .Y(memrd_comb) );
  MUX2X1 U1809 ( .D0(n825), .D1(temp[0]), .S(n1974), .Y(N12824) );
  NAND21X1 U1810 ( .B(n706), .A(n705), .Y(n1571) );
  OA2222XL U1811 ( .A(n788), .B(n1516), .C(n703), .D(n167), .E(n2176), .F(n959), .G(n68), .H(n2470), .Y(n705) );
  AO2222XL U1812 ( .A(alu_out[0]), .B(n913), .C(n196), .D(n702), .E(n740), .F(
        pc_o[0]), .G(n739), .H(pc_i[0]), .Y(n706) );
  INVX1 U1813 ( .A(n742), .Y(n702) );
  NAND21X1 U1814 ( .B(n718), .A(n716), .Y(n1579) );
  OA2222XL U1815 ( .A(n788), .B(n2199), .C(n167), .D(n2434), .E(n2176), .F(
        n946), .G(n697), .H(n715), .Y(n716) );
  AO2222XL U1816 ( .A(alu_out[2]), .B(n913), .C(n196), .D(n714), .E(n740), .F(
        pc_o[2]), .G(pc_i[2]), .H(n739), .Y(n718) );
  NAND21X1 U1817 ( .B(n728), .A(n726), .Y(n1585) );
  OA2222XL U1818 ( .A(n788), .B(n725), .C(n167), .D(n2332), .E(n2176), .F(n936), .G(n697), .H(n2468), .Y(n726) );
  AO2222XL U1819 ( .A(alu_out[4]), .B(n913), .C(n196), .D(n724), .E(n740), .F(
        pc_o[4]), .G(pc_i[4]), .H(n739), .Y(n728) );
  INVX1 U1820 ( .A(n722), .Y(n724) );
  NAND21X1 U1821 ( .B(n738), .A(n736), .Y(n1634) );
  OA2222XL U1822 ( .A(n788), .B(n2208), .C(n2283), .D(n167), .E(n2176), .F(
        n926), .G(n68), .H(n735), .Y(n736) );
  AO2222XL U1823 ( .A(alu_out[6]), .B(n913), .C(n195), .D(n734), .E(n740), .F(
        pc_o[6]), .G(pc_i[6]), .H(n739), .Y(n738) );
  INVX1 U1824 ( .A(n712), .Y(n734) );
  NAND21X1 U1825 ( .B(n713), .A(n711), .Y(n1557) );
  OA2222XL U1826 ( .A(n788), .B(n2197), .C(n2433), .D(n167), .E(n2176), .F(
        n952), .G(n68), .H(n2469), .Y(n711) );
  AO2222XL U1827 ( .A(alu_out[1]), .B(n913), .C(n195), .D(n710), .E(n740), .F(
        pc_o[1]), .G(n739), .H(pc_i[1]), .Y(n713) );
  INVX1 U1828 ( .A(n737), .Y(n710) );
  NAND21X1 U1829 ( .B(n723), .A(n721), .Y(n1593) );
  OA2222XL U1830 ( .A(n788), .B(n2195), .C(n167), .D(n2400), .E(n2176), .F(
        n941), .G(n68), .H(n720), .Y(n721) );
  AO2222XL U1831 ( .A(alu_out[3]), .B(n913), .C(n195), .D(n719), .E(n740), .F(
        pc_o[3]), .G(pc_i[3]), .H(n739), .Y(n723) );
  NAND21X1 U1832 ( .B(n733), .A(n731), .Y(n1621) );
  OA2222XL U1833 ( .A(n788), .B(n730), .C(n167), .D(n2315), .E(n2176), .F(n931), .G(n697), .H(n2467), .Y(n731) );
  AO2222XL U1834 ( .A(alu_out[5]), .B(n913), .C(n1449), .D(n729), .E(n740), 
        .F(memaddr[5]), .G(pc_i[5]), .H(n739), .Y(n733) );
  INVX1 U1835 ( .A(n717), .Y(n729) );
  ENOX1 U1836 ( .A(n612), .B(n2191), .C(N13336), .D(n2191), .Y(n2135) );
  MUX2X1 U1837 ( .D0(pc_o[14]), .D1(n1594), .S(n260), .Y(memaddr_comb[14]) );
  AO2222XL U1838 ( .A(alu_out[14]), .B(n101), .C(n906), .D(n196), .E(pc_i[14]), 
        .F(n168), .G(n670), .H(temp[6]), .Y(n907) );
  MUX2X1 U1839 ( .D0(mempsrd), .D1(n677), .S(n260), .Y(mempsrd_comb) );
  AO21X1 U1840 ( .B(n676), .C(n1600), .A(n1601), .Y(n677) );
  AO22X1 U1841 ( .A(divtempreg[0]), .B(N13343), .C(N13337), .D(n2191), .Y(n184) );
  AO22X1 U1842 ( .A(divtempreg[1]), .B(N13343), .C(N13338), .D(n2191), .Y(n185) );
  AO21X1 U1843 ( .B(n1551), .C(n1627), .A(n288), .Y(n1674) );
  OAI31XL U1844 ( .A(n287), .B(instr[3]), .C(n2324), .D(n2185), .Y(n288) );
  OA222X1 U1845 ( .A(n1784), .B(n102), .C(n1785), .D(n2373), .E(n2410), .F(
        n2389), .Y(n287) );
  AOI221XL U1846 ( .A(instr[2]), .B(n2172), .C(n979), .D(n2407), .E(n974), .Y(
        n1784) );
  XNOR2XL U1847 ( .A(acc[3]), .B(n1376), .Y(N11544) );
  OAI21X1 U1848 ( .B(n1377), .C(n2400), .A(n1378), .Y(N11525) );
  AO2222XL U1849 ( .A(alu_out[15]), .B(n101), .C(n908), .D(n195), .E(pc_i[15]), 
        .F(n168), .G(n670), .H(temp[7]), .Y(n924) );
  OAI22X1 U1850 ( .A(n2317), .B(n645), .C(n145), .D(n15), .Y(N12856) );
  XNOR2XL U1851 ( .A(acc[2]), .B(n1376), .Y(N11543) );
  OAI21X1 U1852 ( .B(n1377), .C(n2434), .A(n2438), .Y(N11524) );
  OAI21BBX1 U1853 ( .A(n583), .B(n584), .C(n585), .Y(
        add_1_root_add_5140_2_carry[2]) );
  NAND41X1 U1854 ( .D(n1417), .A(n1418), .B(n1419), .C(n1420), .Y(n832) );
  AOI22X1 U1855 ( .A(n1372), .B(acc[3]), .C(n2182), .D(ramdatao[7]), .Y(n1420)
         );
  AOI222XL U1856 ( .A(c), .B(n1055), .C(n2304), .D(n612), .E(multemp2[1]), .F(
        n1044), .Y(n1418) );
  OAI21BX1 U1857 ( .C(temp2_comb[7]), .B(n1427), .A(n1428), .Y(n1417) );
  AO21X1 U1858 ( .B(n2010), .C(n1515), .A(n675), .Y(n1601) );
  GEN2XL U1859 ( .D(n674), .E(n496), .C(n2354), .B(n673), .A(n672), .Y(n675)
         );
  AND2X1 U1860 ( .A(cs_run), .B(phase[0]), .Y(n673) );
  INVX1 U1861 ( .A(n668), .Y(n674) );
  NAND21X1 U1862 ( .B(n661), .A(n659), .Y(n1702) );
  MUX2X1 U1863 ( .D0(cs_run), .D1(n1518), .S(codefetch_s), .Y(n661) );
  MUX2X1 U1864 ( .D0(n658), .D1(n657), .S(n1701), .Y(n659) );
  INVX1 U1865 ( .A(state[0]), .Y(n658) );
  MUX2X1 U1866 ( .D0(pc_o[15]), .D1(n1595), .S(n260), .Y(memaddr_comb[15]) );
  NAND3X1 U1867 ( .A(n1453), .B(n1454), .C(n1455), .Y(n831) );
  AOI22X1 U1868 ( .A(acc[2]), .B(n1372), .C(n2182), .D(ramdatao[6]), .Y(n1453)
         );
  AOI222XL U1869 ( .A(n2481), .B(n2180), .C(n2304), .D(n2369), .E(multemp1_0_), 
        .F(n1044), .Y(n1454) );
  AOI221XL U1870 ( .A(acc[5]), .B(n2178), .C(n2179), .D(acc[4]), .E(n1456), 
        .Y(n1455) );
  AO22X1 U1871 ( .A(divtempreg[2]), .B(N13343), .C(N13339), .D(n2191), .Y(n186) );
  NOR2X1 U1872 ( .A(n1726), .B(dec_accop[9]), .Y(n1610) );
  NAND21X1 U1873 ( .B(n748), .A(n747), .Y(n1574) );
  OA2222XL U1874 ( .A(n788), .B(n2209), .C(n746), .D(n167), .E(n2176), .F(n917), .G(n68), .H(n2466), .Y(n747) );
  AO2222XL U1875 ( .A(alu_out[7]), .B(n913), .C(n196), .D(n741), .E(n740), .F(
        pc_o[7]), .G(pc_i[7]), .H(n739), .Y(n748) );
  INVX1 U1876 ( .A(n704), .Y(n741) );
  NAND21X1 U1877 ( .B(n836), .A(n835), .Y(n1578) );
  OA2222XL U1878 ( .A(n2422), .B(n896), .C(n699), .D(n1436), .E(n2414), .F(
        n870), .G(n881), .H(n834), .Y(n835) );
  AO2222XL U1879 ( .A(n1948), .B(pc_i[8]), .C(alu_out[8]), .D(n101), .E(n670), 
        .F(temp[0]), .G(n2476), .H(n2175), .Y(n836) );
  INVX1 U1880 ( .A(p2[0]), .Y(n834) );
  NAND21X1 U1881 ( .B(n866), .A(n838), .Y(n1576) );
  OA2222XL U1882 ( .A(n2423), .B(n896), .C(n684), .D(n1436), .E(n2415), .F(
        n870), .G(n881), .H(n837), .Y(n838) );
  AO2222XL U1883 ( .A(n1948), .B(pc_i[9]), .C(alu_out[9]), .D(n101), .E(
        temp[1]), .F(n670), .G(instr[6]), .H(n2175), .Y(n866) );
  INVX1 U1884 ( .A(p2[1]), .Y(n837) );
  NAND21X1 U1885 ( .B(n869), .A(n868), .Y(n1577) );
  OA2222XL U1886 ( .A(n42), .B(n896), .C(n678), .D(n1436), .E(n870), .F(n2316), 
        .G(n881), .H(n867), .Y(n868) );
  AO2222XL U1887 ( .A(pc_i[10]), .B(n1948), .C(alu_out[10]), .D(n101), .E(
        temp[2]), .F(n670), .G(instr[7]), .H(n2175), .Y(n869) );
  INVX1 U1888 ( .A(p2[2]), .Y(n867) );
  INVX1 U1889 ( .A(n1609), .Y(n2438) );
  GEN2XL U1890 ( .D(acc[3]), .E(n1495), .C(ac), .B(n2452), .A(n2451), .Y(n1609) );
  INVX1 U1891 ( .A(n1492), .Y(n2452) );
  AOI221XL U1892 ( .A(n2449), .B(temp2_comb[0]), .C(dec_accop[5]), .D(n1610), 
        .E(n2451), .Y(n1611) );
  NAND3X1 U1893 ( .A(dec_accop[6]), .B(n2454), .C(n1610), .Y(n1378) );
  NAND2X1 U1894 ( .A(n1483), .B(n1484), .Y(n830) );
  AOI221XL U1895 ( .A(acc[1]), .B(n1372), .C(n2182), .D(ramdatao[5]), .E(n1497), .Y(n1483) );
  AOI221XL U1896 ( .A(acc[4]), .B(n2178), .C(n2179), .D(acc[3]), .E(n1485), 
        .Y(n1484) );
  OAI222XL U1897 ( .A(n612), .B(n2306), .C(acc[5]), .D(n1368), .E(n1498), .F(
        n2369), .Y(n1497) );
  OAI222XL U1898 ( .A(n1457), .B(n2283), .C(n1458), .D(n2369), .E(n1459), .F(
        n1460), .Y(n1456) );
  AOI221XL U1899 ( .A(n2305), .B(n2369), .C(acc[6]), .D(n1371), .E(n1370), .Y(
        n1457) );
  AOI21X1 U1900 ( .B(n2305), .C(n2283), .A(n2262), .Y(n1458) );
  XNOR2XL U1901 ( .A(n1461), .B(n1424), .Y(n1460) );
  OAI222XL U1902 ( .A(n1486), .B(n2315), .C(n1487), .D(n2334), .E(n1459), .F(
        n1488), .Y(n1485) );
  AOI221XL U1903 ( .A(n2305), .B(n2334), .C(acc[5]), .D(n1371), .E(n1370), .Y(
        n1486) );
  AOI21X1 U1904 ( .B(n2305), .C(n2315), .A(n2262), .Y(n1487) );
  XNOR2XL U1905 ( .A(n1489), .B(n1465), .Y(n1488) );
  AOI222XL U1906 ( .A(n2179), .B(acc[5]), .C(n1421), .D(n2181), .E(acc[6]), 
        .F(n2178), .Y(n1419) );
  XOR2X1 U1907 ( .A(n1081), .B(n1080), .Y(n1421) );
  OR2X1 U1908 ( .A(dec_accop[8]), .B(dec_accop[10]), .Y(n1726) );
  INVX1 U1909 ( .A(n626), .Y(n466) );
  NAND41X1 U1910 ( .D(n625), .A(n1391), .B(n1388), .C(n1390), .Y(n626) );
  AOI22X1 U1911 ( .A(pc_o[15]), .B(n391), .C(pc_i[7]), .D(n392), .Y(n1388) );
  AOI222XL U1912 ( .A(pc_i[15]), .B(n2086), .C(pc_o[7]), .D(n2145), .E(n2159), 
        .F(temp2_comb[7]), .Y(n1391) );
  NAND42X1 U1913 ( .C(dec_accop[6]), .D(dec_accop[16]), .A(n1725), .B(n1728), 
        .Y(n1376) );
  NOR2X1 U1914 ( .A(dec_accop[8]), .B(dec_accop[7]), .Y(n1728) );
  AO22X1 U1915 ( .A(divtempreg[3]), .B(N13343), .C(N13340), .D(n2191), .Y(n187) );
  AO22X1 U1916 ( .A(divtempreg[4]), .B(N13343), .C(N13341), .D(n2191), .Y(n188) );
  INVX1 U1917 ( .A(acc[1]), .Y(n2459) );
  XNOR2XL U1918 ( .A(n1376), .B(acc[0]), .Y(n1614) );
  XNOR2XL U1919 ( .A(n1079), .B(n1041), .Y(n1068) );
  NOR2X1 U1920 ( .A(dec_accop[10]), .B(dec_accop[9]), .Y(n1079) );
  NAND2X1 U1921 ( .A(n1522), .B(n1523), .Y(n829) );
  AOI221XL U1922 ( .A(n1372), .B(acc[0]), .C(n2182), .D(ramdatao[4]), .E(n1529), .Y(n1522) );
  AOI221XL U1923 ( .A(acc[3]), .B(n2178), .C(acc[2]), .D(n2179), .E(n1524), 
        .Y(n1523) );
  OAI222XL U1924 ( .A(n2369), .B(n2306), .C(acc[4]), .D(n1368), .E(n1498), .F(
        n2334), .Y(n1529) );
  NAND3X1 U1925 ( .A(n1052), .B(n1053), .C(n1054), .Y(n820) );
  OAI211X1 U1926 ( .C(dec_cop[0]), .D(n1060), .A(n151), .B(n1037), .Y(n1053)
         );
  AOI221XL U1927 ( .A(n1055), .B(n69), .C(n1056), .D(acc[7]), .E(n1057), .Y(
        n1054) );
  AOI21X1 U1928 ( .B(n1068), .C(n2303), .A(n1069), .Y(n1052) );
  NAND3X1 U1929 ( .A(n1610), .B(n2454), .C(dec_accop[18]), .Y(n1492) );
  INVX1 U1930 ( .A(acc[2]), .Y(n2458) );
  OAI222XL U1931 ( .A(n1525), .B(n2332), .C(n1526), .D(n2335), .E(n1459), .F(
        n1527), .Y(n1524) );
  AOI221XL U1932 ( .A(n2305), .B(n2335), .C(acc[4]), .D(n1371), .E(n1370), .Y(
        n1525) );
  AOI21X1 U1933 ( .B(n2305), .C(n2332), .A(n2262), .Y(n1526) );
  XNOR2XL U1934 ( .A(n1528), .B(n2336), .Y(n1527) );
  NOR2X1 U1935 ( .A(dec_accop[5]), .B(dec_accop[18]), .Y(n1725) );
  INVX1 U1936 ( .A(dec_accop[5]), .Y(n2454) );
  XNOR2XL U1937 ( .A(n1727), .B(n1376), .Y(n1612) );
  NAND2X1 U1938 ( .A(c), .B(n1726), .Y(n1727) );
  XNOR2XL U1939 ( .A(n1376), .B(acc[1]), .Y(n584) );
  AO22X1 U1940 ( .A(divtempreg[5]), .B(N13343), .C(N13342), .D(n2191), .Y(n189) );
  INVX1 U1941 ( .A(n600), .Y(n469) );
  NAND41X1 U1942 ( .D(n599), .A(n1440), .B(n1437), .C(n1439), .Y(n600) );
  AOI22X1 U1943 ( .A(memaddr[6]), .B(n2145), .C(pc_i[6]), .D(n392), .Y(n1437)
         );
  AOI222XL U1944 ( .A(pc_i[14]), .B(n2086), .C(pc_o[14]), .D(n391), .E(n2159), 
        .F(temp2_comb[6]), .Y(n1440) );
  NOR43XL U1945 ( .B(n1369), .C(n1723), .D(n1719), .A(dec_accop[15]), .Y(n1035) );
  NAND21X1 U1946 ( .B(dec_accop[7]), .A(n1610), .Y(n1723) );
  NOR32XL U1947 ( .B(n1369), .C(dec_accop[18]), .A(n1051), .Y(n1038) );
  NAND32X1 U1948 ( .B(n1615), .C(n413), .A(n412), .Y(n826) );
  OAI222XL U1949 ( .A(n2446), .B(n2306), .C(acc[1]), .D(n1368), .E(n1498), .F(
        n2458), .Y(n1615) );
  OA222X1 U1950 ( .A(n411), .B(n2334), .C(N13343), .D(n1047), .E(n1430), .F(
        n2415), .Y(n412) );
  AO21X1 U1951 ( .B(acc[0]), .C(n2178), .A(n1604), .Y(n413) );
  NOR32XL U1952 ( .B(n1352), .C(ramsfraddr[6]), .A(n851), .Y(n1375) );
  AOI21X1 U1953 ( .B(n2449), .C(temp2_comb[4]), .A(n2451), .Y(n1468) );
  NAND4X1 U1954 ( .A(n1939), .B(n1940), .C(n1941), .D(n1942), .Y(n1923) );
  NAND4X1 U1955 ( .A(n1931), .B(n1932), .C(n1933), .D(n1934), .Y(n1925) );
  NAND4X1 U1956 ( .A(n1935), .B(n1936), .C(n1937), .D(n1938), .Y(n1924) );
  AO222X1 U1957 ( .A(n391), .B(pc_o[12]), .C(pc_i[12]), .D(n2086), .E(n1531), 
        .F(n2320), .Y(n467) );
  XOR2X1 U1958 ( .A(n1502), .B(n1532), .Y(n1531) );
  XNOR2XL U1959 ( .A(n1503), .B(n2149), .Y(n1532) );
  AOI211X1 U1960 ( .C(n151), .D(dec_accop[17]), .A(n849), .B(n1714), .Y(n1037)
         );
  OR2X1 U1961 ( .A(n1715), .B(n2307), .Y(n1714) );
  INVX1 U1962 ( .A(n153), .Y(n2172) );
  AND2X1 U1963 ( .A(ramsfrwe), .B(ramsfraddr[7]), .Y(n1352) );
  NAND3X1 U1964 ( .A(n1586), .B(n1587), .C(n1588), .Y(n827) );
  AOI22X1 U1965 ( .A(n1372), .B(acc[6]), .C(n2182), .D(ramdatao[2]), .Y(n1586)
         );
  AOI222XL U1966 ( .A(acc[3]), .B(n2180), .C(n1044), .D(acc[4]), .E(
        adder_out[2]), .F(n2181), .Y(n1587) );
  AOI221XL U1967 ( .A(n2179), .B(acc[0]), .C(n2304), .D(n2458), .E(n1589), .Y(
        n1588) );
  NOR2X1 U1968 ( .A(ramsfraddr[4]), .B(ramsfraddr[3]), .Y(n859) );
  INVX1 U1969 ( .A(n2475), .Y(n2436) );
  INVX1 U1970 ( .A(ramsfraddr[1]), .Y(n2440) );
  AOI21X1 U1971 ( .B(n150), .C(dec_accop[1]), .A(n2327), .Y(n1717) );
  NAND3X1 U1972 ( .A(n859), .B(n1375), .C(ramsfraddr[5]), .Y(n1430) );
  AND4X1 U1973 ( .A(n1914), .B(n1915), .C(n1912), .D(n1913), .Y(n324) );
  AOI22X1 U1974 ( .A(rn_reg[180]), .B(n117), .C(rn_reg[212]), .D(n97), .Y(
        n1915) );
  AOI22X1 U1975 ( .A(rn_reg[244]), .B(n58), .C(rn_reg[132]), .D(n65), .Y(n1914) );
  AOI22X1 U1976 ( .A(rn_reg[164]), .B(n79), .C(rn_reg[196]), .D(n135), .Y(
        n1913) );
  NAND3X1 U1977 ( .A(n1562), .B(n1563), .C(n1564), .Y(n828) );
  AOI22X1 U1978 ( .A(n1372), .B(acc[7]), .C(n2182), .D(ramdatao[3]), .Y(n1562)
         );
  AOI222XL U1979 ( .A(acc[4]), .B(n2180), .C(n1044), .D(acc[5]), .E(
        adder_out[3]), .F(n2181), .Y(n1563) );
  AOI221XL U1980 ( .A(acc[1]), .B(n2179), .C(n2304), .D(n2446), .E(n1565), .Y(
        n1564) );
  INVX1 U1981 ( .A(ramsfraddr[0]), .Y(n2444) );
  INVX1 U1982 ( .A(ramsfraddr[2]), .Y(n2443) );
  NAND2X1 U1983 ( .A(dec_accop[13]), .B(n1369), .Y(n1365) );
  NAND2X1 U1984 ( .A(n2479), .B(n2049), .Y(n2040) );
  OAI21X1 U1985 ( .B(instr[2]), .C(n1781), .A(n2048), .Y(n2049) );
  OAI222XL U1986 ( .A(n1566), .B(n2400), .C(n1567), .D(n2446), .E(n1568), .F(
        n2458), .Y(n1565) );
  AOI221XL U1987 ( .A(n2305), .B(n2446), .C(acc[3]), .D(n1371), .E(n1370), .Y(
        n1566) );
  AOI21X1 U1988 ( .B(n2305), .C(n2400), .A(n2262), .Y(n1567) );
  OAI222XL U1989 ( .A(n1590), .B(n2434), .C(n1591), .D(n2458), .E(n1568), .F(
        n2459), .Y(n1589) );
  AOI221XL U1990 ( .A(n2305), .B(n2458), .C(acc[2]), .D(n1371), .E(n1370), .Y(
        n1590) );
  AOI21X1 U1991 ( .B(n2305), .C(n2434), .A(n2262), .Y(n1591) );
  OAI222XL U1992 ( .A(n1605), .B(n2433), .C(n1606), .D(n2459), .E(n1459), .F(
        n1607), .Y(n1604) );
  XOR2X1 U1993 ( .A(n1608), .B(n584), .Y(n1607) );
  AOI221XL U1994 ( .A(n88), .B(n2459), .C(acc[1]), .D(n1371), .E(n1370), .Y(
        n1605) );
  AOI21X1 U1995 ( .B(n88), .C(n2433), .A(n2262), .Y(n1606) );
  AOI211X1 U1996 ( .C(n151), .D(dec_accop[6]), .A(n1710), .B(n1711), .Y(n1712)
         );
  AOI21X1 U1997 ( .B(rn_reg[99]), .C(n112), .A(n1814), .Y(n1927) );
  AOI32X1 U1998 ( .A(n1429), .B(n1430), .C(acc[0]), .D(n2481), .E(n1431), .Y(
        n1428) );
  OAI21X1 U1999 ( .B(temp2_comb[7]), .C(n1365), .A(n1432), .Y(n1431) );
  AOI21X1 U2000 ( .B(rn_reg[228]), .C(n112), .A(n1832), .Y(n1912) );
  INVX1 U2001 ( .A(temp2_comb[1]), .Y(n2433) );
  NAND4X1 U2002 ( .A(n1927), .B(n1928), .C(n1929), .D(n1930), .Y(n1926) );
  AOI22X1 U2003 ( .A(rn_reg[35]), .B(n79), .C(rn_reg[67]), .D(n135), .Y(n1928)
         );
  AOI22X1 U2004 ( .A(rn_reg[51]), .B(n117), .C(rn_reg[83]), .D(n97), .Y(n1930)
         );
  AOI22X1 U2005 ( .A(rn_reg[115]), .B(n58), .C(rn_reg[3]), .D(n65), .Y(n1929)
         );
  NOR32XL U2006 ( .B(n1369), .C(dec_accop[2]), .A(dec_accop[13]), .Y(n1372) );
  AO222X1 U2007 ( .A(n330), .B(n329), .C(n328), .D(n327), .E(n406), .F(n2256), 
        .Y(n931) );
  AND4X1 U2008 ( .A(n1889), .B(n1890), .C(n1887), .D(n1888), .Y(n329) );
  AND4X1 U2009 ( .A(n1897), .B(n1898), .C(n1895), .D(n1896), .Y(n327) );
  NOR21XL U2010 ( .B(dec_accop[0]), .A(n149), .Y(n1429) );
  NAND4X1 U2011 ( .A(n1833), .B(n1834), .C(n1835), .D(n1836), .Y(n1798) );
  NAND4X1 U2012 ( .A(n1815), .B(n1816), .C(n1817), .D(n1818), .Y(n1800) );
  NAND4X1 U2013 ( .A(n1828), .B(n1829), .C(n1830), .D(n1831), .Y(n1799) );
  XNOR2XL U2014 ( .A(n1376), .B(acc[4]), .Y(n1467) );
  OAI221X1 U2015 ( .A(n2309), .B(n483), .C(n1347), .D(n2310), .E(n1348), .Y(
        n1345) );
  AOI33X1 U2016 ( .A(n2427), .B(n1347), .C(ramdatao[2]), .D(n484), .E(n2396), 
        .F(n2482), .Y(n1348) );
  OAI221X1 U2017 ( .A(n2394), .B(n483), .C(n1347), .D(n2395), .E(n1349), .Y(
        n1344) );
  AOI33X1 U2018 ( .A(n2427), .B(n1347), .C(ramdatao[1]), .D(n484), .E(n2396), 
        .F(dps[1]), .Y(n1349) );
  NOR2X1 U2019 ( .A(n2408), .B(n2475), .Y(n1738) );
  NOR21XL U2020 ( .B(dec_accop[4]), .A(n149), .Y(n1729) );
  OAI22X1 U2021 ( .A(n2414), .B(n1151), .C(n2426), .D(n1229), .Y(
        dpl_current[0]) );
  AND4X1 U2022 ( .A(n1230), .B(n1231), .C(n1232), .D(n1233), .Y(n1229) );
  AOI22X1 U2023 ( .A(n1163), .B(dpl_reg[48]), .C(n1164), .D(dpl_reg[56]), .Y(
        n1230) );
  AOI22X1 U2024 ( .A(n1161), .B(dpl_reg[32]), .C(n1162), .D(dpl_reg[40]), .Y(
        n1231) );
  NOR2X1 U2025 ( .A(n2475), .B(n2474), .Y(n765) );
  NOR2X1 U2026 ( .A(n2387), .B(n2479), .Y(n776) );
  NOR42XL U2027 ( .C(accactv), .D(n1709), .A(n1710), .B(dec_accop[6]), .Y(
        n1371) );
  NOR2X1 U2028 ( .A(n1711), .B(n2308), .Y(n1709) );
  NOR2X1 U2029 ( .A(n2411), .B(n153), .Y(n1690) );
  INVX1 U2030 ( .A(n2479), .Y(n2417) );
  AOI21X1 U2031 ( .B(n151), .C(dec_accop[18]), .A(n1051), .Y(n1716) );
  NOR2X1 U2032 ( .A(n2417), .B(n2480), .Y(n1014) );
  INVX1 U2033 ( .A(n2474), .Y(n2408) );
  INVX1 U2034 ( .A(n2480), .Y(n2387) );
  NOR2X1 U2035 ( .A(n2478), .B(instr[2]), .Y(n808) );
  OAI21X1 U2036 ( .B(n1722), .C(n149), .A(n1719), .Y(n1051) );
  NOR3XL U2037 ( .A(n2450), .B(dec_accop[7]), .C(dec_accop[15]), .Y(n1722) );
  NOR2X1 U2038 ( .A(n2417), .B(n2478), .Y(n2048) );
  NOR2X1 U2039 ( .A(n2386), .B(n2478), .Y(n1791) );
  MUX2BXL U2040 ( .D0(n1368), .D1(n1707), .S(acc[0]), .Y(n299) );
  OAI21X1 U2041 ( .B(temp2_comb[0]), .C(n1365), .A(n1432), .Y(n1707) );
  NAND4X1 U2042 ( .A(n2184), .B(n1543), .C(n953), .D(n2009), .Y(n1837) );
  AOI21X1 U2043 ( .B(n1693), .C(phase[1]), .A(n1686), .Y(n2009) );
  AND4X1 U2044 ( .A(n1365), .B(n1366), .C(n1367), .D(n1368), .Y(n1071) );
  AOI21X1 U2045 ( .B(dec_accop[14]), .C(n1369), .A(n1370), .Y(n1367) );
  NOR4XL U2046 ( .A(n1371), .B(n1372), .C(n1373), .D(n1374), .Y(n1366) );
  NOR3XL U2047 ( .A(ramsfraddr[0]), .B(ramsfraddr[2]), .C(n2440), .Y(n864) );
  ENOX1 U2048 ( .A(n1844), .B(n2415), .C(sp[1]), .D(n1844), .Y(N12770) );
  INVX1 U2049 ( .A(acc[5]), .Y(n2334) );
  INVX1 U2050 ( .A(acc[6]), .Y(n2369) );
  INVX1 U2051 ( .A(n876), .Y(n1479) );
  GEN2XL U2052 ( .D(n2079), .E(n2398), .C(test_so), .B(n2080), .A(n2081), .Y(
        n876) );
  NAND21X1 U2053 ( .B(n2079), .A(ckcon[6]), .Y(n2080) );
  AOI222XL U2054 ( .A(ckcon[6]), .B(n2397), .C(ckcon[4]), .D(n2328), .E(
        ckcon[5]), .F(n2329), .Y(n2081) );
  NAND3X1 U2055 ( .A(n1369), .B(n1719), .C(dec_accop[15]), .Y(n1368) );
  AND4X1 U2056 ( .A(n1885), .B(n1886), .C(n1876), .D(n1877), .Y(n330) );
  AOI22X1 U2057 ( .A(rn_reg[117]), .B(n59), .C(rn_reg[5]), .D(n66), .Y(n1885)
         );
  AOI22X1 U2058 ( .A(rn_reg[53]), .B(n118), .C(rn_reg[85]), .D(n98), .Y(n1886)
         );
  AOI22X1 U2059 ( .A(rn_reg[37]), .B(n80), .C(rn_reg[69]), .D(n136), .Y(n1877)
         );
  AND4X1 U2060 ( .A(n2025), .B(n2026), .C(n2023), .D(n2024), .Y(n293) );
  AOI22X1 U2061 ( .A(rn_reg[240]), .B(n59), .C(rn_reg[128]), .D(n66), .Y(n2025) );
  AOI22X1 U2062 ( .A(rn_reg[176]), .B(n118), .C(rn_reg[208]), .D(n98), .Y(
        n2026) );
  AOI22X1 U2063 ( .A(rn_reg[160]), .B(n80), .C(rn_reg[192]), .D(n136), .Y(
        n2024) );
  AND4X1 U2064 ( .A(n1961), .B(n1962), .C(n1959), .D(n1960), .Y(n320) );
  AOI22X1 U2065 ( .A(rn_reg[242]), .B(n59), .C(rn_reg[130]), .D(n66), .Y(n1961) );
  AOI22X1 U2066 ( .A(rn_reg[178]), .B(n118), .C(rn_reg[210]), .D(n98), .Y(
        n1962) );
  AOI22X1 U2067 ( .A(rn_reg[162]), .B(n80), .C(rn_reg[194]), .D(n136), .Y(
        n1960) );
  AND4X1 U2068 ( .A(n1987), .B(n1988), .C(n1985), .D(n1986), .Y(n408) );
  AOI22X1 U2069 ( .A(rn_reg[177]), .B(n118), .C(rn_reg[209]), .D(n98), .Y(
        n1988) );
  AOI22X1 U2070 ( .A(rn_reg[161]), .B(n80), .C(rn_reg[193]), .D(n136), .Y(
        n1986) );
  AOI22X1 U2071 ( .A(rn_reg[241]), .B(n59), .C(rn_reg[129]), .D(n66), .Y(n1987) );
  AND4X1 U2072 ( .A(n1893), .B(n1894), .C(n1891), .D(n1892), .Y(n328) );
  AOI22X1 U2073 ( .A(rn_reg[245]), .B(n59), .C(rn_reg[133]), .D(n66), .Y(n1893) );
  AOI22X1 U2074 ( .A(rn_reg[181]), .B(n118), .C(rn_reg[213]), .D(n98), .Y(
        n1894) );
  AOI22X1 U2075 ( .A(rn_reg[165]), .B(n80), .C(rn_reg[197]), .D(n136), .Y(
        n1892) );
  NOR2X1 U2076 ( .A(n2447), .B(ramsfraddr[3]), .Y(n862) );
  AOI21X1 U2077 ( .B(n2449), .C(temp2_comb[6]), .A(n1462), .Y(n1423) );
  OAI22X1 U2078 ( .A(n2415), .B(n1151), .C(n2426), .D(n1222), .Y(
        dpl_current[1]) );
  AND4X1 U2079 ( .A(n1223), .B(n1224), .C(n1225), .D(n1226), .Y(n1222) );
  AOI22X1 U2080 ( .A(n1163), .B(dpl_reg[49]), .C(n1164), .D(dpl_reg[57]), .Y(
        n1223) );
  AOI22X1 U2081 ( .A(n1161), .B(dpl_reg[33]), .C(n1162), .D(dpl_reg[41]), .Y(
        n1224) );
  OAI22X1 U2082 ( .A(n2316), .B(n1151), .C(n2426), .D(n1215), .Y(
        dpl_current[2]) );
  AND4X1 U2083 ( .A(n1216), .B(n1217), .C(n1218), .D(n1219), .Y(n1215) );
  AOI22X1 U2084 ( .A(n1163), .B(dpl_reg[50]), .C(n1164), .D(dpl_reg[58]), .Y(
        n1216) );
  AOI22X1 U2085 ( .A(n1161), .B(dpl_reg[34]), .C(n1162), .D(dpl_reg[42]), .Y(
        n1217) );
  INVX1 U2086 ( .A(ramsfraddr[5]), .Y(n2445) );
  INVX1 U2087 ( .A(ramsfraddr[4]), .Y(n2447) );
  AOI222XL U2088 ( .A(rn_reg[91]), .B(n77), .C(rn_reg[27]), .D(n115), .E(
        rn_reg[59]), .F(n95), .Y(n1934) );
  AOI222XL U2089 ( .A(rn_reg[219]), .B(n77), .C(rn_reg[155]), .D(n115), .E(
        rn_reg[187]), .F(n95), .Y(n1942) );
  INVX1 U2090 ( .A(ramsfraddr[6]), .Y(n2441) );
  AOI21X1 U2091 ( .B(n2449), .C(temp2_comb[5]), .A(n1462), .Y(n1463) );
  OAI21X1 U2092 ( .B(n1491), .C(n1492), .A(n1378), .Y(n1462) );
  AOI211X1 U2093 ( .C(n2481), .D(n1493), .A(c), .B(n1494), .Y(n1491) );
  NAND2X1 U2094 ( .A(n2334), .B(n2369), .Y(n1493) );
  NOR43XL U2095 ( .B(n1495), .C(n2481), .D(acc[3]), .A(n2335), .Y(n1494) );
  AOI22X1 U2096 ( .A(rn_reg[243]), .B(n58), .C(rn_reg[131]), .D(n65), .Y(n1937) );
  AOI22X1 U2097 ( .A(rn_reg[123]), .B(n139), .C(rn_reg[11]), .D(n99), .Y(n1933) );
  AOI22X1 U2098 ( .A(rn_reg[251]), .B(n139), .C(rn_reg[139]), .D(n99), .Y(
        n1941) );
  AOI22X1 U2099 ( .A(rn_reg[43]), .B(n141), .C(rn_reg[75]), .D(n119), .Y(n1932) );
  AOI22X1 U2100 ( .A(rn_reg[107]), .B(n81), .C(rn_reg[19]), .D(n137), .Y(n1931) );
  AOI22X1 U2101 ( .A(rn_reg[235]), .B(n81), .C(rn_reg[147]), .D(n137), .Y(
        n1939) );
  AOI21X1 U2102 ( .B(rn_reg[227]), .C(n112), .A(n1832), .Y(n1935) );
  AOI21X1 U2103 ( .B(rn_reg[103]), .C(n112), .A(n1814), .Y(n1803) );
  AOI21X1 U2104 ( .B(rn_reg[231]), .C(n112), .A(n1832), .Y(n1828) );
  AOI222XL U2105 ( .A(rn_reg[220]), .B(n77), .C(rn_reg[156]), .D(n115), .E(
        rn_reg[188]), .F(n95), .Y(n1919) );
  AOI222XL U2106 ( .A(rn_reg[92]), .B(n77), .C(rn_reg[28]), .D(n115), .E(
        rn_reg[60]), .F(n95), .Y(n1911) );
  AOI222XL U2107 ( .A(rn_reg[217]), .B(n78), .C(rn_reg[153]), .D(n116), .E(
        rn_reg[185]), .F(n96), .Y(n1992) );
  AOI222XL U2108 ( .A(rn_reg[89]), .B(n78), .C(rn_reg[25]), .D(n116), .E(
        rn_reg[57]), .F(n96), .Y(n1984) );
  NOR2X1 U2109 ( .A(n2040), .B(n2480), .Y(n2046) );
  NOR2X1 U2110 ( .A(n2360), .B(n2480), .Y(n2045) );
  AOI221XL U2111 ( .A(n88), .B(n612), .C(n1371), .D(n2481), .E(n1370), .Y(
        n1427) );
  AOI221XL U2112 ( .A(acc[0]), .B(n1371), .C(n2448), .D(n88), .E(n1370), .Y(
        n1708) );
  INVX1 U2113 ( .A(waitcnt_1_), .Y(n2329) );
  INVX1 U2114 ( .A(temp2_comb[3]), .Y(n2400) );
  AOI22X1 U2115 ( .A(rn_reg[172]), .B(n141), .C(rn_reg[204]), .D(n119), .Y(
        n1917) );
  AOI22X1 U2116 ( .A(n1157), .B(dpl_reg[0]), .C(n1158), .D(dpl_reg[8]), .Y(
        n1233) );
  AOI22X1 U2117 ( .A(n1157), .B(dpl_reg[1]), .C(n1158), .D(dpl_reg[9]), .Y(
        n1226) );
  AOI22X1 U2118 ( .A(n1157), .B(dpl_reg[2]), .C(n1158), .D(dpl_reg[10]), .Y(
        n1219) );
  AOI22X1 U2119 ( .A(rn_reg[236]), .B(n81), .C(rn_reg[148]), .D(n137), .Y(
        n1916) );
  AOI22X1 U2120 ( .A(n1159), .B(dpl_reg[16]), .C(n1160), .D(dpl_reg[24]), .Y(
        n1232) );
  AOI22X1 U2121 ( .A(n1159), .B(dpl_reg[17]), .C(n1160), .D(dpl_reg[25]), .Y(
        n1225) );
  AOI21X1 U2122 ( .B(rn_reg[100]), .C(n112), .A(n1814), .Y(n1904) );
  AOI21X1 U2123 ( .B(rn_reg[224]), .C(n113), .A(n1832), .Y(n2023) );
  AOI21X1 U2124 ( .B(rn_reg[96]), .C(n113), .A(n1814), .Y(n2014) );
  AOI21X1 U2125 ( .B(rn_reg[226]), .C(n113), .A(n1832), .Y(n1959) );
  AOI21X1 U2126 ( .B(rn_reg[225]), .C(n113), .A(n1832), .Y(n1985) );
  AOI21X1 U2127 ( .B(rn_reg[97]), .C(n113), .A(n1814), .Y(n1977) );
  AOI21X1 U2128 ( .B(rn_reg[229]), .C(n113), .A(n1832), .Y(n1891) );
  AOI21X1 U2129 ( .B(rn_reg[101]), .C(n113), .A(n1814), .Y(n1876) );
  INVX1 U2130 ( .A(temp2_comb[2]), .Y(n2434) );
  INVX1 U2131 ( .A(n636), .Y(n892) );
  NAND21X1 U2132 ( .B(n2003), .A(n635), .Y(n636) );
  OAI222XL U2133 ( .A(n1795), .B(n2444), .C(n1090), .D(n2312), .E(n2268), .F(
        n1796), .Y(n2003) );
  AOI22X1 U2134 ( .A(n2002), .B(instr[0]), .C(n2321), .D(n634), .Y(n635) );
  AOI22X1 U2135 ( .A(ckcon[0]), .B(n2328), .C(ckcon[1]), .D(n2329), .Y(n2078)
         );
  NAND2X1 U2136 ( .A(ramdatao[3]), .B(n2427), .Y(n1347) );
  NAND4X1 U2137 ( .A(dec_cop[3]), .B(n1074), .C(n1037), .D(accactv), .Y(n1058)
         );
  AOI31X1 U2138 ( .A(n1070), .B(n1071), .C(n1072), .D(n2455), .Y(n1069) );
  AOI31X1 U2139 ( .A(n1076), .B(n1074), .C(n1077), .D(n2327), .Y(n1070) );
  NOR42XL U2140 ( .C(n1058), .D(n1059), .A(n1038), .B(n1073), .Y(n1072) );
  AOI211X1 U2141 ( .C(dec_cop[7]), .D(n151), .A(n2244), .B(n849), .Y(n1077) );
  NAND2X1 U2142 ( .A(dps[3]), .B(n484), .Y(n483) );
  INVX1 U2143 ( .A(waitcnt_0_), .Y(n2328) );
  NAND4X1 U2144 ( .A(n1803), .B(n1804), .C(n1805), .D(n1806), .Y(n1801) );
  AOI22X1 U2145 ( .A(rn_reg[119]), .B(n58), .C(rn_reg[7]), .D(n65), .Y(n1805)
         );
  AOI22X1 U2146 ( .A(rn_reg[39]), .B(n79), .C(rn_reg[71]), .D(n135), .Y(n1804)
         );
  AOI22X1 U2147 ( .A(rn_reg[55]), .B(n117), .C(rn_reg[87]), .D(n97), .Y(n1806)
         );
  NOR2X1 U2148 ( .A(n2329), .B(ckcon[5]), .Y(n2079) );
  INVX1 U2149 ( .A(test_so), .Y(n2397) );
  INVX1 U2150 ( .A(n877), .Y(n1477) );
  OAI221X1 U2151 ( .A(ckcon[2]), .B(n2397), .C(memwr), .D(memrd), .E(n2076), 
        .Y(n877) );
  OAI22X1 U2152 ( .A(n2077), .B(n2078), .C(test_so), .D(n2330), .Y(n2076) );
  NOR2X1 U2153 ( .A(ckcon[1]), .B(n2329), .Y(n2077) );
  NOR32XL U2154 ( .B(dec_accop[6]), .C(accactv), .A(n1711), .Y(n1373) );
  NOR2X1 U2155 ( .A(n2479), .B(n2480), .Y(n1015) );
  NAND4X1 U2156 ( .A(n1861), .B(n1862), .C(n1863), .D(n1864), .Y(n1845) );
  NAND4X1 U2157 ( .A(n1853), .B(n1854), .C(n1855), .D(n1856), .Y(n1847) );
  NAND4X1 U2158 ( .A(n1857), .B(n1858), .C(n1859), .D(n1860), .Y(n1846) );
  AOI22X1 U2159 ( .A(n484), .B(dps[0]), .C(n2427), .D(ramdatao[0]), .Y(n1101)
         );
  INVX1 U2160 ( .A(n2477), .Y(n2170) );
  NAND21X1 U2161 ( .B(mempswr), .A(n693), .Y(n280) );
  ENOX1 U2162 ( .A(n1844), .B(n2435), .C(sp[3]), .D(n1844), .Y(N12772) );
  ENOX1 U2163 ( .A(n1844), .B(n2316), .C(sp[2]), .D(n1844), .Y(N12771) );
  NOR2X1 U2164 ( .A(n2477), .B(instr[5]), .Y(n819) );
  NOR2X1 U2165 ( .A(n2436), .B(instr[5]), .Y(n1777) );
  XNOR2XL U2166 ( .A(n2387), .B(ramsfraddr[0]), .Y(n2036) );
  NOR2X1 U2167 ( .A(n2170), .B(instr[2]), .Y(n1766) );
  NOR2X1 U2168 ( .A(n25), .B(n2477), .Y(n979) );
  INVX1 U2169 ( .A(acc[4]), .Y(n2335) );
  NAND3X1 U2170 ( .A(n1369), .B(dec_accop[17]), .C(n1720), .Y(n1047) );
  NOR3XL U2171 ( .A(n1051), .B(dec_accop[18]), .C(n849), .Y(n1720) );
  INVX1 U2172 ( .A(ramdatao[3]), .Y(n2435) );
  NAND2X1 U2173 ( .A(phase[2]), .B(n1976), .Y(n697) );
  AOI221XL U2174 ( .A(n443), .B(n2320), .C(n2145), .D(pc_o[2]), .E(n442), .Y(
        n444) );
  AO21X1 U2175 ( .B(temp2_comb[2]), .C(n2159), .A(n1592), .Y(n442) );
  XOR3X1 U2176 ( .A(n2149), .B(n441), .C(n11), .Y(n443) );
  AO222X1 U2177 ( .A(n391), .B(pc_o[10]), .C(n2086), .D(pc_i[10]), .E(n392), 
        .F(pc_i[2]), .Y(n1592) );
  OAI22X1 U2178 ( .A(n2435), .B(n1151), .C(n2426), .D(n1205), .Y(n2141) );
  AND4X1 U2179 ( .A(n1206), .B(n1207), .C(n1208), .D(n1209), .Y(n1205) );
  AOI22X1 U2180 ( .A(n1163), .B(dpl_reg[51]), .C(n1164), .D(dpl_reg[59]), .Y(
        n1206) );
  AOI22X1 U2181 ( .A(n1161), .B(dpl_reg[35]), .C(n1162), .D(dpl_reg[43]), .Y(
        n1207) );
  OAI31XL U2182 ( .A(dec_accop[13]), .B(dec_accop[2]), .C(dec_accop[14]), .D(
        n150), .Y(n1719) );
  AOI222XL U2183 ( .A(rn_reg[94]), .B(n78), .C(rn_reg[30]), .D(n116), .E(
        rn_reg[62]), .F(n96), .Y(n1856) );
  AOI222XL U2184 ( .A(rn_reg[222]), .B(n78), .C(rn_reg[158]), .D(n116), .E(
        rn_reg[190]), .F(n96), .Y(n1864) );
  AOI222XL U2185 ( .A(rn_reg[95]), .B(n77), .C(rn_reg[31]), .D(n115), .E(
        rn_reg[63]), .F(n95), .Y(n1818) );
  AOI222XL U2186 ( .A(rn_reg[223]), .B(n77), .C(rn_reg[159]), .D(n115), .E(
        rn_reg[191]), .F(n95), .Y(n1836) );
  INVX1 U2187 ( .A(ramdatao[4]), .Y(n2169) );
  AOI22X1 U2188 ( .A(rn_reg[179]), .B(n117), .C(rn_reg[211]), .D(n97), .Y(
        n1938) );
  AOI22X1 U2189 ( .A(rn_reg[183]), .B(n117), .C(rn_reg[215]), .D(n97), .Y(
        n1831) );
  AOI22X1 U2190 ( .A(rn_reg[247]), .B(n58), .C(rn_reg[135]), .D(n65), .Y(n1830) );
  AOI22X1 U2191 ( .A(rn_reg[127]), .B(n139), .C(rn_reg[15]), .D(n99), .Y(n1817) );
  AOI22X1 U2192 ( .A(rn_reg[255]), .B(n139), .C(rn_reg[143]), .D(n99), .Y(
        n1835) );
  INVX1 U2193 ( .A(phase[1]), .Y(n2361) );
  AOI22X1 U2194 ( .A(rn_reg[163]), .B(n79), .C(rn_reg[195]), .D(n135), .Y(
        n1936) );
  AOI22X1 U2195 ( .A(rn_reg[171]), .B(n141), .C(rn_reg[203]), .D(n119), .Y(
        n1940) );
  AOI22X1 U2196 ( .A(rn_reg[167]), .B(n79), .C(rn_reg[199]), .D(n135), .Y(
        n1829) );
  AOI22X1 U2197 ( .A(rn_reg[47]), .B(n141), .C(rn_reg[79]), .D(n119), .Y(n1816) );
  AOI22X1 U2198 ( .A(rn_reg[175]), .B(n141), .C(rn_reg[207]), .D(n119), .Y(
        n1834) );
  NAND2X1 U2199 ( .A(dec_accop[3]), .B(n151), .Y(n1718) );
  AOI22X1 U2200 ( .A(rn_reg[111]), .B(n81), .C(rn_reg[23]), .D(n137), .Y(n1815) );
  AOI22X1 U2201 ( .A(rn_reg[239]), .B(n81), .C(rn_reg[151]), .D(n137), .Y(
        n1833) );
  AOI21X1 U2202 ( .B(rn_reg[102]), .C(n113), .A(n1814), .Y(n1849) );
  AOI21X1 U2203 ( .B(rn_reg[230]), .C(n113), .A(n1832), .Y(n1857) );
  AOI222XL U2204 ( .A(rn_reg[216]), .B(n78), .C(rn_reg[152]), .D(n116), .E(
        rn_reg[184]), .F(n96), .Y(n2044) );
  AOI222XL U2205 ( .A(rn_reg[88]), .B(n78), .C(rn_reg[24]), .D(n116), .E(
        rn_reg[56]), .F(n96), .Y(n2022) );
  AOI222XL U2206 ( .A(rn_reg[218]), .B(n78), .C(rn_reg[154]), .D(n116), .E(
        rn_reg[186]), .F(n96), .Y(n1966) );
  AOI222XL U2207 ( .A(rn_reg[221]), .B(n78), .C(rn_reg[157]), .D(n116), .E(
        rn_reg[189]), .F(n96), .Y(n1898) );
  AOI222XL U2208 ( .A(rn_reg[93]), .B(n78), .C(rn_reg[29]), .D(n116), .E(
        rn_reg[61]), .F(n96), .Y(n1890) );
  AOI31X1 U2209 ( .A(n2161), .B(n1737), .C(phase[1]), .D(n1016), .Y(n2006) );
  NAND3X1 U2210 ( .A(n2440), .B(n2443), .C(ramsfraddr[0]), .Y(n853) );
  AOI22X1 U2211 ( .A(rn_reg[36]), .B(n79), .C(rn_reg[68]), .D(n135), .Y(n1905)
         );
  AOI22X1 U2212 ( .A(rn_reg[44]), .B(n141), .C(rn_reg[76]), .D(n119), .Y(n1909) );
  AOI22X1 U2213 ( .A(rn_reg[32]), .B(n80), .C(rn_reg[64]), .D(n136), .Y(n2015)
         );
  AOI22X1 U2214 ( .A(rn_reg[168]), .B(n142), .C(rn_reg[200]), .D(n120), .Y(
        n2042) );
  AOI22X1 U2215 ( .A(rn_reg[40]), .B(n142), .C(rn_reg[72]), .D(n120), .Y(n2020) );
  AOI22X1 U2216 ( .A(rn_reg[33]), .B(n80), .C(rn_reg[65]), .D(n136), .Y(n1978)
         );
  AOI22X1 U2217 ( .A(rn_reg[169]), .B(n142), .C(rn_reg[201]), .D(n120), .Y(
        n1990) );
  AOI22X1 U2218 ( .A(rn_reg[41]), .B(n142), .C(rn_reg[73]), .D(n120), .Y(n1982) );
  AOI22X1 U2219 ( .A(rn_reg[173]), .B(n142), .C(rn_reg[205]), .D(n120), .Y(
        n1896) );
  AOI22X1 U2220 ( .A(rn_reg[45]), .B(n142), .C(rn_reg[77]), .D(n120), .Y(n1888) );
  AOI22X1 U2221 ( .A(n1157), .B(dpl_reg[3]), .C(n1158), .D(dpl_reg[11]), .Y(
        n1209) );
  AOI22X1 U2222 ( .A(rn_reg[108]), .B(n81), .C(rn_reg[20]), .D(n137), .Y(n1908) );
  AOI22X1 U2223 ( .A(rn_reg[232]), .B(n82), .C(rn_reg[144]), .D(n138), .Y(
        n2041) );
  AOI22X1 U2224 ( .A(rn_reg[104]), .B(n82), .C(rn_reg[16]), .D(n138), .Y(n2019) );
  AOI22X1 U2225 ( .A(rn_reg[233]), .B(n82), .C(rn_reg[145]), .D(n138), .Y(
        n1989) );
  AOI22X1 U2226 ( .A(rn_reg[105]), .B(n82), .C(rn_reg[17]), .D(n138), .Y(n1981) );
  AOI22X1 U2227 ( .A(rn_reg[237]), .B(n82), .C(rn_reg[149]), .D(n138), .Y(
        n1895) );
  AOI22X1 U2228 ( .A(rn_reg[109]), .B(n82), .C(rn_reg[21]), .D(n138), .Y(n1887) );
  AOI22X1 U2229 ( .A(n1159), .B(dpl_reg[18]), .C(n1160), .D(dpl_reg[26]), .Y(
        n1218) );
  AOI22X1 U2230 ( .A(n1159), .B(dpl_reg[19]), .C(n1160), .D(dpl_reg[27]), .Y(
        n1208) );
  AOI22X1 U2231 ( .A(rn_reg[116]), .B(n58), .C(rn_reg[4]), .D(n65), .Y(n1906)
         );
  AOI22X1 U2232 ( .A(rn_reg[252]), .B(n139), .C(rn_reg[140]), .D(n99), .Y(
        n1918) );
  AOI22X1 U2233 ( .A(rn_reg[124]), .B(n139), .C(rn_reg[12]), .D(n99), .Y(n1910) );
  AOI22X1 U2234 ( .A(rn_reg[112]), .B(n59), .C(rn_reg[0]), .D(n66), .Y(n2016)
         );
  AOI22X1 U2235 ( .A(rn_reg[248]), .B(n140), .C(rn_reg[136]), .D(n100), .Y(
        n2043) );
  AOI22X1 U2236 ( .A(rn_reg[120]), .B(n140), .C(rn_reg[8]), .D(n100), .Y(n2021) );
  AOI22X1 U2237 ( .A(rn_reg[113]), .B(n59), .C(rn_reg[1]), .D(n66), .Y(n1979)
         );
  AOI22X1 U2238 ( .A(rn_reg[249]), .B(n140), .C(rn_reg[137]), .D(n100), .Y(
        n1991) );
  AOI22X1 U2239 ( .A(rn_reg[121]), .B(n140), .C(rn_reg[9]), .D(n100), .Y(n1983) );
  AOI22X1 U2240 ( .A(rn_reg[253]), .B(n140), .C(rn_reg[141]), .D(n100), .Y(
        n1897) );
  AOI22X1 U2241 ( .A(rn_reg[52]), .B(n117), .C(rn_reg[84]), .D(n97), .Y(n1907)
         );
  AOI22X1 U2242 ( .A(rn_reg[48]), .B(n118), .C(rn_reg[80]), .D(n98), .Y(n2017)
         );
  AOI22X1 U2243 ( .A(rn_reg[49]), .B(n118), .C(rn_reg[81]), .D(n98), .Y(n1980)
         );
  AOI21X1 U2244 ( .B(rn_reg[98]), .C(n113), .A(n1814), .Y(n1951) );
  NAND2X1 U2245 ( .A(dec_accop[11]), .B(accactv), .Y(n1713) );
  INVX1 U2246 ( .A(interrupt), .Y(n2168) );
  INVX1 U2247 ( .A(n2324), .Y(n254) );
  INVX1 U2248 ( .A(phase[0]), .Y(n2324) );
  NAND4X1 U2249 ( .A(n1849), .B(n1850), .C(n1851), .D(n1852), .Y(n1848) );
  AOI22X1 U2250 ( .A(rn_reg[38]), .B(n80), .C(rn_reg[70]), .D(n136), .Y(n1850)
         );
  AOI22X1 U2251 ( .A(rn_reg[54]), .B(n118), .C(rn_reg[86]), .D(n98), .Y(n1852)
         );
  AOI22X1 U2252 ( .A(rn_reg[118]), .B(n59), .C(rn_reg[6]), .D(n66), .Y(n1851)
         );
  INVX1 U2253 ( .A(ckcon[6]), .Y(n2398) );
  INVX1 U2254 ( .A(dps[3]), .Y(n2396) );
  INVX1 U2255 ( .A(ckcon[2]), .Y(n2330) );
  INVX1 U2256 ( .A(rs[0]), .Y(n2395) );
  INVX1 U2257 ( .A(rs[1]), .Y(n2310) );
  MUX2AXL U2258 ( .D0(pmw), .D1(n2169), .S(n487), .Y(n2011) );
  NOR43XL U2259 ( .B(n2165), .C(n2166), .D(n641), .A(n839), .Y(n642) );
  INVX1 U2260 ( .A(phase[5]), .Y(n641) );
  NAND3X1 U2261 ( .A(n255), .B(n2275), .C(n252), .Y(n839) );
  NAND21X1 U2262 ( .B(n640), .A(n639), .Y(n620) );
  AOI222XL U2263 ( .A(n2088), .B(phase[0]), .C(n662), .D(phase[4]), .E(n638), 
        .F(phase[1]), .Y(n639) );
  AO21X1 U2264 ( .B(n2089), .C(phase[2]), .A(n2090), .Y(n640) );
  OAI2B11X1 U2265 ( .D(n2103), .C(n51), .A(n2104), .B(n2105), .Y(n2088) );
  OAI22X1 U2269 ( .A(n880), .B(n2113), .C(n2114), .D(n2424), .Y(n609) );
  AOI22X1 U2270 ( .A(ckcon[7]), .B(n496), .C(ckcon[3]), .D(n2011), .Y(n2113)
         );
  AOI22X1 U2271 ( .A(n496), .B(ramdatao[7]), .C(ramdatao[3]), .D(n2011), .Y(
        n2114) );
  AND2X1 U2272 ( .A(dec_accop[16]), .B(accactv), .Y(n849) );
  AO222X1 U2273 ( .A(n23), .B(pc_o[10]), .C(n21), .D(n1577), .E(pc_ini[10]), 
        .F(n269), .Y(N490) );
  AO222X1 U2274 ( .A(n24), .B(pc_o[9]), .C(n22), .D(n1576), .E(pc_ini[9]), .F(
        n269), .Y(N489) );
  AO222X1 U2275 ( .A(n23), .B(pc_o[8]), .C(n21), .D(n1578), .E(pc_ini[8]), .F(
        n269), .Y(N488) );
  AO222X1 U2276 ( .A(n24), .B(pc_o[7]), .C(n22), .D(n1574), .E(pc_ini[7]), .F(
        n269), .Y(N487) );
  AO222X1 U2277 ( .A(n23), .B(memaddr[6]), .C(n21), .D(n1634), .E(pc_ini[6]), 
        .F(n269), .Y(N486) );
  AO222X1 U2278 ( .A(n24), .B(memaddr[5]), .C(n22), .D(n1621), .E(pc_ini[5]), 
        .F(n269), .Y(N485) );
  AO222X1 U2279 ( .A(n23), .B(pc_o[4]), .C(n21), .D(n1585), .E(pc_ini[4]), .F(
        n269), .Y(N484) );
  AO222X1 U2280 ( .A(n24), .B(pc_o[3]), .C(n22), .D(n1593), .E(pc_ini[3]), .F(
        n273), .Y(N483) );
  AO222X1 U2281 ( .A(n23), .B(pc_o[2]), .C(n21), .D(n1579), .E(pc_ini[2]), .F(
        n272), .Y(N482) );
  AO222X1 U2282 ( .A(n24), .B(pc_o[1]), .C(n22), .D(n1557), .E(pc_ini[1]), .F(
        n273), .Y(N481) );
  AO222X1 U2283 ( .A(n23), .B(pc_o[0]), .C(n21), .D(n1571), .E(pc_ini[0]), .F(
        n271), .Y(N480) );
  AOI22AXL U2284 ( .A(n1692), .B(phase[1]), .D(n1997), .C(phase[0]), .Y(n1945)
         );
  NOR4XL U2285 ( .A(n1998), .B(n1692), .C(n1691), .D(n1999), .Y(n1997) );
  NAND2X1 U2286 ( .A(n2000), .B(n1768), .Y(n1998) );
  AOI32X1 U2287 ( .A(n2479), .B(n2377), .C(n1026), .D(n2001), .E(n2407), .Y(
        n2000) );
  XNOR2XL U2288 ( .A(n1376), .B(n2481), .Y(n1422) );
  ENOX1 U2289 ( .A(n134), .B(n2169), .C(sp[4]), .D(n134), .Y(N12773) );
  AND3X1 U2290 ( .A(dec_accop[1]), .B(n151), .C(n1364), .Y(n1055) );
  INVX1 U2291 ( .A(ramdatao[1]), .Y(n2415) );
  AO21X1 U2292 ( .B(waitstaten), .C(n1663), .A(n273), .Y(N520) );
  MUX2X1 U2293 ( .D0(p2sel), .D1(n1662), .S(n1661), .Y(n1663) );
  AO22X1 U2294 ( .A(n215), .B(n1595), .C(pc_ini[15]), .D(n271), .Y(N495) );
  AO22X1 U2295 ( .A(n214), .B(n1594), .C(pc_ini[14]), .D(n271), .Y(N494) );
  AO22X1 U2296 ( .A(n214), .B(n1575), .C(pc_ini[13]), .D(n271), .Y(N493) );
  AO22X1 U2297 ( .A(n214), .B(n1580), .C(pc_ini[12]), .D(n271), .Y(N492) );
  AO22X1 U2298 ( .A(n214), .B(n1581), .C(pc_ini[11]), .D(n271), .Y(N491) );
  NOR2X1 U2299 ( .A(n1111), .B(n2482), .Y(n207) );
  NOR2X1 U2300 ( .A(n1110), .B(n2482), .Y(n205) );
  NOR2X1 U2301 ( .A(n1109), .B(n2482), .Y(n208) );
  NOR2X1 U2302 ( .A(n1109), .B(n2482), .Y(n516) );
  OAI22X1 U2303 ( .A(n2169), .B(n1151), .C(n2426), .D(n1193), .Y(n2142) );
  AND4X1 U2304 ( .A(n1194), .B(n1195), .C(n1196), .D(n1197), .Y(n1193) );
  AOI22X1 U2305 ( .A(n1163), .B(dpl_reg[52]), .C(n1164), .D(dpl_reg[60]), .Y(
        n1194) );
  AOI22X1 U2306 ( .A(n1161), .B(dpl_reg[36]), .C(n1162), .D(dpl_reg[44]), .Y(
        n1195) );
  OAI22X1 U2307 ( .A(n2256), .B(n1151), .C(n2426), .D(n1183), .Y(
        dpl_current[5]) );
  AND4X1 U2308 ( .A(n1184), .B(n1185), .C(n1186), .D(n1187), .Y(n1183) );
  AOI22X1 U2309 ( .A(n1163), .B(dpl_reg[53]), .C(n1164), .D(dpl_reg[61]), .Y(
        n1184) );
  AOI22X1 U2310 ( .A(n1161), .B(dpl_reg[37]), .C(n1162), .D(dpl_reg[45]), .Y(
        n1185) );
  NAND2X1 U2311 ( .A(dps[0]), .B(n2390), .Y(n1110) );
  NAND2X1 U2312 ( .A(dps[1]), .B(n2392), .Y(n1109) );
  INVX1 U2313 ( .A(ramdatao[2]), .Y(n2316) );
  INVX1 U2314 ( .A(ramsfraddr[3]), .Y(n2432) );
  NAND2X1 U2315 ( .A(n2382), .B(phase[1]), .Y(n1758) );
  OAI221X1 U2316 ( .A(n2474), .B(n1785), .C(n2386), .D(n2347), .E(n2100), .Y(
        n757) );
  GEN2XL U2317 ( .D(instr[4]), .E(n609), .C(n2408), .B(n2381), .A(instr[2]), 
        .Y(n2100) );
  AOI22X1 U2318 ( .A(rn_reg[182]), .B(n118), .C(rn_reg[214]), .D(n98), .Y(
        n1860) );
  AOI22X1 U2319 ( .A(n515), .B(dph_reg[4]), .C(n208), .D(dph_reg[20]), .Y(n566) );
  AOI22X1 U2320 ( .A(n207), .B(dpl_reg[4]), .C(n516), .D(dpl_reg[20]), .Y(n534) );
  AOI22X1 U2321 ( .A(n20), .B(dph_reg[5]), .C(n18), .D(dph_reg[21]), .Y(n562)
         );
  AOI22X1 U2322 ( .A(rn_reg[246]), .B(n59), .C(rn_reg[134]), .D(n66), .Y(n1859) );
  AOI22X1 U2323 ( .A(rn_reg[126]), .B(n140), .C(rn_reg[14]), .D(n100), .Y(
        n1855) );
  AOI22X1 U2324 ( .A(rn_reg[254]), .B(n140), .C(rn_reg[142]), .D(n100), .Y(
        n1863) );
  AOI22X1 U2325 ( .A(n205), .B(dph_reg[12]), .C(n206), .D(dph_reg[28]), .Y(
        n565) );
  AOI21X1 U2326 ( .B(n2449), .C(temp2_comb[7]), .A(n2451), .Y(n1080) );
  AOI22X1 U2327 ( .A(rn_reg[166]), .B(n80), .C(rn_reg[198]), .D(n136), .Y(
        n1858) );
  AOI22X1 U2328 ( .A(rn_reg[46]), .B(n142), .C(rn_reg[78]), .D(n120), .Y(n1854) );
  AOI22X1 U2329 ( .A(rn_reg[174]), .B(n142), .C(rn_reg[206]), .D(n120), .Y(
        n1862) );
  AOI22X1 U2330 ( .A(n202), .B(dph_reg[36]), .C(n204), .D(dph_reg[52]), .Y(
        n564) );
  AOI22X1 U2331 ( .A(rn_reg[110]), .B(n82), .C(rn_reg[22]), .D(n138), .Y(n1853) );
  AOI22X1 U2332 ( .A(rn_reg[238]), .B(n82), .C(rn_reg[150]), .D(n138), .Y(
        n1861) );
  AOI222XL U2333 ( .A(rn_reg[90]), .B(n78), .C(rn_reg[26]), .D(n116), .E(
        rn_reg[58]), .F(n96), .Y(n1958) );
  OAI221X1 U2334 ( .A(n2210), .B(n1706), .C(n1705), .D(n1704), .E(n275), .Y(
        n1878) );
  INVX1 U2335 ( .A(newinstrlock), .Y(n2210) );
  OAI22AX1 U2336 ( .D(idle), .C(n1660), .A(n2163), .B(n1704), .Y(n1879) );
  INVX1 U2337 ( .A(dps[1]), .Y(n2390) );
  AOI22X1 U2338 ( .A(rn_reg[34]), .B(n80), .C(rn_reg[66]), .D(n136), .Y(n1952)
         );
  AOI22X1 U2339 ( .A(rn_reg[170]), .B(n142), .C(rn_reg[202]), .D(n120), .Y(
        n1964) );
  AOI22X1 U2340 ( .A(rn_reg[42]), .B(n142), .C(rn_reg[74]), .D(n120), .Y(n1956) );
  AOI22X1 U2341 ( .A(n1157), .B(dpl_reg[4]), .C(n1158), .D(dpl_reg[12]), .Y(
        n1197) );
  AOI22X1 U2342 ( .A(n1157), .B(dpl_reg[5]), .C(n1158), .D(dpl_reg[13]), .Y(
        n1187) );
  AOI22X1 U2343 ( .A(rn_reg[234]), .B(n82), .C(rn_reg[146]), .D(n138), .Y(
        n1963) );
  AOI22X1 U2344 ( .A(rn_reg[106]), .B(n82), .C(rn_reg[18]), .D(n138), .Y(n1955) );
  AOI22X1 U2345 ( .A(n1159), .B(dpl_reg[20]), .C(n1160), .D(dpl_reg[28]), .Y(
        n1196) );
  AOI22X1 U2346 ( .A(rn_reg[114]), .B(n59), .C(rn_reg[2]), .D(n66), .Y(n1953)
         );
  AOI22X1 U2347 ( .A(rn_reg[250]), .B(n140), .C(rn_reg[138]), .D(n100), .Y(
        n1965) );
  AOI22X1 U2348 ( .A(rn_reg[122]), .B(n140), .C(rn_reg[10]), .D(n100), .Y(
        n1957) );
  AOI22X1 U2349 ( .A(rn_reg[125]), .B(n140), .C(rn_reg[13]), .D(n100), .Y(
        n1889) );
  AOI22X1 U2350 ( .A(rn_reg[50]), .B(n118), .C(rn_reg[82]), .D(n98), .Y(n1954)
         );
  INVX1 U2351 ( .A(dps[0]), .Y(n2392) );
  INVX1 U2352 ( .A(mempsrd), .Y(n693) );
  OAI21AX1 U2353 ( .B(n2093), .C(n2094), .A(n755), .Y(n2089) );
  AOI22X1 U2354 ( .A(n751), .B(n752), .C(n1733), .D(n776), .Y(n2093) );
  AOI32X1 U2355 ( .A(n979), .B(n2436), .C(interrupt), .D(n2475), .E(n757), .Y(
        n2094) );
  INVX1 U2356 ( .A(dec_accop[12]), .Y(n2308) );
  INVX1 U2357 ( .A(ramwe), .Y(n2263) );
  NAND21X1 U2358 ( .B(instr[5]), .A(n2157), .Y(n343) );
  NAND21X1 U2359 ( .B(n2475), .A(n1336), .Y(n2356) );
  NOR4XL U2360 ( .A(n1774), .B(n1775), .C(n778), .D(n591), .Y(n1773) );
  AO2222XL U2361 ( .A(n2144), .B(n2157), .C(n1669), .D(n1738), .E(n2147), .F(
        n1777), .G(n1780), .H(n2189), .Y(n1774) );
  OAI22X1 U2362 ( .A(n1763), .B(n2342), .C(instr[0]), .D(n1776), .Y(n1775) );
  AO21X1 U2363 ( .B(n367), .C(N345), .A(n1411), .Y(n418) );
  NAND32X1 U2364 ( .B(n2476), .C(n928), .A(n2144), .Y(n317) );
  NAND21X1 U2365 ( .B(n1542), .A(n1530), .Y(n451) );
  OAI22X1 U2366 ( .A(n1679), .B(n257), .C(n1680), .D(n2324), .Y(n1530) );
  AOI22X1 U2367 ( .A(n775), .B(instr[3]), .C(n1681), .D(n1682), .Y(n1680) );
  AOI32X1 U2368 ( .A(n1683), .B(instr[0]), .C(n775), .D(n764), .E(n1684), .Y(
        n1679) );
  NOR42XL U2369 ( .C(ramsfraddr[3]), .D(n1114), .A(ramsfraddr[4]), .B(n856), 
        .Y(n880) );
  OR2X1 U2370 ( .A(memwr), .B(memrd), .Y(n278) );
  AOI222XL U2371 ( .A(dptr_inc[8]), .B(n148), .C(n1247), .D(dph_current[0]), 
        .E(n1022), .F(temp[0]), .Y(n699) );
  AOI222XL U2372 ( .A(dptr_inc[9]), .B(n148), .C(n1247), .D(dph_current[1]), 
        .E(n1022), .F(temp[1]), .Y(n684) );
  INVX1 U2373 ( .A(n2482), .Y(n2293) );
  OAI31XL U2374 ( .A(n2111), .B(n2416), .C(n152), .D(n2112), .Y(n662) );
  NAND4X1 U2375 ( .A(n608), .B(n1015), .C(instr[4]), .D(n609), .Y(n2112) );
  AOI32X1 U2376 ( .A(n1682), .B(n609), .C(n1766), .D(n974), .E(instr[7]), .Y(
        n2111) );
  NOR2X1 U2377 ( .A(n2417), .B(n2477), .Y(n792) );
  INVX1 U2378 ( .A(n2478), .Y(n2171) );
  NOR2X1 U2379 ( .A(n2430), .B(n2474), .Y(n781) );
  NOR2X1 U2380 ( .A(n25), .B(n2478), .Y(n1683) );
  INVX1 U2381 ( .A(acc[0]), .Y(n2448) );
  NOR2X1 U2382 ( .A(n2407), .B(n153), .Y(n980) );
  INVX1 U2383 ( .A(acc[3]), .Y(n2446) );
  NOR2X1 U2384 ( .A(n2436), .B(n2474), .Y(n982) );
  NOR2X1 U2385 ( .A(n1111), .B(n2482), .Y(n515) );
  NOR2X1 U2386 ( .A(n1107), .B(n2482), .Y(n206) );
  NAND4X1 U2387 ( .A(phase[0]), .B(n808), .C(n1995), .D(n2387), .Y(n1755) );
  OAI222XL U2388 ( .A(n2479), .B(n1792), .C(n1996), .D(n2417), .E(n610), .F(
        n2412), .Y(n1995) );
  AOI21X1 U2389 ( .B(n2474), .C(n2172), .A(n1738), .Y(n1996) );
  OAI22X1 U2390 ( .A(n2255), .B(n1151), .C(n2426), .D(n1170), .Y(n2143) );
  AND4X1 U2391 ( .A(n1171), .B(n1172), .C(n1173), .D(n1174), .Y(n1170) );
  AOI22X1 U2392 ( .A(n1163), .B(dpl_reg[54]), .C(n1164), .D(dpl_reg[62]), .Y(
        n1171) );
  AOI22X1 U2393 ( .A(n1161), .B(dpl_reg[38]), .C(n1162), .D(dpl_reg[46]), .Y(
        n1172) );
  NAND3X1 U2394 ( .A(instr[5]), .B(n2387), .C(n792), .Y(n2056) );
  NAND2X1 U2395 ( .A(dps[1]), .B(dps[0]), .Y(n1107) );
  INVX1 U2396 ( .A(b[0]), .Y(n2464) );
  INVX1 U2397 ( .A(b[1]), .Y(n2463) );
  NAND3X1 U2398 ( .A(ramsfraddr[1]), .B(ramsfraddr[2]), .C(ramsfraddr[0]), .Y(
        n857) );
  AOI22X1 U2399 ( .A(dpc_tab[0]), .B(n515), .C(dpc_tab[12]), .D(n208), .Y(
        n1327) );
  AOI22X1 U2400 ( .A(dpc_tab[4]), .B(n207), .C(dpc_tab[16]), .D(n208), .Y(
        n1100) );
  AOI22X1 U2401 ( .A(dpc_tab[5]), .B(n515), .C(dpc_tab[17]), .D(n18), .Y(n1096) );
  AOI22X1 U2402 ( .A(n20), .B(dph_reg[3]), .C(n516), .D(dph_reg[19]), .Y(n570)
         );
  AOI22X1 U2403 ( .A(n207), .B(dpl_reg[0]), .C(n208), .D(dpl_reg[16]), .Y(n550) );
  AOI22X1 U2404 ( .A(n515), .B(dph_reg[0]), .C(n208), .D(dph_reg[16]), .Y(n582) );
  AOI22X1 U2405 ( .A(n207), .B(dph_reg[6]), .C(n516), .D(dph_reg[22]), .Y(n558) );
  AOI22X1 U2406 ( .A(n515), .B(dpl_reg[6]), .C(n208), .D(dpl_reg[22]), .Y(n526) );
  AOI22X1 U2407 ( .A(n515), .B(dpl_reg[7]), .C(n18), .D(dpl_reg[23]), .Y(n514)
         );
  AOI22X1 U2408 ( .A(n515), .B(dpl_reg[5]), .C(n18), .D(dpl_reg[21]), .Y(n530)
         );
  AOI22X1 U2409 ( .A(n515), .B(dph_reg[2]), .C(n208), .D(dph_reg[18]), .Y(n574) );
  AOI22X1 U2410 ( .A(n515), .B(dpl_reg[2]), .C(n208), .D(dpl_reg[18]), .Y(n542) );
  NOR2X1 U2411 ( .A(dec_cop[1]), .B(n1061), .Y(n1060) );
  AOI32X1 U2412 ( .A(n1062), .B(n1063), .C(n1064), .D(N11584), .E(n1065), .Y(
        n1061) );
  OAI21BBX1 U2413 ( .A(n2251), .B(dec_cop[7]), .C(n2455), .Y(n1063) );
  OAI21BBX1 U2414 ( .A(c), .B(dec_cop[4]), .C(n1066), .Y(n1065) );
  NOR2X1 U2415 ( .A(n2448), .B(n2463), .Y(N14337) );
  AOI22X1 U2416 ( .A(n205), .B(dpl_reg[8]), .C(n206), .D(dpl_reg[24]), .Y(n549) );
  AOI22X1 U2417 ( .A(n53), .B(dph_reg[8]), .C(n49), .D(dph_reg[24]), .Y(n581)
         );
  AOI22X1 U2418 ( .A(n205), .B(dph_reg[14]), .C(n206), .D(dph_reg[30]), .Y(
        n557) );
  AOI22X1 U2419 ( .A(n205), .B(dpl_reg[14]), .C(n206), .D(dpl_reg[30]), .Y(
        n525) );
  AOI22X1 U2420 ( .A(n205), .B(dpl_reg[12]), .C(n206), .D(dpl_reg[28]), .Y(
        n533) );
  AOI22X1 U2421 ( .A(n1), .B(dph_reg[13]), .C(n2), .D(dph_reg[29]), .Y(n561)
         );
  AOI22X1 U2422 ( .A(n1), .B(dpl_reg[13]), .C(n2), .D(dpl_reg[29]), .Y(n529)
         );
  AOI22X1 U2423 ( .A(n205), .B(dph_reg[10]), .C(n206), .D(dph_reg[26]), .Y(
        n573) );
  AOI22X1 U2424 ( .A(n205), .B(dpl_reg[10]), .C(n206), .D(dpl_reg[26]), .Y(
        n541) );
  AOI22X1 U2425 ( .A(n201), .B(dph_reg[35]), .C(n203), .D(dph_reg[51]), .Y(
        n568) );
  AOI22X1 U2426 ( .A(n519), .B(dpl_reg[32]), .C(n520), .D(dpl_reg[48]), .Y(
        n548) );
  AOI22X1 U2427 ( .A(n201), .B(dph_reg[32]), .C(n203), .D(dph_reg[48]), .Y(
        n580) );
  AOI22X1 U2428 ( .A(n201), .B(dph_reg[38]), .C(n203), .D(dph_reg[54]), .Y(
        n556) );
  AOI22X1 U2429 ( .A(n519), .B(dpl_reg[38]), .C(n520), .D(dpl_reg[54]), .Y(
        n524) );
  AOI22X1 U2430 ( .A(n201), .B(dpl_reg[36]), .C(n203), .D(dpl_reg[52]), .Y(
        n532) );
  AOI22X1 U2431 ( .A(n519), .B(dph_reg[37]), .C(n520), .D(dph_reg[53]), .Y(
        n560) );
  AOI22X1 U2432 ( .A(n202), .B(dpl_reg[37]), .C(n204), .D(dpl_reg[53]), .Y(
        n528) );
  AOI22X1 U2433 ( .A(n519), .B(dph_reg[34]), .C(n520), .D(dph_reg[50]), .Y(
        n572) );
  AOI22X1 U2434 ( .A(n202), .B(dpl_reg[34]), .C(n204), .D(dpl_reg[50]), .Y(
        n540) );
  AOI22X1 U2435 ( .A(n521), .B(dpl_reg[40]), .C(n522), .D(dpl_reg[56]), .Y(
        n547) );
  AOI22X1 U2436 ( .A(n197), .B(dph_reg[46]), .C(n199), .D(dph_reg[62]), .Y(
        n555) );
  AOI22X1 U2437 ( .A(n521), .B(dpl_reg[46]), .C(n522), .D(dpl_reg[62]), .Y(
        n523) );
  AOI22X1 U2438 ( .A(n198), .B(dph_reg[44]), .C(n200), .D(dph_reg[60]), .Y(
        n563) );
  AOI22X1 U2439 ( .A(n521), .B(dph_reg[45]), .C(n522), .D(dph_reg[61]), .Y(
        n559) );
  NOR2X1 U2440 ( .A(n2171), .B(n2477), .Y(n2053) );
  OAI21X1 U2441 ( .B(N11584), .C(n2251), .A(c), .Y(n1062) );
  NAND3X1 U2442 ( .A(n1015), .B(n2477), .C(n2156), .Y(n1023) );
  AOI32X1 U2443 ( .A(n1777), .B(instr[4]), .C(n1336), .D(n792), .E(n1026), .Y(
        n1776) );
  AOI22X1 U2444 ( .A(n1157), .B(dpl_reg[6]), .C(n1158), .D(dpl_reg[14]), .Y(
        n1174) );
  AOI21X1 U2445 ( .B(accactv), .C(n1078), .A(n2307), .Y(n1076) );
  OR4X1 U2446 ( .A(dec_accop[17]), .B(dec_accop[1]), .C(dec_accop[4]), .D(
        dec_cop[6]), .Y(n1078) );
  AOI22X1 U2447 ( .A(n1159), .B(dpl_reg[21]), .C(n1160), .D(dpl_reg[29]), .Y(
        n1186) );
  AOI22X1 U2448 ( .A(n1159), .B(dpl_reg[22]), .C(n1160), .D(dpl_reg[30]), .Y(
        n1173) );
  NAND4X1 U2449 ( .A(n1324), .B(n1325), .C(n1326), .D(n1327), .Y(dpc[0]) );
  AOI22X1 U2450 ( .A(dpc_tab[30]), .B(n521), .C(dpc_tab[42]), .D(n522), .Y(
        n1324) );
  AOI22X1 U2451 ( .A(dpc_tab[6]), .B(n205), .C(dpc_tab[18]), .D(n206), .Y(
        n1326) );
  AOI22X1 U2452 ( .A(dpc_tab[24]), .B(n519), .C(dpc_tab[36]), .D(n520), .Y(
        n1325) );
  AOI22X1 U2453 ( .A(phase[0]), .B(n761), .C(n259), .D(n618), .Y(n745) );
  NAND31X1 U2454 ( .C(n767), .A(n2345), .B(n762), .Y(n761) );
  NAND4X1 U2455 ( .A(n1097), .B(n1098), .C(n1099), .D(n1100), .Y(dpc[4]) );
  AOI22X1 U2456 ( .A(dpc_tab[34]), .B(n198), .C(dpc_tab[46]), .D(n200), .Y(
        n1097) );
  AOI22X1 U2457 ( .A(dpc_tab[10]), .B(n205), .C(dpc_tab[22]), .D(n206), .Y(
        n1099) );
  AOI22X1 U2458 ( .A(dpc_tab[28]), .B(n202), .C(dpc_tab[40]), .D(n204), .Y(
        n1098) );
  NAND4X1 U2459 ( .A(n1093), .B(n1094), .C(n1095), .D(n1096), .Y(dpc[5]) );
  AOI22X1 U2460 ( .A(dpc_tab[35]), .B(n521), .C(dpc_tab[47]), .D(n522), .Y(
        n1093) );
  AOI22X1 U2461 ( .A(dpc_tab[11]), .B(n1), .C(dpc_tab[23]), .D(n2), .Y(n1095)
         );
  AOI22X1 U2462 ( .A(dpc_tab[29]), .B(n519), .C(dpc_tab[41]), .D(n520), .Y(
        n1094) );
  NAND4X1 U2463 ( .A(n511), .B(n512), .C(n513), .D(n514), .Y(dpl[7]) );
  AOI22X1 U2464 ( .A(n197), .B(dpl_reg[47]), .C(n199), .D(dpl_reg[63]), .Y(
        n511) );
  AOI22X1 U2465 ( .A(n1), .B(dpl_reg[15]), .C(n2), .D(dpl_reg[31]), .Y(n513)
         );
  AOI22X1 U2466 ( .A(n201), .B(dpl_reg[39]), .C(n203), .D(dpl_reg[55]), .Y(
        n512) );
  OAI31XL U2467 ( .A(n304), .B(n303), .C(n2382), .D(phase[1]), .Y(n381) );
  INVX1 U2468 ( .A(n589), .Y(n304) );
  INVX1 U2469 ( .A(n587), .Y(n303) );
  NAND42X1 U2470 ( .C(n2159), .D(n286), .A(n1759), .B(n1760), .Y(n1650) );
  NAND3X1 U2471 ( .A(n1770), .B(intcall), .C(n1733), .Y(n1759) );
  INVX1 U2472 ( .A(n1758), .Y(n286) );
  AOI22X1 U2473 ( .A(phase[1]), .B(n1761), .C(phase[0]), .D(n1762), .Y(n1760)
         );
  AO222X1 U2474 ( .A(dph_current[3]), .B(n1247), .C(n1022), .D(temp[3]), .E(
        dptr_inc[11]), .F(n148), .Y(n871) );
  AO222X1 U2475 ( .A(dph_current[4]), .B(n1247), .C(n1022), .D(temp[4]), .E(
        dptr_inc[12]), .F(n148), .Y(n899) );
  AO222X1 U2476 ( .A(dph_current[5]), .B(n1247), .C(n1022), .D(temp[5]), .E(
        dptr_inc[13]), .F(n148), .Y(n904) );
  OR2X1 U2477 ( .A(n2480), .B(n610), .Y(n344) );
  NAND42X1 U2478 ( .C(n1739), .D(n2340), .A(phase[1]), .B(n2183), .Y(n1507) );
  OR3XL U2479 ( .A(instr[4]), .B(n2352), .C(n776), .Y(n668) );
  NAND32X1 U2480 ( .B(ramsfraddr[7]), .C(n2325), .A(n14), .Y(n1508) );
  OAI21X1 U2481 ( .B(dec_cop[3]), .C(dec_cop[4]), .A(accactv), .Y(n1075) );
  AOI222XL U2482 ( .A(dptr_inc[10]), .B(n148), .C(n1247), .D(dph_current[2]), 
        .E(n1022), .F(temp[2]), .Y(n678) );
  AOI22X1 U2483 ( .A(n2436), .B(n2476), .C(instr[4]), .D(n765), .Y(n1792) );
  NAND43X1 U2484 ( .B(n782), .C(n2116), .D(n2115), .A(n1652), .Y(n638) );
  OAI222XL U2485 ( .A(n1748), .B(n2340), .C(n2110), .D(n2385), .E(n610), .F(
        n2412), .Y(n2116) );
  OAI211X1 U2486 ( .C(n2479), .D(n2118), .A(n2119), .B(n2120), .Y(n2115) );
  AOI211X1 U2487 ( .C(n2121), .D(n980), .A(n777), .B(n1999), .Y(n2120) );
  NAND3X1 U2488 ( .A(n2048), .B(n2480), .C(n1766), .Y(n911) );
  AOI21X1 U2489 ( .B(n151), .C(dec_cop[1]), .A(n2241), .Y(n1074) );
  NAND2X1 U2490 ( .A(n1336), .B(n1337), .Y(n1102) );
  OAI21X1 U2491 ( .B(n791), .C(n810), .A(n1338), .Y(n1337) );
  NAND4X1 U2492 ( .A(n752), .B(n259), .C(n1015), .D(n105), .Y(n1338) );
  NOR2X1 U2493 ( .A(n2172), .B(n2477), .Y(n822) );
  NAND2X1 U2494 ( .A(n2479), .B(n2477), .Y(n610) );
  NAND4X1 U2495 ( .A(n1328), .B(n1329), .C(n1330), .D(n1331), .Y(dpc[2]) );
  AOI22X1 U2496 ( .A(dpc_tab[32]), .B(n198), .C(dpc_tab[44]), .D(n200), .Y(
        n1328) );
  AOI22X1 U2497 ( .A(dpc_tab[8]), .B(n53), .C(dpc_tab[20]), .D(n49), .Y(n1330)
         );
  AOI22X1 U2498 ( .A(dpc_tab[26]), .B(n202), .C(dpc_tab[38]), .D(n204), .Y(
        n1329) );
  OAI22X1 U2499 ( .A(n1786), .B(n2324), .C(n590), .D(n257), .Y(n1627) );
  NOR4XL U2500 ( .A(n1787), .B(n1788), .C(n2382), .D(n1789), .Y(n1786) );
  AO2222XL U2501 ( .A(n2189), .B(n2407), .C(n1014), .D(n1026), .E(n1737), .F(
        n2383), .G(n974), .H(n1791), .Y(n1787) );
  OAI22X1 U2502 ( .A(n2476), .B(n2342), .C(n1790), .D(n2357), .Y(n1788) );
  OAI22X1 U2503 ( .A(n2257), .B(n1151), .C(n2426), .D(n1152), .Y(
        dpl_current[7]) );
  AND4X1 U2504 ( .A(n1153), .B(n1154), .C(n1155), .D(n1156), .Y(n1152) );
  AOI22X1 U2505 ( .A(n1163), .B(dpl_reg[55]), .C(n1164), .D(dpl_reg[63]), .Y(
        n1153) );
  AOI22X1 U2506 ( .A(n1161), .B(dpl_reg[39]), .C(n1162), .D(dpl_reg[47]), .Y(
        n1154) );
  AND2XL U2507 ( .A(sfroe_r), .B(n262), .Y(sfroe) );
  AOI31X1 U2508 ( .A(n2479), .B(n753), .C(n758), .D(n964), .Y(n986) );
  NAND4X1 U2509 ( .A(n1332), .B(n1333), .C(n1334), .D(n1335), .Y(dpc[1]) );
  AOI22X1 U2510 ( .A(dpc_tab[31]), .B(n198), .C(dpc_tab[43]), .D(n200), .Y(
        n1332) );
  AOI22X1 U2511 ( .A(dpc_tab[25]), .B(n202), .C(dpc_tab[37]), .D(n204), .Y(
        n1333) );
  AOI22X1 U2512 ( .A(dpc_tab[7]), .B(n53), .C(dpc_tab[19]), .D(n49), .Y(n1334)
         );
  NOR3XL U2513 ( .A(n2347), .B(n2478), .C(n2388), .Y(n1754) );
  AOI22X1 U2514 ( .A(n609), .B(phase[3]), .C(n259), .D(n2253), .Y(n791) );
  NAND2X1 U2515 ( .A(dec_cop[2]), .B(accactv), .Y(n1066) );
  AOI221XL U2516 ( .A(n978), .B(n979), .C(n974), .D(n2476), .E(n1747), .Y(
        n1745) );
  OAI33XL U2517 ( .A(n2408), .B(n2476), .C(n2347), .D(n2436), .E(n1748), .F(
        n26), .Y(n1747) );
  AOI22X1 U2518 ( .A(dpc_tab[1]), .B(n207), .C(dpc_tab[13]), .D(n516), .Y(
        n1335) );
  AOI22X1 U2519 ( .A(dpc_tab[3]), .B(n20), .C(dpc_tab[15]), .D(n516), .Y(n1106) );
  AOI22X1 U2520 ( .A(dpc_tab[2]), .B(n20), .C(dpc_tab[14]), .D(n516), .Y(n1331) );
  AOI22X1 U2521 ( .A(n207), .B(dpl_reg[1]), .C(n18), .D(dpl_reg[17]), .Y(n546)
         );
  AOI22X1 U2522 ( .A(n515), .B(dph_reg[1]), .C(n18), .D(dph_reg[17]), .Y(n578)
         );
  AOI22X1 U2523 ( .A(n207), .B(dpl_reg[3]), .C(n18), .D(dpl_reg[19]), .Y(n538)
         );
  AOI22X1 U2524 ( .A(n20), .B(dph_reg[7]), .C(n516), .D(dph_reg[23]), .Y(n554)
         );
  NOR2X1 U2525 ( .A(n2347), .B(n2475), .Y(n974) );
  AOI22X1 U2526 ( .A(n1), .B(dpl_reg[9]), .C(n2), .D(dpl_reg[25]), .Y(n545) );
  AOI22X1 U2527 ( .A(n1), .B(dph_reg[9]), .C(n2), .D(dph_reg[25]), .Y(n577) );
  AOI22X1 U2528 ( .A(n1), .B(dpl_reg[11]), .C(n2), .D(dpl_reg[27]), .Y(n537)
         );
  AOI22X1 U2529 ( .A(n53), .B(dph_reg[15]), .C(n49), .D(dph_reg[31]), .Y(n553)
         );
  AOI22X1 U2530 ( .A(n201), .B(dpl_reg[33]), .C(n203), .D(dpl_reg[49]), .Y(
        n544) );
  AOI22X1 U2531 ( .A(n519), .B(dpl_reg[35]), .C(n520), .D(dpl_reg[51]), .Y(
        n536) );
  AOI22X1 U2532 ( .A(n202), .B(dph_reg[39]), .C(n204), .D(dph_reg[55]), .Y(
        n552) );
  NOR2X1 U2533 ( .A(n2404), .B(n2478), .Y(n1733) );
  NAND3X1 U2534 ( .A(ramsfraddr[2]), .B(n2444), .C(ramsfraddr[1]), .Y(n856) );
  OAI211X1 U2535 ( .C(n2403), .D(n2340), .A(n1768), .B(n1769), .Y(n1761) );
  INVX1 U2536 ( .A(n1684), .Y(n2403) );
  AOI32X1 U2537 ( .A(n1770), .B(interrupt), .C(n1733), .D(n1690), .E(n1771), 
        .Y(n1769) );
  ENOX1 U2538 ( .A(n2343), .B(n102), .C(n2171), .D(n2144), .Y(n1771) );
  AOI32X1 U2539 ( .A(n2475), .B(n2387), .C(n819), .D(n1014), .E(n2430), .Y(
        n1790) );
  AOI22X1 U2540 ( .A(n1157), .B(dpl_reg[7]), .C(n1158), .D(dpl_reg[15]), .Y(
        n1156) );
  GEN2XL U2541 ( .D(n1730), .E(n296), .C(n2361), .B(n1732), .A(n2182), .Y(n400) );
  AOI32X1 U2542 ( .A(n1733), .B(n758), .C(phase[3]), .D(phase[2]), .E(n1734), 
        .Y(n1732) );
  NAND41X1 U2543 ( .D(n778), .A(n2375), .B(n1021), .C(n1735), .Y(n1734) );
  AOI31X1 U2544 ( .A(n776), .B(instr[2]), .C(n2161), .D(n809), .Y(n1735) );
  OAI21X1 U2545 ( .B(n1745), .C(n44), .A(n1746), .Y(n1744) );
  NAND4X1 U2546 ( .A(n765), .B(n2379), .C(n44), .D(n25), .Y(n1746) );
  NAND4X1 U2547 ( .A(n1103), .B(n1104), .C(n1105), .D(n1106), .Y(dpc[3]) );
  AOI22X1 U2548 ( .A(dpc_tab[33]), .B(n197), .C(dpc_tab[45]), .D(n199), .Y(
        n1103) );
  AOI22X1 U2549 ( .A(dpc_tab[9]), .B(n53), .C(dpc_tab[21]), .D(n49), .Y(n1105)
         );
  AOI22X1 U2550 ( .A(dpc_tab[27]), .B(n201), .C(dpc_tab[39]), .D(n203), .Y(
        n1104) );
  OAI211X1 U2551 ( .C(n1763), .D(n51), .A(n1764), .B(n1765), .Y(n1762) );
  AOI22X1 U2552 ( .A(n766), .B(n752), .C(n1681), .D(instr[6]), .Y(n1765) );
  AOI31X1 U2553 ( .A(n1690), .B(n1014), .C(n1766), .D(n175), .Y(n1764) );
  INVX1 U2554 ( .A(temp2_comb[6]), .Y(n2283) );
  INVX1 U2555 ( .A(temp2_comb[4]), .Y(n2332) );
  INVX1 U2556 ( .A(temp2_comb[5]), .Y(n2315) );
  AO222X1 U2557 ( .A(dph_current[6]), .B(n1247), .C(n1022), .D(temp[6]), .E(
        dptr_inc[14]), .F(n148), .Y(n906) );
  INVX1 U2558 ( .A(ramdatao[0]), .Y(n2414) );
  OAI22X1 U2559 ( .A(n2414), .B(n1248), .C(n2425), .D(n1339), .Y(
        dph_current[0]) );
  AND4X1 U2560 ( .A(n1340), .B(n1341), .C(n1342), .D(n1343), .Y(n1339) );
  AOI22X1 U2561 ( .A(n1163), .B(dph_reg[48]), .C(n1164), .D(dph_reg[56]), .Y(
        n1340) );
  AOI22X1 U2562 ( .A(n1161), .B(dph_reg[32]), .C(n1162), .D(dph_reg[40]), .Y(
        n1341) );
  AND2X1 U2563 ( .A(dec_cop[5]), .B(n151), .Y(n1067) );
  INVX1 U2564 ( .A(phase[2]), .Y(n2275) );
  INVX1 U2565 ( .A(n2481), .Y(n612) );
  AOI32X1 U2566 ( .A(n781), .B(n758), .C(instr[1]), .D(n982), .E(n1681), .Y(
        n1730) );
  OAI21X1 U2567 ( .B(n2431), .C(n2095), .A(n2096), .Y(n755) );
  GEN2XL U2568 ( .D(n2388), .E(n2384), .C(instr[7]), .B(n2171), .A(n2099), .Y(
        n2095) );
  GEN2XL U2569 ( .D(instr[0]), .E(n56), .C(n2097), .B(n1785), .A(n2098), .Y(
        n2096) );
  AOI21X1 U2570 ( .B(instr[7]), .C(instr[4]), .A(n808), .Y(n2099) );
  MUX2AXL U2571 ( .D0(n2459), .D1(temp[1]), .S(n1150), .Y(n181) );
  AOI21X1 U2572 ( .B(n2170), .C(n2475), .A(n1781), .Y(n2110) );
  AOI22AXL U2573 ( .A(n2106), .B(n2107), .D(n2108), .C(n2071), .Y(n2105) );
  OAI222XL U2574 ( .A(interrupt), .B(n2407), .C(n1766), .D(n2474), .E(n2480), 
        .F(n2402), .Y(n2107) );
  OAI21X1 U2575 ( .B(n2388), .C(n2409), .A(n2109), .Y(n2106) );
  AOI33X1 U2576 ( .A(n1683), .B(n2417), .C(n1682), .D(n2189), .E(n2474), .F(
        n2476), .Y(n2109) );
  NOR3XL U2577 ( .A(n285), .B(instr[4]), .C(n2410), .Y(n804) );
  AOI22X1 U2578 ( .A(n1157), .B(dph_reg[0]), .C(n1158), .D(dph_reg[8]), .Y(
        n1343) );
  AOI32X1 U2579 ( .A(n2479), .B(n808), .C(n1780), .D(n980), .E(n2171), .Y(
        n2098) );
  AOI22X1 U2580 ( .A(n1159), .B(dpl_reg[23]), .C(n1160), .D(dpl_reg[31]), .Y(
        n1155) );
  NOR2X1 U2581 ( .A(n2172), .B(n2474), .Y(n978) );
  AOI22X1 U2582 ( .A(n2157), .B(instr[5]), .C(n1336), .D(n1777), .Y(n2118) );
  NOR2X1 U2583 ( .A(n2475), .B(instr[5]), .Y(n1780) );
  INVX1 U2584 ( .A(c), .Y(n2455) );
  INVX1 U2585 ( .A(temp[3]), .Y(n2264) );
  INVX1 U2586 ( .A(temp2_comb[0]), .Y(n703) );
  INVX1 U2587 ( .A(temp[4]), .Y(n2265) );
  NOR2X1 U2588 ( .A(n2478), .B(n2347), .Y(n2121) );
  INVX1 U2589 ( .A(dec_cop[6]), .Y(n2251) );
  NAND21X1 U2590 ( .B(N343), .A(N344), .Y(n2274) );
  NAND2X1 U2591 ( .A(N343), .B(N344), .Y(n2272) );
  NAND21X1 U2592 ( .B(N344), .A(N343), .Y(n488) );
  OR2X1 U2593 ( .A(N343), .B(N344), .Y(n2273) );
  AO222X1 U2594 ( .A(n1247), .B(dph_current[7]), .C(n1022), .D(temp[7]), .E(
        dptr_inc[15]), .F(n148), .Y(n908) );
  OAI22X1 U2595 ( .A(n2257), .B(n1248), .C(n2425), .D(n1249), .Y(
        dph_current[7]) );
  AND4X1 U2596 ( .A(n1250), .B(n1251), .C(n1252), .D(n1253), .Y(n1249) );
  AOI21BBXL U2597 ( .B(n2101), .C(n2102), .A(n2478), .Y(n751) );
  XNOR2XL U2598 ( .A(n2417), .B(n2408), .Y(n2101) );
  XNOR2XL U2599 ( .A(n2408), .B(n2480), .Y(n2102) );
  OAI22X1 U2600 ( .A(n2415), .B(n1248), .C(n2425), .D(n1315), .Y(
        dph_current[1]) );
  AND4X1 U2601 ( .A(n1316), .B(n1317), .C(n1318), .D(n1319), .Y(n1315) );
  AOI22X1 U2602 ( .A(n86), .B(dph_reg[49]), .C(n104), .D(dph_reg[57]), .Y(
        n1316) );
  AOI22X1 U2603 ( .A(n123), .B(dph_reg[33]), .C(n147), .D(dph_reg[41]), .Y(
        n1317) );
  INVX1 U2604 ( .A(temp[1]), .Y(n2269) );
  OAI32X1 U2605 ( .A(n813), .B(n591), .C(n804), .D(n803), .E(n2254), .Y(n812)
         );
  INVX1 U2606 ( .A(n813), .Y(n2254) );
  OAI22X1 U2607 ( .A(n814), .B(n815), .C(n816), .D(n817), .Y(n813) );
  OAI21X1 U2608 ( .B(n2335), .C(n2273), .A(N345), .Y(n817) );
  INVX1 U2609 ( .A(ramsfraddr[7]), .Y(n2173) );
  AOI22X1 U2610 ( .A(n103), .B(dph_reg[1]), .C(n85), .D(dph_reg[9]), .Y(n1319)
         );
  AOI22X1 U2611 ( .A(n1159), .B(dph_reg[16]), .C(n1160), .D(dph_reg[24]), .Y(
        n1342) );
  AOI22X1 U2612 ( .A(n146), .B(dph_reg[17]), .C(n122), .D(dph_reg[25]), .Y(
        n1318) );
  INVX1 U2613 ( .A(n1741), .Y(n2183) );
  AOI221XL U2614 ( .A(instr[7]), .B(n821), .C(n2377), .D(instr[6]), .E(n1742), 
        .Y(n1741) );
  OAI211X1 U2615 ( .C(instr[7]), .D(instr[5]), .A(n2110), .B(n2411), .Y(n2103)
         );
  INVX1 U2616 ( .A(temp[7]), .Y(n2271) );
  NOR2X1 U2617 ( .A(n105), .B(instr[5]), .Y(n821) );
  INVX1 U2618 ( .A(temp[0]), .Y(n2268) );
  INVX1 U2619 ( .A(temp[5]), .Y(n2266) );
  INVX1 U2620 ( .A(memaddr[1]), .Y(n2437) );
  INVX1 U2621 ( .A(memaddr[2]), .Y(n2420) );
  NAND21X1 U2622 ( .B(n344), .A(c), .Y(n345) );
  MUX2X1 U2623 ( .D0(n2146), .D1(n2145), .S(pc_o[1]), .Y(n414) );
  OAI22X1 U2624 ( .A(n2435), .B(n1248), .C(n2425), .D(n1293), .Y(
        dph_current[3]) );
  AND4X1 U2625 ( .A(n1294), .B(n1295), .C(n1296), .D(n1297), .Y(n1293) );
  AOI22X1 U2626 ( .A(n86), .B(dph_reg[51]), .C(n104), .D(dph_reg[59]), .Y(
        n1294) );
  AOI22X1 U2627 ( .A(n123), .B(dph_reg[35]), .C(n147), .D(dph_reg[43]), .Y(
        n1295) );
  OAI22X1 U2628 ( .A(n2316), .B(n1248), .C(n2425), .D(n1304), .Y(
        dph_current[2]) );
  AND4X1 U2629 ( .A(n1305), .B(n1306), .C(n1307), .D(n1308), .Y(n1304) );
  AOI22X1 U2630 ( .A(n86), .B(dph_reg[50]), .C(n104), .D(dph_reg[58]), .Y(
        n1305) );
  AOI22X1 U2631 ( .A(n123), .B(dph_reg[34]), .C(n147), .D(dph_reg[42]), .Y(
        n1306) );
  AOI21X1 U2632 ( .B(n1976), .C(instr[4]), .A(israccess), .Y(n182) );
  OAI21X1 U2633 ( .B(instr[4]), .C(n2168), .A(n102), .Y(n759) );
  AOI22X1 U2634 ( .A(n103), .B(dph_reg[2]), .C(n85), .D(dph_reg[10]), .Y(n1308) );
  AOI22X1 U2635 ( .A(n103), .B(dph_reg[3]), .C(n85), .D(dph_reg[11]), .Y(n1297) );
  AOI22X1 U2636 ( .A(n146), .B(dph_reg[18]), .C(n122), .D(dph_reg[26]), .Y(
        n1307) );
  AOI22X1 U2637 ( .A(n146), .B(dph_reg[19]), .C(n122), .D(dph_reg[27]), .Y(
        n1296) );
  INVX1 U2638 ( .A(temp[2]), .Y(n2270) );
  INVX1 U2639 ( .A(N345), .Y(n2167) );
  INVX1 U2640 ( .A(temp[6]), .Y(n2267) );
  OAI22X1 U2641 ( .A(n2169), .B(n1248), .C(n2425), .D(n1282), .Y(
        dph_current[4]) );
  AND4X1 U2642 ( .A(n1283), .B(n1284), .C(n1285), .D(n1286), .Y(n1282) );
  AOI22X1 U2643 ( .A(n86), .B(dph_reg[52]), .C(n104), .D(dph_reg[60]), .Y(
        n1283) );
  AOI22X1 U2644 ( .A(n123), .B(dph_reg[36]), .C(n147), .D(dph_reg[44]), .Y(
        n1284) );
  OAI22X1 U2645 ( .A(n2256), .B(n1248), .C(n2425), .D(n1272), .Y(
        dph_current[5]) );
  AND4X1 U2646 ( .A(n1273), .B(n1274), .C(n1275), .D(n1276), .Y(n1272) );
  AOI22X1 U2648 ( .A(n86), .B(dph_reg[53]), .C(n104), .D(dph_reg[61]), .Y(
        n1273) );
  AOI22X1 U2649 ( .A(n123), .B(dph_reg[37]), .C(n147), .D(dph_reg[45]), .Y(
        n1274) );
  INVX1 U2650 ( .A(ramdatao[5]), .Y(n2256) );
  NAND2X1 U2651 ( .A(n777), .B(phase[0]), .Y(n696) );
  INVX1 U2652 ( .A(ramdatao[6]), .Y(n2255) );
  INVX1 U2653 ( .A(phase[3]), .Y(n2166) );
  AOI22X1 U2654 ( .A(n103), .B(dph_reg[4]), .C(n85), .D(dph_reg[12]), .Y(n1286) );
  AOI22X1 U2655 ( .A(n103), .B(dph_reg[5]), .C(n85), .D(dph_reg[13]), .Y(n1276) );
  AOI22X1 U2656 ( .A(n146), .B(dph_reg[20]), .C(n122), .D(dph_reg[28]), .Y(
        n1285) );
  AOI22X1 U2657 ( .A(n146), .B(dph_reg[21]), .C(n122), .D(dph_reg[29]), .Y(
        n1275) );
  INVX1 U2658 ( .A(memaddr[9]), .Y(n2423) );
  MUX2X1 U2659 ( .D0(ramsfraddr[7]), .D1(n1651), .S(n261), .Y(
        ramsfraddr_comb[7]) );
  NAND32X1 U2660 ( .B(p2sel), .C(n1434), .A(n833), .Y(n881) );
  OR2X1 U2661 ( .A(state[1]), .B(state[2]), .Y(n1677) );
  NAND32X1 U2662 ( .B(p2sel), .C(n690), .A(n833), .Y(n870) );
  NAND21X1 U2663 ( .B(state[0]), .A(n1701), .Y(n1545) );
  INVX1 U2664 ( .A(memaddr[4]), .Y(n2371) );
  AO2222XL U2665 ( .A(n1359), .B(b[2]), .C(n1360), .D(multemp2[4]), .E(n1361), 
        .F(n2366), .G(n2429), .H(n240), .Y(N12479) );
  INVX1 U2666 ( .A(n845), .Y(n2366) );
  AO2222XL U2667 ( .A(n1359), .B(b[3]), .C(n1360), .D(multemp2[5]), .E(n1361), 
        .F(n2365), .G(n2429), .H(n237), .Y(N12480) );
  INVX1 U2668 ( .A(n844), .Y(n2365) );
  OAI22X1 U2669 ( .A(n2255), .B(n1248), .C(n2425), .D(n1258), .Y(
        dph_current[6]) );
  AND4X1 U2670 ( .A(n1259), .B(n1260), .C(n1261), .D(n1262), .Y(n1258) );
  AOI22X1 U2671 ( .A(n86), .B(dph_reg[54]), .C(n104), .D(dph_reg[62]), .Y(
        n1259) );
  AOI22X1 U2672 ( .A(n123), .B(dph_reg[38]), .C(n147), .D(dph_reg[46]), .Y(
        n1260) );
  OAI22XL U2673 ( .A(n987), .B(n1639), .C(n1002), .D(n272), .Y(N12716) );
  AOI221XL U2674 ( .A(n993), .B(memaddr[10]), .C(ramdatai[2]), .D(n994), .E(
        n1003), .Y(n1002) );
  OAI22X1 U2675 ( .A(n2279), .B(n2199), .C(n437), .D(n2280), .Y(n1003) );
  OAI22XL U2676 ( .A(n987), .B(n1646), .C(n992), .D(n271), .Y(N12720) );
  AOI221XL U2677 ( .A(n993), .B(pc_o[14]), .C(ramdatai[6]), .D(n994), .E(n995), 
        .Y(n992) );
  OAI22X1 U2678 ( .A(n2279), .B(n2208), .C(n2252), .D(n2280), .Y(n995) );
  OAI22XL U2679 ( .A(n987), .B(n1649), .C(n1000), .D(n272), .Y(N12717) );
  AOI221XL U2680 ( .A(n993), .B(pc_o[11]), .C(ramdatai[3]), .D(n994), .E(n1001), .Y(n1000) );
  OAI22X1 U2681 ( .A(n2279), .B(n2195), .C(n2259), .D(n2280), .Y(n1001) );
  AOI22X1 U2682 ( .A(n103), .B(dph_reg[6]), .C(n85), .D(dph_reg[14]), .Y(n1262) );
  AOI22X1 U2683 ( .A(n146), .B(dph_reg[22]), .C(n122), .D(dph_reg[30]), .Y(
        n1261) );
  INVX1 U2684 ( .A(phase[4]), .Y(n2165) );
  AND2XL U2685 ( .A(phase0_ff), .B(n262), .Y(newinstr) );
  AO2222XL U2686 ( .A(n2429), .B(n248), .C(n1359), .D(b[0]), .E(n1360), .F(
        multemp2[2]), .G(n1361), .H(n2368), .Y(N12477) );
  INVX1 U2687 ( .A(n847), .Y(n2368) );
  AO2222XL U2688 ( .A(n2429), .B(n244), .C(n1359), .D(b[1]), .E(n1360), .F(
        multemp2[3]), .G(n1361), .H(n2367), .Y(N12478) );
  INVX1 U2689 ( .A(n846), .Y(n2367) );
  AO2222XL U2690 ( .A(n2429), .B(n234), .C(n1359), .D(b[4]), .E(n1360), .F(
        multemp2[6]), .G(n1361), .H(n2364), .Y(N12481) );
  INVX1 U2691 ( .A(n843), .Y(n2364) );
  AO2222XL U2692 ( .A(n2429), .B(n228), .C(n1359), .D(b[6]), .E(n1360), .F(
        multemp2[8]), .G(n1361), .H(n2362), .Y(N12483) );
  INVX1 U2693 ( .A(n840), .Y(n2362) );
  AO2222XL U2694 ( .A(n1359), .B(b[5]), .C(n1360), .D(multemp2[7]), .E(n2429), 
        .F(n231), .G(n1361), .H(n2363), .Y(N12482) );
  INVX1 U2695 ( .A(n842), .Y(n2363) );
  NAND3X1 U2696 ( .A(ramsfraddr[3]), .B(ramsfraddr[4]), .C(n858), .Y(n863) );
  NAND3X1 U2697 ( .A(ramsfraddr[3]), .B(n2447), .C(n858), .Y(n860) );
  INVX1 U2698 ( .A(ramdatao[7]), .Y(n2257) );
  OAI221X1 U2699 ( .A(n834), .B(n1350), .C(n690), .D(n2207), .E(n275), .Y(
        N12485) );
  OAI221X1 U2700 ( .A(n2245), .B(n1350), .C(n690), .D(n2201), .E(n275), .Y(
        N12491) );
  INVX1 U2701 ( .A(p2[6]), .Y(n2245) );
  OAI221X1 U2702 ( .A(n837), .B(n1350), .C(n2206), .D(n690), .E(n275), .Y(
        N12486) );
  OAI221X1 U2703 ( .A(n867), .B(n1350), .C(n2205), .D(n690), .E(n275), .Y(
        N12487) );
  OAI221X1 U2704 ( .A(n2240), .B(n1350), .C(n690), .D(n2203), .E(n274), .Y(
        N12489) );
  INVX1 U2705 ( .A(p2[4]), .Y(n2240) );
  OAI221X1 U2706 ( .A(n2238), .B(n1350), .C(n690), .D(n2200), .E(n274), .Y(
        N12492) );
  INVX1 U2707 ( .A(p2[7]), .Y(n2238) );
  OAI221X1 U2708 ( .A(n2246), .B(n1350), .C(n2204), .D(n690), .E(n274), .Y(
        N12488) );
  INVX1 U2709 ( .A(p2[3]), .Y(n2246) );
  OAI221X1 U2710 ( .A(n2239), .B(n1350), .C(n2202), .D(n690), .E(n274), .Y(
        N12490) );
  INVX1 U2711 ( .A(p2[5]), .Y(n2239) );
  OAI22X1 U2712 ( .A(n2200), .B(n1353), .C(n1354), .D(n1355), .Y(N12484) );
  AOI21X1 U2713 ( .B(b[7]), .C(n1356), .A(n1357), .Y(n1354) );
  OAI33XL U2714 ( .A(n2212), .B(n2306), .C(n2213), .D(n2211), .E(n1358), .F(
        n1047), .Y(n1357) );
  AOI22X1 U2715 ( .A(N13353), .B(n189), .C(N13352), .D(n2190), .Y(n1358) );
  OAI22X1 U2716 ( .A(n943), .B(n216), .C(n918), .D(n2198), .Y(N12725) );
  AOI211X1 U2717 ( .C(n915), .D(ramdatai[2]), .A(n944), .B(n945), .Y(n943) );
  AO2222XL U2718 ( .A(n921), .B(temp[2]), .C(n919), .D(pc_i[10]), .E(n920), 
        .F(temp2_comb[2]), .G(n2314), .H(pc_o[2]), .Y(n944) );
  OAI22X1 U2719 ( .A(n946), .B(n2323), .C(n437), .D(n942), .Y(n945) );
  AOI22X1 U2720 ( .A(n103), .B(dph_reg[7]), .C(n85), .D(dph_reg[15]), .Y(n1253) );
  AOI22X1 U2721 ( .A(n146), .B(dph_reg[23]), .C(n122), .D(dph_reg[31]), .Y(
        n1252) );
  AOI22X1 U2722 ( .A(n86), .B(dph_reg[55]), .C(n104), .D(dph_reg[63]), .Y(
        n1250) );
  AOI22X1 U2723 ( .A(n123), .B(dph_reg[39]), .C(n147), .D(dph_reg[47]), .Y(
        n1251) );
  ENOX1 U2724 ( .A(n1027), .B(n2201), .C(n1028), .D(n1048), .Y(N12706) );
  OAI22BX1 U2725 ( .B(ac), .A(n1049), .D(n1035), .C(n1050), .Y(n1048) );
  AND3X1 U2726 ( .A(n1039), .B(n1034), .C(n1051), .Y(n1049) );
  AOI32X1 U2727 ( .A(n2460), .B(n2453), .C(N11555), .D(dec_accop[10]), .E(
        n2399), .Y(n1050) );
  ENOX1 U2728 ( .A(n485), .B(n2206), .C(f1), .D(n485), .Y(n1883) );
  ENOX1 U2729 ( .A(n486), .B(n2205), .C(gf0), .D(n486), .Y(n1881) );
  NOR2X1 U2730 ( .A(n269), .B(n487), .Y(n486) );
  ENOX1 U2731 ( .A(n485), .B(n2202), .C(f0), .D(n485), .Y(n1882) );
  NAND2X1 U2732 ( .A(n1112), .B(dps[2]), .Y(n1108) );
  INVX1 U2733 ( .A(stop_r), .Y(n2164) );
  NOR32XL U2734 ( .B(n211), .C(n792), .A(n2070), .Y(N10566) );
  NAND3X1 U2735 ( .A(n808), .B(instr[0]), .C(n1742), .Y(n2070) );
  OA21X1 U2736 ( .B(n1618), .C(n1617), .A(n215), .Y(N10562) );
  AO21X1 U2737 ( .B(n2084), .C(n259), .A(n2085), .Y(n1618) );
  OAI21BBX1 U2738 ( .A(n2083), .B(n620), .C(n2073), .Y(n1617) );
  AOI31X1 U2739 ( .A(n255), .B(n2275), .C(n252), .D(n2348), .Y(n2085) );
  NOR32XL U2740 ( .B(n212), .C(n254), .A(newinstrlock), .Y(N689) );
  OAI21X1 U2741 ( .B(n850), .C(n1671), .A(n274), .Y(N13324) );
  NOR2X1 U2742 ( .A(n849), .B(finishmul), .Y(n850) );
  AND2X1 U2743 ( .A(state[2]), .B(n214), .Y(N590) );
  AND2X1 U2744 ( .A(state[1]), .B(n214), .Y(N589) );
  INVX1 U2745 ( .A(n1513), .Y(n1757) );
  NAND32X1 U2746 ( .B(instr[5]), .C(n219), .A(n749), .Y(n1513) );
  AOI21X1 U2747 ( .B(n1584), .C(n1583), .A(n1671), .Y(N12726) );
  AOI221XL U2748 ( .A(n2314), .B(pc_o[3]), .C(n915), .D(ramdatai[3]), .E(n1582), .Y(n1584) );
  AOI221XL U2749 ( .A(n919), .B(pc_i[11]), .C(temp2_comb[3]), .D(n920), .E(
        n940), .Y(n1583) );
  OAI21BBX1 U2750 ( .A(intvect[0]), .B(n2145), .C(n937), .Y(n1582) );
  AOI21X1 U2751 ( .B(n1599), .C(n1598), .A(n1671), .Y(N12727) );
  AOI221XL U2752 ( .A(n2314), .B(pc_o[4]), .C(n915), .D(ramdatai[4]), .E(n1597), .Y(n1599) );
  AOI221XL U2753 ( .A(pc_i[12]), .B(n919), .C(temp2_comb[4]), .D(n920), .E(
        n935), .Y(n1598) );
  OAI21BBX1 U2754 ( .A(intvect[1]), .B(n2145), .C(n932), .Y(n1597) );
  AOI21X1 U2755 ( .B(n1626), .C(n1625), .A(n1671), .Y(N12728) );
  AOI221XL U2756 ( .A(pc_i[13]), .B(n919), .C(temp2_comb[5]), .D(n920), .E(
        n930), .Y(n1625) );
  AOI221XL U2757 ( .A(n2314), .B(pc_o[5]), .C(n915), .D(ramdatai[5]), .E(n1624), .Y(n1626) );
  OAI22X1 U2758 ( .A(n931), .B(n2323), .C(n730), .D(n918), .Y(n930) );
  AOI21X1 U2759 ( .B(n1637), .C(n1636), .A(n221), .Y(N12729) );
  AOI221XL U2760 ( .A(pc_i[14]), .B(n919), .C(temp2_comb[6]), .D(n920), .E(
        n925), .Y(n1636) );
  AOI221XL U2761 ( .A(n2314), .B(pc_o[6]), .C(n915), .D(ramdatai[6]), .E(n1635), .Y(n1637) );
  OAI22X1 U2762 ( .A(n926), .B(n2323), .C(n2208), .D(n918), .Y(n925) );
  AOI21X1 U2763 ( .B(n1658), .C(n1656), .A(n218), .Y(N12730) );
  AOI221XL U2764 ( .A(n919), .B(pc_i[15]), .C(n920), .D(temp2_comb[7]), .E(
        n916), .Y(n1656) );
  AOI221XL U2765 ( .A(n2314), .B(pc_o[7]), .C(n915), .D(ramdatai[7]), .E(n1654), .Y(n1658) );
  OAI22X1 U2766 ( .A(n917), .B(n2323), .C(n2209), .D(n918), .Y(n916) );
  INVX1 U2767 ( .A(idle_r), .Y(n2163) );
  INVX1 U2768 ( .A(memaddr[8]), .Y(n2422) );
  AOI21X1 U2769 ( .B(n2397), .C(n872), .A(n873), .Y(N12976) );
  NAND2X1 U2770 ( .A(waitcnt_0_), .B(waitcnt_1_), .Y(n872) );
  NOR2X1 U2771 ( .A(waitcnt_0_), .B(n873), .Y(N12974) );
  NAND43X1 U2772 ( .B(n785), .C(n750), .D(n2445), .A(n1351), .Y(n690) );
  INVX1 U2773 ( .A(n859), .Y(n785) );
  NOR2X1 U2774 ( .A(ramsfraddr[6]), .B(n851), .Y(n1351) );
  AO21X1 U2775 ( .B(d_hold), .C(n656), .A(cpu_resume_fff), .Y(n1521) );
  INVX1 U2776 ( .A(cpu_hold), .Y(n656) );
  INVX1 U2777 ( .A(memaddr[11]), .Y(n2418) );
  AOI22X1 U2778 ( .A(acc[6]), .B(N13353), .C(N13345), .D(n2190), .Y(n847) );
  OAI21BBX1 U2779 ( .A(intvect[3]), .B(n2145), .C(n922), .Y(n1635) );
  AOI22X1 U2780 ( .A(n921), .B(temp[6]), .C(n2326), .D(n831), .Y(n922) );
  OAI21BBX1 U2781 ( .A(intvect[2]), .B(n2145), .C(n927), .Y(n1624) );
  AOI22X1 U2782 ( .A(n921), .B(temp[5]), .C(n2326), .D(n830), .Y(n927) );
  OAI21BBX1 U2783 ( .A(intvect[4]), .B(n2145), .C(n912), .Y(n1654) );
  AOI22X1 U2784 ( .A(n921), .B(temp[7]), .C(n2326), .D(n832), .Y(n912) );
  INVX1 U2785 ( .A(temp2_comb[7]), .Y(n746) );
  AOI32X1 U2786 ( .A(n1033), .B(n1034), .C(n1035), .D(ov), .E(n1036), .Y(n1032) );
  NAND42X1 U2787 ( .C(n1037), .D(n1038), .A(n1039), .B(n1034), .Y(n1036) );
  XOR2X1 U2788 ( .A(n1040), .B(n1041), .Y(n1033) );
  AOI21BBXL U2789 ( .B(N345), .C(n2139), .A(n1411), .Y(n183) );
  AOI22X1 U2790 ( .A(n921), .B(temp[4]), .C(n2326), .D(n829), .Y(n932) );
  MUX2AXL U2791 ( .D0(n126), .D1(n2264), .S(n1150), .Y(n1903) );
  AOI221X1 U2792 ( .A(n1179), .B(n55), .C(pc_i[4]), .D(n1139), .E(n1188), .Y(
        n1119) );
  AO222X1 U2793 ( .A(n1138), .B(n1189), .C(pc_o[4]), .D(n1190), .E(n50), .F(
        n1181), .Y(n1188) );
  OAI221X1 U2794 ( .A(n36), .B(n1146), .C(n1191), .D(n1144), .E(n1192), .Y(
        n1190) );
  AOI221X1 U2795 ( .A(n1165), .B(n71), .C(pc_i[6]), .D(n1139), .E(n1166), .Y(
        n1118) );
  AO222X1 U2796 ( .A(n1145), .B(n2232), .C(pc_o[6]), .D(n1167), .E(n1143), .F(
        n2231), .Y(n1166) );
  OAI221X1 U2797 ( .A(n29), .B(n1146), .C(n1168), .D(n1144), .E(n1169), .Y(
        n1167) );
  AOI221X1 U2798 ( .A(n50), .B(n1268), .C(pc_i[11]), .D(n1139), .E(n2227), .Y(
        n1237) );
  INVX1 U2799 ( .A(n1287), .Y(n2227) );
  AOI221XL U2800 ( .A(n1280), .B(n2232), .C(pc_o[11]), .D(n1288), .E(n1289), 
        .Y(n1287) );
  NOR4XL U2801 ( .A(pc_o[11]), .B(n42), .C(n2235), .D(n1281), .Y(n1289) );
  OAI211X1 U2802 ( .C(pc_o[10]), .D(n2235), .A(n1290), .B(n1291), .Y(n1288) );
  AOI22X1 U2803 ( .A(n2232), .B(n1292), .C(n2231), .D(pc_o[10]), .Y(n1291) );
  OAI211X1 U2804 ( .C(pc_o[8]), .D(n2235), .A(n1312), .B(n1313), .Y(n1310) );
  AOI22X1 U2805 ( .A(n2232), .B(n1314), .C(n2231), .D(pc_o[8]), .Y(n1313) );
  AOI221X1 U2806 ( .A(n50), .B(n1303), .C(pc_i[9]), .D(n1139), .E(n2229), .Y(
        n1238) );
  INVX1 U2807 ( .A(n1309), .Y(n2229) );
  AOI221XL U2808 ( .A(n1301), .B(n2232), .C(pc_o[9]), .D(n1310), .E(n1311), 
        .Y(n1309) );
  NOR4XL U2809 ( .A(pc_o[9]), .B(n2422), .C(n2235), .D(n1302), .Y(n1311) );
  NOR2X1 U2810 ( .A(n2448), .B(n2462), .Y(N14339) );
  NOR2X1 U2811 ( .A(n2448), .B(n2461), .Y(N14340) );
  NOR2X1 U2812 ( .A(n2448), .B(n2456), .Y(N14341) );
  NOR2X1 U2813 ( .A(n2448), .B(n2457), .Y(N14342) );
  NOR2X1 U2814 ( .A(n2448), .B(n2465), .Y(N14338) );
  NOR2X1 U2815 ( .A(n2448), .B(n2442), .Y(N14343) );
  OA222X1 U2816 ( .A(n1241), .B(n15), .C(pc_o[15]), .D(n1242), .E(n2284), .F(
        n2234), .Y(n1235) );
  INVX1 U2817 ( .A(pc_i[15]), .Y(n2284) );
  INVX1 U2818 ( .A(n1139), .Y(n2234) );
  AOI32X1 U2819 ( .A(n71), .B(pc_o[14]), .C(n1243), .D(n1244), .E(n38), .Y(
        n1242) );
  MUX2AXL U2820 ( .D0(n2335), .D1(temp[4]), .S(n1150), .Y(n1517) );
  MUX2AXL U2821 ( .D0(n2334), .D1(temp[5]), .S(n1150), .Y(n1478) );
  AOI221X1 U2822 ( .A(n1137), .B(n71), .C(pc_i[7]), .D(n1139), .E(n1140), .Y(
        n1116) );
  AO222X1 U2823 ( .A(n2286), .B(n50), .C(pc_o[7]), .D(n1141), .E(n1142), .F(
        n2232), .Y(n1140) );
  INVX1 U2824 ( .A(n1147), .Y(n2286) );
  OAI221X1 U2825 ( .A(n1143), .B(n1144), .C(n1145), .D(n1146), .E(n2233), .Y(
        n1141) );
  AOI222XL U2826 ( .A(n1245), .B(pc_o[14]), .C(n38), .D(n1254), .E(pc_i[14]), 
        .F(n1139), .Y(n1236) );
  AO21X1 U2827 ( .B(n1243), .C(n1138), .A(n1244), .Y(n1254) );
  INVX1 U2828 ( .A(n1198), .Y(n2223) );
  OAI211X1 U2829 ( .C(n1199), .D(n2235), .A(n1200), .B(n1201), .Y(n1198) );
  AOI22X1 U2830 ( .A(n50), .B(n1191), .C(n93), .D(pc_i[3]), .Y(n1201) );
  AOI32X1 U2831 ( .A(n2421), .B(n36), .C(n2232), .D(pc_o[3]), .E(n1202), .Y(
        n1200) );
  INVX1 U2832 ( .A(n1263), .Y(n2224) );
  OAI211X1 U2833 ( .C(n1264), .D(n31), .A(n1265), .B(n1266), .Y(n1263) );
  NAND4X1 U2834 ( .A(n1269), .B(n71), .C(pc_o[12]), .D(n31), .Y(n1265) );
  AOI21X1 U2835 ( .B(n93), .C(pc_i[13]), .A(n1244), .Y(n1266) );
  OAI32X1 U2836 ( .A(n1267), .B(pc_o[13]), .C(n1146), .D(n1144), .E(n1256), 
        .Y(n1244) );
  MUX2BXL U2837 ( .D0(acc[6]), .D1(n2267), .S(n1150), .Y(n190) );
  INVX1 U2838 ( .A(n1175), .Y(n2222) );
  OAI2B11X1 U2839 ( .D(n1176), .C(n2235), .A(n1177), .B(n1178), .Y(n1175) );
  AOI22X1 U2840 ( .A(n50), .B(n1168), .C(n1139), .D(pc_i[5]), .Y(n1178) );
  AOI32X1 U2841 ( .A(n1179), .B(n29), .C(n2232), .D(pc_o[5]), .E(n1180), .Y(
        n1177) );
  AOI22X1 U2842 ( .A(n921), .B(temp[3]), .C(n2326), .D(n828), .Y(n937) );
  AOI221X1 U2843 ( .A(n2419), .B(n71), .C(pc_i[2]), .D(n1139), .E(n2221), .Y(
        n1120) );
  INVX1 U2844 ( .A(n1210), .Y(n2221) );
  AOI221XL U2845 ( .A(n1211), .B(n2231), .C(pc_o[2]), .D(n1212), .E(n1213), 
        .Y(n1210) );
  AOI21X1 U2846 ( .B(n1204), .C(n1214), .A(n1146), .Y(n1213) );
  NAND21X1 U2847 ( .B(n1677), .A(state[0]), .Y(n1603) );
  AOI222XL U2848 ( .A(n1212), .B(pc_o[1]), .C(n2437), .D(n1220), .E(pc_i[1]), 
        .F(n1139), .Y(n1121) );
  OAI21X1 U2849 ( .B(n1146), .C(pc_o[0]), .A(n1221), .Y(n1220) );
  INVX1 U2850 ( .A(n1320), .Y(n2230) );
  AO2222XL U2851 ( .A(n93), .B(pc_i[8]), .C(n2289), .D(n55), .E(pc_o[8]), .F(
        n1321), .G(n1322), .H(n2422), .Y(n1320) );
  INVX1 U2852 ( .A(n1314), .Y(n2289) );
  OAI22X1 U2853 ( .A(n2235), .B(n1302), .C(n1144), .D(n1147), .Y(n1322) );
  INVX1 U2854 ( .A(n1298), .Y(n2228) );
  AO2222XL U2855 ( .A(n93), .B(pc_i[10]), .C(n2290), .D(n55), .E(pc_o[10]), 
        .F(n1299), .G(n1300), .H(n42), .Y(n1298) );
  INVX1 U2856 ( .A(n1292), .Y(n2290) );
  OAI22X1 U2857 ( .A(n2235), .B(n1281), .C(n1144), .D(n2288), .Y(n1300) );
  INVX1 U2858 ( .A(n1277), .Y(n2226) );
  AO2222XL U2859 ( .A(n93), .B(pc_i[12]), .C(n2291), .D(n55), .E(pc_o[12]), 
        .F(n1278), .G(n1279), .H(n27), .Y(n1277) );
  OAI22X1 U2860 ( .A(n2235), .B(n2292), .C(n45), .D(n2287), .Y(n1279) );
  OAI21X1 U2861 ( .B(n1280), .C(n62), .A(n1271), .Y(n1278) );
  INVX1 U2862 ( .A(b[3]), .Y(n2462) );
  INVX1 U2863 ( .A(b[2]), .Y(n2465) );
  MUX2AXL U2864 ( .D0(n2458), .D1(temp[2]), .S(n1150), .Y(n191) );
  NAND3X1 U2865 ( .A(pc_o[5]), .B(n1442), .C(pc_o[4]), .Y(n1323) );
  NAND2X1 U2866 ( .A(pc_o[2]), .B(pc_o[1]), .Y(n1214) );
  INVX1 U2867 ( .A(pdmode), .Y(n2162) );
  XNOR2XL U2868 ( .A(n1323), .B(memaddr[6]), .Y(n1165) );
  XNOR2XL U2869 ( .A(n1499), .B(memaddr[5]), .Y(n1176) );
  NAND2X1 U2870 ( .A(pc_o[4]), .B(n1442), .Y(n1499) );
  NOR3XL U2871 ( .A(pc_o[4]), .B(pc_o[3]), .C(n1204), .Y(n1179) );
  NOR3XL U2872 ( .A(memaddr[10]), .B(pc_o[11]), .C(n2288), .Y(n1268) );
  NOR3XL U2873 ( .A(pc_o[8]), .B(pc_o[9]), .C(n1147), .Y(n1303) );
  INVX1 U2874 ( .A(b[4]), .Y(n2461) );
  NOR3XL U2875 ( .A(memaddr[6]), .B(pc_o[5]), .C(n2370), .Y(n1145) );
  NOR2X1 U2876 ( .A(pc_o[2]), .B(pc_o[1]), .Y(n1203) );
  NOR2X1 U2877 ( .A(n1314), .B(pc_o[9]), .Y(n1301) );
  NOR2X1 U2878 ( .A(n1292), .B(pc_o[11]), .Y(n1280) );
  NAND32X1 U2879 ( .B(n1302), .C(n2422), .A(pc_o[9]), .Y(n1281) );
  NAND32X1 U2880 ( .B(n1323), .C(n40), .A(pc_o[6]), .Y(n1302) );
  NOR42XL U2881 ( .C(n1008), .D(n254), .A(n2319), .B(n986), .Y(n989) );
  INVX1 U2882 ( .A(b[5]), .Y(n2456) );
  INVX1 U2883 ( .A(b[6]), .Y(n2457) );
  NOR4XL U2884 ( .A(b[2]), .B(b[1]), .C(b[0]), .D(n1047), .Y(n1046) );
  AOI22X1 U2885 ( .A(n920), .B(temp2_comb[1]), .C(n919), .D(pc_i[9]), .Y(n954)
         );
  AOI22X1 U2886 ( .A(n920), .B(temp2_comb[0]), .C(n919), .D(pc_i[8]), .Y(n963)
         );
  OAI211X1 U2887 ( .C(n1017), .D(n253), .A(n2355), .B(n1018), .Y(n990) );
  INVX1 U2888 ( .A(n1022), .Y(n2355) );
  AOI22X1 U2889 ( .A(n259), .B(n1019), .C(n965), .D(phase[2]), .Y(n1018) );
  NOR3XL U2890 ( .A(n767), .B(n318), .C(n783), .Y(n1017) );
  NAND2X1 U2891 ( .A(n2185), .B(n1009), .Y(n994) );
  NAND4X1 U2892 ( .A(n2279), .B(n259), .C(n1010), .D(n2173), .Y(n1009) );
  AOI21X1 U2893 ( .B(phase[0]), .C(n2354), .A(n692), .Y(n961) );
  OAI21X1 U2894 ( .B(n1012), .C(n2356), .A(n1013), .Y(n1010) );
  AOI22X1 U2895 ( .A(n1014), .B(n105), .C(n2476), .D(n54), .Y(n1012) );
  AOI22X1 U2896 ( .A(n259), .B(n964), .C(phase[2]), .D(n965), .Y(n962) );
  NAND3X1 U2897 ( .A(n1008), .B(ramsfraddr[7]), .C(n1011), .Y(n987) );
  NOR3XL U2898 ( .A(n256), .B(n270), .C(n2353), .Y(n1011) );
  INVX1 U2899 ( .A(b[7]), .Y(n2442) );
  OAI21X1 U2900 ( .B(n980), .C(n981), .A(instr[3]), .Y(n976) );
  OAI31XL U2901 ( .A(n968), .B(n969), .C(n970), .D(phase[0]), .Y(n942) );
  OAI22X1 U2902 ( .A(n2388), .B(n2410), .C(n971), .D(n2431), .Y(n970) );
  OAI31XL U2903 ( .A(n2411), .B(n105), .C(n285), .D(n973), .Y(n969) );
  OAI211X1 U2904 ( .C(n975), .D(n25), .A(n976), .B(n977), .Y(n968) );
  NAND4X1 U2905 ( .A(n974), .B(instr[5]), .C(n51), .D(n102), .Y(n973) );
  AOI211X1 U2906 ( .C(n254), .D(n2082), .A(n915), .B(n967), .Y(n2073) );
  OAI21BBX1 U2907 ( .A(n1754), .B(n753), .C(n2372), .Y(n2082) );
  NAND3X1 U2908 ( .A(n862), .B(n1375), .C(ramsfraddr[5]), .Y(n1353) );
  INVX1 U2909 ( .A(finishdiv), .Y(n2211) );
  INVX1 U2910 ( .A(finishmul), .Y(n2212) );
  NOR3XL U2911 ( .A(b[5]), .B(b[7]), .C(b[6]), .Y(n1045) );
  OAI22AX1 U2912 ( .D(ckcon[1]), .C(n878), .A(n2415), .B(n879), .Y(N12966) );
  OAI22AX1 U2913 ( .D(ckcon[5]), .C(n878), .A(n2256), .B(n879), .Y(N12970) );
  OAI22AX1 U2914 ( .D(ckcon[4]), .C(n878), .A(n2169), .B(n879), .Y(N12969) );
  OAI22AX1 U2915 ( .D(ckcon[0]), .C(n878), .A(n2414), .B(n879), .Y(N12965) );
  OAI22AX1 U2916 ( .D(ckcon[3]), .C(n878), .A(n2435), .B(n879), .Y(N12968) );
  OAI22AX1 U2917 ( .D(ckcon[7]), .C(n878), .A(n2257), .B(n879), .Y(N12972) );
  NAND2X1 U2918 ( .A(dec_accop[9]), .B(n2460), .Y(n1034) );
  AND2X1 U2919 ( .A(cpu_resume_ff1), .B(n264), .Y(N13380) );
  INVX1 U2920 ( .A(dec_accop[10]), .Y(n2460) );
  INVX1 U2921 ( .A(dec_accop[9]), .Y(n2453) );
  NAND2X1 U2922 ( .A(dec_accop[17]), .B(accactv), .Y(n1510) );
  INVX1 U2923 ( .A(stop), .Y(n1676) );
  NAND3X1 U2924 ( .A(ramsfraddr[2]), .B(n2440), .C(ramsfraddr[0]), .Y(n855) );
  NAND3X1 U2925 ( .A(n2444), .B(n2440), .C(ramsfraddr[2]), .Y(n854) );
  INVX1 U2926 ( .A(mempswr), .Y(n2331) );
  BUFX3 U2927 ( .A(pc_o[6]), .Y(memaddr[6]) );
  BUFX3 U2928 ( .A(memaddr[4]), .Y(pc_o[4]) );
  BUFX3 U2929 ( .A(memaddr[2]), .Y(pc_o[2]) );
  MUX2X1 U2930 ( .D0(memaddr[5]), .D1(n1621), .S(n155), .Y(memaddr_comb[5]) );
  INVXL U2931 ( .A(n433), .Y(n436) );
  AO2222XL U2932 ( .A(ramdatao[7]), .B(n172), .C(n924), .D(n923), .E(n173), 
        .F(p2[7]), .G(n914), .H(pc_o[15]), .Y(n1595) );
  AO2222XL U2933 ( .A(ramdatao[6]), .B(n172), .C(n907), .D(n923), .E(n173), 
        .F(p2[6]), .G(n914), .H(pc_o[14]), .Y(n1594) );
  AO2222XL U2934 ( .A(ramdatao[5]), .B(n172), .C(n905), .D(n923), .E(n173), 
        .F(p2[5]), .G(n914), .H(pc_o[13]), .Y(n1575) );
  AO2222XL U2935 ( .A(n172), .B(ramdatao[4]), .C(n903), .D(n923), .E(n173), 
        .F(p2[4]), .G(n914), .H(pc_o[12]), .Y(n1580) );
  AO2222XL U2936 ( .A(ramdatao[3]), .B(n172), .C(n898), .D(n923), .E(n173), 
        .F(p2[3]), .G(n914), .H(pc_o[11]), .Y(n1581) );
  OA21XL U2937 ( .B(n1703), .C(n1702), .A(n1701), .Y(n1706) );
  NAND21XL U2938 ( .B(pdmode), .A(n1703), .Y(n1622) );
  INVXL U2939 ( .A(n1703), .Y(n1705) );
  INVXL U2940 ( .A(n455), .Y(n462) );
  AO222XL U2941 ( .A(n2150), .B(ramdatai[5]), .C(n2151), .D(sfrdatai[5]), .E(
        n2152), .F(n2087), .Y(n1445) );
  OAI22XL U2942 ( .A(n987), .B(n1647), .C(n996), .D(n272), .Y(N12719) );
  OAI211XL U2943 ( .C(n1647), .D(n938), .A(n503), .B(n502), .Y(n504) );
  OAI21BBXL U2944 ( .A(n1445), .B(n1444), .C(n2149), .Y(n1446) );
  XNOR2XL U2945 ( .A(n1445), .B(n1501), .Y(n1500) );
  INVX1 U2946 ( .A(n1383), .Y(n1397) );
  OAI22X1 U2947 ( .A(n355), .B(n1649), .C(n354), .D(n720), .Y(n1383) );
  OAI211XL U2948 ( .C(n1648), .D(n938), .A(n475), .B(n473), .Y(n1476) );
  OAI22XL U2949 ( .A(n987), .B(n1648), .C(n998), .D(n271), .Y(N12718) );
  AOI222XL U2950 ( .A(n2150), .B(ramdatai[4]), .C(n2151), .D(sfrdatai[4]), .E(
        n2152), .F(n2136), .Y(n1503) );
  OA21XL U2951 ( .B(n507), .C(n482), .A(n481), .Y(n489) );
  AOI22XL U2952 ( .A(n2153), .B(n827), .C(sfrdatai[2]), .D(n2155), .Y(n1569)
         );
  NAND21XL U2953 ( .B(n216), .A(n1555), .Y(n1554) );
  NAND21XL U2954 ( .B(n1555), .A(n211), .Y(n1556) );
  NAND21XL U2955 ( .B(n1555), .A(n896), .Y(n914) );
  OA21XL U2956 ( .B(n507), .C(n455), .A(n481), .Y(n457) );
  NAND42X1 U2957 ( .C(n379), .D(n378), .A(n377), .B(n376), .Y(n380) );
  AO2222X1 U2958 ( .A(n482), .B(n357), .C(n455), .D(n352), .E(n351), .F(n614), 
        .G(n356), .H(n506), .Y(n358) );
  AO2222X1 U2959 ( .A(n352), .B(n364), .C(n356), .D(n433), .E(n351), .F(n1383), 
        .G(n416), .H(n357), .Y(n359) );
endmodule


module mcu51_cpu_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module mcu51_cpu_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
endmodule


module mcu51_cpu_a0_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
endmodule


module mcu51_cpu_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n10), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n13), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n17), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n14), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  INVX1 U1 ( .A(B[2]), .Y(n17) );
  INVX1 U2 ( .A(B[3]), .Y(n13) );
  INVX1 U3 ( .A(B[4]), .Y(n12) );
  INVX1 U4 ( .A(B[5]), .Y(n10) );
  INVX1 U5 ( .A(B[1]), .Y(n14) );
  NAND21X1 U6 ( .B(n15), .A(n16), .Y(carry[1]) );
  INVX1 U7 ( .A(A[0]), .Y(n16) );
  INVX1 U8 ( .A(B[6]), .Y(n11) );
  AOI21X1 U9 ( .B(carry[7]), .C(A[7]), .A(n9), .Y(DIFF[8]) );
  AOI21BBXL U10 ( .B(A[7]), .C(carry[7]), .A(B[7]), .Y(n9) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U12 ( .A(B[0]), .Y(n15) );
endmodule


module mcu51_cpu_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [8:1] carry;

  FAD1X1 U2_7 ( .A(A[7]), .B(n11), .CI(carry[7]), .CO(carry[8]), .SO(DIFF[7])
         );
  FAD1X1 U2_6 ( .A(A[6]), .B(n13), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n14), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n18), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  INVX1 U1 ( .A(carry[8]), .Y(DIFF[8]) );
  INVX1 U2 ( .A(B[7]), .Y(n11) );
  INVX1 U3 ( .A(B[2]), .Y(n18) );
  INVX1 U4 ( .A(B[3]), .Y(n15) );
  INVX1 U5 ( .A(B[4]), .Y(n14) );
  INVX1 U6 ( .A(B[5]), .Y(n12) );
  INVX1 U7 ( .A(B[6]), .Y(n13) );
  INVX1 U8 ( .A(B[1]), .Y(n16) );
  NAND21X1 U9 ( .B(n17), .A(n10), .Y(carry[1]) );
  INVX1 U10 ( .A(A[0]), .Y(n10) );
  INVX1 U11 ( .A(B[0]), .Y(n17) );
  XOR2X1 U12 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module mcu51_cpu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [15:1] carry;

  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  INVX1 U1 ( .A(B[0]), .Y(n2) );
  NOR21XL U2 ( .B(A[0]), .A(n2), .Y(carry[1]) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mpb_a0 ( i_rd, i_wr, wdat0, wdat1, addr0, addr1, r_i2c_attr, esfrm_oe, 
        esfrm_we, sfrack, esfrm_wdat, esfrm_adr, mcu_esfr_rdat, delay_rdat, 
        delay_rrdy, esfrm_rrdy, esfrm_rdat, channel_sel, r_pg0_sel, dma_w, 
        dma_r, dma_addr, dma_wdat, dma_ack, memaddr, memaddr_c, memwr, memrd, 
        memrd_c, cpurst, memdatao, memack, hit_xd, hit_xr, hit_ps, hit_ps_c, 
        idat_r, idat_w, idat_adr, idat_wdat, iram_ce, xram_ce, regx_re, 
        iram_we, xram_we, regx_we, iram_a, xram_a, iram_d, xram_d, iram_rdat, 
        xram_rdat, regx_rdat, bist_en, bist_wr, bist_adr, bist_wdat, bist_xram, 
        mclk, srstz, test_si, test_so, test_se );
  input [1:0] i_rd;
  input [1:0] i_wr;
  input [7:0] wdat0;
  input [7:0] wdat1;
  input [7:0] addr0;
  input [7:0] addr1;
  output [7:0] esfrm_wdat;
  output [6:0] esfrm_adr;
  input [7:0] mcu_esfr_rdat;
  input [7:0] delay_rdat;
  output [7:0] esfrm_rdat;
  input [3:0] r_pg0_sel;
  input [10:0] dma_addr;
  input [7:0] dma_wdat;
  input [15:0] memaddr;
  input [15:0] memaddr_c;
  input [7:0] memdatao;
  input [7:0] idat_adr;
  input [7:0] idat_wdat;
  output [10:0] iram_a;
  output [10:0] xram_a;
  output [7:0] iram_d;
  output [7:0] xram_d;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  input [7:0] regx_rdat;
  input [10:0] bist_adr;
  input [7:0] bist_wdat;
  input r_i2c_attr, delay_rrdy, channel_sel, dma_w, dma_r, memwr, memrd,
         memrd_c, cpurst, idat_r, idat_w, bist_en, bist_wr, bist_xram, mclk,
         srstz, test_si, test_se;
  output esfrm_oe, esfrm_we, sfrack, esfrm_rrdy, dma_ack, memack, hit_xd,
         hit_xr, hit_ps, hit_ps_c, iram_ce, xram_ce, regx_re, iram_we, xram_we,
         regx_we, test_so;
  wire   pg0_rdwait, pg0_wrwait, N44, N45, r_pg0_rdrdy, N46, xram_rdsel_0_,
         n55, n91, n110, n112, n114, n128, n129, n130, n132, n133, n134, n136,
         n137, n140, n142, n143, n144, n145, n146, n147, n148, n149, n150, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n111, n113, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n131,
         n135, n138, n139, n141, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229;

  SDFFRQX1 r_pg0_rdrdy_reg ( .D(N46), .SIN(pg0_wrwait), .SMC(test_se), .C(mclk), .XR(srstz), .Q(r_pg0_rdrdy) );
  SDFFRQX1 xram_rdsel_reg_1_ ( .D(n224), .SIN(xram_rdsel_0_), .SMC(test_se), 
        .C(mclk), .XR(srstz), .Q(test_so) );
  SDFFRQX1 xram_rdsel_reg_0_ ( .D(n225), .SIN(n3), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(xram_rdsel_0_) );
  SDFFRQX1 pg0_rdwait_reg ( .D(N45), .SIN(test_si), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(pg0_rdwait) );
  SDFFRQX1 pg0_wrwait_reg ( .D(N44), .SIN(pg0_rdwait), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(pg0_wrwait) );
  INVX2 U3 ( .A(i_rd[1]), .Y(n31) );
  OAI31X1 U4 ( .A(r_i2c_attr), .B(n30), .C(n209), .D(n29), .Y(n219) );
  INVX1 U5 ( .A(n222), .Y(n32) );
  NOR2X1 U6 ( .A(n21), .B(cpurst), .Y(memack) );
  NAND2X1 U7 ( .A(n12), .B(n209), .Y(n214) );
  NAND21X1 U8 ( .B(n208), .A(n207), .Y(n213) );
  INVX1 U9 ( .A(n213), .Y(esfrm_oe) );
  AO21X1 U10 ( .B(n208), .C(n207), .A(pg0_rdwait), .Y(n222) );
  OAI2B11X1 U11 ( .D(dma_addr[5]), .C(n127), .A(n158), .B(n95), .Y(xram_a[5])
         );
  AND3X1 U12 ( .A(n13), .B(n14), .C(n15), .Y(n97) );
  OAI2B11X1 U13 ( .D(dma_addr[1]), .C(n127), .A(n138), .B(n87), .Y(xram_a[1])
         );
  AND3X1 U14 ( .A(n17), .B(n18), .C(n19), .Y(n94) );
  OAI211X1 U15 ( .C(n86), .D(n123), .A(n131), .B(n85), .Y(xram_a[0]) );
  OA33X1 U16 ( .A(n181), .B(n215), .C(n180), .D(bist_en), .E(n173), .F(n172), 
        .Y(n1) );
  INVX1 U17 ( .A(n180), .Y(n2) );
  BUFX3 U18 ( .A(r_pg0_rdrdy), .Y(n3) );
  INVX1 U19 ( .A(n170), .Y(n4) );
  INVX1 U20 ( .A(n217), .Y(n5) );
  BUFX3 U21 ( .A(bist_en), .Y(n6) );
  OR2X1 U22 ( .A(i_wr[0]), .B(i_wr[1]), .Y(n210) );
  NAND2X1 U23 ( .A(r_pg0_sel[2]), .B(n27), .Y(n25) );
  INVX1 U24 ( .A(n25), .Y(n7) );
  INVX1 U25 ( .A(n25), .Y(n8) );
  NAND42X1 U26 ( .C(n93), .D(n92), .A(n90), .B(n89), .Y(xram_a[3]) );
  BUFX3 U27 ( .A(bist_en), .Y(n183) );
  INVX1 U28 ( .A(n183), .Y(n9) );
  INVX1 U29 ( .A(n183), .Y(n10) );
  INVX1 U30 ( .A(n183), .Y(n11) );
  INVX1 U31 ( .A(n214), .Y(esfrm_we) );
  OA21X1 U32 ( .B(n212), .C(n211), .A(n210), .Y(n12) );
  NAND2XL U33 ( .A(n116), .B(esfrm_adr[6]), .Y(n14) );
  INVX1 U34 ( .A(n121), .Y(n103) );
  INVX1 U35 ( .A(n125), .Y(n105) );
  NAND2X1 U36 ( .A(memaddr[6]), .B(n105), .Y(n13) );
  NAND2X2 U37 ( .A(memaddr_c[6]), .B(n103), .Y(n15) );
  OA21X1 U38 ( .B(n154), .C(n123), .A(n16), .Y(n89) );
  NAND2X1 U39 ( .A(memaddr_c[3]), .B(n103), .Y(n16) );
  NAND2X1 U40 ( .A(memaddr_c[4]), .B(n103), .Y(n19) );
  NAND2X1 U41 ( .A(memaddr[4]), .B(n105), .Y(n17) );
  NAND2XL U42 ( .A(n116), .B(esfrm_adr[4]), .Y(n18) );
  INVXL U43 ( .A(n163), .Y(esfrm_adr[6]) );
  INVXL U44 ( .A(n86), .Y(esfrm_adr[0]) );
  AO22XL U45 ( .A(idat_adr[0]), .B(n185), .C(n168), .D(esfrm_adr[0]), .Y(n135)
         );
  OAI221XL U46 ( .A(n160), .B(n180), .C(n170), .D(n159), .E(n158), .Y(
        iram_a[5]) );
  AO22XL U47 ( .A(idat_adr[2]), .B(n185), .C(n168), .D(esfrm_adr[2]), .Y(n151)
         );
  OAI221XL U48 ( .A(n163), .B(n180), .C(n170), .D(n162), .E(n161), .Y(
        iram_a[6]) );
  OAI221XL U49 ( .A(n157), .B(n180), .C(n170), .D(n156), .E(n155), .Y(
        iram_a[4]) );
  OAI221XL U50 ( .A(n154), .B(n180), .C(n170), .D(n153), .E(n152), .Y(
        iram_a[3]) );
  OAI21BXL U51 ( .C(n204), .B(n110), .A(n187), .Y(regx_we) );
  INVXL U52 ( .A(n210), .Y(n30) );
  INVXL U53 ( .A(n157), .Y(esfrm_adr[4]) );
  OAI2B11X1 U54 ( .D(dma_addr[4]), .C(n127), .A(n155), .B(n94), .Y(xram_a[4])
         );
  INVX1 U55 ( .A(n177), .Y(n82) );
  INVX1 U56 ( .A(n123), .Y(n116) );
  INVX1 U57 ( .A(n170), .Y(n185) );
  INVX1 U58 ( .A(n180), .Y(n168) );
  INVX1 U59 ( .A(n127), .Y(n106) );
  INVX4 U60 ( .A(n28), .Y(n96) );
  NAND21X2 U61 ( .B(i_wr[1]), .A(n31), .Y(n28) );
  INVX1 U62 ( .A(n81), .Y(n84) );
  INVX1 U63 ( .A(n44), .Y(n60) );
  NAND32X1 U64 ( .B(bist_en), .C(n84), .A(n43), .Y(n44) );
  AND3X1 U65 ( .A(n201), .B(n200), .C(n199), .Y(n193) );
  NAND21X1 U66 ( .B(bist_en), .A(n177), .Y(n83) );
  NAND21X1 U67 ( .B(bist_en), .A(n82), .Y(n123) );
  OR2X1 U68 ( .A(bist_en), .B(n43), .Y(n63) );
  NAND21X1 U69 ( .B(bist_en), .A(n223), .Y(n180) );
  INVX1 U70 ( .A(n217), .Y(n216) );
  INVX1 U71 ( .A(n221), .Y(n223) );
  NAND21X1 U72 ( .B(bist_en), .A(n221), .Y(n170) );
  NAND21X1 U73 ( .B(n11), .A(bist_wdat[0]), .Y(n65) );
  NAND21X1 U74 ( .B(n11), .A(bist_wdat[1]), .Y(n67) );
  NAND21X1 U75 ( .B(n11), .A(bist_wdat[4]), .Y(n73) );
  NAND21X1 U76 ( .B(n10), .A(bist_wdat[2]), .Y(n69) );
  NAND21X1 U77 ( .B(n10), .A(bist_wdat[3]), .Y(n71) );
  NAND21X1 U78 ( .B(n10), .A(bist_wdat[6]), .Y(n77) );
  NAND21X1 U79 ( .B(n218), .A(n217), .Y(n220) );
  NAND32X1 U80 ( .B(n82), .C(n81), .A(n11), .Y(n127) );
  INVX1 U81 ( .A(n42), .Y(n61) );
  NAND32X1 U82 ( .B(n6), .C(n81), .A(n43), .Y(n42) );
  NAND31X1 U83 ( .C(n6), .A(n189), .B(n205), .Y(n197) );
  OA21X1 U84 ( .B(idat_adr[4]), .C(idat_adr[3]), .A(idat_adr[5]), .Y(n129) );
  NAND21X1 U85 ( .B(n219), .A(n32), .Y(n171) );
  INVX1 U86 ( .A(n154), .Y(esfrm_adr[3]) );
  INVX1 U87 ( .A(n160), .Y(esfrm_adr[5]) );
  INVX1 U88 ( .A(n52), .Y(esfrm_wdat[3]) );
  OR2X1 U89 ( .A(idat_r), .B(idat_w), .Y(n221) );
  OR3XL U90 ( .A(n84), .B(n26), .C(n83), .Y(n125) );
  NAND32X1 U91 ( .B(n84), .C(n83), .A(n26), .Y(n121) );
  AO21X1 U92 ( .B(n191), .C(n178), .A(n225), .Y(n81) );
  INVX1 U93 ( .A(memaddr_c[11]), .Y(n201) );
  INVX1 U94 ( .A(memaddr_c[13]), .Y(n199) );
  INVX1 U95 ( .A(memaddr_c[12]), .Y(n200) );
  NAND5XL U96 ( .A(n20), .B(n202), .C(n201), .D(n200), .E(n199), .Y(n203) );
  INVX1 U97 ( .A(memaddr_c[7]), .Y(n202) );
  NAND21X1 U98 ( .B(memaddr_c[9]), .A(n109), .Y(n190) );
  INVX1 U99 ( .A(memaddr_c[8]), .Y(n109) );
  NAND21X1 U100 ( .B(n80), .A(n79), .Y(iram_d[7]) );
  AO22X1 U101 ( .A(idat_wdat[7]), .B(n185), .C(n168), .D(esfrm_wdat[7]), .Y(
        n80) );
  NOR2X1 U102 ( .A(memaddr_c[10]), .B(n190), .Y(n20) );
  INVX1 U103 ( .A(idat_adr[6]), .Y(n162) );
  INVX1 U104 ( .A(idat_adr[4]), .Y(n156) );
  INVX1 U105 ( .A(idat_adr[3]), .Y(n153) );
  NAND21X1 U106 ( .B(n135), .A(n131), .Y(iram_a[0]) );
  NAND21X1 U107 ( .B(n139), .A(n138), .Y(iram_a[1]) );
  AO22X1 U108 ( .A(idat_adr[1]), .B(n185), .C(n168), .D(esfrm_adr[1]), .Y(n139) );
  NAND21X1 U109 ( .B(n151), .A(n141), .Y(iram_a[2]) );
  INVX1 U110 ( .A(idat_adr[5]), .Y(n159) );
  AOI211X1 U111 ( .C(memaddr_c[10]), .D(n190), .A(memaddr_c[14]), .B(
        memaddr_c[15]), .Y(n192) );
  NAND21X1 U112 ( .B(n78), .A(n77), .Y(iram_d[6]) );
  AO22X1 U113 ( .A(idat_wdat[6]), .B(n185), .C(n168), .D(esfrm_wdat[6]), .Y(
        n78) );
  NAND21X1 U114 ( .B(n76), .A(n75), .Y(iram_d[5]) );
  AO22X1 U115 ( .A(idat_wdat[5]), .B(n185), .C(n168), .D(esfrm_wdat[5]), .Y(
        n76) );
  NAND21X1 U116 ( .B(n74), .A(n73), .Y(iram_d[4]) );
  AO22X1 U117 ( .A(idat_wdat[4]), .B(n185), .C(n168), .D(esfrm_wdat[4]), .Y(
        n74) );
  NAND21X1 U118 ( .B(n72), .A(n71), .Y(iram_d[3]) );
  AO22X1 U119 ( .A(idat_wdat[3]), .B(n185), .C(n168), .D(esfrm_wdat[3]), .Y(
        n72) );
  NAND4X1 U120 ( .A(memaddr_c[14]), .B(memaddr_c[13]), .C(memaddr_c[15]), .D(
        n114), .Y(n112) );
  AND3X1 U121 ( .A(memaddr_c[12]), .B(memaddr_c[11]), .C(memaddr_c[7]), .Y(
        n114) );
  NOR43XL U122 ( .B(n225), .C(n187), .D(n186), .A(n112), .Y(n188) );
  AND4X1 U123 ( .A(memaddr_c[9]), .B(memaddr_c[10]), .C(memaddr_c[8]), .D(n224), .Y(n186) );
  NAND21X1 U124 ( .B(n181), .A(n7), .Y(n187) );
  NAND21X1 U125 ( .B(n70), .A(n69), .Y(iram_d[2]) );
  AO22X1 U126 ( .A(idat_wdat[2]), .B(n4), .C(n168), .D(esfrm_wdat[2]), .Y(n70)
         );
  INVX1 U127 ( .A(memaddr_c[9]), .Y(n120) );
  NAND21X1 U128 ( .B(n66), .A(n65), .Y(iram_d[0]) );
  AO22X1 U129 ( .A(idat_wdat[0]), .B(n185), .C(n168), .D(esfrm_wdat[0]), .Y(
        n66) );
  NAND21X1 U130 ( .B(n68), .A(n67), .Y(iram_d[1]) );
  AO22X1 U131 ( .A(idat_wdat[1]), .B(n4), .C(n2), .D(esfrm_wdat[1]), .Y(n68)
         );
  INVX1 U132 ( .A(n110), .Y(hit_xr) );
  INVX1 U133 ( .A(n46), .Y(esfrm_wdat[0]) );
  INVX1 U134 ( .A(hit_xd), .Y(n172) );
  INVX1 U135 ( .A(n48), .Y(esfrm_wdat[1]) );
  NAND21X1 U136 ( .B(n7), .A(n215), .Y(n217) );
  OAI211X1 U137 ( .C(n55), .D(n229), .A(n1), .B(n197), .Y(xram_we) );
  NAND2X1 U138 ( .A(bist_wr), .B(n6), .Y(n55) );
  INVX1 U139 ( .A(n191), .Y(n224) );
  INVX1 U140 ( .A(n124), .Y(n27) );
  INVX1 U141 ( .A(n64), .Y(esfrm_wdat[7]) );
  INVX1 U142 ( .A(n57), .Y(esfrm_wdat[5]) );
  INVX1 U143 ( .A(n54), .Y(esfrm_wdat[4]) );
  INVX1 U144 ( .A(n50), .Y(esfrm_wdat[2]) );
  INVX1 U145 ( .A(n59), .Y(esfrm_wdat[6]) );
  NAND21XL U146 ( .B(esfrm_oe), .A(n140), .Y(esfrm_rrdy) );
  AO21X1 U147 ( .B(idat_w), .C(n185), .A(n184), .Y(iram_we) );
  OAI33XL U148 ( .A(bist_xram), .B(n10), .C(n182), .D(n181), .E(n217), .F(n180), .Y(n184) );
  INVX1 U149 ( .A(bist_wr), .Y(n182) );
  INVX1 U150 ( .A(idat_adr[7]), .Y(n165) );
  NAND21X1 U151 ( .B(n10), .A(bist_wdat[5]), .Y(n75) );
  INVX1 U152 ( .A(n215), .Y(n218) );
  INVX1 U153 ( .A(n179), .Y(n205) );
  NAND32X1 U154 ( .B(n198), .C(n178), .A(n177), .Y(n179) );
  AO21X1 U155 ( .B(test_so), .C(n206), .A(n205), .Y(dma_ack) );
  INVX1 U156 ( .A(n228), .Y(n101) );
  AOI31X1 U157 ( .A(idat_adr[4]), .B(idat_adr[6]), .C(idat_adr[5]), .D(
        idat_adr[7]), .Y(n130) );
  INVX1 U158 ( .A(n91), .Y(n100) );
  AO21X1 U159 ( .B(n176), .C(n175), .A(n174), .Y(n189) );
  NAND21X1 U160 ( .B(n127), .A(dma_addr[3]), .Y(n90) );
  INVX1 U161 ( .A(n152), .Y(n92) );
  AND2X1 U162 ( .A(memaddr[3]), .B(n105), .Y(n93) );
  MUX2IXL U163 ( .D0(addr1[3]), .D1(addr0[3]), .S(n96), .Y(n154) );
  INVX1 U164 ( .A(r_i2c_attr), .Y(n211) );
  MUX2IXL U165 ( .D0(addr1[0]), .D1(addr0[0]), .S(n96), .Y(n86) );
  MUX2IXL U166 ( .D0(addr1[4]), .D1(addr0[4]), .S(n96), .Y(n157) );
  MUX2IXL U167 ( .D0(addr1[6]), .D1(addr0[6]), .S(n96), .Y(n163) );
  MUX2IXL U168 ( .D0(addr1[5]), .D1(addr0[5]), .S(n96), .Y(n160) );
  AOI222XL U169 ( .A(dma_addr[0]), .B(n106), .C(memaddr_c[0]), .D(n103), .E(
        memaddr[0]), .F(n105), .Y(n85) );
  AOI222XL U170 ( .A(memaddr[1]), .B(n105), .C(n116), .D(esfrm_adr[1]), .E(
        memaddr_c[1]), .F(n103), .Y(n87) );
  INVX1 U171 ( .A(pg0_wrwait), .Y(n29) );
  AOI222XL U172 ( .A(memaddr[5]), .B(n105), .C(n116), .D(esfrm_adr[5]), .E(
        memaddr_c[5]), .F(n103), .Y(n95) );
  AOI21X1 U173 ( .B(test_so), .C(xram_rdsel_0_), .A(n204), .Y(n21) );
  OAI2B11X1 U174 ( .D(dma_addr[6]), .C(n127), .A(n161), .B(n97), .Y(xram_a[6])
         );
  MUX2XL U175 ( .D0(addr1[1]), .D1(addr0[1]), .S(n96), .Y(esfrm_adr[1]) );
  MUX2XL U176 ( .D0(addr1[2]), .D1(addr0[2]), .S(n96), .Y(esfrm_adr[2]) );
  GEN3XL U177 ( .F(xram_rdsel_0_), .G(n36), .E(n35), .D(n37), .C(n82), .B(n34), 
        .A(n198), .Y(n191) );
  INVX1 U178 ( .A(dma_r), .Y(n35) );
  OAI211X1 U179 ( .C(dma_r), .D(memrd_c), .A(xram_rdsel_0_), .B(n33), .Y(n34)
         );
  AND2X1 U180 ( .A(n178), .B(n36), .Y(n33) );
  INVX1 U181 ( .A(n41), .Y(n225) );
  MUX3X1 U182 ( .D0(n38), .D1(n24), .D2(n181), .S0(xram_rdsel_0_), .S1(test_so), .Y(n39) );
  INVX1 U183 ( .A(n198), .Y(n40) );
  NAND21X1 U184 ( .B(dma_w), .A(memrd_c), .Y(n37) );
  NOR2X1 U185 ( .A(dma_r), .B(n37), .Y(n24) );
  OAI211X1 U186 ( .C(n46), .D(n63), .A(n65), .B(n45), .Y(xram_d[0]) );
  AOI22X1 U187 ( .A(dma_wdat[0]), .B(n61), .C(memdatao[0]), .D(n60), .Y(n45)
         );
  AOI211X1 U188 ( .C(memaddr_c[14]), .D(n203), .A(memaddr_c[15]), .B(cpurst), 
        .Y(hit_ps_c) );
  OAI211X1 U189 ( .C(n120), .D(n121), .A(n119), .B(n118), .Y(xram_a[9]) );
  AOI31X1 U190 ( .A(n116), .B(r_pg0_sel[2]), .C(n212), .D(iram_a[9]), .Y(n119)
         );
  OA22X1 U191 ( .A(n125), .B(n117), .C(n127), .D(n175), .Y(n118) );
  NAND32X1 U192 ( .B(n2), .C(n4), .A(n167), .Y(iram_a[8]) );
  OAI221X1 U193 ( .A(n113), .B(n123), .C(n10), .D(n167), .E(n111), .Y(
        xram_a[8]) );
  INVX1 U194 ( .A(bist_adr[8]), .Y(n167) );
  OAI221X1 U195 ( .A(n180), .B(n166), .C(n170), .D(n165), .E(n164), .Y(
        iram_a[7]) );
  OAI211X1 U196 ( .C(n166), .D(n123), .A(n164), .B(n107), .Y(xram_a[7]) );
  INVX1 U197 ( .A(r_pg0_sel[0]), .Y(n166) );
  OAI2B11X1 U198 ( .D(n128), .C(n170), .A(n180), .B(n169), .Y(iram_a[10]) );
  OAI211X1 U199 ( .C(n174), .D(n127), .A(n169), .B(n126), .Y(xram_a[10]) );
  OAI211X1 U200 ( .C(n129), .D(idat_adr[6]), .A(n130), .B(channel_sel), .Y(
        n128) );
  OAI211X1 U201 ( .C(n224), .D(n1), .A(n197), .B(n196), .Y(xram_ce) );
  MUX3IX1 U202 ( .D0(n195), .D1(n194), .D2(bist_xram), .S0(n225), .S1(bist_en), 
        .Y(n196) );
  AND2X1 U203 ( .A(n224), .B(n189), .Y(n195) );
  AO21X1 U204 ( .B(n193), .C(n192), .A(n191), .Y(n194) );
  OAI211X1 U205 ( .C(r_pg0_sel[1]), .D(r_pg0_sel[0]), .A(r_pg0_sel[2]), .B(
        r_pg0_sel[3]), .Y(n212) );
  OA222X1 U206 ( .A(n125), .B(n228), .C(n124), .D(n123), .E(n122), .F(n121), 
        .Y(n126) );
  INVX1 U207 ( .A(memaddr_c[10]), .Y(n122) );
  AOI211X1 U208 ( .C(memaddr[14]), .D(n136), .A(memaddr[15]), .B(cpurst), .Y(
        hit_ps) );
  NAND4X1 U209 ( .A(n226), .B(n228), .C(n91), .D(n137), .Y(n136) );
  NOR3XL U210 ( .A(memaddr[12]), .B(memaddr[7]), .C(memaddr[13]), .Y(n137) );
  AOI222XL U211 ( .A(dma_addr[7]), .B(n106), .C(n105), .D(n104), .E(n103), .F(
        n102), .Y(n107) );
  OAI31XL U212 ( .A(n101), .B(n100), .C(n99), .D(n98), .Y(n104) );
  AO21X1 U213 ( .B(channel_sel), .C(n20), .A(memaddr_c[7]), .Y(n102) );
  INVX1 U214 ( .A(channel_sel), .Y(n99) );
  NOR2X1 U215 ( .A(memaddr[8]), .B(memaddr[9]), .Y(n91) );
  INVX1 U216 ( .A(memaddr[10]), .Y(n228) );
  OAI211X1 U217 ( .C(n54), .D(n63), .A(n73), .B(n53), .Y(xram_d[4]) );
  AOI22X1 U218 ( .A(dma_wdat[4]), .B(n61), .C(memdatao[4]), .D(n60), .Y(n53)
         );
  OAI211X1 U219 ( .C(n64), .D(n63), .A(n79), .B(n62), .Y(xram_d[7]) );
  AOI22X1 U220 ( .A(dma_wdat[7]), .B(n61), .C(memdatao[7]), .D(n60), .Y(n62)
         );
  INVX1 U221 ( .A(memaddr[11]), .Y(n226) );
  OA222X1 U222 ( .A(n127), .B(n176), .C(n109), .D(n121), .E(n125), .F(n108), 
        .Y(n111) );
  INVX1 U223 ( .A(memaddr[8]), .Y(n108) );
  OAI211X1 U224 ( .C(n48), .D(n63), .A(n67), .B(n47), .Y(xram_d[1]) );
  AOI22X1 U225 ( .A(dma_wdat[1]), .B(n61), .C(memdatao[1]), .D(n60), .Y(n47)
         );
  OAI211X1 U226 ( .C(n59), .D(n63), .A(n77), .B(n58), .Y(xram_d[6]) );
  AOI22X1 U227 ( .A(dma_wdat[6]), .B(n61), .C(memdatao[6]), .D(n60), .Y(n58)
         );
  OAI211X1 U228 ( .C(n57), .D(n63), .A(n75), .B(n56), .Y(xram_d[5]) );
  AOI22X1 U229 ( .A(dma_wdat[5]), .B(n61), .C(memdatao[5]), .D(n60), .Y(n56)
         );
  OAI211X1 U230 ( .C(n50), .D(n63), .A(n69), .B(n49), .Y(xram_d[2]) );
  AOI22X1 U231 ( .A(dma_wdat[2]), .B(n61), .C(memdatao[2]), .D(n60), .Y(n49)
         );
  OAI211X1 U232 ( .C(n52), .D(n63), .A(n71), .B(n51), .Y(xram_d[3]) );
  AOI22X1 U233 ( .A(dma_wdat[3]), .B(n61), .C(memdatao[3]), .D(n60), .Y(n51)
         );
  INVX1 U234 ( .A(memaddr[12]), .Y(n227) );
  NAND4X1 U235 ( .A(memaddr[11]), .B(memaddr[7]), .C(n132), .D(n133), .Y(n110)
         );
  NOR43XL U236 ( .B(memaddr[15]), .C(memaddr[13]), .D(memaddr[14]), .A(n227), 
        .Y(n133) );
  AND3X1 U237 ( .A(memaddr[8]), .B(memaddr[9]), .C(memaddr[10]), .Y(n132) );
  NOR4XL U238 ( .A(memaddr[14]), .B(memaddr[15]), .C(memaddr[13]), .D(n134), 
        .Y(hit_xd) );
  OAI211X1 U239 ( .C(n228), .D(n91), .A(n227), .B(n226), .Y(n134) );
  NOR21XL U240 ( .B(delay_rrdy), .A(r_pg0_rdrdy), .Y(n143) );
  AO222XL U241 ( .A(mcu_esfr_rdat[7]), .B(n140), .C(r_pg0_rdrdy), .D(n142), 
        .E(delay_rdat[7]), .F(n143), .Y(esfrm_rdat[7]) );
  AO222X1 U242 ( .A(xram_rdat[7]), .B(n218), .C(iram_rdat[7]), .D(n216), .E(
        regx_rdat[7]), .F(n8), .Y(n142) );
  AO21X1 U243 ( .B(r_pg0_sel[1]), .C(n27), .A(n7), .Y(n215) );
  NAND2X1 U244 ( .A(n212), .B(r_pg0_sel[3]), .Y(n124) );
  NOR2X1 U245 ( .A(delay_rrdy), .B(r_pg0_rdrdy), .Y(n140) );
  AO222X1 U246 ( .A(xram_rdat[2]), .B(n218), .C(iram_rdat[2]), .D(n216), .E(
        regx_rdat[2]), .F(n8), .Y(n148) );
  AO222X1 U247 ( .A(xram_rdat[4]), .B(n218), .C(iram_rdat[4]), .D(n216), .E(
        regx_rdat[4]), .F(n8), .Y(n146) );
  AO222X1 U248 ( .A(xram_rdat[5]), .B(n218), .C(iram_rdat[5]), .D(n216), .E(
        regx_rdat[5]), .F(n8), .Y(n145) );
  MUX2BXL U249 ( .D0(n198), .D1(bist_xram), .S(n6), .Y(iram_ce) );
  AO222XL U250 ( .A(mcu_esfr_rdat[6]), .B(n140), .C(r_pg0_rdrdy), .D(n144), 
        .E(delay_rdat[6]), .F(n143), .Y(esfrm_rdat[6]) );
  AO222X1 U251 ( .A(xram_rdat[6]), .B(n218), .C(iram_rdat[6]), .D(n216), .E(
        regx_rdat[6]), .F(n8), .Y(n144) );
  AO222XL U252 ( .A(mcu_esfr_rdat[3]), .B(n140), .C(r_pg0_rdrdy), .D(n147), 
        .E(delay_rdat[3]), .F(n143), .Y(esfrm_rdat[3]) );
  AO222X1 U253 ( .A(xram_rdat[3]), .B(n218), .C(iram_rdat[3]), .D(n216), .E(
        regx_rdat[3]), .F(n8), .Y(n147) );
  AO222XL U254 ( .A(mcu_esfr_rdat[1]), .B(n140), .C(r_pg0_rdrdy), .D(n149), 
        .E(delay_rdat[1]), .F(n143), .Y(esfrm_rdat[1]) );
  AO222X1 U255 ( .A(xram_rdat[1]), .B(n218), .C(iram_rdat[1]), .D(n216), .E(
        regx_rdat[1]), .F(n8), .Y(n149) );
  AO222XL U256 ( .A(mcu_esfr_rdat[0]), .B(n140), .C(n3), .D(n150), .E(
        delay_rdat[0]), .F(n143), .Y(esfrm_rdat[0]) );
  AO222X1 U257 ( .A(xram_rdat[0]), .B(n218), .C(iram_rdat[0]), .D(n216), .E(
        regx_rdat[0]), .F(n8), .Y(n150) );
  NAND21X1 U258 ( .B(n9), .A(bist_adr[3]), .Y(n152) );
  NAND21X1 U259 ( .B(n11), .A(bist_adr[1]), .Y(n138) );
  NAND21X1 U260 ( .B(n10), .A(bist_adr[2]), .Y(n141) );
  NAND21X1 U261 ( .B(n11), .A(bist_adr[0]), .Y(n131) );
  NAND21X1 U262 ( .B(n10), .A(bist_adr[5]), .Y(n158) );
  NAND21X1 U263 ( .B(n10), .A(bist_adr[6]), .Y(n161) );
  NAND21X1 U264 ( .B(n11), .A(bist_adr[4]), .Y(n155) );
  INVX1 U265 ( .A(test_so), .Y(n36) );
  NOR2X1 U266 ( .A(memrd), .B(memwr), .Y(n26) );
  NAND21X1 U267 ( .B(n11), .A(bist_wdat[7]), .Y(n79) );
  INVX1 U268 ( .A(n115), .Y(iram_a[9]) );
  NAND21X1 U269 ( .B(n11), .A(bist_adr[9]), .Y(n115) );
  NAND21X1 U270 ( .B(n10), .A(bist_adr[10]), .Y(n169) );
  NAND21X1 U271 ( .B(n11), .A(bist_adr[7]), .Y(n164) );
  INVX1 U272 ( .A(memaddr[7]), .Y(n98) );
  INVX1 U273 ( .A(memaddr[9]), .Y(n117) );
  INVX1 U274 ( .A(r_pg0_sel[1]), .Y(n113) );
  INVX1 U275 ( .A(xram_rdsel_0_), .Y(n206) );
  INVX1 U276 ( .A(bist_xram), .Y(n229) );
  INVX1 U277 ( .A(dma_w), .Y(n178) );
  INVX1 U278 ( .A(dma_addr[10]), .Y(n174) );
  INVX1 U279 ( .A(dma_addr[8]), .Y(n176) );
  INVX1 U280 ( .A(dma_addr[9]), .Y(n175) );
  AO21XL U281 ( .B(n216), .C(n171), .A(n221), .Y(n198) );
  NAND21XL U282 ( .B(n5), .A(n171), .Y(n177) );
  AND3XL U283 ( .A(n219), .B(n221), .C(n220), .Y(N44) );
  INVXL U284 ( .A(n219), .Y(n181) );
  AND3XL U285 ( .A(n221), .B(n222), .C(n220), .Y(N45) );
  OA21XL U286 ( .B(n223), .C(n8), .A(n222), .Y(N46) );
  AO21XL U287 ( .B(n8), .C(n222), .A(n188), .Y(regx_re) );
  OAI211XL U288 ( .C(n24), .D(n222), .A(n40), .B(n39), .Y(n41) );
  NAND21XL U289 ( .B(n222), .A(n82), .Y(n38) );
  NAND21XL U290 ( .B(n216), .A(n219), .Y(n43) );
  INVX1 U291 ( .A(n173), .Y(n204) );
  NAND43X1 U292 ( .B(dma_r), .C(dma_w), .D(n171), .A(memwr), .Y(n173) );
  MUX2IX2 U293 ( .D0(addr1[7]), .D1(addr0[7]), .S(n96), .Y(n208) );
  AND2XL U294 ( .A(n214), .B(n213), .Y(sfrack) );
  AO222XL U295 ( .A(mcu_esfr_rdat[5]), .B(n140), .C(r_pg0_rdrdy), .D(n145), 
        .E(delay_rdat[5]), .F(n143), .Y(esfrm_rdat[5]) );
  AO222XL U296 ( .A(mcu_esfr_rdat[4]), .B(n140), .C(r_pg0_rdrdy), .D(n146), 
        .E(delay_rdat[4]), .F(n143), .Y(esfrm_rdat[4]) );
  MUX2IXL U297 ( .D0(wdat0[5]), .D1(wdat1[5]), .S(i_wr[1]), .Y(n57) );
  MUX2IXL U298 ( .D0(wdat0[2]), .D1(wdat1[2]), .S(i_wr[1]), .Y(n50) );
  MUX2IXL U299 ( .D0(wdat0[4]), .D1(wdat1[4]), .S(i_wr[1]), .Y(n54) );
  MUX2IXL U300 ( .D0(wdat0[6]), .D1(wdat1[6]), .S(i_wr[1]), .Y(n59) );
  MUX2IXL U301 ( .D0(wdat0[7]), .D1(wdat1[7]), .S(i_wr[1]), .Y(n64) );
  MUX2IXL U302 ( .D0(wdat0[1]), .D1(wdat1[1]), .S(i_wr[1]), .Y(n48) );
  MUX2IXL U303 ( .D0(wdat0[0]), .D1(wdat1[0]), .S(i_wr[1]), .Y(n46) );
  MUX2IXL U304 ( .D0(wdat0[3]), .D1(wdat1[3]), .S(i_wr[1]), .Y(n52) );
  NAND21XL U305 ( .B(i_rd[0]), .A(n31), .Y(n207) );
  AOI222XL U306 ( .A(memaddr[2]), .B(n105), .C(n116), .D(esfrm_adr[2]), .E(
        memaddr_c[2]), .F(n103), .Y(n88) );
  AO222XL U307 ( .A(mcu_esfr_rdat[2]), .B(n140), .C(r_pg0_rdrdy), .D(n148), 
        .E(delay_rdat[2]), .F(n143), .Y(esfrm_rdat[2]) );
  INVX2 U308 ( .A(n208), .Y(n209) );
  OAI2B11X4 U309 ( .D(dma_addr[2]), .C(n127), .A(n141), .B(n88), .Y(xram_a[2])
         );
endmodule


module ATO0008KX8MX180LBX4DA ( A, CSB, CLK, PGM, RE, TWLB, VSS, VDD, VDDP, SAP, 
        Q );
  input [15:0] A;
  input [1:0] TWLB;
  input [1:0] SAP;
  output [7:0] Q;
  input CSB, CLK, PGM, RE, VSS, VDD, VDDP;


endmodule


module MSL18B_1536X8_RW10TM4_16 ( DO, CK, CSB, OEB, WEB, A, DI );
  output [7:0] DO;
  input [10:0] A;
  input [7:0] DI;
  input CK, CSB, OEB, WEB;


endmodule


module IOBMURUDA_A1 ( PAD, IE, DI, OE, DO, PU, PD, ANA_R, RSTB_5, VB, ANA_P );
  input IE, OE, DO, PU, PD, RSTB_5, VB, ANA_P;
  output DI, ANA_R;
  inout PAD;


endmodule


module IOBMURUDA_A0 ( PAD, IE, DI, OE, DO, PU, PD, ANA_R, RSTB_5, VB );
  input IE, OE, DO, PU, PD, RSTB_5, VB;
  output DI, ANA_R;
  inout PAD;


endmodule


module IODMURUDA_A0 ( PAD, IE, DI, OE, DO, PU, PD, ANA_R, RSTB_5, VB );
  input IE, OE, DO, PU, PD, RSTB_5, VB;
  output DI, ANA_R;
  inout PAD;


endmodule


module anatop_1127a0 ( CC1, CC2, DP, DN, VFB, CSP, CSN, COM, LG, SW, HG, BST, 
        GATE, VDRV, BST_SET, DCM_SEL, HGOFF, HGLGOFF, HGON, LGON, ENDRV, FSW, 
        EN_OSC, MAXDS, EN_GM, EN_ODLDO, EN_IBUK, RP_SEL, RP1_EN, RP2_EN, 
        VCONN1_EN, VCONN2_EN, SGP, S20U, S100U, TX_EN, TX_DAT, CC_SEL, TRA, 
        TFA, LSR, RX_DAT, RX_SQL, SEL_RX_TH, DAC1_EN, DPDN_SHORT, DP_2V7_EN, 
        DN_2V7_EN, DP_0P6V_EN, DN_0P6V_EN, DP_DWN_EN, DN_DWN_EN, PWR_I, DAC3, 
        DAC1, CV2, LFOSC_ENB, VO_DISCHG, DISCHG_SEL, CMP_SEL_VO10, 
        CMP_SEL_VO20, CMP_SEL_GP1, CMP_SEL_GP2, CMP_SEL_GP3, CMP_SEL_GP4, 
        CMP_SEL_GP5, CMP_SEL_VIN20, CMP_SEL_TS, CMP_SEL_IS, CMP_SEL_CC2, 
        CMP_SEL_CC1, CMP_SEL_CC2_4, CMP_SEL_CC1_4, CMP_SEL_DP, CMP_SEL_DP_3, 
        CMP_SEL_DN, CMP_SEL_DN_3, OCP_EN, CS_EN, COMP_O, CCI2C_EN, UVP_SEL, TM, 
        V5OCP, RSTB, DAC0, SLEEP, OSC_LOW, OSC_STOP, PWRDN, VPP_ZERO, OSC_O, 
        RD_DET, IMP_OSC, DRP_OSC, STB_RP, RD_ENB, PWREN, OCP, SCP, UVP, 
        LDO3P9V, VPP_SEL, CC1_DOB, CC2_DOB, CC1_DI, CC2_DI, ANTI_INRUSH, OTPI, 
        OVP_SEL, OVP, DN_COMP, DP_COMP, DPDN_VTH, DPDEN, DPDO, DPIE, DNDEN, 
        DNDO, DNIE, DUMMY_IN, CP_CLKX2, SEL_CONST_OVP, LP_EN, DNCHK_EN, IRP_EN, 
        CCBFEN, REGTRM, AD_RST, AD_HOLD, DN_FAULT, SEL_CCGAIN, VFB_SW, CPV_SEL, 
        CLAMPV_EN, HVNG_CPEN, PWREN_HOLD, OCP_SEL, OCP_80M, OCP_160M, OPTO1, 
        OPTO2, VPP_OTP, VDD_OTP, RSTB_5, V1P1, TS_ANA_R, GP5_ANA_R, GP4_ANA_R, 
        GP3_ANA_R, GP2_ANA_R, GP1_ANA_R, TS_ANA_P, GP5_ANA_P, GP4_ANA_P, 
        GP3_ANA_P, GP2_ANA_P, GP1_ANA_P );
  input [1:0] FSW;
  input [1:0] RP_SEL;
  input [5:1] SGP;
  input [7:0] PWR_I;
  input [5:0] DAC3;
  input [9:0] DAC1;
  input [3:0] TM;
  input [10:0] DAC0;
  input [1:0] OVP_SEL;
  input [7:0] DUMMY_IN;
  input [55:0] REGTRM;
  input BST_SET, DCM_SEL, HGOFF, HGLGOFF, HGON, LGON, ENDRV, EN_OSC, MAXDS,
         EN_GM, EN_ODLDO, EN_IBUK, RP1_EN, RP2_EN, VCONN1_EN, VCONN2_EN, S20U,
         S100U, TX_EN, TX_DAT, CC_SEL, TRA, TFA, LSR, SEL_RX_TH, DAC1_EN,
         DPDN_SHORT, DP_2V7_EN, DN_2V7_EN, DP_0P6V_EN, DN_0P6V_EN, DP_DWN_EN,
         DN_DWN_EN, CV2, LFOSC_ENB, VO_DISCHG, DISCHG_SEL, CMP_SEL_VO10,
         CMP_SEL_VO20, CMP_SEL_GP1, CMP_SEL_GP2, CMP_SEL_GP3, CMP_SEL_GP4,
         CMP_SEL_GP5, CMP_SEL_VIN20, CMP_SEL_TS, CMP_SEL_IS, CMP_SEL_CC2,
         CMP_SEL_CC1, CMP_SEL_CC2_4, CMP_SEL_CC1_4, CMP_SEL_DP, CMP_SEL_DP_3,
         CMP_SEL_DN, CMP_SEL_DN_3, OCP_EN, CS_EN, CCI2C_EN, UVP_SEL, SLEEP,
         OSC_LOW, OSC_STOP, PWRDN, VPP_ZERO, STB_RP, RD_ENB, PWREN, LDO3P9V,
         VPP_SEL, CC1_DOB, CC2_DOB, ANTI_INRUSH, DPDN_VTH, DPDEN, DPDO, DPIE,
         DNDEN, DNDO, DNIE, CP_CLKX2, SEL_CONST_OVP, LP_EN, DNCHK_EN, IRP_EN,
         CCBFEN, AD_RST, AD_HOLD, SEL_CCGAIN, VFB_SW, CPV_SEL, CLAMPV_EN,
         HVNG_CPEN, PWREN_HOLD, OCP_SEL, TS_ANA_R, GP5_ANA_R, GP4_ANA_R,
         GP3_ANA_R, GP2_ANA_R, GP1_ANA_R;
  output RX_DAT, RX_SQL, COMP_O, V5OCP, RSTB, OSC_O, RD_DET, IMP_OSC, DRP_OSC,
         OCP, SCP, UVP, CC1_DI, CC2_DI, OTPI, OVP, DN_COMP, DP_COMP, DN_FAULT,
         OCP_80M, OCP_160M, OPTO1, OPTO2, VPP_OTP, VDD_OTP, RSTB_5, V1P1,
         TS_ANA_P, GP5_ANA_P, GP4_ANA_P, GP3_ANA_P, GP2_ANA_P, GP1_ANA_P;
  inout CC1,  CC2,  DP,  DN,  VFB,  CSP,  CSN,  COM,  LG,  SW,  HG,  BST, 
     GATE,  VDRV;


endmodule

