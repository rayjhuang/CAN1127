module anatop_1127a0 ( VBUS, CC1, CC2, DP, DN, VFB, IFB, ISENP, ISENN, OCDRV, 
        GATE_A, GATE_B, RP_SEL, RP1_EN, RP2_EN, VCONN1_EN, VCONN2_EN, GP3_20U, 
        GP4_20U, GP5_20U, S20UB, S100UB, TX_EN, TX_DAT, CC_SEL, TRA, TFA, 
        RX_D_PK, RX_D_49, RX_SQL, CCBIAS, CCLEVEL, CV_ENB, CC_ENB, DAC1_EN, 
        DPDN_SHORT, DP_2V7_EN, DN_2V7_EN, DP_0P6V_EN, DN_0P6V_EN, DP_DWN_EN, 
        DN_DWN_EN, PWR_I, DAC3, DAC1, CV2, CS_DIR, LFOSC_ENB, VIN_DISCHG_EN, 
        VBUS_DISCHG_EN, DISCHG_SEL, T3A, CC_FT, CMP_SEL_GP3, CMP_SEL_GP4, 
        CMP_SEL_GP5, CMP_SEL_VIN20, CMP_SEL_DI, CMP_SEL_DV, CMP_SEL_T, 
        CMP_SEL_VIN, CMP_SEL_IS, CMP_SEL_VBUS, CMP_SEL_CC2, CMP_SEL_CC1, 
        CMP_SEL_CC2_4, CMP_SEL_CC1_4, CMP_SEL_DN, CMP_SEL_DP, OCP_EN, CS_EN, 
        COMP_O, CCI2C_EN, UVP_SEL, TM, V5OCP, RSTB, RSTB_5, V1P1, DAC0, SLEEP, 
        OSC_LOW, OSC_STOP, PWRDN, VPP_ZERO, OCDRV_ENZ, OSC_O, RD_DET, STB_OVP, 
        IMP_OSC, DRP_OSC, STB_RP, RD_ENB, PWREN_A, PWREN_B, OCP, SCP, UVP, 
        LDO3P9V, VPP_SEL, VPP_OTP, VDD_OTP, CC1_DOB, CC2_DOB, CC1_DI, CC2_DI, 
        ANTI_INRUSH, IFB_CUT, OTPI, CF, CC_PROT, OVP_SEL, OVP, TX_DRV0, 
        DN_COMP, DP_COMP, DPDN_VTH, DPDEN, DPDO, DPIE, DNDEN, DNDO, DNIE, IDEN, 
        IDDO, IDIN, DUMMY_IN, REGTRM, AD_RST, AD_HOLD, DN_FAULT, VBUS_400K, 
        SEL_CCGAIN, SEL_OCDRV, SEL_FB, CPV_SEL, CLAMPV_EN, HVNG_CPEN, 
        PWREN_HOLD, OCP_SEL, IDAC_EN, IDAC_SEN, OCP_80M, OCP_160M, OPTO1, 
        OPTO2, TS_ANA_R, GP5_ANA_R, GP4_ANA_R, GP3_ANA_R, TS_ANA_P, GP5_ANA_P, 
        GP4_ANA_P, GP3_ANA_P );
  input [1:0] RP_SEL;
  input [7:0] PWR_I;
  input [5:0] DAC3;
  input [9:0] DAC1;
  input [3:0] TM;
  input [10:0] DAC0;
  input [1:0] OVP_SEL;
  input [7:0] DUMMY_IN;
  input [47:0] REGTRM;
  input VFB, IFB, ISENP, ISENN, RP1_EN, RP2_EN, VCONN1_EN, VCONN2_EN, GP3_20U,
         GP4_20U, GP5_20U, S20UB, S100UB, TX_EN, TX_DAT, CC_SEL, TRA, TFA,
         CCBIAS, CCLEVEL, CV_ENB, CC_ENB, DAC1_EN, DPDN_SHORT, DP_2V7_EN,
         DN_2V7_EN, DP_0P6V_EN, DN_0P6V_EN, DP_DWN_EN, DN_DWN_EN, CV2, CS_DIR,
         LFOSC_ENB, VIN_DISCHG_EN, VBUS_DISCHG_EN, DISCHG_SEL, T3A, CC_FT,
         CMP_SEL_GP3, CMP_SEL_GP4, CMP_SEL_GP5, CMP_SEL_VIN20, CMP_SEL_DI,
         CMP_SEL_DV, CMP_SEL_T, CMP_SEL_VIN, CMP_SEL_IS, CMP_SEL_VBUS,
         CMP_SEL_CC2, CMP_SEL_CC1, CMP_SEL_CC2_4, CMP_SEL_CC1_4, CMP_SEL_DN,
         CMP_SEL_DP, OCP_EN, CS_EN, CCI2C_EN, UVP_SEL, SLEEP, OSC_LOW,
         OSC_STOP, PWRDN, VPP_ZERO, OCDRV_ENZ, STB_RP, RD_ENB, PWREN_A,
         PWREN_B, LDO3P9V, VPP_SEL, CC1_DOB, CC2_DOB, ANTI_INRUSH, IFB_CUT,
         CC_PROT, TX_DRV0, DPDN_VTH, DPDEN, DPDO, DPIE, DNDEN, DNDO, DNIE,
         IDEN, IDDO, AD_RST, AD_HOLD, VBUS_400K, SEL_CCGAIN, SEL_OCDRV, SEL_FB,
         CPV_SEL, CLAMPV_EN, HVNG_CPEN, PWREN_HOLD, OCP_SEL, IDAC_EN, IDAC_SEN,
         TS_ANA_R, GP5_ANA_R, GP4_ANA_R, GP3_ANA_R;
  output OCDRV, GATE_A, GATE_B, RX_D_PK, RX_D_49, RX_SQL, COMP_O, V5OCP, RSTB,
         RSTB_5, V1P1, OSC_O, RD_DET, STB_OVP, IMP_OSC, DRP_OSC, OCP, SCP, UVP,
         VPP_OTP, VDD_OTP, CC1_DI, CC2_DI, OTPI, CF, OVP, DN_COMP, DP_COMP,
         IDIN, DN_FAULT, OCP_80M, OCP_160M, OPTO1, OPTO2, TS_ANA_P, GP5_ANA_P,
         GP4_ANA_P, GP3_ANA_P;
  inout VBUS,  CC1,  CC2,  DP,  DN;

reg r_rstz=0;
assign RSTB = r_rstz;

endmodule

