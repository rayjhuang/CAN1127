
module chiptop_1127a0 ( CSP, CSN, VFB, COMP, SW, BST, VDRV, LG, HG, GATE, DP, 
        DN, CC1, CC2, TST, GPIO_TS, SCL, SDA, GPIO1, GPIO2, GPIO3, GPIO4, 
        GPIO5 );
  input TST;
  output LG, HG, GATE;
  inout CSP,  CSN,  VFB,  COMP,  SW,  BST,  VDRV,  DP,  DN,  CC1,  CC2, 
     GPIO_TS,  SCL,  SDA,  GPIO1,  GPIO2,  GPIO3,  GPIO4,  GPIO5;
  wire   SRAM_WEB, SRAM_CEB, SRAM_OEB, PWREN_HOLD, RD_ENB, STB_RP, DRP_OSC,
         IMP_OSC, TX_EN, TX_DAT, RX_DAT, RX_SQL, DAC1_EN, AD_RST, AD_HOLD,
         COMP_O, CCI2C_EN, RSTB, SLEEP, OSC_LOW, OSC_STOP, PWRDN, VPP_0V,
         VPP_SEL, LDO3P9V, OSC_O, RD_DET, OCP_SEL, CC1_DOB, CC2_DOB, CC1_DI,
         CC2_DI, DP_COMP, DN_COMP, DN_FAULT, LFOSC_ENB, VPP_OTP, IO_RSTB5,
         V1P1, ANAP_TS, TS_ANA_R, ANAP_GP1, GP1_ANA_R, ANAP_GP2, GP2_ANA_R,
         ANAP_GP3, GP3_ANA_R, ANAP_GP4, GP4_ANA_R, ANAP_GP5, GP5_ANA_R, DI_TST,
         DI_TS, SRAM_CLK, PMEM_RE, PMEM_PGM, PMEM_CSB, do_ccctl_0_,
         do_srcctl_0, tm_atpg, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17;
  wire   [10:0] SRAM_A;
  wire   [7:0] SRAM_D;
  wire   [7:0] ANAOPT;
  wire   [1:0] FSW;
  wire   [1:0] RP_EN;
  wire   [1:0] VCONN_EN;
  wire   [17:0] SAMPL_SEL;
  wire   [4:0] DUMMY_IN;
  wire   [55:0] REGTRM;
  wire   [7:0] PWR_I;
  wire   [1:0] OVP_SEL;
  wire   [1:0] CC_SLOPE;
  wire   [5:0] DAC3_V;
  wire   [10:0] DAC0;
  wire   [3:0] ANA_TM;
  wire   [9:0] DAC1;
  wire   [1:0] RP_SEL;
  wire   [1:0] IE_GPIO;
  wire   [6:0] DI_GPIO;
  wire   [6:0] OE_GPIO;
  wire   [6:0] DO_GPIO;
  wire   [6:0] PU_GPIO;
  wire   [6:0] PD_GPIO;
  wire   [3:0] DO_TS;
  wire   [1:0] PMEM_CLK;
  wire   [7:0] PMEM_Q1;
  wire   [7:0] PMEM_Q0;
  wire   [1:0] PMEM_SAP;
  wire   [1:0] PMEM_TWLB;
  wire   [15:0] PMEM_A;
  wire   [7:0] bck_regx0;
  wire   [7:2] bck_regx1;
  wire   [7:2] do_xana1;
  wire   [7:0] do_xana0;
  wire   [3:0] do_regx_xtm;
  wire   [5:2] do_cvctl;
  wire   [3:0] do_vooc;
  wire   [5:0] do_dpdm;
  wire   [5:4] do_srcctl;
  wire   [7:0] do_cctrx;
  wire   [5:0] di_xanav;
  wire   [5:0] srci;
  tri   CSP;
  tri   CSN;
  tri   VFB;
  tri   COMP;
  tri   SW;
  tri   BST;
  tri   VDRV;
  tri   DP;
  tri   DN;
  tri   CC1;
  tri   CC2;
  tri   TST;
  tri   GPIO_TS;
  tri   SCL;
  tri   SDA;
  tri   GPIO1;
  tri   GPIO2;
  tri   GPIO3;
  tri   GPIO4;
  tri   GPIO5;
  tri   [7:0] xdat_o;

  anatop_1127a0 U0_ANALOG_TOP ( .CC1(CC1), .CC2(CC2), .DP(DP), .DN(DN), .VFB(
        VFB), .CSP(CSP), .CSN(CSN), .COMP(COMP), .SW(SW), .BST(BST), .VDRV(
        VDRV), .LG(LG), .HG(HG), .GATE(GATE), .BST_SET(bck_regx0[0]), 
        .DCM_SEL(bck_regx0[1]), .HGOFF(bck_regx0[2]), .HGON(bck_regx0[4]), 
        .LGOFF(bck_regx0[3]), .LGON(bck_regx0[5]), .EN_DRV(bck_regx0[6]), 
        .FSW(FSW), .EN_OSC(bck_regx1[2]), .MAXDS(bck_regx1[3]), .EN_GM(
        bck_regx1[4]), .EN_ODLDO(bck_regx1[5]), .EN_IBUK(bck_regx1[6]), 
        .EN_CP(do_srcctl_0), .EXT_CP(bck_regx1[7]), .INT_CP(bck_regx0[7]), 
        .ANTI_INRUSH(do_cvctl[5]), .PWREN_HOLD(PWREN_HOLD), .RP_SEL(RP_SEL), 
        .RP1_EN(RP_EN[0]), .RP2_EN(RP_EN[1]), .VCONN1_EN(VCONN_EN[0]), 
        .VCONN2_EN(VCONN_EN[1]), .SGP({do_cctrx[0], do_regx_xtm}), .S20U(
        do_cctrx[1]), .S100U(do_cctrx[2]), .TX_EN(TX_EN), .TX_DAT(TX_DAT), 
        .CC_SEL(do_ccctl_0_), .TRA(do_cctrx[4]), .TFA(do_cctrx[5]), .LSR(
        do_cctrx[6]), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .SEL_RX_TH(do_cctrx[7]), .DAC1_EN(DAC1_EN), .DPDN_SHORT(do_dpdm[0]), .DP_2V7_EN(do_dpdm[4]), 
        .DN_2V7_EN(do_dpdm[3]), .DP_0P6V_EN(do_xana1[3]), .DN_0P6V_EN(
        do_xana1[2]), .DP_DWN_EN(do_dpdm[2]), .DN_DWN_EN(do_dpdm[1]), 
        .CC_SLOPE(CC_SLOPE), .DAC2(PWR_I), .DAC3(DAC3_V), .DAC1(DAC1), .CV2(
        do_xana0[0]), .LFOSC_ENB(LFOSC_ENB), .VO_DISCHG(do_srcctl[4]), 
        .DISCHG_SEL(do_srcctl[5]), .CMP_SEL_VO10(SAMPL_SEL[1]), .CMP_SEL_VO20(
        SAMPL_SEL[10]), .CMP_SEL_GP1(SAMPL_SEL[17]), .CMP_SEL_GP2(
        SAMPL_SEL[16]), .CMP_SEL_GP3(SAMPL_SEL[15]), .CMP_SEL_GP4(
        SAMPL_SEL[14]), .CMP_SEL_GP5(SAMPL_SEL[13]), .CMP_SEL_VIN20(
        SAMPL_SEL[0]), .CMP_SEL_TS(SAMPL_SEL[3]), .CMP_SEL_IS(SAMPL_SEL[2]), 
        .CMP_SEL_CC2(SAMPL_SEL[7]), .CMP_SEL_CC1(SAMPL_SEL[6]), 
        .CMP_SEL_CC2_4(SAMPL_SEL[12]), .CMP_SEL_CC1_4(SAMPL_SEL[11]), 
        .CMP_SEL_DP(SAMPL_SEL[4]), .CMP_SEL_DP_3(SAMPL_SEL[8]), .CMP_SEL_DN(
        SAMPL_SEL[5]), .CMP_SEL_DN_3(SAMPL_SEL[9]), .OCP_EN(do_cvctl[2]), 
        .COMP_O(COMP_O), .CCI2C_EN(CCI2C_EN), .UVP_SEL(do_xana0[7]), .TM(
        ANA_TM), .V5OCP(srci[4]), .RSTB(RSTB), .DAC0(DAC0), .SLEEP(SLEEP), 
        .OSC_LOW(OSC_LOW), .OSC_STOP(OSC_STOP), .PWRDN(PWRDN), .VPP_ZERO(
        VPP_0V), .OSC_O(OSC_O), .RD_DET(RD_DET), .IMP_OSC(IMP_OSC), .DRP_OSC(
        DRP_OSC), .STB_RP(STB_RP), .RD_ENB(RD_ENB), .OCP(srci[1]), .SCP(
        srci[3]), .UVP(srci[0]), .LDO3P9V(LDO3P9V), .VPP_SEL(VPP_SEL), 
        .CC1_DOB(CC1_DOB), .CC2_DOB(CC2_DOB), .CC1_DI(CC1_DI), .CC2_DI(CC2_DI), 
        .OTPI(srci[5]), .OVP_SEL(OVP_SEL), .OVP(srci[2]), .DN_COMP(DN_COMP), 
        .DP_COMP(DP_COMP), .DPDN_VTH(do_xana0[5]), .DPDEN(do_vooc[3]), .DPDO(
        do_vooc[2]), .DPIE(do_dpdm[5]), .DNDEN(do_vooc[1]), .DNDO(do_vooc[0]), 
        .DNIE(do_dpdm[5]), .CP_CLKX2(ANAOPT[7]), .SEL_CONST_OVP(ANAOPT[6]), 
        .LP_EN(ANAOPT[5]), .DNCHK_EN(ANAOPT[3]), .IRP_EN(ANAOPT[2]), .CCFBEN(
        ANAOPT[0]), .REGTRM(REGTRM), .AD_RST(AD_RST), .AD_HOLD(AD_HOLD), 
        .DN_FAULT(DN_FAULT), .SEL_CCGAIN(do_xana0[3]), .VFB_SWB(do_xana0[1]), 
        .CPVSEL(do_xana1[6]), .CLAMPV_EN(do_xana1[5]), .HVNG_CPEN(do_xana1[7]), 
        .OCP_SEL(OCP_SEL), .OCP_80M(di_xanav[1]), .OCP_160M(di_xanav[0]), 
        .DMY_OUT(di_xanav[5:2]), .DMY_IN(DUMMY_IN), .VPP_OTP(VPP_OTP), 
        .RSTB_5(IO_RSTB5), .V1P1(V1P1), .TS_ANA_R(TS_ANA_R), .GP5_ANA_R(
        GP5_ANA_R), .GP4_ANA_R(GP4_ANA_R), .GP3_ANA_R(GP3_ANA_R), .GP2_ANA_R(
        GP2_ANA_R), .GP1_ANA_R(GP1_ANA_R), .TS_ANA_P(ANAP_TS), .GP5_ANA_P(
        ANAP_GP5), .GP4_ANA_P(ANAP_GP4), .GP3_ANA_P(ANAP_GP3), .GP2_ANA_P(
        ANAP_GP2), .GP1_ANA_P(ANAP_GP1) );
  IODMURUDA_A0 PAD_SCL ( .DO(DO_GPIO[0]), .IE(IE_GPIO[1]), .OE(OE_GPIO[0]), 
        .PD(PD_GPIO[0]), .PU(PU_GPIO[0]), .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(
        SCL), .ANA_R(), .DI(DI_GPIO[0]) );
  IODMURUDA_A0 PAD_SDA ( .DO(DO_GPIO[1]), .IE(IE_GPIO[1]), .OE(OE_GPIO[1]), 
        .PD(PD_GPIO[1]), .PU(PU_GPIO[1]), .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(
        SDA), .ANA_R(), .DI(DI_GPIO[1]) );
  IOBMURUDA_A0 PAD_TST ( .DO(1'b0), .IE(1'b1), .OE(1'b0), .PD(1'b1), .PU(1'b0), 
        .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(TST), .ANA_R(), .DI(DI_TST) );
  IOBMURUDA_A1 PAD_GPIO1 ( .ANA_P(ANAP_GP1), .DO(DO_GPIO[2]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[2]), .PD(PD_GPIO[2]), .PU(PU_GPIO[2]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO1), .ANA_R(GP1_ANA_R), .DI(DI_GPIO[2]) );
  IOBMURUDA_A1 PAD_GPIO2 ( .ANA_P(ANAP_GP2), .DO(DO_GPIO[3]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[3]), .PD(PD_GPIO[3]), .PU(PU_GPIO[3]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO2), .ANA_R(GP2_ANA_R), .DI(DI_GPIO[3]) );
  IOBMURUDA_A1 PAD_GPIO3 ( .ANA_P(ANAP_GP3), .DO(DO_GPIO[4]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[4]), .PD(PD_GPIO[4]), .PU(PU_GPIO[4]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO3), .ANA_R(GP3_ANA_R), .DI(DI_GPIO[4]) );
  IOBMURUDA_A1 PAD_GPIO4 ( .ANA_P(ANAP_GP4), .DO(DO_GPIO[5]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[5]), .PD(PD_GPIO[5]), .PU(PU_GPIO[5]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO4), .ANA_R(GP4_ANA_R), .DI(DI_GPIO[5]) );
  IOBMURUDA_A1 PAD_GPIO5 ( .ANA_P(ANAP_GP5), .DO(DO_GPIO[6]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[6]), .PD(PD_GPIO[6]), .PU(PU_GPIO[6]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO5), .ANA_R(GP5_ANA_R), .DI(DI_GPIO[6]) );
  IOBMURUDA_A1 PAD_GPIO_TS ( .ANA_P(ANAP_TS), .DO(DO_TS[3]), .IE(IE_GPIO[0]), 
        .OE(DO_TS[2]), .PD(DO_TS[0]), .PU(DO_TS[1]), .RSTB_5(IO_RSTB5), .VB(
        V1P1), .PAD(GPIO_TS), .ANA_R(TS_ANA_R), .DI(DI_TS) );
  MSL18B_1536X8_RW10TM4_16_20221107 U0_SRAM ( .A(SRAM_A), .DI(SRAM_D), .DO(
        xdat_o), .CK(SRAM_CLK), .WEB(SRAM_WEB), .CSB(SRAM_CEB), .OEB(SRAM_OEB)
         );
  ATO0008KX8MX180LBX4DA U0_CODE_0_ ( .A(PMEM_A), .TWLB(PMEM_TWLB), .Q(PMEM_Q0), 
        .SAP(PMEM_SAP), .CSB(PMEM_CSB), .CLK(PMEM_CLK[0]), .PGM(PMEM_PGM), 
        .RE(PMEM_RE), .VDDP(VPP_OTP), .VDD(), .VSS() );
  ATO0008KX8MX180LBX4DA U0_CODE_1_ ( .A(PMEM_A), .TWLB(PMEM_TWLB), .Q(PMEM_Q1), 
        .SAP(PMEM_SAP), .CSB(PMEM_CSB), .CLK(PMEM_CLK[1]), .PGM(PMEM_PGM), 
        .RE(PMEM_RE), .VDDP(VPP_OTP), .VDD(), .VSS() );
  core_a0 U0_CORE ( .SRCI(srci), .XANAV(di_xanav), .BCK_REGX({bck_regx1, FSW, 
        bck_regx0}), .ANA_REGX({do_xana1[7:5], SYNOPSYS_UNCONNECTED_1, 
        do_xana1[3:2], SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        do_xana0[7], SYNOPSYS_UNCONNECTED_4, do_xana0[5], 
        SYNOPSYS_UNCONNECTED_5, do_xana0[3], SYNOPSYS_UNCONNECTED_6, 
        do_xana0[1:0]}), .LFOSC_ENB(LFOSC_ENB), .STB_RP(STB_RP), .RD_ENB(
        RD_ENB), .OCP_SEL(OCP_SEL), .PWREN_HOLD(PWREN_HOLD), .CC1_DI(CC1_DI), 
        .CC2_DI(CC2_DI), .DRP_OSC(DRP_OSC), .IMP_OSC(IMP_OSC), .CC1_DOB(
        CC1_DOB), .CC2_DOB(CC2_DOB), .DAC1_EN(DAC1_EN), .SH_RST(AD_RST), 
        .SH_HOLD(AD_HOLD), .LDO3P9V(LDO3P9V), .XTM(do_regx_xtm), .DO_CVCTL({
        OVP_SEL, do_cvctl[5], SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        do_cvctl[2], SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10}), 
        .DO_CCTRX({do_cctrx[7:4], SYNOPSYS_UNCONNECTED_11, do_cctrx[2:0]}), 
        .DO_SRCCTL({CC_SLOPE, do_srcctl, VCONN_EN, SYNOPSYS_UNCONNECTED_12, 
        do_srcctl_0}), .DO_CCCTL({RP_EN, RP_SEL, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, do_ccctl_0_}), 
        .DO_DAC0(DAC0), .DO_DPDN(do_dpdm), .DO_VOOC(do_vooc), .DO_PWR_I(PWR_I), 
        .PMEM_A(PMEM_A), .PMEM_Q0(PMEM_Q0), .PMEM_Q1(PMEM_Q1), .PMEM_TWLB(
        PMEM_TWLB), .PMEM_SAP(PMEM_SAP), .PMEM_CLK(PMEM_CLK), .PMEM_CSB(
        PMEM_CSB), .PMEM_RE(PMEM_RE), .PMEM_PGM(PMEM_PGM), .VPP_SEL(VPP_SEL), 
        .VPP_0V(VPP_0V), .SRAM_WEB(SRAM_WEB), .SRAM_CEB(SRAM_CEB), .SRAM_OEB(
        SRAM_OEB), .SRAM_CLK(SRAM_CLK), .SRAM_A(SRAM_A), .SRAM_D(SRAM_D), 
        .SRAM_RDAT(xdat_o), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .RD_DET(RD_DET), 
        .TX_DAT(TX_DAT), .TX_EN(TX_EN), .OSC_STOP(OSC_STOP), .OSC_LOW(OSC_LOW), 
        .SLEEP(SLEEP), .PWRDN(PWRDN), .OCDRV_ENZ(), .DAC1_V(DAC1), .SAMPL_SEL(
        SAMPL_SEL), .DAC1_COMP(COMP_O), .CCI2C_EN(CCI2C_EN), .ANA_TM(ANA_TM), 
        .DM_FAULT(DN_FAULT), .DM_COMP(DN_COMP), .DP_COMP(DP_COMP), .DI_GPIO(
        DI_GPIO), .DO_GPIO(DO_GPIO), .OE_GPIO(OE_GPIO), .GPIO_PU(PU_GPIO), 
        .GPIO_PD(PD_GPIO), .GPIO_IE(IE_GPIO), .DO_TS(DO_TS), .DI_TS(DI_TS), 
        .REGTRM(REGTRM), .ANAOPT({ANAOPT[7:5], SYNOPSYS_UNCONNECTED_16, 
        ANAOPT[3:2], SYNOPSYS_UNCONNECTED_17, ANAOPT[0]}), .DUMMY_IN(DUMMY_IN), 
        .DAC3_V(DAC3_V), .i_clk(OSC_O), .i_rstz(RSTB), .atpg_en(tm_atpg), 
        .di_tst(DI_TST), .tm_atpg(tm_atpg) );
endmodule


module core_a0 ( SRCI, XANAV, BCK_REGX, ANA_REGX, LFOSC_ENB, STB_RP, RD_ENB, 
        OCP_SEL, PWREN_HOLD, CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, CC1_DOB, 
        CC2_DOB, DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, XTM, DO_CVCTL, DO_CCTRX, 
        DO_SRCCTL, DO_CCCTL, DO_DAC0, DO_DPDN, DO_VOOC, DO_PWR_I, PMEM_A, 
        PMEM_Q0, PMEM_Q1, PMEM_TWLB, PMEM_SAP, PMEM_CLK, PMEM_CSB, PMEM_RE, 
        PMEM_PGM, VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, 
        SRAM_A, SRAM_D, SRAM_RDAT, RX_DAT, RX_SQL, RD_DET, TX_DAT, TX_EN, 
        OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, DAC1_V, SAMPL_SEL, 
        DAC1_COMP, CCI2C_EN, ANA_TM, DM_FAULT, DM_COMP, DP_COMP, DI_GPIO, 
        DO_GPIO, OE_GPIO, GPIO_PU, GPIO_PD, GPIO_IE, DO_TS, DI_TS, REGTRM, 
        ANAOPT, DUMMY_IN, DAC3_V, i_clk, i_rstz, atpg_en, di_tst, tm_atpg );
  input [5:0] SRCI;
  input [5:0] XANAV;
  output [15:0] BCK_REGX;
  output [15:0] ANA_REGX;
  output [3:0] XTM;
  output [7:0] DO_CVCTL;
  output [7:0] DO_CCTRX;
  output [7:0] DO_SRCCTL;
  output [7:0] DO_CCCTL;
  output [10:0] DO_DAC0;
  output [5:0] DO_DPDN;
  output [3:0] DO_VOOC;
  output [7:0] DO_PWR_I;
  output [15:0] PMEM_A;
  input [7:0] PMEM_Q0;
  input [7:0] PMEM_Q1;
  output [1:0] PMEM_TWLB;
  output [1:0] PMEM_SAP;
  output [1:0] PMEM_CLK;
  output [10:0] SRAM_A;
  output [7:0] SRAM_D;
  input [7:0] SRAM_RDAT;
  output [9:0] DAC1_V;
  output [17:0] SAMPL_SEL;
  output [3:0] ANA_TM;
  input [6:0] DI_GPIO;
  output [6:0] DO_GPIO;
  output [6:0] OE_GPIO;
  output [6:0] GPIO_PU;
  output [6:0] GPIO_PD;
  output [1:0] GPIO_IE;
  output [3:0] DO_TS;
  output [55:0] REGTRM;
  output [7:0] ANAOPT;
  output [4:0] DUMMY_IN;
  output [5:0] DAC3_V;
  input CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, RX_DAT, RX_SQL, RD_DET, DAC1_COMP,
         DM_FAULT, DM_COMP, DP_COMP, DI_TS, i_clk, i_rstz, atpg_en, di_tst;
  output LFOSC_ENB, STB_RP, RD_ENB, OCP_SEL, PWREN_HOLD, CC1_DOB, CC2_DOB,
         DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, PMEM_CSB, PMEM_RE, PMEM_PGM,
         VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, TX_DAT,
         TX_EN, OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, CCI2C_EN, tm_atpg;
  wire   N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N268, n675, n676, n677, n678, n679, aswclk, detclk, tclk_sel, s_clk,
         aswkup, x_clk, t_di_gpio4, t_pmem_clk, pmem_csb, t_pmem_csb,
         r_osc_gate, t_osc_gate, g_clk, xram_ce, iram_ce, sram_en, r_i2c_attr,
         esfrm_oe, esfrm_we, sfrack, ictlr_psrack, esfrm_rrdy, memwr, memrd,
         memrd_c, memack, o_cpurst, hit_xd, hit_xr, hit_ps, hit_ps_c,
         mcu_ram_r, mcu_ram_w, regx_re, iram_we, xram_we, regx_we, bist_en,
         bist_wr, srstz, prl_cany0w, prl_cany0r, mempsrd, r_bclk_sel,
         r_hold_mcu, t0_intr, fcp_intr, dpdm_urx, s0_rxdoe, mcuo_scl, mcuo_sda,
         mempsack, mempswr, mempsrd_c, sfr_w, sfr_r, ictlr_psack, ictlr_inc,
         set_hold, bkpt_hold, bkpt_ena, r_psrd, r_pswr, prl_cany0, prl_c0set,
         pmem_pgm, pmem_re, we_twlb, r_otp_wpls, pwrdn_rst, r_otp_pwdn_en,
         ramacc, frc_lg_on, gating_pwr, cc1_di, cc2_di, r_sleep, ps_pwrdn,
         r_pwrdn, r_ocdrv_enz, r_osc_stop, r_pwrv_upd, r_otpi_gate, r_fcpre,
         r_fortxdat, r_fortxrdy, r_fortxen, r_gpio_tm, pid_goidle, pid_gobusy,
         bus_idle, sse_idle, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop,
         r_unlock, r_first, r_last, r_fiforst, r_set_cpmsgid, r_txendk,
         r_txshrt, r_auto_discard, r_dat_portrole, r_dat_datarole, r_pshords,
         r_discard, r_strtch, r_i2c_ninc, r_i2c_fwnak, r_i2c_fwack,
         hwi2c_stretch, i2c_ev_6_, i2c_ev_3, i2c_ev_2, prl_discard,
         prl_GCTxDone, pff_obsd, pff_empty, pff_full, ptx_ack, clk_1p0m,
         clk_500, prstz, sse_rdrdy, upd_rdrdy, sse_prefetch, slvo_sda, slvo_re,
         slvo_early, dm_comp, dp_comp, di_sqlch, ptx_cc, ptx_oe, sh_rst,
         sh_hold, fcp_oe, fcp_do, sdischg_duty, clk_100k, r_bck2_2_, r_imp_osc,
         clk_500k, r_vpp_en, r_vpp0v_en, di_ts, di_aswk_0, r_xana_23,
         r_xana_19, r_xana_18, divff_o1, clk_50k, do_opt_1, do_opt_0, N448,
         o_dodat0_15_, o_dodat5_2_, N568, N569, N570, N571, N572, N575, N576,
         N577, N578, N579, N580, N581, N582, N583, N584, N593, N594, N595,
         N596, N598, N599, N600, N601, N603, N606, N607, N608, N627, N628,
         N629, N630, N632, N633, N634, N635, N637, N640, N641, N642, N1478,
         N1483, net8853, n28, n29, n30, n76, n117, n123, n126, n128, n129,
         n131, n133, n135, n137, n138, n140, n147, n160, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n181, n182, n183,
         n184, n186, n188, n190, n192, n193, n195, n197, n199, n200, n214,
         n217, n218, n220, n223, n224, n226, n227, n229, n230, n232, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n254, n255, n258, n259, n260, n261,
         n264, n265, n266, n267, n270, n271, n272, n273, n274, n277, n278,
         n279, n282, n283, n287, n288, n289, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n444, n445, n447, n472, n493, n494, n495, n496, n497, n498,
         n504, n505, n506, n508, n509, n510, n511, sll_232_2_A_0_, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n41, n42, n44, n45, n46, n47, n48, n49, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n118, n119, n120, n121,
         n122, n124, n125, n127, n130, n132, n134, n136, n139, n141, n143,
         n144, n146, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n161, n162, n163, n164, n165, n166, n167, n168,
         n180, n185, n187, n189, n191, n194, n196, n198, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n215,
         n216, n219, n221, n222, n225, n228, n231, n233, n234, n252, n253,
         n256, n257, n262, n263, n268, n269, n275, n276, n280, n281, n284,
         n285, n286, n290, n291, n357, n393, n443, n446, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n499, n500, n501,
         n502, n503, n507, n512, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109;
  wire   [9:0] aswclk_ps;
  wire   [9:0] detclk_ps;
  wire   [1:0] pmem_clk;
  wire   [7:0] sse_wdat;
  wire   [7:0] prx_fifowdat;
  wire   [7:0] sse_adr;
  wire   [7:0] prl_cany0adr;
  wire   [7:0] esfrm_wdat;
  wire   [6:0] esfrm_adr;
  wire   [7:0] mcu_esfrrdat;
  wire   [7:0] delay_inst;
  wire   [7:0] esfrm_rdat;
  wire   [3:0] r_pg0_sel;
  wire   [15:0] memaddr;
  wire   [15:0] memaddr_c;
  wire   [7:0] memdatao;
  wire   [7:0] idat_adr;
  wire   [7:0] idat_wdat;
  wire   [10:0] iram_a;
  wire   [10:0] xram_a;
  wire   [7:0] iram_d;
  wire   [7:0] xram_d;
  wire   [1:0] sram_rdat;
  wire   [7:0] regx_rdat;
  wire   [10:0] bist_adr;
  wire   [7:0] bist_wdat;
  wire   [7:0] memdatai;
  wire   [7:0] ictlr_inst;
  wire   [15:0] mcu_pc;
  wire   [22:16] mcu_dbgpo;
  wire   [3:2] sfr_intr;
  wire   [7:0] exint;
  wire   [7:0] ff_p0;
  wire   [6:0] do_p0;
  wire   [7:0] sfr_rdat;
  wire   [7:0] sfr_wdat;
  wire   [6:0] sfr_adr;
  wire   [14:0] bkpt_pc;
  wire   [14:0] r_inst_ofs;
  wire   [7:0] pmem_q0;
  wire   [7:0] pmem_q1;
  wire   [1:0] pmem_twlb;
  wire   [1:0] wd_twlb;
  wire   [1:0] r_sqlch;
  wire   [3:2] r_ccrx;
  wire   [1:0] r_rxdb_opt;
  wire   [7:4] r_pwrctl;
  wire   [5:2] di_pro;
  wire   [1:0] lg_pulse_len;
  wire   [7:0] r_srcctl;
  wire   [7:0] r_dpdmctl;
  wire   [11:0] r_fw_pwrv;
  wire   [5:0] r_cvcwr;
  wire   [15:0] r_cvofs;
  wire   [7:0] r_cctrx;
  wire   [7:0] r_ccctl;
  wire   [6:0] r_fcpwr;
  wire   [7:0] fcp_r_dat;
  wire   [7:0] fcp_r_sta;
  wire   [7:0] fcp_r_msk;
  wire   [7:0] fcp_r_ctl;
  wire   [7:0] fcp_r_crc;
  wire   [7:0] fcp_r_acc;
  wire   [7:0] fcp_r_tui;
  wire   [7:0] r_accctl;
  wire   [7:5] r_comp_opt;
  wire   [14:0] sfr_dacwr;
  wire   [17:0] r_dac_en;
  wire   [17:0] r_sar_en;
  wire   [7:0] r_isofs;
  wire   [7:0] r_adofs;
  wire   [7:0] dac_r_ctl;
  wire   [7:0] dac_r_cmpsta;
  wire   [17:0] dac_r_comp;
  wire   [143:0] dac_r_vs;
  wire   [5:0] x_daclsb;
  wire   [6:0] REVID;
  wire   [6:0] r_pu_gpio;
  wire   [6:0] r_pd_gpio;
  wire   [6:0] r_gpio_oe;
  wire   [1:0] r_gpio_ie;
  wire   [55:0] r_regtrm;
  wire   [3:0] r_ana_tm;
  wire   [7:0] i2c_ltbuf;
  wire   [7:0] i2c_lt_ofs;
  wire   [4:0] r_txnumk;
  wire   [1:0] r_auto_gdcrc;
  wire   [1:0] r_spec;
  wire   [1:0] r_dat_spec;
  wire   [6:0] r_txauto;
  wire   [6:0] r_rxords_ena;
  wire   [7:1] r_i2c_deva;
  wire   [2:0] prl_cpmsgid;
  wire   [1:0] pff_ack;
  wire   [7:0] pff_rdat;
  wire   [15:0] pff_rxpart;
  wire   [5:0] pff_ptr;
  wire   [6:0] prx_setsta;
  wire   [1:0] prx_rst;
  wire   [4:0] prx_rcvinf;
  wire   [5:0] prx_adpn;
  wire   [3:0] prx_fsm;
  wire   [2:0] ptx_fsm;
  wire   [3:0] prl_fsm;
  wire   [3:0] slvo_ev;
  wire   [1:0] r_i2cslv_route;
  wire   [5:4] r_i2crout;
  wire   [1:0] r_i2cmcu_route;
  wire   [18:17] upd_dbgpo;
  wire   [7:0] r_dacwdat;
  wire   [17:8] wr_dacv;
  wire   [10:7] r_dacwr;
  wire   [17:0] dacmux_sel;
  wire   [3:0] comp_smpl;
  wire   [7:0] r_cvcwdat;
  wire   [7:0] r_sdischg;
  wire   [7:0] r_vcomp;
  wire   [7:0] r_idacsh;
  wire   [7:0] r_cvofsx;
  wire   [7:0] r_xtm;
  wire   [6:0] bist_r_ctl;
  wire   [1:0] regx_hitbst;
  wire   [7:0] bist_r_dat;
  wire   [1:0] regx_wrpwm;
  wire   [15:0] r_pwm;
  wire   [1:0] r_sap;
  wire   [3:0] lt_gpi;
  wire   [6:0] r_do_ts;
  wire   [3:0] r_dpdo_sel;
  wire   [3:0] r_dndo_sel;
  wire   [4:2] di_aswk;
  wire   [7:0] r_bck0;
  wire   [7:0] r_bck1;
  wire   [15:0] r_xana;
  wire   [5:0] di_xanav;
  wire   [7:0] r_aopt;
  wire   [6:0] di_gpio;
  wire   [7:6] do_opt;
  wire   [1:0] pwm_o;
  wire   [15:0] d_dodat;
  wire   [3:0] r_lt_gpi;
  tri   [7:0] SRAM_RDAT;

  CKBUFX1 U0_ASWCLK_BUF_0_ ( .A(aswclk_ps[0]), .Y(aswclk_ps[1]) );
  CKBUFX1 U0_ASWCLK_BUF_1_ ( .A(aswclk_ps[1]), .Y(aswclk_ps[2]) );
  CKBUFX1 U0_ASWCLK_BUF_2_ ( .A(aswclk_ps[2]), .Y(aswclk_ps[3]) );
  CKBUFX1 U0_ASWCLK_BUF_3_ ( .A(aswclk_ps[3]), .Y(aswclk_ps[4]) );
  CKBUFX1 U0_ASWCLK_BUF_4_ ( .A(aswclk_ps[4]), .Y(aswclk_ps[5]) );
  CKBUFX1 U0_ASWCLK_BUF_5_ ( .A(aswclk_ps[5]), .Y(aswclk_ps[6]) );
  CKBUFX1 U0_ASWCLK_BUF_6_ ( .A(aswclk_ps[6]), .Y(aswclk_ps[7]) );
  CKBUFX1 U0_ASWCLK_BUF_7_ ( .A(aswclk_ps[7]), .Y(aswclk_ps[8]) );
  CKBUFX1 U0_ASWCLK_BUF_8_ ( .A(aswclk_ps[8]), .Y(aswclk_ps[9]) );
  CKBUFX1 U0_ASWCLK_BUF_9_ ( .A(aswclk_ps[9]), .Y(aswclk) );
  CKBUFX1 U0_DETCLK_BUF_0_ ( .A(detclk_ps[0]), .Y(detclk_ps[1]) );
  CKBUFX1 U0_DETCLK_BUF_1_ ( .A(detclk_ps[1]), .Y(detclk_ps[2]) );
  CKBUFX1 U0_DETCLK_BUF_2_ ( .A(detclk_ps[2]), .Y(detclk_ps[3]) );
  CKBUFX1 U0_DETCLK_BUF_3_ ( .A(detclk_ps[3]), .Y(detclk_ps[4]) );
  CKBUFX1 U0_DETCLK_BUF_4_ ( .A(detclk_ps[4]), .Y(detclk_ps[5]) );
  CKBUFX1 U0_DETCLK_BUF_5_ ( .A(detclk_ps[5]), .Y(detclk_ps[6]) );
  CKBUFX1 U0_DETCLK_BUF_6_ ( .A(detclk_ps[6]), .Y(detclk_ps[7]) );
  CKBUFX1 U0_DETCLK_BUF_7_ ( .A(detclk_ps[7]), .Y(detclk_ps[8]) );
  CKBUFX1 U0_DETCLK_BUF_8_ ( .A(detclk_ps[8]), .Y(detclk_ps[9]) );
  CKBUFX1 U0_DETCLK_BUF_9_ ( .A(detclk_ps[9]), .Y(detclk) );
  AND2X1 U0_SCAN_EN ( .A(DI_GPIO[2]), .B(n107), .Y() );
  CKMUX2X1 U0_CLK_MUX ( .D0(i_clk), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(s_clk)
         );
  CKMUX2X1 U0_DCLKMUX ( .D0(RD_DET), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        detclk_ps[0]) );
  CKMUX2X1 U0_ACLKMUX ( .D0(aswkup), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        aswclk_ps[0]) );
  CKBUFX1 U0_MCK_BUF ( .A(i_clk), .Y(x_clk) );
  CKBUFX1 U0_TCK_BUF ( .A(DI_GPIO[4]), .Y(t_di_gpio4) );
  CKBUFX1 U0_BUF_NEG0 ( .A(pmem_clk[0]), .Y(t_pmem_clk) );
  CKBUFX1 U0_BUF_NEG1 ( .A(pmem_csb), .Y(t_pmem_csb) );
  CKBUFX1 U0_BUF_NEG2 ( .A(r_osc_gate), .Y(t_osc_gate) );
  CLKDLX1 U0_MCLK_ICG ( .CK(s_clk), .E(n644), .SE(n136), .ECK(g_clk) );
  CLKDLX1 U0_SRAM_ICG ( .CK(g_clk), .E(sram_en), .SE(n136), .ECK(SRAM_CLK) );
  INVX1 U0_REVIDZ_0_ ( .A(1'b0), .Y(REVID[0]) );
  INVX1 U0_REVIDZ_1_ ( .A(1'b1), .Y(REVID[1]) );
  INVX1 U0_REVIDZ_2_ ( .A(1'b1), .Y(REVID[2]) );
  INVX1 U0_REVIDZ_3_ ( .A(1'b1), .Y(REVID[3]) );
  INVX1 U0_REVIDZ_4_ ( .A(1'b0), .Y(REVID[4]) );
  INVX1 U0_REVIDZ_5_ ( .A(1'b0), .Y(REVID[5]) );
  INVX1 U0_REVIDZ_6_ ( .A(1'b1), .Y(REVID[6]) );
  mpb_a0 u0_mpb ( .i_rd({prl_cany0r, n76}), .i_wr({prl_cany0w, i2c_ev_3}), 
        .wdat0(sse_wdat), .wdat1(prx_fifowdat), .addr0(sse_adr), .addr1(
        prl_cany0adr), .r_i2c_attr(r_i2c_attr), .esfrm_oe(esfrm_oe), 
        .esfrm_we(esfrm_we), .sfrack(sfrack), .esfrm_wdat(esfrm_wdat), 
        .esfrm_adr(esfrm_adr), .mcu_esfr_rdat(mcu_esfrrdat), .delay_rdat(
        delay_inst), .delay_rrdy(ictlr_psrack), .esfrm_rrdy(esfrm_rrdy), 
        .esfrm_rdat(esfrm_rdat), .channel_sel(1'b0), .r_pg0_sel(r_pg0_sel), 
        .dma_w(1'b0), .dma_r(1'b0), .dma_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_wdat({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_ack(), .memaddr(memaddr), 
        .memaddr_c(memaddr_c), .memwr(memwr), .memrd(memrd), .memrd_c(memrd_c), 
        .cpurst(o_cpurst), .memdatao(memdatao), .memack(memack), .hit_xd(
        hit_xd), .hit_xr(hit_xr), .hit_ps(hit_ps), .hit_ps_c(hit_ps_c), 
        .idat_r(mcu_ram_r), .idat_w(mcu_ram_w), .idat_adr(idat_adr), 
        .idat_wdat(idat_wdat), .iram_ce(iram_ce), .xram_ce(xram_ce), .regx_re(
        regx_re), .iram_we(iram_we), .xram_we(xram_we), .regx_we(regx_we), 
        .iram_a(iram_a), .xram_a(xram_a), .iram_d(iram_d), .xram_d(xram_d), 
        .iram_rdat({n129, n131, n133, n135, n138, n140, sram_rdat}), 
        .xram_rdat({n129, n131, n133, n135, n138, n140, sram_rdat}), 
        .regx_rdat({n14, regx_rdat[6:0]}), .bist_en(n38), .bist_wr(bist_wr), 
        .bist_adr(bist_adr), .bist_wdat(bist_wdat), .bist_xram(1'b0), .mclk(
        g_clk), .srstz(srstz) );
  mcu51_a0 u0_mcu ( .bclki2c(r_bclk_sel), .pc_ini({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .slp2wakeup(1'b0), .r_hold_mcu(r_hold_mcu), .wdt_slow(1'b0), .wdtov({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}), .mdubsy(), .cs_run(), 
        .t0_intr(t0_intr), .clki2c(g_clk), .clkmdu(g_clk), .clkur0(g_clk), 
        .clktm0(g_clk), .clktm1(g_clk), .clkwdt(g_clk), .i2c_autoack(1'b0), 
        .i2c_con_ens1(), .clkcpu(g_clk), .clkper(g_clk), .reset(n84), .ro(
        o_cpurst), .port0i({n4, di_gpio[6:4], n137, di_gpio[2:0]}), .exint_9(
        fcp_intr), .exint({exint[7:4], n30, n29, exint[1:0]}), .clkcpuen(), 
        .clkperen(), .port0o({SYNOPSYS_UNCONNECTED_3, do_p0}), .port0ff(ff_p0), 
        .rxd0o(do_opt[7]), .txd0(do_opt[6]), .rxd0i(dpdm_urx), .rxd0oe(
        s0_rxdoe), .scli(n509), .sdai(n511), .sclo(mcuo_scl), .sdao(mcuo_sda), 
        .waitstaten(), .mempsack(mempsack), .memack(memack), .memdatai(
        memdatai), .memdatao(memdatao), .memaddr(memaddr), .mempswr(mempswr), 
        .mempsrd(mempsrd), .memwr(memwr), .memrd(memrd), .memdatao_comb({
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11}), .memaddr_comb(
        memaddr_c), .mempswr_comb(), .mempsrd_comb(mempsrd_c), .memwr_comb(), 
        .memrd_comb(memrd_c), .ramdatai({n129, n131, n133, n135, n138, n140, 
        sram_rdat}), .ramdatao(idat_wdat), .ramaddr(idat_adr), .ramwe(
        mcu_ram_w), .ramoe(mcu_ram_r), .dbgpo({SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, mcu_dbgpo, mcu_pc}), 
        .sfrack(sfrack), .sfrdatai(sfr_rdat), .sfrdatao(sfr_wdat), .sfraddr(
        sfr_adr), .sfrwe(sfr_w), .sfroe(sfr_r), .esfrm_wrdata(esfrm_wdat), 
        .esfrm_addr(esfrm_adr), .esfrm_we(esfrm_we), .esfrm_oe(esfrm_oe), 
        .esfrm_rddata(mcu_esfrrdat) );
  ictlr_a0 u0_ictlr ( .bkpt_ena(bkpt_ena), .bkpt_pc(bkpt_pc), .memaddr_c({
        memaddr_c[14:7], n27, n33, n21, n31, n24, n13, n25}), .memaddr(
        memaddr[14:0]), .mcu_psr_c(mempsrd_c), .mcu_psw(mempswr), .hit_ps_c(
        hit_ps_c), .hit_ps(hit_ps), .mempsack(ictlr_psack), .memdatao(memdatao), .o_set_hold(set_hold), .o_bkp_hold(bkpt_hold), .o_ofs_inc(ictlr_inc), 
        .o_inst(ictlr_inst), .d_inst(delay_inst), .sfr_psrack(ictlr_psrack), 
        .sfr_psofs(r_inst_ofs), .sfr_psr(r_psrd), .sfr_psw(r_pswr), .dw_rst(
        prl_c0set), .dw_ena(prl_cany0), .sfr_wdat({n80, n78, n75, n72, n70, 
        n67, n64, n61}), .pmem_pgm(pmem_pgm), .pmem_re(pmem_re), .pmem_csb(
        pmem_csb), .pmem_clk(pmem_clk), .pmem_a(PMEM_A), .pmem_q0(pmem_q0), 
        .pmem_q1(pmem_q1), .pmem_twlb(pmem_twlb), .wd_twlb(wd_twlb), .we_twlb(
        we_twlb), .pwrdn_rst(pwrdn_rst), .r_pwdn_en(r_otp_pwdn_en), .r_multi(
        r_otp_wpls), .r_hold_mcu(r_hold_mcu), .clk(g_clk), .srst(o_cpurst) );
  regbank_a0 u0_regbank ( .srci({di_pro[5], n531, n532, di_pro[2], n126, n128}), .lg_pulse_len(lg_pulse_len), .dm_fault(n117), .cc1_di(cc1_di), .cc2_di(
        cc2_di), .di_rd_det(di_aswk[2]), .i_tmrf(t0_intr), .i_vcbyval(r_xtm[4]), .dnchk_en(o_dodat5_2_), .r_pwrv_upd(r_pwrv_upd), .aswkup(aswkup), 
        .lg_dischg(frc_lg_on), .gating_pwr(gating_pwr), .ps_pwrdn(ps_pwrdn), 
        .r_sleep(r_sleep), .r_pwrdn(r_pwrdn), .r_ocdrv_enz(r_ocdrv_enz), 
        .r_osc_stop(r_osc_stop), .r_osc_lo(o_dodat0_15_), .r_osc_gate(
        r_osc_gate), .r_fw_pwrv(r_fw_pwrv), .r_cvcwr(r_cvcwr[1:0]), .r_cvofs(
        r_cvofs), .r_otpi_gate(r_otpi_gate), .r_pwrctl(r_pwrctl), .r_pwr_i(
        DO_PWR_I), .r_cvctl(DO_CVCTL), .r_srcctl(r_srcctl), .r_dpdmctl(
        r_dpdmctl), .r_ccrx({r_sqlch, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, r_ccrx, r_rxdb_opt}), .r_cctrx(r_cctrx), 
        .r_ccctl(r_ccctl), .r_fcpwr(r_fcpwr), .r_fcpre(r_fcpre), .fcp_r_dat(
        fcp_r_dat), .fcp_r_sta(fcp_r_sta), .fcp_r_msk(fcp_r_msk), .fcp_r_ctl(
        fcp_r_ctl), .fcp_r_crc(fcp_r_crc), .fcp_r_acc(fcp_r_acc), .fcp_r_tui(
        fcp_r_tui), .r_accctl(r_accctl), .r_bclk_sel(r_bclk_sel), .r_dacwr(
        sfr_dacwr), .r_dac_en({r_dac_en[7:4], n49, r_dac_en[2:0]}), .r_sar_en(
        r_sar_en[7:0]), .r_adofs({r_adofs[7:6], n48, n47, n42, n46, n45, 
        r_adofs[0]}), .r_isofs(r_isofs), .x_daclsb(x_daclsb), .r_comp_opt({
        r_comp_opt, SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27}), .dac_r_ctl(dac_r_ctl), .dac_r_comp(
        dac_r_comp[7:0]), .dac_r_cmpsta(dac_r_cmpsta), .dac_r_vs(
        dac_r_vs[63:0]), .REVID(REVID), .atpg_en(n104), .sfr_r(sfr_r), .sfr_w(
        sfr_w), .set_hold(set_hold), .bkpt_hold(bkpt_hold), .cpurst(o_cpurst), 
        .sfr_addr({1'b1, sfr_adr}), .sfr_wdat({n80, n78, n74, n72, n69, n66, 
        n63, n60}), .sfr_rdat(sfr_rdat), .ff_p0(ff_p0), .di_p0({n4, 
        di_gpio[6:4], n137, di_gpio[2:0]}), .ictlr_idle(pmem_csb), .ictlr_inc(
        ictlr_inc), .r_inst_ofs(r_inst_ofs), .r_psrd(r_psrd), .r_pswr(r_pswr), 
        .r_fortxdat(r_fortxdat), .r_fortxrdy(r_fortxrdy), .r_fortxen(r_fortxen), .r_ana_tm(r_ana_tm), .r_gpio_tm(r_gpio_tm), .r_gpio_ie(r_gpio_ie), 
        .r_gpio_oe(r_gpio_oe), .r_gpio_pu(r_pu_gpio), .r_gpio_pd(r_pd_gpio), 
        .r_gpio_s0({N268, N267, N266}), .r_gpio_s1({N265, N264, N263}), 
        .r_gpio_s2({N262, N261, N260}), .r_gpio_s3({N259, N258, N257}), 
        .r_regtrm(r_regtrm), .i_pc(mcu_pc), .i_goidle(pid_goidle), .i_gobusy(
        pid_gobusy), .i_i2c_idle(sse_idle), .bus_idle(bus_idle), .i2c_stretch(
        hwi2c_stretch), .i_i2c_rwbuf(sse_wdat), .i_i2c_ltbuf(i2c_ltbuf), 
        .i_i2c_ofs(i2c_lt_ofs), .o_intr({exint[6], sfr_intr, exint[5:4]}), 
        .r_auto_gdcrc(r_auto_gdcrc), .r_exist1st(r_exist1st), .r_ordrs4(
        r_ordrs4), .r_fifopsh(r_fifopsh), .r_fifopop(r_fifopop), .r_unlock(
        r_unlock), .r_first(r_first), .r_last(r_last), .r_fiforst(r_fiforst), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_txendk(r_txendk), .r_txnumk(r_txnumk), .r_txshrt(r_txshrt), .r_auto_discard(r_auto_discard), .r_hold_mcu(r_hold_mcu), .r_txauto(r_txauto), .r_rxords_ena(r_rxords_ena), .r_spec(r_spec), 
        .r_dat_spec(r_dat_spec), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_discard(r_discard), .r_pshords(
        r_pshords), .r_pg0_sel(r_pg0_sel), .r_strtch(r_strtch), .r_i2c_attr(
        r_i2c_attr), .r_i2c_ninc(r_i2c_ninc), .r_hwi2c_en(), .r_i2c_fwnak(
        r_i2c_fwnak), .r_i2c_fwack(r_i2c_fwack), .r_i2c_deva(r_i2c_deva), 
        .i2c_ev({n76, i2c_ev_6_, slvo_ev[3:2], i2c_ev_3, i2c_ev_2, 
        slvo_ev[1:0]}), .prl_c0set(prl_c0set), .prl_cany0(prl_cany0), 
        .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_cpmsgid(
        prl_cpmsgid), .pff_ack(pff_ack), .prx_rst(prx_rst), .pff_obsd(pff_obsd), .pff_full(pff_full), .pff_empty(pff_empty), .ptx_ack(ptx_ack), .pff_ptr(
        pff_ptr), .prx_adpn(prx_adpn), .pff_rdat(pff_rdat), .pff_rxpart(
        pff_rxpart), .prx_rcvinf(prx_rcvinf), .ptx_fsm(ptx_fsm), .prx_fsm(
        prx_fsm), .prl_fsm(prl_fsm), .prx_setsta(prx_setsta), .clk_1p0m(
        clk_1p0m), .clk_500(clk_500), .clk(g_clk), .xrstz(i_rstz), .xclk(s_clk), .dbgpo({SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59}), .srstz(srstz), 
        .prstz(prstz) );
  i2cslv_a0 u0_i2cslv ( .i_sda(n510), .i_scl(n508), .o_sda(slvo_sda), .i_deva(
        r_i2c_deva), .i_inc(n28), .i_fwnak(r_i2c_fwnak), .i_fwack(r_i2c_fwack), 
        .o_we(i2c_ev_3), .o_re(slvo_re), .o_r_early(slvo_early), .o_idle(
        sse_idle), .o_dec(), .o_busev(slvo_ev), .o_ofs(sse_adr), .o_lt_ofs(
        i2c_lt_ofs), .o_wdat(sse_wdat), .o_lt_buf(i2c_ltbuf), .o_dbgpo({
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67}), .i_rdat(esfrm_rdat), .i_rd_mem(sse_rdrdy), .i_clk(g_clk), .i_rstz(n83), .i_prefetch(sse_prefetch)
         );
  updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 u0_updphy ( .i_cc(n58), .i_cc_49(n123), 
        .i_sqlch(di_sqlch), .r_sqlch(r_sqlch), .r_adprx_en(r_ccrx[3]), 
        .r_adp2nd(r_ccrx[2]), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), 
        .r_fifopsh(r_fifopsh), .r_fifopop(r_fifopop), .r_fiforst(r_fiforst), 
        .r_unlock(r_unlock), .r_first(r_first), .r_last(r_last), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_rdy(upd_rdrdy), .r_wdat({sfr_wdat[7], 
        n78, n75, n72, n70, n67, n64, n61}), .r_rdat(esfrm_rdat), .r_txnumk(
        r_txnumk), .r_txendk(r_txendk), .r_txshrt(r_txshrt), .r_auto_discard(
        r_auto_discard), .r_txauto(r_txauto), .r_rxords_ena(r_rxords_ena), 
        .r_spec(r_spec), .r_dat_spec(r_dat_spec), .r_auto_gdcrc(r_auto_gdcrc), 
        .r_rxdb_opt(r_rxdb_opt), .r_pshords(r_pshords), .r_dat_portrole(
        r_dat_portrole), .r_dat_datarole(r_dat_datarole), .r_discard(r_discard), .pid_goidle(pid_goidle), .pid_gobusy(pid_gobusy), .pff_ack(pff_ack), 
        .pff_rdat(pff_rdat), .pff_rxpart(pff_rxpart), .prx_rcvinf(prx_rcvinf), 
        .pff_obsd(pff_obsd), .pff_ptr(pff_ptr), .pff_empty(pff_empty), 
        .pff_full(pff_full), .ptx_ack(ptx_ack), .ptx_cc(ptx_cc), .ptx_oe(
        ptx_oe), .prx_setsta(prx_setsta), .prx_rst(prx_rst), .prl_c0set(
        prl_c0set), .prl_cany0(prl_cany0), .prl_cany0r(prl_cany0r), 
        .prl_cany0w(prl_cany0w), .prl_discard(prl_discard), .prl_GCTxDone(
        prl_GCTxDone), .prl_cany0adr(prl_cany0adr), .prl_cpmsgid(prl_cpmsgid), 
        .prx_fifowdat(prx_fifowdat), .ptx_fsm(ptx_fsm), .prl_fsm(prl_fsm), 
        .prx_fsm(prx_fsm), .prx_adpn(prx_adpn), .dbgpo({
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, upd_dbgpo, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97}), .clk(g_clk), 
        .srstz(prstz) );
  dacmux_a0 u0_dacmux ( .clk(g_clk), .srstz(n82), .i_comp(n4), .r_comp_opt(
        r_comp_opt), .r_wdat(r_dacwdat), .r_adofs(r_adofs), .r_isofs(r_isofs), 
        .r_wr({r_dacwr[10], n23, r_dacwr[8:7], sfr_dacwr[14:8]}), .dacv_wr({
        n15, n11, n37, n22, n17, n32, n18, wr_dacv[10], n36, n34, 
        sfr_dacwr[7:0]}), .o_dacv(dac_r_vs), .o_shrst(sh_rst), .o_hold(sh_hold), .o_dac1(DAC1_V), .o_daci_sel(dacmux_sel), .o_dat(dac_r_comp), .r_dac_en(
        r_dac_en), .r_sar_en(r_sar_en), .o_dactl(dac_r_ctl), .o_cmpsta(
        dac_r_cmpsta), .x_daclsb(x_daclsb), .o_intr(exint[7]), .o_smpl({
        SYNOPSYS_UNCONNECTED_98, comp_smpl}) );
  fcp_a0 u0_fcp ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(1'b0), .intr(
        fcp_intr), .tx_en(fcp_oe), .tx_dat(fcp_do), .r_dat(fcp_r_dat), .r_sta(
        fcp_r_sta), .r_ctl(fcp_r_ctl), .r_msk(fcp_r_msk), .r_crc(fcp_r_crc), 
        .r_acc(fcp_r_acc), .r_dpdmsta(r_accctl), .r_wdat({n80, n78, n75, n72, 
        n70, n67, n64, n61}), .r_wr(r_fcpwr), .r_re(r_fcpre), .clk(g_clk), 
        .srstz(n83), .r_tui(fcp_r_tui) );
  cvctl_a0 u0_cvctl ( .r_cvcwr(r_cvcwr), .wdat(r_cvcwdat), .r_sdischg(
        r_sdischg), .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), .r_cvofsx(r_cvofsx), .r_cvofs(r_cvofs), .sdischg_duty(sdischg_duty), .r_hlsb_en(r_pwrctl[4]), 
        .r_hlsb_sel(r_pwrctl[5]), .r_hlsb_freq(r_xtm[5]), .r_hlsb_duty(
        r_xtm[6]), .r_fw_pwrv(r_fw_pwrv), .r_dac0(DO_DAC0), .r_dac3(DAC3_V), 
        .clk_100k(clk_100k), .clk(g_clk), .srstz(n83) );
  regx_a0 u0_regx ( .regx_r(regx_re), .regx_w(regx_we), .di_drposc(di_aswk_0), 
        .di_imposc(di_aswk[4]), .di_rd_det(di_aswk[2]), .clk_500k(clk_500k), 
        .r_imp_osc(r_imp_osc), .regx_addr(xram_a[6:0]), .regx_wdat({
        xram_d[7:1], n85}), .regx_rdat(regx_rdat), .regx_hitbst(regx_hitbst), 
        .regx_wrpwm(regx_wrpwm), .regx_wrcvc({r_cvcwr[2], r_cvcwr[5:3]}), 
        .r_sdischg(r_sdischg), .r_bistctl(bist_r_ctl), .r_bistdat(bist_r_dat), 
        .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), .r_cvofsx(r_cvofsx), .r_pwm(
        r_pwm), .regx_wrdac({wr_dacv[17:16], r_dacwr[10:9], wr_dacv[15:8], 
        r_dacwr[8:7]}), .dac_r_vs(dac_r_vs[143:64]), .dac_comp(
        dac_r_comp[17:8]), .r_dac_en(r_dac_en[17:8]), .r_sar_en(r_sar_en[17:8]), .r_aopt(r_aopt), .r_xtm(r_xtm), .r_adummyi({SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, DUMMY_IN}), 
        .r_bck0(r_bck0), .r_bck1(r_bck1), .r_bck2({SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, r_bck2_2_, 
        lg_pulse_len}), .r_i2crout({r_i2crout, r_i2cmcu_route, r_i2cslv_route}), .r_xana({r_xana_23, SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, r_xana_19, r_xana_18, OCP_SEL, PWREN_HOLD, 
        r_xana}), .di_xanav(di_xanav), .lt_gpi(lt_gpi), .di_tst(di_tst), 
        .bkpt_pc(bkpt_pc), .bkpt_ena(bkpt_ena), .we_twlb(we_twlb), .r_vpp_en(
        r_vpp_en), .r_vpp0v_en(r_vpp0v_en), .r_otp_pwdn_en(r_otp_pwdn_en), 
        .r_otp_wpls(r_otp_wpls), .wd_twlb(wd_twlb), .r_sap(r_sap), .r_twlb(
        pmem_twlb), .upd_pwrv(r_pwrv_upd), .ramacc(ramacc), .sse_idle(sse_idle), .bus_idle(bus_idle), .r_do_ts(r_do_ts), .r_dpdo_sel(r_dpdo_sel), 
        .r_dndo_sel(r_dndo_sel), .di_ts(di_ts), .detclk(detclk), .aswclk(
        aswclk), .atpg_en(n107), .di_aswk({di_aswk[4], n117, di_aswk[2], 1'b0, 
        di_aswk_0}), .clk(g_clk), .rrstz(n82) );
  srambist_a0 u0_srambist ( .clk(g_clk), .srstz(n83), .reg_hit(regx_hitbst), 
        .reg_w(regx_we), .reg_r(regx_re), .reg_wdat({xram_d[7:1], n85}), 
        .iram_rdat({n129, n131, n133, n135, n138, n140, sram_rdat}), 
        .xram_rdat({n129, n131, n133, n135, n138, n140, sram_rdat}), .bist_en(
        bist_en), .bist_xram(), .bist_wr(bist_wr), .bist_adr(bist_adr), 
        .bist_wdat(bist_wdat), .o_bistctl(bist_r_ctl), .o_bistdat(bist_r_dat)
         );
  divclk_a0 u0_divclk ( .mclk(g_clk), .srstz(n83), .atpg_en(n87), .clk_1p0m(
        clk_1p0m), .clk_500k(clk_500k), .clk_100k(clk_100k), .clk_50k(clk_50k), 
        .clk_500(clk_500), .divff_o1(divff_o1), .divff_o2() );
  glpwm_a0_0 u0_pwm_0_ ( .clk(g_clk), .rstz(n83), .clk_base(clk_50k), .we(
        regx_wrpwm[0]), .wdat({xram_d[7:1], n85}), .r_pwm(r_pwm[7:0]), .pwm_o(
        pwm_o[0]) );
  glpwm_a0_1 u0_pwm_1_ ( .clk(g_clk), .rstz(n82), .clk_base(clk_50k), .we(
        regx_wrpwm[1]), .wdat({xram_d[7:1], n85}), .r_pwm(r_pwm[15:8]), 
        .pwm_o(pwm_o[1]) );
  SNPS_CLOCK_GATE_HIGH_core_a0 clk_gate_d_dodat_reg ( .CLK(g_clk), .EN(N568), 
        .ENCLK(net8853), .TE(1'b0) );
  DLNQX1 r_lt_gpi_reg_1_ ( .D(DI_GPIO[2]), .XG(i_rstz), .Q(r_lt_gpi[1]) );
  DLNQX1 r_lt_gpi_reg_0_ ( .D(DI_GPIO[3]), .XG(i_rstz), .Q(r_lt_gpi[0]) );
  DLNQX1 r_lt_gpi_reg_2_ ( .D(DI_GPIO[1]), .XG(i_rstz), .Q(r_lt_gpi[2]) );
  DLNQX1 r_lt_gpi_reg_3_ ( .D(DI_GPIO[0]), .XG(i_rstz), .Q(r_lt_gpi[3]) );
  DFFQX1 d_dodat_reg_10_ ( .D(N1483), .C(net8853), .Q(d_dodat[10]) );
  DFFQX1 d_dodat_reg_9_ ( .D(N575), .C(net8853), .Q(d_dodat[9]) );
  DFFQX1 d_dodat_reg_11_ ( .D(N1478), .C(net8853), .Q(d_dodat[11]) );
  DFFQX1 d_dodat_reg_12_ ( .D(N572), .C(net8853), .Q(d_dodat[12]) );
  DFFQX1 d_dodat_reg_14_ ( .D(N570), .C(net8853), .Q(d_dodat[14]) );
  DFFQX1 d_dodat_reg_8_ ( .D(N576), .C(net8853), .Q(d_dodat[8]) );
  DFFQX1 d_dodat_reg_15_ ( .D(N569), .C(net8853), .Q(d_dodat[15]) );
  DFFQX1 d_dodat_reg_13_ ( .D(N571), .C(net8853), .Q(d_dodat[13]) );
  DFFQX1 d_dodat_reg_1_ ( .D(N583), .C(net8853), .Q(d_dodat[1]) );
  DFFQX1 d_dodat_reg_2_ ( .D(N582), .C(net8853), .Q(d_dodat[2]) );
  DFFQX1 d_dodat_reg_3_ ( .D(N581), .C(net8853), .Q(d_dodat[3]) );
  DFFQX1 d_dodat_reg_0_ ( .D(N584), .C(net8853), .Q(d_dodat[0]) );
  DFFQX1 d_dodat_reg_5_ ( .D(N579), .C(net8853), .Q(d_dodat[5]) );
  DFFQX1 d_dodat_reg_6_ ( .D(N578), .C(net8853), .Q(d_dodat[6]) );
  DFFQX1 d_dodat_reg_4_ ( .D(N580), .C(net8853), .Q(d_dodat[4]) );
  DFFQX1 d_dodat_reg_7_ ( .D(N577), .C(net8853), .Q(d_dodat[7]) );
  NAND42X4 U3 ( .C(n275), .D(n269), .A(n56), .B(n268), .Y(DO_GPIO[4]) );
  AND2X1 U4 ( .A(n476), .B(n59), .Y(sse_prefetch) );
  NAND4X1 U5 ( .A(r_pg0_sel[2]), .B(r_pg0_sel[3]), .C(n475), .D(n474), .Y(n59)
         );
  INVX1 U6 ( .A(r_pg0_sel[0]), .Y(n475) );
  INVX1 U7 ( .A(r_pg0_sel[1]), .Y(n474) );
  INVX2 U8 ( .A(wr_dacv[15]), .Y(n465) );
  INVX1 U9 ( .A(sse_adr[7]), .Y(n476) );
  OAI211X1 U10 ( .C(n522), .D(n491), .A(n516), .B(n490), .Y(memdatai[2]) );
  AO21X1 U11 ( .B(SRAM_RDAT[7]), .C(n139), .A(n484), .Y(n129) );
  OR2X1 U12 ( .A(slvo_early), .B(slvo_re), .Y(n76) );
  NAND21X1 U13 ( .B(n470), .A(n20), .Y(n471) );
  NOR2X1 U14 ( .A(n521), .B(n522), .Y(n1) );
  INVX1 U15 ( .A(n471), .Y(n473) );
  AO2222XL U16 ( .A(cc2_di), .B(n537), .C(prx_rcvinf[4]), .D(n222), .E(
        r_vpp_en), .F(n639), .G(comp_smpl[0]), .H(n640), .Y(n233) );
  OAI211X1 U17 ( .C(n522), .D(n501), .A(n516), .B(n500), .Y(memdatai[4]) );
  NOR2X1 U18 ( .A(n520), .B(n519), .Y(n2) );
  INVX1 U19 ( .A(n518), .Y(n3) );
  OR3X4 U20 ( .A(n1), .B(n2), .C(n3), .Y(memdatai[7]) );
  INVX1 U21 ( .A(n129), .Y(n520) );
  MUX2IX2 U22 ( .D0(n86), .D1(n62), .S(n468), .Y(r_dacwdat[0]) );
  AO21X1 U23 ( .B(DAC1_COMP), .C(n119), .A(n648), .Y(n4) );
  MUX2IX1 U24 ( .D0(n552), .D1(di_gpio[0]), .S(n193), .Y(n5) );
  MUX2IX1 U25 ( .D0(n555), .D1(di_gpio[0]), .S(n184), .Y(n6) );
  AOI21X1 U26 ( .B(N603), .C(n204), .A(n191), .Y(n7) );
  BUFX2 U27 ( .A(xram_ce), .Y(n8) );
  INVX1 U28 ( .A(xram_d[4]), .Y(n26) );
  INVXL U29 ( .A(n679), .Y(n9) );
  INVX24 U30 ( .A(n9), .Y(PMEM_PGM) );
  NOR21XL U31 ( .B(pmem_pgm), .A(atpg_en), .Y(n679) );
  BUFXL U32 ( .A(wr_dacv[16]), .Y(n11) );
  BUFXL U33 ( .A(n463), .Y(n12) );
  BUFXL U34 ( .A(memaddr_c[1]), .Y(n13) );
  INVX1 U35 ( .A(regx_rdat[7]), .Y(n521) );
  INVXL U36 ( .A(n521), .Y(n14) );
  INVX3 U37 ( .A(wr_dacv[14]), .Y(n464) );
  BUFXL U38 ( .A(wr_dacv[17]), .Y(n15) );
  BUFXL U39 ( .A(xram_a[3]), .Y(n16) );
  INVXL U40 ( .A(n12), .Y(n17) );
  INVX2 U41 ( .A(wr_dacv[13]), .Y(n463) );
  BUFXL U42 ( .A(wr_dacv[11]), .Y(n18) );
  INVXL U43 ( .A(n469), .Y(n19) );
  INVXL U44 ( .A(n19), .Y(n20) );
  BUFXL U45 ( .A(memaddr_c[4]), .Y(n21) );
  INVXL U46 ( .A(n464), .Y(n22) );
  NAND43X2 U47 ( .B(r_dacwr[8]), .C(wr_dacv[8]), .D(r_dacwr[7]), .A(n467), .Y(
        n470) );
  NOR3X2 U48 ( .A(n466), .B(wr_dacv[10]), .C(wr_dacv[9]), .Y(n467) );
  BUFXL U49 ( .A(r_dacwr[9]), .Y(n23) );
  BUFXL U50 ( .A(memaddr_c[2]), .Y(n24) );
  BUFXL U51 ( .A(memaddr_c[0]), .Y(n25) );
  MUX2IX1 U52 ( .D0(n73), .D1(n26), .S(n471), .Y(r_dacwdat[4]) );
  INVX1 U53 ( .A(r_dacwr[10]), .Y(n461) );
  BUFXL U54 ( .A(memaddr_c[6]), .Y(n27) );
  BUFXL U55 ( .A(memaddr_c[3]), .Y(n31) );
  BUFXL U56 ( .A(wr_dacv[12]), .Y(n32) );
  BUFXL U57 ( .A(memaddr_c[5]), .Y(n33) );
  BUFXL U58 ( .A(wr_dacv[8]), .Y(n34) );
  INVXL U59 ( .A(wr_dacv[9]), .Y(n35) );
  INVX1 U60 ( .A(n35), .Y(n36) );
  NAND43X1 U61 ( .B(wr_dacv[17]), .C(r_dacwr[9]), .D(wr_dacv[16]), .A(n461), 
        .Y(n462) );
  INVXL U62 ( .A(n465), .Y(n37) );
  OR2X2 U63 ( .A(wr_dacv[11]), .B(wr_dacv[12]), .Y(n466) );
  BUFX3 U64 ( .A(bist_en), .Y(n38) );
  BUFX3 U65 ( .A(iram_ce), .Y(n39) );
  BUFX3 U66 ( .A(n676), .Y(PMEM_TWLB[0]) );
  NOR21XL U67 ( .B(pmem_twlb[0]), .A(n132), .Y(n676) );
  INVX1 U68 ( .A(n150), .Y(n41) );
  BUFXL U69 ( .A(r_adofs[3]), .Y(n42) );
  BUFX3 U70 ( .A(n675), .Y(PMEM_TWLB[1]) );
  NOR21XL U71 ( .B(pmem_twlb[1]), .A(n130), .Y(n675) );
  INVX1 U72 ( .A(n149), .Y(n44) );
  BUFXL U73 ( .A(r_adofs[1]), .Y(n45) );
  BUFXL U74 ( .A(r_adofs[2]), .Y(n46) );
  BUFXL U75 ( .A(r_adofs[4]), .Y(n47) );
  BUFXL U76 ( .A(r_adofs[5]), .Y(n48) );
  BUFX3 U77 ( .A(r_dac_en[3]), .Y(n49) );
  BUFX4 U78 ( .A(n678), .Y(PMEM_SAP[0]) );
  NOR21XL U79 ( .B(r_sap[0]), .A(n134), .Y(n678) );
  BUFX4 U80 ( .A(n677), .Y(PMEM_SAP[1]) );
  NOR21XL U81 ( .B(r_sap[1]), .A(n134), .Y(n677) );
  NAND42X1 U82 ( .C(n215), .D(n53), .A(n213), .B(n212), .Y(DO_GPIO[5]) );
  AO2222XL U83 ( .A(r_accctl[4]), .B(n446), .C(n58), .D(n443), .E(comp_smpl[3]), .F(n640), .G(n537), .H(TX_DAT), .Y(n454) );
  XOR2XL U84 ( .A(DO_GPIO[6]), .B(n289), .Y(n457) );
  NOR4XL U85 ( .A(r_cvcwr[3]), .B(r_cvcwr[2]), .C(r_cvcwr[5]), .D(r_cvcwr[4]), 
        .Y(n160) );
  XOR3X1 U86 ( .A(n52), .B(DO_GPIO[5]), .C(n57), .Y(N579) );
  XNOR2XL U87 ( .A(SRAM_D[1]), .B(SRAM_A[5]), .Y(n52) );
  INVXL U88 ( .A(n86), .Y(n85) );
  AOI21AX1 U89 ( .B(ictlr_inst[7]), .C(n517), .A(n516), .Y(n518) );
  INVXL U90 ( .A(regx_rdat[6]), .Y(n515) );
  INVXL U91 ( .A(regx_rdat[3]), .Y(n499) );
  INVXL U92 ( .A(regx_rdat[4]), .Y(n501) );
  INVX1 U93 ( .A(regx_rdat[2]), .Y(n491) );
  OAI222XL U94 ( .A(n147), .B(n654), .C(n451), .D(n180), .E(n449), .F(n168), 
        .Y(n53) );
  XNOR3X1 U95 ( .A(n277), .B(n278), .C(n54), .Y(N580) );
  XNOR2XL U96 ( .A(DO_GPIO[4]), .B(n279), .Y(n54) );
  XNOR3X1 U97 ( .A(n270), .B(n271), .C(n55), .Y(N581) );
  XNOR2XL U98 ( .A(DO_GPIO[3]), .B(n272), .Y(n55) );
  OAI22AXL U99 ( .D(xram_d[0]), .C(n160), .A(n565), .B(n62), .Y(r_cvcwdat[0])
         );
  AND2XL U100 ( .A(n76), .B(n476), .Y(i2c_ev_6_) );
  AO2222XL U101 ( .A(do_p0[6]), .B(n357), .C(n531), .D(n535), .E(mcu_dbgpo[16]), .F(n291), .G(n290), .H(r_ccctl[0]), .Y(n455) );
  AO2222XL U102 ( .A(n532), .B(n285), .C(mcu_dbgpo[17]), .D(n284), .E(n123), 
        .F(n281), .G(n280), .H(n4), .Y(n456) );
  AOI222XL U103 ( .A(n256), .B(n126), .C(n290), .D(n619), .E(upd_dbgpo[18]), 
        .F(n443), .Y(n56) );
  NOR21XL U104 ( .B(r_aopt[1]), .A(n97), .Y(ANAOPT[1]) );
  NOR21XL U105 ( .B(r_aopt[4]), .A(n97), .Y(ANAOPT[4]) );
  NOR21XL U106 ( .B(r_xana[12]), .A(n99), .Y(ANA_REGX[12]) );
  NOR21XL U107 ( .B(r_xana[2]), .A(n100), .Y(ANA_REGX[2]) );
  NOR21XL U108 ( .B(r_xana[4]), .A(n101), .Y(ANA_REGX[4]) );
  NOR21XL U109 ( .B(r_xana[6]), .A(n101), .Y(ANA_REGX[6]) );
  NOR21XL U110 ( .B(r_xana[8]), .A(n103), .Y(ANA_REGX[8]) );
  NOR21XL U111 ( .B(r_xana[9]), .A(n103), .Y(ANA_REGX[9]) );
  NOR21XL U112 ( .B(r_ccctl[1]), .A(n100), .Y(DO_CCCTL[1]) );
  NOR21XL U113 ( .B(r_ccctl[2]), .A(n100), .Y(DO_CCCTL[2]) );
  NOR21XL U114 ( .B(r_ccctl[3]), .A(n101), .Y(DO_CCCTL[3]) );
  NOR21XL U115 ( .B(r_cctrx[3]), .A(n100), .Y(DO_CCTRX[3]) );
  INVX1 U116 ( .A(n225), .Y(n357) );
  INVX1 U117 ( .A(n497), .Y(n205) );
  INVX1 U118 ( .A(n160), .Y(n565) );
  INVX1 U119 ( .A(n141), .Y(n94) );
  INVX1 U120 ( .A(n112), .Y(n93) );
  INVX1 U121 ( .A(n112), .Y(n92) );
  INVX1 U122 ( .A(n111), .Y(n91) );
  INVX1 U123 ( .A(n111), .Y(n90) );
  INVX1 U124 ( .A(n112), .Y(n96) );
  INVX1 U125 ( .A(n111), .Y(n89) );
  INVX1 U126 ( .A(n110), .Y(n95) );
  INVX1 U127 ( .A(n127), .Y(n88) );
  INVX1 U128 ( .A(n115), .Y(n102) );
  INVX1 U129 ( .A(n114), .Y(n97) );
  INVX1 U130 ( .A(n114), .Y(n99) );
  INVX1 U131 ( .A(n114), .Y(n101) );
  INVX1 U132 ( .A(n113), .Y(n100) );
  INVX1 U133 ( .A(n116), .Y(n98) );
  INVX1 U134 ( .A(n113), .Y(n103) );
  INVX1 U135 ( .A(n110), .Y(n87) );
  INVX1 U136 ( .A(n114), .Y(n106) );
  INVX1 U137 ( .A(n113), .Y(n105) );
  INVX1 U138 ( .A(n110), .Y(n104) );
  INVX1 U139 ( .A(n113), .Y(n107) );
  INVX1 U140 ( .A(n71), .Y(n69) );
  INVX1 U141 ( .A(n519), .Y(n507) );
  NAND21X1 U142 ( .B(n356), .A(n556), .Y(n225) );
  NAND21X1 U143 ( .B(n222), .A(n221), .Y(n497) );
  INVX1 U144 ( .A(fcp_oe), .Y(n450) );
  INVX1 U145 ( .A(n256), .Y(n219) );
  NAND2X1 U146 ( .A(n139), .B(sram_en), .Y(SRAM_CEB) );
  INVX1 U147 ( .A(n84), .Y(n82) );
  INVX1 U148 ( .A(n65), .Y(n64) );
  INVX1 U149 ( .A(n81), .Y(n80) );
  INVX1 U150 ( .A(n68), .Y(n67) );
  INVX1 U151 ( .A(n71), .Y(n70) );
  INVX1 U152 ( .A(n77), .Y(n75) );
  INVX1 U153 ( .A(n73), .Y(n72) );
  INVX1 U154 ( .A(n62), .Y(n60) );
  INVX1 U155 ( .A(n68), .Y(n66) );
  INVX1 U156 ( .A(n65), .Y(n63) );
  INVX1 U157 ( .A(n77), .Y(n74) );
  INVX1 U158 ( .A(n79), .Y(n78) );
  INVX1 U159 ( .A(n62), .Y(n61) );
  NOR2X1 U160 ( .A(n106), .B(n577), .Y(OSC_STOP) );
  NOR2X1 U161 ( .A(n106), .B(n576), .Y(OSC_LOW) );
  INVX1 U162 ( .A(n84), .Y(n83) );
  INVX1 U163 ( .A(n136), .Y(n109) );
  INVX1 U164 ( .A(n134), .Y(n110) );
  INVX1 U165 ( .A(n134), .Y(n114) );
  INVX1 U166 ( .A(n134), .Y(n112) );
  INVX1 U167 ( .A(n132), .Y(n111) );
  INVX1 U168 ( .A(n134), .Y(n113) );
  INVX1 U169 ( .A(n132), .Y(n119) );
  INVX1 U170 ( .A(n132), .Y(n120) );
  INVX1 U171 ( .A(n130), .Y(n122) );
  INVX1 U172 ( .A(atpg_en), .Y(n125) );
  INVX1 U173 ( .A(n130), .Y(n124) );
  INVX1 U174 ( .A(n130), .Y(n121) );
  INVX1 U175 ( .A(n132), .Y(n116) );
  INVX1 U176 ( .A(n130), .Y(n115) );
  INVX1 U177 ( .A(atpg_en), .Y(n118) );
  INVX1 U178 ( .A(atpg_en), .Y(n127) );
  NAND21X1 U179 ( .B(hit_xr), .A(n485), .Y(n519) );
  INVX1 U180 ( .A(sfr_wdat[3]), .Y(n71) );
  INVX1 U181 ( .A(sfr_wdat[4]), .Y(n73) );
  INVX1 U182 ( .A(sfr_wdat[0]), .Y(n62) );
  XNOR2XL U183 ( .A(n282), .B(n283), .Y(n57) );
  NAND43X1 U184 ( .B(n290), .C(n291), .D(n446), .A(n451), .Y(n533) );
  NAND43X1 U185 ( .B(n284), .C(n256), .D(n533), .A(n208), .Y(n356) );
  AND4X1 U186 ( .A(n449), .B(n207), .C(n206), .D(n205), .Y(n208) );
  INVX1 U187 ( .A(n640), .Y(n207) );
  INVX1 U188 ( .A(n537), .Y(n206) );
  OR2X1 U189 ( .A(n281), .B(n443), .Y(n222) );
  INVX1 U190 ( .A(n314), .Y(do_opt_0) );
  NAND21X1 U191 ( .B(n535), .A(n536), .Y(n256) );
  XNOR2XL U192 ( .A(n240), .B(SRAM_D[2]), .Y(n289) );
  NAND21X1 U193 ( .B(n534), .A(n7), .Y(n284) );
  NAND21X1 U194 ( .B(n638), .A(n225), .Y(n538) );
  INVX1 U195 ( .A(n280), .Y(n221) );
  INVX1 U196 ( .A(n253), .Y(n451) );
  INVX1 U197 ( .A(n285), .Y(n536) );
  INVX1 U198 ( .A(srstz), .Y(n84) );
  INVX1 U199 ( .A(n639), .Y(n449) );
  INVX1 U200 ( .A(n638), .Y(n556) );
  OR3XL U201 ( .A(n535), .B(n534), .C(n533), .Y(n498) );
  INVX1 U202 ( .A(s0_rxdoe), .Y(n641) );
  INVX1 U203 ( .A(n240), .Y(SRAM_A[6]) );
  INVX1 U204 ( .A(n241), .Y(SRAM_A[3]) );
  OR2X1 U205 ( .A(xram_ce), .B(iram_ce), .Y(sram_en) );
  INVX1 U206 ( .A(o_dodat0_15_), .Y(n576) );
  INVX1 U207 ( .A(n236), .Y(SRAM_D[5]) );
  INVX1 U208 ( .A(n237), .Y(SRAM_D[4]) );
  OAI22X1 U209 ( .A(n160), .B(n567), .C(n65), .D(n565), .Y(r_cvcwdat[1]) );
  OAI22X1 U210 ( .A(n160), .B(n568), .C(n68), .D(n565), .Y(r_cvcwdat[2]) );
  OAI22X1 U211 ( .A(n160), .B(n569), .C(n71), .D(n565), .Y(r_cvcwdat[3]) );
  OAI22X1 U212 ( .A(n160), .B(n571), .C(n79), .D(n565), .Y(r_cvcwdat[6]) );
  OAI22X1 U213 ( .A(n160), .B(n572), .C(n81), .D(n565), .Y(r_cvcwdat[7]) );
  INVX1 U214 ( .A(sfr_wdat[7]), .Y(n81) );
  INVX1 U215 ( .A(sfr_wdat[1]), .Y(n65) );
  INVX1 U216 ( .A(n238), .Y(SRAM_D[0]) );
  INVX1 U217 ( .A(sfr_wdat[6]), .Y(n79) );
  INVX1 U218 ( .A(sfr_wdat[2]), .Y(n68) );
  INVX1 U219 ( .A(sfr_wdat[5]), .Y(n77) );
  INVX1 U220 ( .A(xram_we), .Y(n566) );
  XNOR2XL U221 ( .A(DO_DAC0[0]), .B(DAC3_V[5]), .Y(n282) );
  OAI21X1 U222 ( .B(xram_we), .C(iram_we), .A(n139), .Y(SRAM_WEB) );
  OR2X1 U223 ( .A(iram_we), .B(xram_we), .Y(n340) );
  INVX1 U224 ( .A(r_osc_stop), .Y(n577) );
  NOR2X1 U225 ( .A(n597), .B(n593), .Y(n364) );
  INVX1 U226 ( .A(n379), .Y(n603) );
  NOR2X1 U227 ( .A(n332), .B(n104), .Y(TX_EN) );
  NOR2X1 U228 ( .A(n105), .B(n584), .Y(STB_RP) );
  AOI21X1 U229 ( .B(n596), .C(n592), .A(n107), .Y(CCI2C_EN) );
  NOR2X1 U230 ( .A(n106), .B(n575), .Y(DO_SRCCTL[3]) );
  NOR2X1 U231 ( .A(n105), .B(n574), .Y(DO_SRCCTL[2]) );
  NOR2X1 U232 ( .A(n106), .B(n579), .Y(DO_SRCCTL[0]) );
  NOR2X1 U233 ( .A(n105), .B(n578), .Y(BCK_REGX[2]) );
  NAND21X1 U234 ( .B(n672), .A(n202), .Y(n165) );
  NAND2X1 U235 ( .A(n650), .B(n651), .Y(n670) );
  NAND2X1 U236 ( .A(n647), .B(n646), .Y(n660) );
  NAND2X1 U237 ( .A(n141), .B(n147), .Y(tclk_sel) );
  INVX1 U238 ( .A(n136), .Y(n108) );
  INVX1 U239 ( .A(n139), .Y(n136) );
  INVX1 U240 ( .A(n141), .Y(n132) );
  INVX1 U241 ( .A(n139), .Y(n134) );
  INVX1 U242 ( .A(n141), .Y(n130) );
  INVX1 U243 ( .A(n147), .Y(n151) );
  OAI211X1 U244 ( .C(n522), .D(n515), .A(n516), .B(n512), .Y(memdatai[6]) );
  AOI22X1 U245 ( .A(n507), .B(n131), .C(ictlr_inst[6]), .D(n517), .Y(n512) );
  OAI211X1 U246 ( .C(n522), .D(n499), .A(n516), .B(n492), .Y(memdatai[3]) );
  AOI22X1 U247 ( .A(n507), .B(n138), .C(ictlr_inst[3]), .D(n517), .Y(n492) );
  AOI22X1 U248 ( .A(n507), .B(n140), .C(ictlr_inst[2]), .D(n517), .Y(n490) );
  AOI22X1 U249 ( .A(n507), .B(n135), .C(ictlr_inst[4]), .D(n517), .Y(n500) );
  OAI211X1 U250 ( .C(n522), .D(n503), .A(n516), .B(n502), .Y(memdatai[5]) );
  AOI22X1 U251 ( .A(n507), .B(n133), .C(ictlr_inst[5]), .D(n517), .Y(n502) );
  INVXL U252 ( .A(regx_rdat[5]), .Y(n503) );
  INVX1 U253 ( .A(xram_d[0]), .Y(n86) );
  OAI211X1 U254 ( .C(n522), .D(n489), .A(n516), .B(n488), .Y(memdatai[1]) );
  AOI22X1 U255 ( .A(n507), .B(sram_rdat[1]), .C(ictlr_inst[1]), .D(n517), .Y(
        n488) );
  INVX1 U256 ( .A(regx_rdat[1]), .Y(n489) );
  OAI211X1 U257 ( .C(n522), .D(n487), .A(n516), .B(n486), .Y(memdatai[0]) );
  AOI22X1 U258 ( .A(n507), .B(sram_rdat[0]), .C(ictlr_inst[0]), .D(n517), .Y(
        n486) );
  INVXL U259 ( .A(regx_rdat[0]), .Y(n487) );
  AOI221XL U260 ( .A(n290), .B(TX_DAT), .C(mcu_dbgpo[22]), .D(n291), .E(n209), 
        .Y(n213) );
  OA222X1 U261 ( .A(n221), .B(n211), .C(n576), .D(n7), .E(n210), .F(n219), .Y(
        n212) );
  NAND21X1 U262 ( .B(n517), .A(hit_xr), .Y(n522) );
  INVX1 U263 ( .A(n517), .Y(n485) );
  INVX1 U264 ( .A(n137), .Y(n544) );
  INVX1 U265 ( .A(n550), .Y(n527) );
  XNOR2XL U266 ( .A(n328), .B(n329), .Y(N570) );
  XNOR2XL U267 ( .A(n330), .B(n331), .Y(n329) );
  XNOR2XL U268 ( .A(n333), .B(n334), .Y(n328) );
  XNOR2XL U269 ( .A(DAC1_V[8]), .B(TX_EN), .Y(n330) );
  INVX1 U270 ( .A(n582), .Y(o_dodat5_2_) );
  INVX1 U271 ( .A(di_gpio[2]), .Y(n546) );
  INVX1 U272 ( .A(n126), .Y(n392) );
  INVX1 U273 ( .A(n128), .Y(n543) );
  OAI22X1 U274 ( .A(n379), .B(n543), .C(n378), .D(n392), .Y(n391) );
  OAI22X1 U275 ( .A(n384), .B(n583), .C(n578), .D(n385), .Y(n386) );
  OAI22X1 U276 ( .A(n274), .B(n378), .C(n584), .D(n379), .Y(n377) );
  INVX1 U277 ( .A(r_xana_19), .Y(n584) );
  XOR3X1 U278 ( .A(n287), .B(n288), .C(n457), .Y(N578) );
  XNOR2XL U279 ( .A(DO_DAC0[1]), .B(DAC1_V[0]), .Y(n287) );
  XNOR2XL U280 ( .A(dacmux_sel[6]), .B(DO_PWR_I[6]), .Y(n288) );
  XOR3X1 U281 ( .A(n292), .B(n293), .C(n154), .Y(N577) );
  XNOR2XL U282 ( .A(DO_DAC0[2]), .B(DAC1_V[1]), .Y(n292) );
  XNOR2XL U283 ( .A(dacmux_sel[7]), .B(DO_PWR_I[7]), .Y(n293) );
  XOR2X1 U284 ( .A(n153), .B(n295), .Y(n154) );
  XNOR2XL U285 ( .A(n315), .B(n316), .Y(N572) );
  XNOR2XL U286 ( .A(n317), .B(n318), .Y(n316) );
  XNOR2XL U287 ( .A(n573), .B(n319), .Y(n315) );
  XNOR2XL U288 ( .A(dacmux_sel[12]), .B(DO_DAC0[7]), .Y(n317) );
  AOI222XL U289 ( .A(n182), .B(n190), .C(n5), .D(n183), .E(n593), .F(n192), 
        .Y(n511) );
  INVX1 U290 ( .A(n123), .Y(n393) );
  AOI222XL U291 ( .A(n612), .B(cc1_di), .C(n414), .D(di_sqlch), .E(n613), .F(
        n619), .Y(n430) );
  AOI222XL U292 ( .A(n612), .B(cc2_di), .C(n414), .D(n123), .E(n613), .F(
        TX_DAT), .Y(n421) );
  AOI222XL U293 ( .A(n177), .B(n190), .C(n5), .D(n179), .E(n597), .F(n192), 
        .Y(n510) );
  AOI222XL U294 ( .A(n177), .B(n178), .C(n179), .D(n6), .E(n597), .F(n181), 
        .Y(n508) );
  INVX1 U295 ( .A(di_xanav[0]), .Y(n542) );
  AOI221XL U296 ( .A(n613), .B(di_pro[5]), .C(n612), .D(n4), .E(n422), .Y(n420) );
  OAI22X1 U297 ( .A(n574), .B(n611), .C(n392), .D(n610), .Y(n422) );
  AOI221XL U298 ( .A(n437), .B(dp_comp), .C(n436), .D(dm_comp), .E(n438), .Y(
        n434) );
  ENOX1 U299 ( .A(n581), .B(n439), .C(pwm_o[1]), .D(n587), .Y(n438) );
  AOI221XL U300 ( .A(n414), .B(di_pro[2]), .C(n406), .D(n128), .E(n431), .Y(
        n429) );
  OAI22X1 U301 ( .A(n416), .B(n585), .C(n575), .D(n417), .Y(n431) );
  AOI221XL U302 ( .A(n588), .B(n126), .C(n587), .D(n532), .E(n442), .Y(n441)
         );
  OAI22X1 U303 ( .A(n542), .B(n541), .C(n540), .D(n539), .Y(n442) );
  INVX1 U304 ( .A(n437), .Y(n541) );
  INVX1 U305 ( .A(n436), .Y(n539) );
  INVX1 U306 ( .A(di_xanav[1]), .Y(n540) );
  NOR3XL U307 ( .A(n177), .B(n393), .C(n182), .Y(n58) );
  INVX1 U308 ( .A(n294), .Y(n153) );
  AOI222XL U309 ( .A(n182), .B(n178), .C(n183), .D(n6), .E(n593), .F(n181), 
        .Y(n509) );
  XNOR2XL U310 ( .A(dacmux_sel[4]), .B(DO_PWR_I[4]), .Y(n278) );
  XNOR2XL U311 ( .A(DAC3_V[4]), .B(n238), .Y(n277) );
  XNOR2XL U312 ( .A(dacmux_sel[3]), .B(DO_PWR_I[3]), .Y(n271) );
  XNOR2XL U313 ( .A(DAC3_V[3]), .B(n241), .Y(n270) );
  XNOR2XL U314 ( .A(r_xana_19), .B(r_srcctl[0]), .Y(n318) );
  XNOR2XL U315 ( .A(n583), .B(dacmux_sel[11]), .Y(n353) );
  XNOR2XL U316 ( .A(n351), .B(n352), .Y(N1478) );
  XNOR2XL U317 ( .A(n354), .B(SRAM_D[7]), .Y(n351) );
  XNOR2XL U318 ( .A(DO_DAC0[6]), .B(n353), .Y(n352) );
  XOR2X1 U319 ( .A(DAC1_V[5]), .B(n248), .Y(n354) );
  OA21X1 U320 ( .B(n281), .C(n280), .A(n123), .Y(n257) );
  INVX1 U321 ( .A(di_pro[2]), .Y(n210) );
  INVX1 U322 ( .A(dp_comp), .Y(n211) );
  MUX2XL U323 ( .D0(xram_d[1]), .D1(n64), .S(n473), .Y(r_dacwdat[1]) );
  MUX2XL U324 ( .D0(xram_d[7]), .D1(n80), .S(n473), .Y(r_dacwdat[7]) );
  XOR3X1 U325 ( .A(n266), .B(o_dodat5_2_), .C(n459), .Y(N582) );
  XOR2X1 U326 ( .A(n264), .B(n265), .Y(n459) );
  XNOR2XL U327 ( .A(DO_GPIO[2]), .B(n267), .Y(n266) );
  XNOR2XL U328 ( .A(dacmux_sel[2]), .B(DO_PWR_I[2]), .Y(n265) );
  AOI22BXL U329 ( .B(n536), .A(di_pro[5]), .D(n7), .C(r_osc_stop), .Y(n494) );
  INVX1 U330 ( .A(di_gpio[0]), .Y(n549) );
  INVX1 U331 ( .A(n460), .Y(n481) );
  MUX2XL U332 ( .D0(xram_d[6]), .D1(n78), .S(n473), .Y(r_dacwdat[6]) );
  MUX2XL U333 ( .D0(xram_d[5]), .D1(n75), .S(n473), .Y(r_dacwdat[5]) );
  MUX2XL U334 ( .D0(xram_d[2]), .D1(n67), .S(n473), .Y(r_dacwdat[2]) );
  MUX2XL U335 ( .D0(xram_d[3]), .D1(n70), .S(n473), .Y(r_dacwdat[3]) );
  INVX1 U336 ( .A(pwm_o[0]), .Y(n581) );
  NOR2X1 U337 ( .A(n106), .B(n294), .Y(DO_TS[3]) );
  OAI22X1 U338 ( .A(n598), .B(n361), .C(mcuo_scl), .D(n594), .Y(n314) );
  AO21X1 U339 ( .B(N595), .C(n204), .A(n163), .Y(n443) );
  NOR2X1 U340 ( .A(n659), .B(n658), .Y(N595) );
  AO21X1 U341 ( .B(N629), .C(n202), .A(n479), .Y(n163) );
  NOR2X1 U342 ( .A(n669), .B(n668), .Y(N629) );
  AO21X1 U343 ( .B(N596), .C(n204), .A(n161), .Y(n281) );
  NOR2X1 U344 ( .A(n660), .B(n658), .Y(N596) );
  AO21X1 U345 ( .B(N630), .C(n202), .A(n480), .Y(n161) );
  NOR2X1 U346 ( .A(n670), .B(n668), .Y(N630) );
  NOR21XL U347 ( .B(dacmux_sel[9]), .A(n88), .Y(SAMPL_SEL[9]) );
  NOR21XL U348 ( .B(dacmux_sel[5]), .A(n88), .Y(SAMPL_SEL[5]) );
  NOR21XL U349 ( .B(dacmux_sel[8]), .A(n88), .Y(SAMPL_SEL[8]) );
  NOR21XL U350 ( .B(dacmux_sel[4]), .A(n88), .Y(SAMPL_SEL[4]) );
  NOR21XL U351 ( .B(dacmux_sel[12]), .A(n89), .Y(SAMPL_SEL[12]) );
  NOR21XL U352 ( .B(dacmux_sel[6]), .A(n88), .Y(SAMPL_SEL[6]) );
  NOR21XL U353 ( .B(dacmux_sel[7]), .A(n88), .Y(SAMPL_SEL[7]) );
  NOR21XL U354 ( .B(dacmux_sel[2]), .A(n89), .Y(SAMPL_SEL[2]) );
  NOR21XL U355 ( .B(dacmux_sel[3]), .A(n88), .Y(SAMPL_SEL[3]) );
  NOR21XL U356 ( .B(dacmux_sel[0]), .A(n89), .Y(SAMPL_SEL[0]) );
  NOR21XL U357 ( .B(dacmux_sel[13]), .A(n89), .Y(SAMPL_SEL[13]) );
  NOR21XL U358 ( .B(dacmux_sel[14]), .A(n89), .Y(SAMPL_SEL[14]) );
  NOR21XL U359 ( .B(dacmux_sel[15]), .A(n89), .Y(SAMPL_SEL[15]) );
  NOR21XL U360 ( .B(dacmux_sel[16]), .A(n89), .Y(SAMPL_SEL[16]) );
  NOR21XL U361 ( .B(dacmux_sel[17]), .A(n89), .Y(SAMPL_SEL[17]) );
  NOR21XL U362 ( .B(dacmux_sel[1]), .A(n89), .Y(SAMPL_SEL[1]) );
  NAND21X1 U363 ( .B(n663), .A(n204), .Y(n157) );
  OAI221X1 U364 ( .A(n674), .B(n158), .C(n664), .D(n157), .E(n175), .Y(n446)
         );
  AND2X1 U365 ( .A(dacmux_sel[11]), .B(n108), .Y(SAMPL_SEL[11]) );
  INVX1 U366 ( .A(n235), .Y(n117) );
  NOR2X1 U367 ( .A(n105), .B(n617), .Y(SAMPL_SEL[10]) );
  INVX1 U368 ( .A(n244), .Y(SRAM_A[0]) );
  INVX1 U369 ( .A(n243), .Y(SRAM_A[1]) );
  AO21X1 U370 ( .B(N598), .C(n204), .A(n203), .Y(n280) );
  NOR2X1 U371 ( .A(n664), .B(n661), .Y(N598) );
  AO21X1 U372 ( .B(N632), .C(n202), .A(n482), .Y(n203) );
  NOR2X1 U373 ( .A(n674), .B(n671), .Y(N632) );
  AO21X1 U374 ( .B(N600), .C(n44), .A(n198), .Y(n285) );
  NOR2X1 U375 ( .A(n661), .B(n660), .Y(N600) );
  AO21X1 U376 ( .B(N634), .C(n202), .A(n484), .Y(n198) );
  NOR2X1 U377 ( .A(n671), .B(n670), .Y(N634) );
  AO21X1 U378 ( .B(N606), .C(n204), .A(n167), .Y(n253) );
  NOR2X1 U379 ( .A(n664), .B(n657), .Y(N606) );
  AO21X1 U380 ( .B(N640), .C(n202), .A(n166), .Y(n167) );
  NOR2X1 U381 ( .A(n674), .B(n667), .Y(N640) );
  OAI221X1 U382 ( .A(n670), .B(n158), .C(n660), .D(n157), .E(n173), .Y(n640)
         );
  OAI221X1 U383 ( .A(n671), .B(n165), .C(n661), .D(n164), .E(n460), .Y(n537)
         );
  OAI221X1 U384 ( .A(n667), .B(n165), .C(n657), .D(n164), .E(n172), .Y(n639)
         );
  XOR3X1 U385 ( .A(DO_PWR_I[0]), .B(n255), .C(n143), .Y(N584) );
  XNOR2XL U386 ( .A(dacmux_sel[16]), .B(dacmux_sel[0]), .Y(n255) );
  XOR2X1 U387 ( .A(SRAM_A[0]), .B(n254), .Y(n143) );
  XNOR2XL U388 ( .A(DO_GPIO[0]), .B(DAC3_V[0]), .Y(n254) );
  XOR3X1 U389 ( .A(n258), .B(n259), .C(n146), .Y(N583) );
  XNOR2XL U390 ( .A(DO_PWR_I[1]), .B(DO_GPIO[1]), .Y(n258) );
  XNOR2XL U391 ( .A(dacmux_sel[1]), .B(dacmux_sel[17]), .Y(n259) );
  XOR2X1 U392 ( .A(SRAM_A[1]), .B(n260), .Y(n146) );
  AO21X1 U393 ( .B(N601), .C(n204), .A(n185), .Y(n290) );
  NOR2X1 U394 ( .A(n663), .B(n662), .Y(N601) );
  AO21X1 U395 ( .B(N635), .C(n202), .A(n648), .Y(n185) );
  NOR2X1 U396 ( .A(n673), .B(n672), .Y(N635) );
  AO21X1 U397 ( .B(N608), .C(n204), .A(n187), .Y(n291) );
  NOR2X1 U398 ( .A(n660), .B(n657), .Y(N608) );
  AO21X1 U399 ( .B(N642), .C(n202), .A(n252), .Y(n187) );
  NOR2X1 U400 ( .A(n670), .B(n667), .Y(N642) );
  NAND21X1 U401 ( .B(n483), .A(n196), .Y(n535) );
  AOI22X1 U402 ( .A(N599), .B(n44), .C(N633), .D(n202), .Y(n196) );
  NOR2X1 U403 ( .A(n671), .B(n669), .Y(N633) );
  NOR2X1 U404 ( .A(n661), .B(n659), .Y(N599) );
  NAND21X1 U405 ( .B(n662), .A(n204), .Y(n164) );
  AO21X1 U406 ( .B(N641), .C(n41), .A(n189), .Y(n534) );
  NOR2X1 U407 ( .A(n669), .B(n667), .Y(N641) );
  AO21X1 U408 ( .B(N607), .C(n204), .A(n216), .Y(n189) );
  NOR2X1 U409 ( .A(n659), .B(n657), .Y(N607) );
  NOR2X1 U410 ( .A(n663), .B(n659), .Y(N603) );
  AO21X1 U411 ( .B(N637), .C(n41), .A(n276), .Y(n191) );
  NOR2X1 U412 ( .A(n106), .B(n250), .Y(OE_GPIO[1]) );
  NOR2X1 U413 ( .A(n106), .B(n251), .Y(OE_GPIO[0]) );
  NOR2X1 U414 ( .A(n105), .B(n247), .Y(OE_GPIO[4]) );
  NOR2X1 U415 ( .A(n106), .B(n248), .Y(OE_GPIO[3]) );
  NOR2X1 U416 ( .A(n106), .B(n249), .Y(OE_GPIO[2]) );
  NAND2X1 U417 ( .A(n245), .B(n111), .Y(OE_GPIO[6]) );
  NAND2X1 U418 ( .A(n246), .B(n109), .Y(OE_GPIO[5]) );
  NOR2X1 U419 ( .A(n104), .B(n618), .Y(SH_RST) );
  INVX1 U420 ( .A(n176), .Y(n648) );
  INVX1 U421 ( .A(n170), .Y(n216) );
  INVX1 U422 ( .A(n169), .Y(n252) );
  INVX1 U423 ( .A(n171), .Y(n166) );
  AO21X1 U424 ( .B(N594), .C(n44), .A(n152), .Y(n638) );
  NOR2X1 U425 ( .A(n662), .B(n658), .Y(N594) );
  AO21X1 U426 ( .B(N627), .C(n41), .A(n151), .Y(n152) );
  NOR2X1 U427 ( .A(n672), .B(n668), .Y(N627) );
  XNOR2XL U428 ( .A(DAC3_V[2]), .B(n242), .Y(n264) );
  XOR2X1 U429 ( .A(n419), .B(SRAM_A[4]), .Y(n279) );
  XNOR2XL U430 ( .A(n239), .B(SRAM_D[3]), .Y(n295) );
  INVX1 U431 ( .A(n305), .Y(do_opt_1) );
  INVX1 U432 ( .A(n172), .Y(n649) );
  INVX1 U433 ( .A(n173), .Y(n286) );
  INVX1 U434 ( .A(n444), .Y(n587) );
  INVX1 U435 ( .A(n439), .Y(n588) );
  INVX1 U436 ( .A(n179), .Y(n598) );
  INVX1 U437 ( .A(n183), .Y(n594) );
  INVX1 U438 ( .A(n174), .Y(n276) );
  AO22X1 U439 ( .A(xram_a[8]), .B(n8), .C(iram_a[8]), .D(n39), .Y(SRAM_A[8])
         );
  AO22XL U440 ( .A(xram_a[5]), .B(xram_ce), .C(iram_a[5]), .D(iram_ce), .Y(
        SRAM_A[5]) );
  AO22X1 U441 ( .A(xram_a[10]), .B(n8), .C(iram_a[10]), .D(n39), .Y(SRAM_A[10]) );
  XNOR2XL U442 ( .A(sram_en), .B(n245), .Y(n333) );
  XNOR2XL U443 ( .A(n306), .B(n307), .Y(N575) );
  XNOR2XL U444 ( .A(n308), .B(n309), .Y(n307) );
  XNOR2XL U445 ( .A(n310), .B(SRAM_A[9]), .Y(n306) );
  XNOR2XL U446 ( .A(DO_DAC0[4]), .B(DAC1_V[3]), .Y(n308) );
  XNOR2XL U447 ( .A(n343), .B(n344), .Y(N1483) );
  XNOR2XL U448 ( .A(DAC1_V[4]), .B(n345), .Y(n344) );
  XNOR2XL U449 ( .A(n346), .B(SRAM_A[10]), .Y(n343) );
  XNOR2XL U450 ( .A(DO_DAC0[5]), .B(n617), .Y(n345) );
  XNOR2XL U451 ( .A(n296), .B(n297), .Y(N576) );
  XNOR2XL U452 ( .A(n298), .B(n299), .Y(n297) );
  XNOR2XL U453 ( .A(n300), .B(SRAM_A[8]), .Y(n296) );
  XNOR2XL U454 ( .A(DO_DAC0[3]), .B(DAC1_V[2]), .Y(n298) );
  INVX1 U455 ( .A(n342), .Y(TX_DAT) );
  INVX1 U456 ( .A(n175), .Y(n156) );
  XOR2X1 U457 ( .A(n249), .B(SRAM_D[6]), .Y(n346) );
  ENOX1 U458 ( .A(n571), .B(n566), .C(iram_d[6]), .D(iram_we), .Y(SRAM_D[6])
         );
  ENOX1 U459 ( .A(n572), .B(n566), .C(iram_we), .D(iram_d[7]), .Y(SRAM_D[7])
         );
  INVX1 U460 ( .A(n239), .Y(SRAM_A[7]) );
  INVX1 U461 ( .A(n242), .Y(SRAM_A[2]) );
  AOI22XL U462 ( .A(xram_d[4]), .B(xram_we), .C(iram_d[4]), .D(iram_we), .Y(
        n237) );
  XNOR2XL U463 ( .A(n236), .B(n250), .Y(n310) );
  XNOR2XL U464 ( .A(n237), .B(n251), .Y(n300) );
  AOI22XL U465 ( .A(xram_d[5]), .B(xram_we), .C(iram_d[5]), .D(iram_we), .Y(
        n236) );
  OAI22X1 U466 ( .A(n160), .B(n570), .C(n77), .D(n565), .Y(r_cvcwdat[5]) );
  INVX1 U467 ( .A(xram_d[5]), .Y(n570) );
  OAI22X1 U468 ( .A(n565), .B(n73), .C(n160), .D(n26), .Y(r_cvcwdat[4]) );
  ENOX1 U469 ( .A(n569), .B(n566), .C(iram_d[3]), .D(iram_we), .Y(SRAM_D[3])
         );
  ENOX1 U470 ( .A(n568), .B(n566), .C(iram_d[2]), .D(iram_we), .Y(SRAM_D[2])
         );
  AOI22X1 U471 ( .A(n85), .B(xram_we), .C(iram_d[0]), .D(iram_we), .Y(n238) );
  XNOR2XL U472 ( .A(o_dodat0_15_), .B(dacmux_sel[15]), .Y(n338) );
  XNOR2XL U473 ( .A(r_srcctl[1]), .B(dacmux_sel[13]), .Y(n324) );
  XNOR2XL U474 ( .A(r_srcctl[2]), .B(dacmux_sel[9]), .Y(n309) );
  XNOR2XL U475 ( .A(r_srcctl[3]), .B(dacmux_sel[8]), .Y(n299) );
  XNOR2XL U476 ( .A(dacmux_sel[14]), .B(DO_DAC0[9]), .Y(n331) );
  XNOR2XL U477 ( .A(dacmux_sel[5]), .B(DO_PWR_I[5]), .Y(n283) );
  XNOR2XL U478 ( .A(n321), .B(n322), .Y(N571) );
  XNOR2XL U479 ( .A(n325), .B(n326), .Y(n321) );
  XNOR2XL U480 ( .A(n323), .B(n324), .Y(n322) );
  XNOR2XL U481 ( .A(n327), .B(n246), .Y(n325) );
  XNOR2XL U482 ( .A(n335), .B(n336), .Y(N569) );
  XNOR2XL U483 ( .A(n339), .B(n340), .Y(n335) );
  XNOR2XL U484 ( .A(n337), .B(n338), .Y(n336) );
  XNOR2XL U485 ( .A(n341), .B(n342), .Y(n339) );
  ENOX1 U486 ( .A(n567), .B(n566), .C(iram_d[1]), .D(iram_we), .Y(SRAM_D[1])
         );
  NOR2X1 U487 ( .A(n106), .B(n573), .Y(DO_VOOC[0]) );
  NOR21XL U488 ( .B(n334), .A(n97), .Y(DO_VOOC[2]) );
  INVX1 U489 ( .A(xram_d[2]), .Y(n568) );
  OAI22X1 U490 ( .A(n596), .B(n361), .C(mcuo_scl), .D(n592), .Y(n504) );
  INVX1 U491 ( .A(xram_d[3]), .Y(n569) );
  INVX1 U492 ( .A(xram_d[1]), .Y(n567) );
  INVX1 U493 ( .A(xram_d[7]), .Y(n572) );
  INVX1 U494 ( .A(xram_d[6]), .Y(n571) );
  INVX1 U495 ( .A(n273), .Y(CC1_DOB) );
  INVX1 U496 ( .A(r_osc_gate), .Y(n644) );
  NOR2X1 U497 ( .A(sh_hold), .B(n618), .Y(N568) );
  INVX1 U498 ( .A(r_srcctl[0]), .Y(n579) );
  OAI22X1 U499 ( .A(n579), .B(n416), .C(n417), .D(n626), .Y(n415) );
  INVX1 U500 ( .A(r_srcctl[3]), .Y(n575) );
  INVX1 U501 ( .A(n182), .Y(n592) );
  INVX1 U502 ( .A(n619), .Y(n332) );
  INVX1 U503 ( .A(n177), .Y(n596) );
  NOR21XL U504 ( .B(n326), .A(n97), .Y(DO_VOOC[1]) );
  NOR21XL U505 ( .B(n341), .A(n97), .Y(DO_VOOC[3]) );
  NAND2X1 U506 ( .A(n624), .B(n605), .Y(n379) );
  OAI22X1 U507 ( .A(n400), .B(n361), .C(mcuo_scl), .D(n401), .Y(n366) );
  OAI32X1 U508 ( .A(n610), .B(n615), .C(n637), .D(n611), .E(n327), .Y(n428) );
  INVX1 U509 ( .A(n267), .Y(n578) );
  INVX1 U510 ( .A(r_srcctl[2]), .Y(n574) );
  INVX1 U511 ( .A(n417), .Y(n613) );
  INVX1 U512 ( .A(n406), .Y(n610) );
  INVX1 U513 ( .A(n414), .Y(n611) );
  INVX1 U514 ( .A(n419), .Y(CC2_DOB) );
  INVX1 U515 ( .A(n416), .Y(n612) );
  INVX1 U516 ( .A(n385), .Y(n606) );
  INVX1 U517 ( .A(n401), .Y(n593) );
  INVX1 U518 ( .A(n384), .Y(n607) );
  INVX1 U519 ( .A(n400), .Y(n597) );
  INVX1 U520 ( .A(n378), .Y(n604) );
  XNOR2XL U521 ( .A(DAC3_V[1]), .B(n261), .Y(n260) );
  NOR2X1 U522 ( .A(n104), .B(n582), .Y(ANAOPT[3]) );
  NOR2X1 U523 ( .A(n104), .B(n327), .Y(ANAOPT[5]) );
  NAND2X1 U524 ( .A(n583), .B(n110), .Y(RD_ENB) );
  NOR21XL U525 ( .B(PWRDN), .A(n615), .Y(VPP_0V) );
  NOR2X1 U526 ( .A(n637), .B(n104), .Y(PWRDN) );
  NOR2X1 U527 ( .A(n105), .B(n261), .Y(DO_SRCCTL[4]) );
  NOR2X1 U528 ( .A(n105), .B(n274), .Y(BCK_REGX[5]) );
  OR2X1 U529 ( .A(sh_hold), .B(n107), .Y(SH_HOLD) );
  NOR2X1 U530 ( .A(n105), .B(n616), .Y(BCK_REGX[4]) );
  NAND2X1 U531 ( .A(n626), .B(n109), .Y(SLEEP) );
  XNOR2XL U532 ( .A(DO_DAC0[8]), .B(DAC1_V[7]), .Y(n323) );
  XNOR2XL U533 ( .A(DO_DAC0[10]), .B(DAC1_V[9]), .Y(n337) );
  XNOR2XL U534 ( .A(DAC1_V[6]), .B(n247), .Y(n319) );
  XNOR2XL U535 ( .A(n273), .B(n274), .Y(n272) );
  NAND21X1 U536 ( .B(n150), .A(N628), .Y(n147) );
  NOR2X1 U537 ( .A(n674), .B(n668), .Y(N628) );
  NOR21XL U538 ( .B(r_srcctl[1]), .A(n98), .Y(DO_SRCCTL[1]) );
  OR2X2 U539 ( .A(pmem_csb), .B(n107), .Y(PMEM_CSB) );
  NAND21X1 U540 ( .B(n673), .A(n202), .Y(n158) );
  INVX1 U541 ( .A(n150), .Y(n202) );
  NAND2X1 U542 ( .A(sll_232_2_A_0_), .B(n653), .Y(N593) );
  NAND2X1 U543 ( .A(n652), .B(n645), .Y(n668) );
  NAND2X1 U544 ( .A(n647), .B(n655), .Y(n659) );
  NAND2X1 U545 ( .A(n650), .B(n665), .Y(n669) );
  NAND2X1 U546 ( .A(n651), .B(n666), .Y(n674) );
  NAND2X1 U547 ( .A(n652), .B(n645), .Y(n658) );
  NAND3X1 U548 ( .A(n655), .B(n656), .C(N593), .Y(n662) );
  NAND3X1 U549 ( .A(n665), .B(n666), .C(sll_232_2_A_0_), .Y(n672) );
  NAND2X1 U550 ( .A(n646), .B(n656), .Y(n664) );
  INVX1 U551 ( .A(atpg_en), .Y(n139) );
  INVX1 U552 ( .A(atpg_en), .Y(n141) );
  NOR2X1 U553 ( .A(n673), .B(n669), .Y(N637) );
  NOR2X1 U554 ( .A(n104), .B(n653), .Y(lt_gpi[0]) );
  INVX1 U555 ( .A(n665), .Y(n651) );
  INVX1 U556 ( .A(n655), .Y(n646) );
  INVX1 U557 ( .A(n656), .Y(n647) );
  INVX1 U558 ( .A(n666), .Y(n650) );
  NAND2X1 U559 ( .A(n636), .B(n108), .Y(OCDRV_ENZ) );
  AOI211X1 U560 ( .C(n357), .D(n263), .A(n262), .B(n257), .Y(n268) );
  AO22X1 U561 ( .A(t_pmem_csb), .B(n639), .C(dm_comp), .D(n253), .Y(n275) );
  AND2X1 U562 ( .A(r_vpp0v_en), .B(ps_pwrdn), .Y(pwrdn_rst) );
  AO222X1 U563 ( .A(slvo_sda), .B(n537), .C(r_dpdmctl[4]), .D(n446), .E(
        comp_smpl[1]), .F(n640), .Y(n269) );
  NAND43X1 U564 ( .B(n456), .C(n455), .D(n454), .A(n453), .Y(DO_GPIO[6]) );
  OA222X1 U565 ( .A(n147), .B(n452), .C(n451), .D(n450), .E(n449), .F(n448), 
        .Y(n453) );
  NAND32X1 U566 ( .B(n234), .C(n233), .A(n231), .Y(DO_GPIO[3]) );
  AOI222XL U567 ( .A(mcu_dbgpo[16]), .B(n284), .C(n228), .D(n538), .E(
        mcu_dbgpo[21]), .F(n533), .Y(n231) );
  OAI22X1 U568 ( .A(n221), .B(n393), .C(n543), .D(n219), .Y(n234) );
  AO2222XL U569 ( .A(n446), .B(r_dpdmctl[6]), .C(upd_dbgpo[17]), .D(n222), .E(
        comp_smpl[2]), .F(n640), .G(n537), .H(n619), .Y(n215) );
  AO21X1 U570 ( .B(mempsrd), .C(hit_ps), .A(n485), .Y(n516) );
  OAI21X1 U571 ( .B(hit_xd), .C(hit_xr), .A(memrd), .Y(n517) );
  AO21X1 U572 ( .B(SRAM_RDAT[0]), .C(n121), .A(n477), .Y(sram_rdat[0]) );
  AO21X1 U573 ( .B(SRAM_RDAT[4]), .C(n108), .A(n481), .Y(n135) );
  AO21X1 U574 ( .B(SRAM_RDAT[5]), .C(n124), .A(n482), .Y(n133) );
  AO21X1 U575 ( .B(SRAM_RDAT[6]), .C(n122), .A(n483), .Y(n131) );
  AO21X1 U576 ( .B(SRAM_RDAT[3]), .C(n124), .A(n480), .Y(n138) );
  AO21X1 U577 ( .B(SRAM_RDAT[1]), .C(n119), .A(n478), .Y(sram_rdat[1]) );
  AO21X1 U578 ( .B(DI_GPIO[3]), .C(n127), .A(n480), .Y(n137) );
  NAND21X1 U579 ( .B(N258), .A(n544), .Y(n550) );
  MUX2X1 U580 ( .D0(di_gpio[0]), .D1(n530), .S(n214), .Y(exint[1]) );
  NAND3X1 U581 ( .A(N266), .B(n634), .C(N268), .Y(n214) );
  MUX2BXL U582 ( .D0(di_gpio[1]), .D1(n529), .S(n217), .Y(n530) );
  NAND3X1 U583 ( .A(N263), .B(n632), .C(N265), .Y(n217) );
  MUX2X1 U584 ( .D0(di_gpio[0]), .D1(n526), .S(n220), .Y(exint[0]) );
  NAND3X1 U585 ( .A(n635), .B(n634), .C(N268), .Y(n220) );
  MUX2X1 U586 ( .D0(di_gpio[1]), .D1(n525), .S(n223), .Y(n526) );
  NAND3X1 U587 ( .A(n633), .B(n632), .C(N265), .Y(n223) );
  MUX2X1 U588 ( .D0(n524), .D1(di_gpio[2]), .S(n224), .Y(n525) );
  NOR3XL U589 ( .A(N260), .B(N261), .C(n629), .Y(n224) );
  NAND21X1 U590 ( .B(n627), .A(n553), .Y(n524) );
  MUX2X1 U591 ( .D0(n528), .D1(n546), .S(n218), .Y(n529) );
  NOR3XL U592 ( .A(n631), .B(N261), .C(n629), .Y(n218) );
  AND3X1 U593 ( .A(n527), .B(N257), .C(N259), .Y(n528) );
  INVX1 U594 ( .A(n523), .Y(n553) );
  NAND21X1 U595 ( .B(N257), .A(n527), .Y(n523) );
  AO21X1 U596 ( .B(SRAM_RDAT[2]), .C(n120), .A(n479), .Y(n140) );
  AO21X1 U597 ( .B(DI_GPIO[1]), .C(n125), .A(n478), .Y(di_gpio[1]) );
  AO21X1 U598 ( .B(DI_GPIO[2]), .C(n121), .A(n479), .Y(di_gpio[2]) );
  AO21X1 U599 ( .B(SRCI[1]), .C(n122), .A(n648), .Y(n126) );
  AO21X1 U600 ( .B(SRCI[0]), .C(n121), .A(n484), .Y(n128) );
  AO21X1 U601 ( .B(IMP_OSC), .C(n120), .A(n483), .Y(di_aswk[4]) );
  OAI21BBX1 U602 ( .A(DRP_OSC), .B(n118), .C(n169), .Y(di_aswk_0) );
  OAI221X1 U603 ( .A(r_dpdo_sel[3]), .B(n367), .C(n368), .D(n600), .E(n369), 
        .Y(n334) );
  NAND4X1 U604 ( .A(n601), .B(n600), .C(n602), .D(n370), .Y(n369) );
  AOI22X1 U605 ( .A(n387), .B(n601), .C(r_dpdo_sel[2]), .D(n388), .Y(n367) );
  AOI22X1 U606 ( .A(n373), .B(n601), .C(r_dpdo_sel[2]), .D(n374), .Y(n368) );
  AND2X1 U607 ( .A(bist_r_ctl[5]), .B(n109), .Y(SRAM_OEB) );
  INVX1 U608 ( .A(r_xana_18), .Y(n583) );
  OAI22X1 U609 ( .A(n381), .B(n602), .C(r_dpdo_sel[1]), .D(n382), .Y(n373) );
  AOI221XL U610 ( .A(n603), .B(pwm_o[0]), .C(n604), .D(pwm_o[1]), .E(n383), 
        .Y(n382) );
  AOI221XL U611 ( .A(n603), .B(di_aswk[2]), .C(r_bck0[3]), .D(n604), .E(n386), 
        .Y(n381) );
  OAI22X1 U612 ( .A(n576), .B(n384), .C(n577), .D(n385), .Y(n383) );
  OAI22X1 U613 ( .A(n375), .B(n602), .C(r_dpdo_sel[1]), .D(n376), .Y(n374) );
  AOI221XL U614 ( .A(r_srcctl[5]), .B(n606), .C(n607), .D(o_dodat5_2_), .E(
        n380), .Y(n375) );
  AOI221XL U615 ( .A(n606), .B(di_aswk_0), .C(n607), .D(di_aswk[4]), .E(n377), 
        .Y(n376) );
  OAI22X1 U616 ( .A(n261), .B(n378), .C(n616), .D(n379), .Y(n380) );
  OAI22X1 U617 ( .A(n389), .B(n602), .C(r_dpdo_sel[1]), .D(n390), .Y(n388) );
  AOI221XL U618 ( .A(n603), .B(n531), .C(n604), .D(di_pro[5]), .E(n394), .Y(
        n389) );
  AOI221XL U619 ( .A(n606), .B(di_pro[2]), .C(n607), .D(n532), .E(n391), .Y(
        n390) );
  OAI22X1 U620 ( .A(n235), .B(n384), .C(n585), .D(n385), .Y(n394) );
  XOR2X1 U621 ( .A(n458), .B(r_aopt[3]), .Y(n582) );
  NAND2X1 U622 ( .A(di_aswk[4]), .B(r_imp_osc), .Y(n458) );
  AO21X1 U623 ( .B(DI_GPIO[0]), .C(n121), .A(n477), .Y(di_gpio[0]) );
  AO21X1 U624 ( .B(RX_DAT), .C(n119), .A(n156), .Y(n123) );
  AO21X1 U625 ( .B(SRCI[5]), .C(n125), .A(n649), .Y(di_pro[5]) );
  AO21X1 U626 ( .B(SRCI[2]), .C(n120), .A(n156), .Y(di_pro[2]) );
  NOR3XL U627 ( .A(N267), .B(N268), .C(N266), .Y(n184) );
  MUX3X1 U628 ( .D0(n554), .D1(di_gpio[2]), .D2(di_gpio[1]), .S0(n188), .S1(
        n186), .Y(n555) );
  NOR3XL U629 ( .A(N267), .B(N268), .C(n635), .Y(n193) );
  MUX3X1 U630 ( .D0(n551), .D1(di_gpio[2]), .D2(di_gpio[1]), .S0(n197), .S1(
        n195), .Y(n552) );
  AO21X1 U631 ( .B(XANAV[0]), .C(n127), .A(n477), .Y(di_xanav[0]) );
  AO21X1 U632 ( .B(SRCI[3]), .C(n120), .A(n276), .Y(n532) );
  AO21X1 U633 ( .B(SRCI[4]), .C(n124), .A(n286), .Y(n531) );
  AO21X1 U634 ( .B(XANAV[1]), .C(n120), .A(n478), .Y(di_xanav[1]) );
  AO21X1 U635 ( .B(CC2_DI), .C(n120), .A(n216), .Y(cc2_di) );
  AOI21X1 U636 ( .B(DM_FAULT), .C(n119), .A(n649), .Y(n235) );
  AOI22AXL U637 ( .A(r_do_ts[6]), .B(n432), .D(r_do_ts[6]), .C(n433), .Y(n294)
         );
  OAI22X1 U638 ( .A(n434), .B(n586), .C(r_do_ts[5]), .D(n435), .Y(n433) );
  OAI22X1 U639 ( .A(n440), .B(n586), .C(r_do_ts[5]), .D(n441), .Y(n432) );
  INVX1 U640 ( .A(r_do_ts[5]), .Y(n586) );
  AO21X1 U641 ( .B(DM_COMP), .C(n122), .A(n252), .Y(dm_comp) );
  OAI21BBX1 U642 ( .A(CC1_DI), .B(n118), .C(n171), .Y(cc1_di) );
  NAND32X1 U643 ( .B(N259), .C(n550), .A(N257), .Y(n551) );
  NAND21X1 U644 ( .B(N259), .A(n553), .Y(n554) );
  OAI21BBX1 U645 ( .A(RX_SQL), .B(n118), .C(n174), .Y(di_sqlch) );
  OAI32X1 U646 ( .A(n605), .B(r_dpdo_sel[1]), .C(n395), .D(n396), .E(n602), 
        .Y(n387) );
  AOI22X1 U647 ( .A(r_dpdmctl[2]), .B(n123), .C(di_sqlch), .D(n624), .Y(n395)
         );
  AOI221XL U648 ( .A(n606), .B(cc1_di), .C(n607), .D(cc2_di), .E(n397), .Y(
        n396) );
  OAI22X1 U649 ( .A(n342), .B(n378), .C(n332), .D(n379), .Y(n397) );
  OAI31XL U650 ( .A(n199), .B(o_cpurst), .C(hit_ps), .D(n200), .Y(mempsack) );
  NOR2X1 U651 ( .A(mempsrd), .B(mempswr), .Y(n199) );
  NAND2X1 U652 ( .A(ictlr_psack), .B(hit_ps), .Y(n200) );
  AOI221XL U653 ( .A(n414), .B(di_aswk[4]), .C(n406), .D(r_vpp_en), .E(n418), 
        .Y(n412) );
  OAI22X1 U654 ( .A(n419), .B(n416), .C(n261), .D(n417), .Y(n418) );
  AOI221XL U655 ( .A(n437), .B(n531), .C(n436), .D(di_pro[5]), .E(n445), .Y(
        n440) );
  ENOX1 U656 ( .A(n235), .B(n444), .C(t_pmem_clk), .D(n588), .Y(n445) );
  AOI22X1 U657 ( .A(n410), .B(n608), .C(r_dndo_sel[3]), .D(n411), .Y(n404) );
  OAI22X1 U658 ( .A(n412), .B(n609), .C(r_dndo_sel[2]), .D(n413), .Y(n411) );
  OAI22X1 U659 ( .A(n420), .B(n609), .C(r_dndo_sel[2]), .D(n421), .Y(n410) );
  AOI221XL U660 ( .A(n406), .B(pwm_o[1]), .C(n414), .D(o_dodat0_15_), .E(n415), 
        .Y(n413) );
  AOI22X1 U661 ( .A(n423), .B(n608), .C(r_dndo_sel[3]), .D(n424), .Y(n403) );
  OAI22X1 U662 ( .A(n425), .B(n609), .C(r_dndo_sel[2]), .D(n426), .Y(n424) );
  OAI22X1 U663 ( .A(n429), .B(n609), .C(r_dndo_sel[2]), .D(n430), .Y(n423) );
  AOI221XL U664 ( .A(r_bck0[4]), .B(n613), .C(n612), .D(CC1_DOB), .E(n428), 
        .Y(n425) );
  INVX1 U665 ( .A(n402), .Y(n573) );
  OAI221X1 U666 ( .A(r_dpdmctl[0]), .B(n403), .C(n404), .D(n625), .E(n405), 
        .Y(n402) );
  INVX1 U667 ( .A(r_dpdmctl[0]), .Y(n625) );
  NAND4X1 U668 ( .A(n406), .B(n407), .C(n609), .D(n608), .Y(n405) );
  AO21X1 U669 ( .B(DP_COMP), .C(n122), .A(n286), .Y(dp_comp) );
  MUX3X1 U670 ( .D0(n547), .D1(n546), .D2(n545), .S0(n232), .S1(n230), .Y(n548) );
  NOR32XL U671 ( .B(N265), .C(N263), .A(n632), .Y(n230) );
  NOR3XL U672 ( .A(n629), .B(n631), .C(n630), .Y(n232) );
  INVX1 U673 ( .A(di_gpio[1]), .Y(n545) );
  OAI22AX1 U674 ( .D(n226), .C(n227), .A(n226), .B(n181), .Y(dpdm_urx) );
  AOI22X1 U675 ( .A(r_i2crout[5]), .B(r_pwrctl[7]), .C(n590), .D(r_pwrctl[6]), 
        .Y(n226) );
  MUX2X1 U676 ( .D0(n549), .D1(n548), .S(n229), .Y(n227) );
  NAND3X1 U677 ( .A(N268), .B(N266), .C(N267), .Y(n229) );
  AND4X1 U678 ( .A(N258), .B(N259), .C(N257), .D(n544), .Y(n547) );
  OAI21BBX1 U679 ( .A(RD_DET), .B(n118), .C(n170), .Y(di_aswk[2]) );
  INVX1 U680 ( .A(n155), .Y(n484) );
  NAND21X1 U681 ( .B(n109), .A(d_dodat[7]), .Y(n155) );
  NAND21X1 U682 ( .B(n111), .A(d_dodat[4]), .Y(n460) );
  INVX1 U683 ( .A(n201), .Y(n482) );
  NAND21X1 U684 ( .B(n141), .A(d_dodat[5]), .Y(n201) );
  INVX1 U685 ( .A(n159), .Y(n480) );
  NAND21X1 U686 ( .B(n113), .A(d_dodat[3]), .Y(n159) );
  OAI22X1 U687 ( .A(dp_comp), .B(n590), .C(r_i2crout[5]), .D(dm_comp), .Y(n181) );
  OAI22X1 U688 ( .A(r_i2crout[5]), .B(dp_comp), .C(dm_comp), .D(n590), .Y(n192) );
  OAI22X1 U689 ( .A(r_i2crout[4]), .B(cc2_di), .C(cc1_di), .D(n591), .Y(n178)
         );
  OAI22X1 U690 ( .A(cc2_di), .B(n591), .C(r_i2crout[4]), .D(cc1_di), .Y(n190)
         );
  NAND4X1 U691 ( .A(n493), .B(n494), .C(n495), .D(n496), .Y(DO_GPIO[2]) );
  AOI22X1 U692 ( .A(n497), .B(di_sqlch), .C(mcu_dbgpo[20]), .D(n498), .Y(n496)
         );
  AOI22X1 U693 ( .A(N448), .B(n538), .C(cc1_di), .D(n537), .Y(n495) );
  AOI22X1 U694 ( .A(n640), .B(n4), .C(t_pmem_clk), .D(n639), .Y(n493) );
  INVX1 U695 ( .A(n194), .Y(n483) );
  NAND21X1 U696 ( .B(n112), .A(d_dodat[6]), .Y(n194) );
  INVX1 U697 ( .A(n144), .Y(n477) );
  NAND21X1 U698 ( .B(n108), .A(d_dodat[0]), .Y(n144) );
  INVX1 U699 ( .A(n162), .Y(n479) );
  NAND21X1 U700 ( .B(n108), .A(d_dodat[2]), .Y(n162) );
  AO21X1 U701 ( .B(DI_GPIO[5]), .C(n125), .A(n482), .Y(di_gpio[5]) );
  AO21X1 U702 ( .B(DI_GPIO[6]), .C(n122), .A(n483), .Y(di_gpio[6]) );
  AO22AXL U703 ( .A(mcu_dbgpo[19]), .B(n534), .C(n357), .D(n472), .Y(n209) );
  XNOR2XL U704 ( .A(pwm_o[1]), .B(do_p0[5]), .Y(n472) );
  INVX1 U705 ( .A(n148), .Y(n478) );
  NAND21X1 U706 ( .B(n114), .A(d_dodat[1]), .Y(n148) );
  OAI21BBX1 U707 ( .A(DI_TS), .B(n115), .C(n171), .Y(di_ts) );
  MUX2X1 U708 ( .D0(n558), .D1(n557), .S(N259), .Y(n228) );
  MUX4X1 U709 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N257), .S1(N258), .Y(n557) );
  MUX4X1 U710 ( .D0(do_opt_0), .D1(do_opt_1), .D2(do_p0[0]), .D3(do_p0[1]), 
        .S0(N257), .S1(N258), .Y(n558) );
  MUX2X1 U711 ( .D0(n560), .D1(n559), .S(N262), .Y(N448) );
  MUX4X1 U712 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N260), .S1(N261), .Y(n559) );
  MUX4X1 U713 ( .D0(do_opt_0), .D1(do_opt_1), .D2(do_p0[0]), .D3(do_p0[1]), 
        .S0(N260), .S1(N261), .Y(n560) );
  XOR2X1 U714 ( .A(do_p0[4]), .B(pwm_o[0]), .Y(n263) );
  AO21X1 U715 ( .B(XANAV[2]), .C(n119), .A(n479), .Y(di_xanav[2]) );
  AO21X1 U716 ( .B(XANAV[3]), .C(n109), .A(n480), .Y(di_xanav[3]) );
  AO21X1 U717 ( .B(XANAV[4]), .C(n127), .A(n481), .Y(di_xanav[4]) );
  AO21X1 U718 ( .B(XANAV[5]), .C(n121), .A(n482), .Y(di_xanav[5]) );
  INVX1 U719 ( .A(n149), .Y(n204) );
  OAI211X1 U720 ( .C(di_tst), .D(r_gpio_tm), .A(i_rstz), .B(n119), .Y(n149) );
  OAI21X1 U721 ( .B(hwi2c_stretch), .C(pmem_pgm), .A(r_strtch), .Y(n361) );
  INVX1 U722 ( .A(dacmux_sel[10]), .Y(n617) );
  MUX2X1 U723 ( .D0(n564), .D1(n563), .S(N268), .Y(DO_GPIO[0]) );
  MUX4X1 U724 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N266), .S1(N267), .Y(n563) );
  MUX4X1 U725 ( .D0(do_opt_0), .D1(do_opt_1), .D2(do_p0[0]), .D3(do_p0[1]), 
        .S0(N266), .S1(N267), .Y(n564) );
  MUX2X1 U726 ( .D0(n562), .D1(n561), .S(N265), .Y(DO_GPIO[1]) );
  MUX4X1 U727 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N263), .S1(N264), .Y(n561) );
  MUX4X1 U728 ( .D0(do_opt_0), .D1(do_opt_1), .D2(do_p0[0]), .D3(do_p0[1]), 
        .S0(N263), .S1(N264), .Y(n562) );
  AND3X1 U729 ( .A(n356), .B(i_rstz), .C(n556), .Y(n320) );
  OAI21X1 U730 ( .B(n347), .C(n320), .A(n302), .Y(n249) );
  NOR21XL U731 ( .B(r_gpio_oe[2]), .A(n348), .Y(n347) );
  AOI221XL U732 ( .A(n314), .B(n631), .C(n349), .D(n629), .E(n350), .Y(n348)
         );
  OAI21X1 U733 ( .B(do_opt_1), .C(n631), .A(n630), .Y(n349) );
  OAI21X1 U734 ( .B(n355), .C(n320), .A(n302), .Y(n248) );
  NOR21XL U735 ( .B(r_gpio_oe[3]), .A(n358), .Y(n355) );
  AOI221XL U736 ( .A(n314), .B(n628), .C(n359), .D(n627), .E(n360), .Y(n358)
         );
  AOI31X1 U737 ( .A(N257), .B(n641), .C(N258), .D(n627), .Y(n360) );
  NAND2X1 U738 ( .A(d_dodat[13]), .B(n103), .Y(n171) );
  NAND2X1 U739 ( .A(d_dodat[14]), .B(n103), .Y(n170) );
  NAND2X1 U740 ( .A(d_dodat[15]), .B(n103), .Y(n169) );
  NAND2X1 U741 ( .A(d_dodat[8]), .B(n104), .Y(n176) );
  NOR3XL U742 ( .A(r_gpio_oe[5]), .B(n638), .C(n320), .Y(n246) );
  NOR3XL U743 ( .A(r_gpio_oe[6]), .B(n638), .C(n320), .Y(n245) );
  NOR2X1 U744 ( .A(r_gpio_oe[4]), .B(n320), .Y(n247) );
  NAND3X1 U745 ( .A(n311), .B(n302), .C(r_gpio_oe[1]), .Y(n250) );
  OAI221X1 U746 ( .A(N265), .B(n312), .C(N263), .D(do_opt_0), .E(n313), .Y(
        n311) );
  OAI31XL U747 ( .A(n632), .B(s0_rxdoe), .C(n633), .D(N265), .Y(n313) );
  AOI21X1 U748 ( .B(N263), .C(n305), .A(N264), .Y(n312) );
  NAND3X1 U749 ( .A(n301), .B(n302), .C(r_gpio_oe[0]), .Y(n251) );
  OAI221X1 U750 ( .A(N268), .B(n303), .C(N266), .D(do_opt_0), .E(n304), .Y(
        n301) );
  OAI31XL U751 ( .A(n634), .B(s0_rxdoe), .C(n635), .D(N268), .Y(n304) );
  AOI21X1 U752 ( .B(N266), .C(n305), .A(N267), .Y(n303) );
  INVX1 U753 ( .A(sh_rst), .Y(n618) );
  OAI22X1 U754 ( .A(slvo_sda), .B(n598), .C(mcuo_sda), .D(n594), .Y(n305) );
  NAND21X1 U755 ( .B(n112), .A(d_dodat[12]), .Y(n172) );
  NAND21X1 U756 ( .B(n127), .A(d_dodat[11]), .Y(n173) );
  NAND21X1 U757 ( .B(n110), .A(d_dodat[9]), .Y(n175) );
  AOI22X1 U758 ( .A(xram_a[7]), .B(xram_ce), .C(iram_a[7]), .D(iram_ce), .Y(
        n239) );
  AOI22XL U759 ( .A(xram_a[2]), .B(xram_ce), .C(iram_a[2]), .D(iram_ce), .Y(
        n242) );
  AO21X1 U760 ( .B(n305), .C(N257), .A(N258), .Y(n359) );
  OA21X1 U761 ( .B(n284), .C(n291), .A(mcu_dbgpo[18]), .Y(n262) );
  NOR2X1 U762 ( .A(n589), .B(r_do_ts[4]), .Y(n436) );
  NOR2X1 U763 ( .A(r_do_ts[3]), .B(r_do_ts[4]), .Y(n437) );
  NOR2X1 U764 ( .A(r_i2cmcu_route[0]), .B(r_i2cmcu_route[1]), .Y(n183) );
  NOR2X1 U765 ( .A(r_i2cslv_route[0]), .B(r_i2cslv_route[1]), .Y(n179) );
  OR2XL U766 ( .A(r_fortxen), .B(ptx_oe), .Y(n619) );
  NAND2X1 U767 ( .A(d_dodat[10]), .B(n104), .Y(n174) );
  NAND2X1 U768 ( .A(r_do_ts[4]), .B(r_do_ts[3]), .Y(n444) );
  NAND2X1 U769 ( .A(r_do_ts[4]), .B(n589), .Y(n439) );
  AOI221XL U770 ( .A(n587), .B(x_clk), .C(divff_o1), .D(n588), .E(n436), .Y(
        n435) );
  INVX1 U771 ( .A(r_do_ts[3]), .Y(n589) );
  AOI31X1 U772 ( .A(N260), .B(n641), .C(N261), .D(n629), .Y(n350) );
  MUX2IX1 U773 ( .D0(ptx_cc), .D1(r_fortxdat), .S(r_fortxrdy), .Y(n342) );
  AO22X1 U774 ( .A(n8), .B(xram_a[9]), .C(n39), .D(iram_a[9]), .Y(SRAM_A[9])
         );
  NOR2X1 U775 ( .A(n595), .B(r_i2cmcu_route[1]), .Y(n182) );
  NOR2X1 U776 ( .A(n599), .B(r_i2cslv_route[1]), .Y(n177) );
  INVX1 U777 ( .A(N259), .Y(n627) );
  INVX1 U778 ( .A(N264), .Y(n632) );
  INVX1 U779 ( .A(N260), .Y(n631) );
  INVX1 U780 ( .A(N266), .Y(n635) );
  INVX1 U781 ( .A(N263), .Y(n633) );
  INVX1 U782 ( .A(N262), .Y(n629) );
  INVX1 U783 ( .A(N267), .Y(n634) );
  INVX1 U784 ( .A(r_i2cmcu_route[0]), .Y(n595) );
  INVX1 U785 ( .A(r_i2cslv_route[0]), .Y(n599) );
  INVX1 U786 ( .A(N261), .Y(n630) );
  INVX1 U787 ( .A(N257), .Y(n628) );
  INVX1 U788 ( .A(pmem_re), .Y(n168) );
  INVX1 U789 ( .A(pmem_pgm), .Y(n448) );
  INVX1 U790 ( .A(fcp_do), .Y(n180) );
  NOR21XL U791 ( .B(r_do_ts[2]), .A(n98), .Y(DO_TS[2]) );
  AOI221XL U792 ( .A(t_osc_gate), .B(n613), .C(n612), .D(n267), .E(n427), .Y(
        n426) );
  OAI22X1 U793 ( .A(n577), .B(n611), .C(n581), .D(n610), .Y(n427) );
  OAI22X1 U794 ( .A(r_i2crout[4]), .B(n504), .C(n591), .D(n505), .Y(n419) );
  NOR21XL U795 ( .B(esfrm_rrdy), .A(prl_cany0), .Y(sse_rdrdy) );
  OAI22X1 U796 ( .A(n591), .B(n504), .C(r_i2crout[4]), .D(n505), .Y(n273) );
  OAI22X1 U797 ( .A(slvo_sda), .B(n596), .C(mcuo_sda), .D(n592), .Y(n505) );
  NAND21X1 U798 ( .B(r_bck0[2]), .A(n506), .Y(n267) );
  NAND21X1 U799 ( .B(r_bck2_2_), .A(gating_pwr), .Y(n506) );
  NOR2X1 U800 ( .A(r_dndo_sel[0]), .B(r_dndo_sel[1]), .Y(n406) );
  NOR2X1 U801 ( .A(n614), .B(r_dndo_sel[1]), .Y(n414) );
  OAI21BBX1 U802 ( .A(r_xtm[7]), .B(n636), .C(r_aopt[5]), .Y(n327) );
  NAND2X1 U803 ( .A(r_dpdmctl[2]), .B(n605), .Y(n378) );
  NAND2X1 U804 ( .A(r_dpdo_sel[0]), .B(r_dpdmctl[2]), .Y(n384) );
  NAND2X1 U805 ( .A(r_dndo_sel[1]), .B(r_dndo_sel[0]), .Y(n416) );
  NAND2X1 U806 ( .A(r_dndo_sel[1]), .B(n614), .Y(n417) );
  NAND2X1 U807 ( .A(r_dpdo_sel[0]), .B(n624), .Y(n385) );
  OAI21X1 U808 ( .B(r_pwrctl[7]), .C(n362), .A(n363), .Y(n341) );
  OAI21X1 U809 ( .B(s0_rxdoe), .C(n590), .A(r_pwrctl[7]), .Y(n363) );
  AOI222XL U810 ( .A(r_dpdmctl[3]), .B(n364), .C(n365), .D(n590), .E(
        r_i2crout[5]), .F(n366), .Y(n362) );
  INVX1 U811 ( .A(r_ocdrv_enz), .Y(n636) );
  INVX1 U812 ( .A(r_pwrdn), .Y(n637) );
  NAND31X1 U813 ( .C(r_otpi_gate), .A(n447), .B(r_srcctl[4]), .Y(n261) );
  NAND21X1 U814 ( .B(sdischg_duty), .A(r_sdischg[6]), .Y(n447) );
  OAI211X1 U815 ( .C(r_pwrctl[6]), .D(n398), .A(n399), .B(n450), .Y(n326) );
  OAI21X1 U816 ( .B(r_i2crout[5]), .C(s0_rxdoe), .A(r_pwrctl[6]), .Y(n399) );
  AOI222XL U817 ( .A(r_dpdmctl[1]), .B(n364), .C(r_i2crout[5]), .D(n365), .E(
        n366), .F(n590), .Y(n398) );
  ENOX1 U818 ( .A(fcp_oe), .B(n408), .C(fcp_do), .D(fcp_oe), .Y(n407) );
  AOI32X1 U819 ( .A(n364), .B(n622), .C(r_dpdmctl[0]), .D(r_pwrctl[6]), .E(
        n409), .Y(n408) );
  INVX1 U820 ( .A(r_pwrctl[6]), .Y(n622) );
  OAI22X1 U821 ( .A(r_i2crout[5]), .B(n643), .C(n590), .D(n642), .Y(n409) );
  NOR2X1 U822 ( .A(frc_lg_on), .B(r_bck0[5]), .Y(n274) );
  INVX1 U823 ( .A(r_dpdo_sel[0]), .Y(n605) );
  INVX1 U824 ( .A(r_dpdmctl[2]), .Y(n624) );
  INVX1 U825 ( .A(r_i2crout[4]), .Y(n591) );
  INVX1 U826 ( .A(r_dndo_sel[0]), .Y(n614) );
  INVX1 U827 ( .A(r_vpp0v_en), .Y(n615) );
  INVX1 U828 ( .A(r_sleep), .Y(n626) );
  AND2X1 U829 ( .A(esfrm_rrdy), .B(prl_cany0), .Y(upd_rdrdy) );
  NAND2X1 U830 ( .A(r_i2cslv_route[1]), .B(n599), .Y(n400) );
  NAND2X1 U831 ( .A(r_i2cmcu_route[1]), .B(n595), .Y(n401) );
  INVX1 U832 ( .A(r_i2crout[5]), .Y(n590) );
  OAI22X1 U833 ( .A(slvo_sda), .B(n400), .C(mcuo_sda), .D(n401), .Y(n365) );
  NOR2X1 U834 ( .A(r_dpdo_sel[0]), .B(n371), .Y(n370) );
  AOI32X1 U835 ( .A(n364), .B(n621), .C(r_dpdmctl[2]), .D(r_pwrctl[7]), .E(
        n372), .Y(n371) );
  INVX1 U836 ( .A(r_pwrctl[7]), .Y(n621) );
  OAI22X1 U837 ( .A(n590), .B(n643), .C(r_i2crout[5]), .D(n642), .Y(n372) );
  INVX1 U838 ( .A(do_opt[6]), .Y(n642) );
  INVX1 U839 ( .A(do_opt[7]), .Y(n643) );
  INVX1 U840 ( .A(r_bck0[4]), .Y(n616) );
  INVX1 U841 ( .A(PWREN_HOLD), .Y(n585) );
  INVX1 U842 ( .A(r_dpdo_sel[1]), .Y(n602) );
  INVX1 U843 ( .A(r_dndo_sel[2]), .Y(n609) );
  INVX1 U844 ( .A(r_dndo_sel[3]), .Y(n608) );
  INVX1 U845 ( .A(r_dpdo_sel[2]), .Y(n601) );
  OR2XL U846 ( .A(mcu_ram_r), .B(mcu_ram_w), .Y(ramacc) );
  INVX1 U847 ( .A(r_dpdo_sel[3]), .Y(n600) );
  NOR21XL U848 ( .B(r_xana[15]), .A(n99), .Y(ANA_REGX[15]) );
  NOR21XL U849 ( .B(r_xana[13]), .A(n98), .Y(ANA_REGX[13]) );
  NOR21XL U850 ( .B(r_xana[14]), .A(n99), .Y(ANA_REGX[14]) );
  NOR21XL U851 ( .B(r_xana[1]), .A(n101), .Y(ANA_REGX[1]) );
  NOR21XL U852 ( .B(r_xana[3]), .A(n102), .Y(ANA_REGX[3]) );
  NOR21XL U853 ( .B(r_regtrm[0]), .A(atpg_en), .Y(REGTRM[0]) );
  NOR21XL U854 ( .B(r_regtrm[1]), .A(n94), .Y(REGTRM[1]) );
  NOR21XL U855 ( .B(r_regtrm[2]), .A(n93), .Y(REGTRM[2]) );
  NOR21XL U856 ( .B(r_regtrm[3]), .A(n96), .Y(REGTRM[3]) );
  NOR21XL U859 ( .B(r_regtrm[4]), .A(n91), .Y(REGTRM[4]) );
  NOR21XL U860 ( .B(r_regtrm[5]), .A(n90), .Y(REGTRM[5]) );
  NOR21XL U861 ( .B(r_regtrm[6]), .A(n90), .Y(REGTRM[6]) );
  NOR21XL U862 ( .B(r_regtrm[7]), .A(n90), .Y(REGTRM[7]) );
  NOR21XL U863 ( .B(r_regtrm[8]), .A(n90), .Y(REGTRM[8]) );
  NOR21XL U864 ( .B(r_regtrm[9]), .A(n89), .Y(REGTRM[9]) );
  NOR21XL U865 ( .B(r_regtrm[10]), .A(n136), .Y(REGTRM[10]) );
  NOR21XL U866 ( .B(r_regtrm[11]), .A(n132), .Y(REGTRM[11]) );
  NOR21XL U867 ( .B(r_regtrm[12]), .A(n130), .Y(REGTRM[12]) );
  NOR21XL U868 ( .B(r_regtrm[13]), .A(n94), .Y(REGTRM[13]) );
  NOR21XL U869 ( .B(r_regtrm[14]), .A(n94), .Y(REGTRM[14]) );
  NOR21XL U870 ( .B(r_regtrm[15]), .A(n94), .Y(REGTRM[15]) );
  NOR21XL U871 ( .B(r_regtrm[16]), .A(n94), .Y(REGTRM[16]) );
  NOR21XL U872 ( .B(r_regtrm[17]), .A(n94), .Y(REGTRM[17]) );
  NOR21XL U873 ( .B(r_regtrm[18]), .A(n94), .Y(REGTRM[18]) );
  NOR21XL U874 ( .B(r_regtrm[19]), .A(n94), .Y(REGTRM[19]) );
  NOR21XL U875 ( .B(r_regtrm[20]), .A(n94), .Y(REGTRM[20]) );
  NOR21XL U876 ( .B(r_regtrm[21]), .A(n94), .Y(REGTRM[21]) );
  NOR21XL U877 ( .B(r_regtrm[22]), .A(n93), .Y(REGTRM[22]) );
  NOR21XL U878 ( .B(r_regtrm[23]), .A(n93), .Y(REGTRM[23]) );
  NOR21XL U879 ( .B(r_regtrm[24]), .A(n93), .Y(REGTRM[24]) );
  NOR21XL U880 ( .B(r_regtrm[25]), .A(n93), .Y(REGTRM[25]) );
  NOR21XL U881 ( .B(r_regtrm[26]), .A(n93), .Y(REGTRM[26]) );
  NOR21XL U882 ( .B(r_regtrm[27]), .A(n93), .Y(REGTRM[27]) );
  NOR21XL U883 ( .B(r_regtrm[28]), .A(n93), .Y(REGTRM[28]) );
  NOR21XL U884 ( .B(r_regtrm[29]), .A(n93), .Y(REGTRM[29]) );
  NOR21XL U885 ( .B(r_regtrm[30]), .A(n93), .Y(REGTRM[30]) );
  NOR21XL U886 ( .B(r_regtrm[31]), .A(n92), .Y(REGTRM[31]) );
  NOR21XL U887 ( .B(r_regtrm[32]), .A(n92), .Y(REGTRM[32]) );
  NOR21XL U888 ( .B(r_regtrm[33]), .A(n92), .Y(REGTRM[33]) );
  NOR21XL U889 ( .B(r_regtrm[34]), .A(n92), .Y(REGTRM[34]) );
  NOR21XL U890 ( .B(r_regtrm[35]), .A(n92), .Y(REGTRM[35]) );
  NOR21XL U891 ( .B(r_regtrm[36]), .A(n92), .Y(REGTRM[36]) );
  NOR21XL U892 ( .B(r_regtrm[37]), .A(n92), .Y(REGTRM[37]) );
  NOR21XL U893 ( .B(r_regtrm[38]), .A(n92), .Y(REGTRM[38]) );
  NOR21XL U894 ( .B(r_regtrm[39]), .A(n92), .Y(REGTRM[39]) );
  NOR21XL U895 ( .B(r_regtrm[40]), .A(n92), .Y(REGTRM[40]) );
  NOR21XL U896 ( .B(r_regtrm[41]), .A(n91), .Y(REGTRM[41]) );
  NOR21XL U897 ( .B(r_regtrm[42]), .A(n91), .Y(REGTRM[42]) );
  NOR21XL U898 ( .B(r_regtrm[43]), .A(n91), .Y(REGTRM[43]) );
  NOR21XL U899 ( .B(r_regtrm[44]), .A(n91), .Y(REGTRM[44]) );
  NOR21XL U900 ( .B(r_regtrm[45]), .A(n91), .Y(REGTRM[45]) );
  NOR21XL U901 ( .B(r_regtrm[46]), .A(n91), .Y(REGTRM[46]) );
  NOR21XL U902 ( .B(r_regtrm[47]), .A(n91), .Y(REGTRM[47]) );
  NOR21XL U903 ( .B(r_regtrm[48]), .A(n91), .Y(REGTRM[48]) );
  NOR21XL U904 ( .B(r_regtrm[49]), .A(n91), .Y(REGTRM[49]) );
  NOR21XL U905 ( .B(r_regtrm[50]), .A(n90), .Y(REGTRM[50]) );
  NOR21XL U906 ( .B(r_regtrm[51]), .A(n90), .Y(REGTRM[51]) );
  NOR21XL U907 ( .B(r_regtrm[52]), .A(n90), .Y(REGTRM[52]) );
  NOR21XL U908 ( .B(r_regtrm[53]), .A(n90), .Y(REGTRM[53]) );
  NOR21XL U909 ( .B(r_regtrm[54]), .A(n90), .Y(REGTRM[54]) );
  NOR21XL U910 ( .B(r_regtrm[55]), .A(n90), .Y(REGTRM[55]) );
  NOR21XL U911 ( .B(r_aopt[0]), .A(n96), .Y(ANAOPT[0]) );
  NOR21XL U912 ( .B(r_aopt[2]), .A(n97), .Y(ANAOPT[2]) );
  NOR21XL U913 ( .B(r_aopt[6]), .A(n97), .Y(ANAOPT[6]) );
  NOR21XL U914 ( .B(r_aopt[7]), .A(n98), .Y(ANAOPT[7]) );
  NOR21XL U915 ( .B(r_accctl[3]), .A(n99), .Y(DO_DPDN[5]) );
  NOR21XL U916 ( .B(r_xana[5]), .A(n98), .Y(ANA_REGX[5]) );
  NOR21XL U917 ( .B(r_vpp_en), .A(n88), .Y(VPP_SEL) );
  NOR21XL U918 ( .B(r_sdischg[7]), .A(n95), .Y(LDO3P9V) );
  NOR21XL U919 ( .B(r_ana_tm[0]), .A(n102), .Y(ANA_TM[0]) );
  NOR21XL U920 ( .B(r_ana_tm[1]), .A(n103), .Y(ANA_TM[1]) );
  NOR21XL U921 ( .B(r_ana_tm[2]), .A(n103), .Y(ANA_TM[2]) );
  NOR21XL U922 ( .B(r_ana_tm[3]), .A(n102), .Y(ANA_TM[3]) );
  NOR21XL U923 ( .B(r_xana[7]), .A(n100), .Y(ANA_REGX[7]) );
  NOR21XL U924 ( .B(r_srcctl[5]), .A(n98), .Y(DO_SRCCTL[5]) );
  NOR21XL U925 ( .B(r_xana_23), .A(n95), .Y(LFOSC_ENB) );
  NOR21XL U926 ( .B(r_xana[0]), .A(n98), .Y(ANA_REGX[0]) );
  NOR21XL U927 ( .B(r_srcctl[6]), .A(n97), .Y(DO_SRCCTL[6]) );
  NOR21XL U928 ( .B(r_srcctl[7]), .A(n98), .Y(DO_SRCCTL[7]) );
  NOR21XL U929 ( .B(r_dpdmctl[4]), .A(n100), .Y(DO_DPDN[1]) );
  NOR21XL U930 ( .B(r_dpdmctl[5]), .A(n99), .Y(DO_DPDN[2]) );
  NOR21XL U931 ( .B(r_xana[10]), .A(n98), .Y(ANA_REGX[10]) );
  NOR21XL U932 ( .B(r_xana[11]), .A(n99), .Y(ANA_REGX[11]) );
  NOR21XL U933 ( .B(r_dpdmctl[7]), .A(n99), .Y(DO_DPDN[4]) );
  NOR21XL U934 ( .B(r_accctl[4]), .A(n99), .Y(DO_DPDN[0]) );
  NOR21XL U935 ( .B(x_daclsb[2]), .A(n101), .Y(DAC1_EN) );
  NOR21XL U936 ( .B(r_cctrx[7]), .A(n100), .Y(DO_CCTRX[7]) );
  NOR21XL U937 ( .B(r_cctrx[6]), .A(n100), .Y(DO_CCTRX[6]) );
  NOR21XL U938 ( .B(r_cctrx[5]), .A(n99), .Y(DO_CCTRX[5]) );
  NOR21XL U939 ( .B(r_cctrx[4]), .A(n100), .Y(DO_CCTRX[4]) );
  NOR21XL U940 ( .B(r_xtm[0]), .A(n88), .Y(XTM[0]) );
  NOR21XL U941 ( .B(r_xtm[1]), .A(n88), .Y(XTM[1]) );
  NOR21XL U942 ( .B(r_xtm[2]), .A(n87), .Y(XTM[2]) );
  NOR21XL U943 ( .B(r_xtm[3]), .A(n87), .Y(XTM[3]) );
  NOR21XL U944 ( .B(r_cctrx[0]), .A(n97), .Y(DO_CCTRX[0]) );
  NOR21XL U945 ( .B(r_ccctl[7]), .A(n99), .Y(DO_CCCTL[7]) );
  NOR21XL U946 ( .B(r_ccctl[6]), .A(n101), .Y(DO_CCCTL[6]) );
  NOR21XL U947 ( .B(r_ccctl[4]), .A(n100), .Y(DO_CCCTL[4]) );
  NOR21XL U948 ( .B(r_ccctl[5]), .A(n101), .Y(DO_CCCTL[5]) );
  NOR21XL U949 ( .B(r_bck0[7]), .A(n102), .Y(BCK_REGX[7]) );
  NOR21XL U950 ( .B(r_bck1[7]), .A(n102), .Y(BCK_REGX[15]) );
  NOR21XL U951 ( .B(r_bck1[6]), .A(n101), .Y(BCK_REGX[14]) );
  NOR21XL U952 ( .B(r_bck1[5]), .A(n103), .Y(BCK_REGX[13]) );
  NOR21XL U953 ( .B(r_bck1[4]), .A(n103), .Y(BCK_REGX[12]) );
  NOR21XL U954 ( .B(r_bck1[3]), .A(n102), .Y(BCK_REGX[11]) );
  NOR21XL U955 ( .B(r_bck1[2]), .A(n103), .Y(BCK_REGX[10]) );
  NOR21XL U956 ( .B(r_bck1[0]), .A(n101), .Y(BCK_REGX[8]) );
  NOR21XL U957 ( .B(r_bck1[1]), .A(n102), .Y(BCK_REGX[9]) );
  NOR21XL U958 ( .B(r_bck0[6]), .A(n102), .Y(BCK_REGX[6]) );
  NOR21XL U959 ( .B(r_bck0[3]), .A(n102), .Y(BCK_REGX[3]) );
  NOR21XL U960 ( .B(r_bck0[1]), .A(n101), .Y(BCK_REGX[1]) );
  NOR21XL U961 ( .B(r_bck0[0]), .A(n102), .Y(BCK_REGX[0]) );
  NOR2X1 U962 ( .A(n105), .B(n623), .Y(DO_DPDN[3]) );
  INVX1 U963 ( .A(r_dpdmctl[6]), .Y(n623) );
  NOR2X1 U964 ( .A(n105), .B(n620), .Y(DO_CCCTL[0]) );
  INVX1 U965 ( .A(r_ccctl[0]), .Y(n620) );
  OR2X1 U966 ( .A(r_cctrx[2]), .B(n107), .Y(DO_CCTRX[2]) );
  OR2X1 U967 ( .A(r_cctrx[1]), .B(n107), .Y(DO_CCTRX[1]) );
  INVX1 U968 ( .A(sfr_intr[2]), .Y(n29) );
  NOR21XL U969 ( .B(i2c_ev_3), .A(sse_adr[7]), .Y(i2c_ev_2) );
  AO21X1 U970 ( .B(PMEM_Q1[7]), .C(n124), .A(n484), .Y(pmem_q1[7]) );
  OAI21BBX1 U971 ( .A(PMEM_Q0[7]), .B(n116), .C(n169), .Y(pmem_q0[7]) );
  AO21X1 U972 ( .B(PMEM_Q1[1]), .C(n122), .A(n478), .Y(pmem_q1[1]) );
  OAI21BBX1 U973 ( .A(PMEM_Q0[1]), .B(n118), .C(n175), .Y(pmem_q0[1]) );
  AO21X1 U974 ( .B(PMEM_Q1[2]), .C(n125), .A(n479), .Y(pmem_q1[2]) );
  OAI21BBX1 U975 ( .A(PMEM_Q0[2]), .B(n116), .C(n174), .Y(pmem_q0[2]) );
  AO21X1 U976 ( .B(PMEM_Q1[3]), .C(n124), .A(n480), .Y(pmem_q1[3]) );
  OAI21BBX1 U977 ( .A(PMEM_Q0[3]), .B(n115), .C(n173), .Y(pmem_q0[3]) );
  AO21X1 U978 ( .B(PMEM_Q1[5]), .C(n127), .A(n482), .Y(pmem_q1[5]) );
  OAI21BBX1 U979 ( .A(PMEM_Q0[5]), .B(n116), .C(n171), .Y(pmem_q0[5]) );
  AO21X1 U980 ( .B(PMEM_Q1[6]), .C(n124), .A(n483), .Y(pmem_q1[6]) );
  OAI21BBX1 U981 ( .A(PMEM_Q0[6]), .B(n115), .C(n170), .Y(pmem_q0[6]) );
  OAI21BBX1 U982 ( .A(PMEM_Q0[4]), .B(n116), .C(n172), .Y(pmem_q0[4]) );
  AO21X1 U983 ( .B(PMEM_Q1[4]), .C(n125), .A(n481), .Y(pmem_q1[4]) );
  AO21X1 U984 ( .B(PMEM_Q1[0]), .C(n121), .A(n477), .Y(pmem_q1[0]) );
  OAI21BBX1 U985 ( .A(PMEM_Q0[0]), .B(n115), .C(n176), .Y(pmem_q0[0]) );
  INVX1 U986 ( .A(sfr_intr[3]), .Y(n30) );
  INVX1 U987 ( .A(r_i2c_ninc), .Y(n28) );
  NOR3XL U988 ( .A(N261), .B(N262), .C(N260), .Y(n188) );
  NOR3XL U989 ( .A(N261), .B(N262), .C(n631), .Y(n197) );
  NOR3XL U990 ( .A(N264), .B(N265), .C(N263), .Y(n186) );
  NOR3XL U991 ( .A(N264), .B(N265), .C(n633), .Y(n195) );
  AO21X1 U992 ( .B(t_di_gpio4), .C(n125), .A(n481), .Y(di_gpio[4]) );
  NOR21X2 U993 ( .B(pmem_re), .A(n136), .Y(PMEM_RE) );
  NOR21X1 U994 ( .B(pmem_clk[1]), .A(n95), .Y(PMEM_CLK[1]) );
  NOR21X1 U995 ( .B(pmem_clk[0]), .A(n95), .Y(PMEM_CLK[0]) );
  NOR21XL U996 ( .B(di_tst), .A(N593), .Y(tm_atpg) );
  NOR21XL U997 ( .B(r_do_ts[1]), .A(n97), .Y(DO_TS[1]) );
  NOR21XL U998 ( .B(r_do_ts[0]), .A(n98), .Y(DO_TS[0]) );
  NOR21XL U999 ( .B(r_pu_gpio[6]), .A(n95), .Y(GPIO_PU[6]) );
  NOR21XL U1000 ( .B(r_pu_gpio[5]), .A(n95), .Y(GPIO_PU[5]) );
  NOR21XL U1001 ( .B(r_pu_gpio[4]), .A(n95), .Y(GPIO_PU[4]) );
  NOR21XL U1002 ( .B(r_pd_gpio[3]), .A(n96), .Y(GPIO_PD[3]) );
  NOR21XL U1003 ( .B(r_pd_gpio[2]), .A(n96), .Y(GPIO_PD[2]) );
  NOR21XL U1004 ( .B(r_pd_gpio[1]), .A(n96), .Y(GPIO_PD[1]) );
  NOR21XL U1005 ( .B(r_pd_gpio[0]), .A(n96), .Y(GPIO_PD[0]) );
  NOR21XL U1006 ( .B(r_pd_gpio[6]), .A(n96), .Y(GPIO_PD[6]) );
  NOR21XL U1007 ( .B(r_pd_gpio[5]), .A(n96), .Y(GPIO_PD[5]) );
  NOR21XL U1008 ( .B(r_pd_gpio[4]), .A(n96), .Y(GPIO_PD[4]) );
  NOR21XL U1009 ( .B(r_pu_gpio[3]), .A(n95), .Y(GPIO_PU[3]) );
  NOR21XL U1010 ( .B(r_pu_gpio[2]), .A(n95), .Y(GPIO_PU[2]) );
  NOR21XL U1011 ( .B(r_pu_gpio[1]), .A(n95), .Y(GPIO_PU[1]) );
  NOR21XL U1012 ( .B(r_pu_gpio[0]), .A(n96), .Y(GPIO_PU[0]) );
  NAND21X1 U1013 ( .B(n107), .A(di_tst), .Y(n150) );
  NOR21XL U1014 ( .B(r_lt_gpi[2]), .A(n87), .Y(lt_gpi[2]) );
  NOR21XL U1015 ( .B(r_lt_gpi[3]), .A(n87), .Y(lt_gpi[3]) );
  NOR21XL U1016 ( .B(r_lt_gpi[1]), .A(n87), .Y(lt_gpi[1]) );
  OR2X1 U1017 ( .A(r_gpio_ie[0]), .B(n107), .Y(GPIO_IE[0]) );
  NOR3XL U1018 ( .A(r_lt_gpi[2]), .B(r_lt_gpi[3]), .C(r_lt_gpi[1]), .Y(
        sll_232_2_A_0_) );
  NAND2X1 U1019 ( .A(r_lt_gpi[0]), .B(sll_232_2_A_0_), .Y(n665) );
  NAND2X1 U1020 ( .A(r_lt_gpi[0]), .B(N593), .Y(n655) );
  NAND2X1 U1021 ( .A(r_lt_gpi[1]), .B(sll_232_2_A_0_), .Y(n666) );
  NAND2X1 U1022 ( .A(r_lt_gpi[1]), .B(N593), .Y(n656) );
  INVX1 U1023 ( .A(r_lt_gpi[3]), .Y(n645) );
  INVX1 U1024 ( .A(r_lt_gpi[2]), .Y(n652) );
  NAND2X1 U1025 ( .A(r_lt_gpi[2]), .B(r_lt_gpi[3]), .Y(n667) );
  NAND2X1 U1026 ( .A(r_lt_gpi[2]), .B(r_lt_gpi[3]), .Y(n657) );
  NAND2X1 U1027 ( .A(r_lt_gpi[2]), .B(n645), .Y(n671) );
  NAND2X1 U1028 ( .A(r_lt_gpi[2]), .B(n645), .Y(n661) );
  OR2X1 U1029 ( .A(r_gpio_ie[1]), .B(n107), .Y(GPIO_IE[1]) );
  NAND2X1 U1030 ( .A(r_lt_gpi[3]), .B(n652), .Y(n673) );
  NAND2X1 U1031 ( .A(r_lt_gpi[3]), .B(n652), .Y(n663) );
  INVX1 U1032 ( .A(r_lt_gpi[0]), .Y(n653) );
  NAND2X1 U1033 ( .A(di_tst), .B(n654), .Y(n302) );
  INVX1 U1034 ( .A(i_rstz), .Y(n654) );
  INVX1 U1035 ( .A(x_clk), .Y(n452) );
  AOI22XL U1036 ( .A(xram_a[6]), .B(xram_ce), .C(iram_a[6]), .D(iram_ce), .Y(
        n240) );
  AO22XL U1037 ( .A(xram_a[4]), .B(xram_ce), .C(iram_a[4]), .D(iram_ce), .Y(
        SRAM_A[4]) );
  AOI22XL U1038 ( .A(xram_a[0]), .B(xram_ce), .C(iram_a[0]), .D(iram_ce), .Y(
        n244) );
  AOI22XL U1039 ( .A(xram_a[1]), .B(xram_ce), .C(iram_a[1]), .D(iram_ce), .Y(
        n243) );
  AOI22XL U1040 ( .A(n16), .B(xram_ce), .C(iram_a[3]), .D(iram_ce), .Y(n241)
         );
  NOR43X2 U1041 ( .B(n465), .C(n463), .D(n464), .A(n462), .Y(n469) );
  NOR21X2 U1042 ( .B(n469), .A(n470), .Y(n468) );
endmodule


module SNPS_CLOCK_GATE_HIGH_core_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_1 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we;
  output pwm_o;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         net8871, n5, n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [6:0] pwmcnt;

  glreg_a0_1 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8871), .TE(1'b0) );
  DFFSQX1 pwmcnt_reg_0_ ( .D(N14), .C(net8871), .XS(n1), .Q(pwmcnt[0]) );
  DFFSQX1 pwmcnt_reg_4_ ( .D(N18), .C(net8871), .XS(n2), .Q(pwmcnt[4]) );
  DFFSQX1 pwmcnt_reg_6_ ( .D(N20), .C(net8871), .XS(n2), .Q(pwmcnt[6]) );
  DFFSQX1 pwmcnt_reg_5_ ( .D(N19), .C(net8871), .XS(n2), .Q(pwmcnt[5]) );
  DFFSQX1 pwmcnt_reg_1_ ( .D(N15), .C(net8871), .XS(n1), .Q(pwmcnt[1]) );
  DFFSQX1 pwmcnt_reg_2_ ( .D(N16), .C(net8871), .XS(n2), .Q(pwmcnt[2]) );
  DFFSQX1 pwmcnt_reg_3_ ( .D(N17), .C(net8871), .XS(n2), .Q(pwmcnt[3]) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  INVX1 U6 ( .A(n12), .Y(n25) );
  INVX1 U7 ( .A(n19), .Y(n26) );
  NAND21X1 U8 ( .B(wdat[7]), .A(we), .Y(n5) );
  INVX1 U9 ( .A(pwmcnt[1]), .Y(n22) );
  INVX1 U10 ( .A(r_pwm[3]), .Y(n24) );
  INVX1 U11 ( .A(r_pwm[2]), .Y(n23) );
  INVX1 U12 ( .A(pwmcnt[5]), .Y(n21) );
  INVX1 U13 ( .A(pwmcnt[6]), .Y(n20) );
  NAND21X1 U14 ( .B(r_pwm[7]), .A(n5), .Y(N13) );
  OAI21BBX1 U15 ( .A(N12), .B(r_pwm[7]), .C(n5), .Y(N20) );
  OAI21BBX1 U16 ( .A(N11), .B(r_pwm[7]), .C(n5), .Y(N19) );
  OAI21BBX1 U17 ( .A(N6), .B(r_pwm[7]), .C(n5), .Y(N14) );
  OAI21BBX1 U18 ( .A(N10), .B(r_pwm[7]), .C(n5), .Y(N18) );
  OAI21BBX1 U19 ( .A(N9), .B(r_pwm[7]), .C(n5), .Y(N17) );
  OAI21BBX1 U20 ( .A(N8), .B(r_pwm[7]), .C(n5), .Y(N16) );
  OAI21BBX1 U21 ( .A(N7), .B(r_pwm[7]), .C(n5), .Y(N15) );
  INVX1 U22 ( .A(pwmcnt[0]), .Y(N6) );
  OR2X1 U23 ( .A(pwmcnt[1]), .B(pwmcnt[0]), .Y(n4) );
  OAI21BBX1 U24 ( .A(pwmcnt[0]), .B(pwmcnt[1]), .C(n4), .Y(N7) );
  OR2X1 U25 ( .A(n4), .B(pwmcnt[2]), .Y(n6) );
  OAI21BBX1 U26 ( .A(n4), .B(pwmcnt[2]), .C(n6), .Y(N8) );
  OR2X1 U27 ( .A(n6), .B(pwmcnt[3]), .Y(n7) );
  OAI21BBX1 U28 ( .A(n6), .B(pwmcnt[3]), .C(n7), .Y(N9) );
  OR2X1 U29 ( .A(n7), .B(pwmcnt[4]), .Y(n8) );
  OAI21BBX1 U30 ( .A(n7), .B(pwmcnt[4]), .C(n8), .Y(N10) );
  XNOR2XL U31 ( .A(n8), .B(pwmcnt[5]), .Y(N11) );
  OR2X1 U32 ( .A(pwmcnt[5]), .B(n8), .Y(n9) );
  XNOR2XL U33 ( .A(pwmcnt[6]), .B(n9), .Y(N12) );
  NOR2X1 U34 ( .A(n20), .B(r_pwm[6]), .Y(n19) );
  OR2X1 U35 ( .A(r_pwm[5]), .B(n21), .Y(n11) );
  NOR32XL U36 ( .B(r_pwm[4]), .C(n11), .A(pwmcnt[4]), .Y(n10) );
  AOI221XL U37 ( .A(r_pwm[6]), .B(n20), .C(r_pwm[5]), .D(n21), .E(n10), .Y(n18) );
  OAI2B11X1 U38 ( .D(pwmcnt[4]), .C(r_pwm[4]), .A(n11), .B(n26), .Y(n17) );
  AND2X1 U39 ( .A(pwmcnt[3]), .B(n24), .Y(n15) );
  OAI32X1 U40 ( .A(n23), .B(pwmcnt[2]), .C(n15), .D(pwmcnt[3]), .E(n24), .Y(
        n12) );
  AOI21BBXL U41 ( .B(n22), .C(r_pwm[1]), .A(pwmcnt[0]), .Y(n13) );
  AOI221XL U42 ( .A(r_pwm[1]), .B(n22), .C(n13), .D(r_pwm[0]), .E(n12), .Y(n14) );
  GEN2XL U43 ( .D(pwmcnt[2]), .E(n23), .C(n15), .B(n25), .A(n14), .Y(n16) );
  OAI22X1 U44 ( .A(n19), .B(n18), .C(n17), .D(n16), .Y(pwm_o) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_1 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net8889;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8889), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net8889), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net8889), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net8889), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net8889), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net8889), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net8889), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net8889), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net8889), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_0 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we;
  output pwm_o;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         net8907, n5, n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [6:0] pwmcnt;

  glreg_a0_0 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8907), .TE(1'b0) );
  DFFSQX1 pwmcnt_reg_6_ ( .D(N20), .C(net8907), .XS(n2), .Q(pwmcnt[6]) );
  DFFSQX1 pwmcnt_reg_2_ ( .D(N16), .C(net8907), .XS(n2), .Q(pwmcnt[2]) );
  DFFSQX1 pwmcnt_reg_0_ ( .D(N14), .C(net8907), .XS(n1), .Q(pwmcnt[0]) );
  DFFSQX1 pwmcnt_reg_4_ ( .D(N18), .C(net8907), .XS(n2), .Q(pwmcnt[4]) );
  DFFSQX1 pwmcnt_reg_5_ ( .D(N19), .C(net8907), .XS(n2), .Q(pwmcnt[5]) );
  DFFSQX1 pwmcnt_reg_1_ ( .D(N15), .C(net8907), .XS(n1), .Q(pwmcnt[1]) );
  DFFSQX1 pwmcnt_reg_3_ ( .D(N17), .C(net8907), .XS(n2), .Q(pwmcnt[3]) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  INVX1 U6 ( .A(n12), .Y(n25) );
  INVX1 U7 ( .A(n19), .Y(n26) );
  NAND21X1 U8 ( .B(wdat[7]), .A(we), .Y(n5) );
  INVX1 U9 ( .A(pwmcnt[1]), .Y(n22) );
  INVX1 U10 ( .A(r_pwm[3]), .Y(n24) );
  INVX1 U11 ( .A(pwmcnt[5]), .Y(n21) );
  INVX1 U12 ( .A(r_pwm[2]), .Y(n23) );
  INVX1 U13 ( .A(pwmcnt[6]), .Y(n20) );
  NAND21X1 U14 ( .B(r_pwm[7]), .A(n5), .Y(N13) );
  OAI21BBX1 U15 ( .A(N12), .B(r_pwm[7]), .C(n5), .Y(N20) );
  OAI21BBX1 U16 ( .A(N11), .B(r_pwm[7]), .C(n5), .Y(N19) );
  OAI21BBX1 U17 ( .A(N6), .B(r_pwm[7]), .C(n5), .Y(N14) );
  OAI21BBX1 U18 ( .A(N10), .B(r_pwm[7]), .C(n5), .Y(N18) );
  OAI21BBX1 U19 ( .A(N9), .B(r_pwm[7]), .C(n5), .Y(N17) );
  OAI21BBX1 U20 ( .A(N8), .B(r_pwm[7]), .C(n5), .Y(N16) );
  OAI21BBX1 U21 ( .A(N7), .B(r_pwm[7]), .C(n5), .Y(N15) );
  INVX1 U22 ( .A(pwmcnt[0]), .Y(N6) );
  OR2X1 U23 ( .A(pwmcnt[1]), .B(pwmcnt[0]), .Y(n4) );
  OAI21BBX1 U24 ( .A(pwmcnt[0]), .B(pwmcnt[1]), .C(n4), .Y(N7) );
  OR2X1 U25 ( .A(n4), .B(pwmcnt[2]), .Y(n6) );
  OAI21BBX1 U26 ( .A(n4), .B(pwmcnt[2]), .C(n6), .Y(N8) );
  OR2X1 U27 ( .A(n6), .B(pwmcnt[3]), .Y(n7) );
  OAI21BBX1 U28 ( .A(n6), .B(pwmcnt[3]), .C(n7), .Y(N9) );
  OR2X1 U29 ( .A(n7), .B(pwmcnt[4]), .Y(n8) );
  OAI21BBX1 U30 ( .A(n7), .B(pwmcnt[4]), .C(n8), .Y(N10) );
  XNOR2XL U31 ( .A(n8), .B(pwmcnt[5]), .Y(N11) );
  OR2X1 U32 ( .A(pwmcnt[5]), .B(n8), .Y(n9) );
  XNOR2XL U33 ( .A(pwmcnt[6]), .B(n9), .Y(N12) );
  NOR2X1 U34 ( .A(n20), .B(r_pwm[6]), .Y(n19) );
  OR2X1 U35 ( .A(r_pwm[5]), .B(n21), .Y(n11) );
  NOR32XL U36 ( .B(r_pwm[4]), .C(n11), .A(pwmcnt[4]), .Y(n10) );
  AOI221XL U37 ( .A(r_pwm[6]), .B(n20), .C(r_pwm[5]), .D(n21), .E(n10), .Y(n18) );
  OAI2B11X1 U38 ( .D(pwmcnt[4]), .C(r_pwm[4]), .A(n11), .B(n26), .Y(n17) );
  AND2X1 U39 ( .A(pwmcnt[3]), .B(n24), .Y(n15) );
  OAI32X1 U40 ( .A(n23), .B(pwmcnt[2]), .C(n15), .D(pwmcnt[3]), .E(n24), .Y(
        n12) );
  AOI21BBXL U41 ( .B(n22), .C(r_pwm[1]), .A(pwmcnt[0]), .Y(n13) );
  AOI221XL U42 ( .A(r_pwm[1]), .B(n22), .C(n13), .D(r_pwm[0]), .E(n12), .Y(n14) );
  GEN2XL U43 ( .D(pwmcnt[2]), .E(n23), .C(n15), .B(n25), .A(n14), .Y(n16) );
  OAI22X1 U44 ( .A(n19), .B(n18), .C(n17), .D(n16), .Y(pwm_o) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_0 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net8925;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8925), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net8925), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net8925), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net8925), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net8925), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net8925), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net8925), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net8925), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net8925), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module divclk_a0 ( mclk, srstz, atpg_en, clk_1p0m, clk_500k, clk_100k, clk_50k, 
        clk_500, divff_o1, divff_o2 );
  input mclk, srstz, atpg_en;
  output clk_1p0m, clk_500k, clk_100k, clk_50k, clk_500, divff_o1, divff_o2;
  wire   div500k_5_2_, div500k_5_0, div1p0m_2, div100k_2, N23, N24, N25, N26,
         N37, N38, N39, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n1, n2, n3, n4, n5, n6, n7, n25, n26,
         n27;
  wire   [2:0] div12;
  wire   [6:0] div50k_100;

  CLKDLX1 U0_D1P0M_ICG ( .CK(mclk), .E(n22), .SE(atpg_en), .ECK(clk_1p0m) );
  CLKDLX1 U0_D500K_ICG ( .CK(clk_1p0m), .E(div1p0m_2), .SE(atpg_en), .ECK(
        clk_500k) );
  CLKDLX1 U0_D100K_ICG ( .CK(clk_500k), .E(n23), .SE(atpg_en), .ECK(clk_100k)
         );
  CLKDLX1 U0_D50K_ICG ( .CK(clk_100k), .E(div100k_2), .SE(atpg_en), .ECK(
        clk_50k) );
  CLKDLX1 U0_D0P5K_ICG ( .CK(clk_50k), .E(n24), .SE(atpg_en), .ECK(clk_500) );
  divclk_a0_DW01_inc_0 add_60 ( .A(div50k_100), .SUM({N52, N51, N50, N49, N48, 
        N47, N46}) );
  DFFRQX1 div1p0m_2_reg ( .D(n6), .C(clk_1p0m), .XR(n1), .Q(div1p0m_2) );
  DFFRQX1 div100k_2_reg ( .D(n27), .C(clk_100k), .XR(n1), .Q(div100k_2) );
  DFFRQX1 div50k_100_reg_6_ ( .D(N59), .C(clk_50k), .XR(n2), .Q(div50k_100[6])
         );
  DFFRQX1 div50k_100_reg_5_ ( .D(N58), .C(clk_50k), .XR(n2), .Q(div50k_100[5])
         );
  DFFRQX1 div50k_100_reg_4_ ( .D(N57), .C(clk_50k), .XR(n2), .Q(div50k_100[4])
         );
  DFFRQX1 div50k_100_reg_1_ ( .D(N54), .C(clk_50k), .XR(n2), .Q(div50k_100[1])
         );
  DFFRQX1 div50k_100_reg_0_ ( .D(N53), .C(clk_50k), .XR(n1), .Q(div50k_100[0])
         );
  DFFRQX1 div50k_100_reg_3_ ( .D(N56), .C(clk_50k), .XR(n2), .Q(div50k_100[3])
         );
  DFFRQX1 div50k_100_reg_2_ ( .D(N55), .C(clk_50k), .XR(n2), .Q(div50k_100[2])
         );
  DFFRQX1 div500k_5_reg_2_ ( .D(N39), .C(clk_500k), .XR(n1), .Q(div500k_5_2_)
         );
  DFFRQX1 div500k_5_reg_1_ ( .D(N38), .C(clk_500k), .XR(n1), .Q(divff_o2) );
  DFFRQX1 div500k_5_reg_0_ ( .D(N37), .C(clk_500k), .XR(n1), .Q(div500k_5_0)
         );
  DFFRQX1 div12_reg_0_ ( .D(N23), .C(mclk), .XR(n1), .Q(div12[0]) );
  DFFRQX1 div12_reg_2_ ( .D(N25), .C(mclk), .XR(n1), .Q(div12[2]) );
  DFFRQX1 div12_reg_1_ ( .D(N24), .C(mclk), .XR(n1), .Q(div12[1]) );
  DFFRQX1 div12_reg_3_ ( .D(N26), .C(mclk), .XR(n1), .Q(divff_o1) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(srstz), .Y(n3) );
  NOR21XL U6 ( .B(n18), .A(n19), .Y(n14) );
  XNOR2XL U7 ( .A(n15), .B(n14), .Y(n12) );
  XNOR2XL U8 ( .A(n10), .B(n12), .Y(N25) );
  NOR2X1 U9 ( .A(n11), .B(n16), .Y(N24) );
  XOR2X1 U10 ( .A(n12), .B(n17), .Y(n16) );
  XNOR2XL U11 ( .A(n18), .B(n19), .Y(n17) );
  NOR21XL U12 ( .B(n10), .A(n11), .Y(N26) );
  NOR21XL U13 ( .B(N51), .A(n24), .Y(N58) );
  NOR21XL U14 ( .B(N50), .A(n24), .Y(N57) );
  NOR21XL U15 ( .B(N49), .A(n24), .Y(N56) );
  NOR21XL U16 ( .B(N48), .A(n24), .Y(N55) );
  NOR21XL U17 ( .B(N47), .A(n24), .Y(N54) );
  XNOR2XL U18 ( .A(divff_o1), .B(n5), .Y(n15) );
  XNOR2XL U19 ( .A(n15), .B(div12[1]), .Y(n19) );
  XNOR2XL U20 ( .A(n13), .B(divff_o1), .Y(n10) );
  NAND2X1 U21 ( .A(n14), .B(n15), .Y(n13) );
  XNOR2XL U22 ( .A(n20), .B(n15), .Y(n18) );
  XNOR2XL U23 ( .A(div12[1]), .B(div12[0]), .Y(n20) );
  INVX1 U24 ( .A(div12[2]), .Y(n5) );
  NOR21XL U25 ( .B(N52), .A(n24), .Y(N59) );
  NOR21XL U26 ( .B(N46), .A(n24), .Y(N53) );
  XNOR2XL U27 ( .A(n21), .B(n4), .Y(N23) );
  XNOR2XL U28 ( .A(divff_o1), .B(div12[2]), .Y(n21) );
  OAI32X1 U29 ( .A(n25), .B(div500k_5_2_), .C(n7), .D(n9), .E(n26), .Y(N39) );
  INVX1 U30 ( .A(div500k_5_0), .Y(n7) );
  AOI21BBXL U31 ( .B(n23), .C(divff_o2), .A(N37), .Y(n9) );
  NOR3XL U32 ( .A(div500k_5_0), .B(divff_o2), .C(n26), .Y(n23) );
  NOR2X1 U33 ( .A(n23), .B(div500k_5_0), .Y(N37) );
  AND4X1 U34 ( .A(div50k_100[5]), .B(div50k_100[1]), .C(div50k_100[6]), .D(n8), 
        .Y(n24) );
  NOR41XL U35 ( .D(div50k_100[0]), .A(div50k_100[4]), .B(div50k_100[3]), .C(
        div50k_100[2]), .Y(n8) );
  NOR4XL U36 ( .A(div12[0]), .B(N23), .C(n4), .D(n5), .Y(n22) );
  INVX1 U37 ( .A(div12[1]), .Y(n4) );
  INVX1 U38 ( .A(div500k_5_2_), .Y(n26) );
  NOR42XL U39 ( .C(divff_o1), .D(div12[2]), .A(n4), .B(div12[0]), .Y(n11) );
  XNOR2XL U40 ( .A(n25), .B(div500k_5_0), .Y(N38) );
  INVX1 U41 ( .A(divff_o2), .Y(n25) );
  INVX1 U42 ( .A(div100k_2), .Y(n27) );
  INVX1 U43 ( .A(div1p0m_2), .Y(n6) );
endmodule


module divclk_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module srambist_a0 ( clk, srstz, reg_hit, reg_w, reg_r, reg_wdat, iram_rdat, 
        xram_rdat, bist_en, bist_xram, bist_wr, bist_adr, bist_wdat, o_bistctl, 
        o_bistdat );
  input [1:0] reg_hit;
  input [7:0] reg_wdat;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  output [10:0] bist_adr;
  output [7:0] bist_wdat;
  output [6:0] o_bistctl;
  output [7:0] o_bistdat;
  input clk, srstz, reg_w, reg_r;
  output bist_en, bist_xram, bist_wr;
  wire   we_1_, bistctl_re, N21, busy_dly, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, r_bistfault, upd_fault, wd_fault, net8943, n30, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n83, n84, n85,
         n86, n87, n88, n89, n90, n92, n94, n105, n106, n107, n108, n109, n110,
         n111, n3, n4, n5, n6, n7, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33,
         n34, n75, n76, n77, n78, n79, n80, n81, n82, n91, n93, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129;
  wire   [1:0] rw_sta;

  glreg_WIDTH1_0 u0_bistfault ( .clk(clk), .arstz(n11), .we(upd_fault), .wdat(
        wd_fault), .rdat(o_bistctl[3]) );
  glreg_WIDTH5_1 u0_bistctl ( .clk(clk), .arstz(n11), .we(n30), .wdat({
        reg_wdat[6:4], reg_wdat[2:1]}), .rdat({o_bistctl[6:4], o_bistctl[2:1]}) );
  glreg_a0_6 u0_bistdat ( .clk(clk), .arstz(n10), .we(we_1_), .wdat(reg_wdat), 
        .rdat(o_bistdat) );
  SNPS_CLOCK_GATE_HIGH_srambist_a0 clk_gate_adr_reg ( .CLK(clk), .EN(N86), 
        .ENCLK(net8943), .TE(1'b0) );
  srambist_a0_DW01_inc_0 add_65 ( .A(bist_adr), .SUM({N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64}) );
  DFFQX1 busy_dly_reg ( .D(o_bistctl[0]), .C(clk), .Q(busy_dly) );
  DFFQX1 r_bistfault_reg ( .D(n110), .C(clk), .Q(r_bistfault) );
  DFFRQX1 bistctl_re_reg ( .D(N21), .C(clk), .XR(n11), .Q(bistctl_re) );
  DFFQX1 rw_sta_reg_1_ ( .D(n121), .C(clk), .Q(rw_sta[1]) );
  DFFQX1 rw_sta_reg_0_ ( .D(n111), .C(clk), .Q(rw_sta[0]) );
  DFFQX1 adr_reg_9_ ( .D(N96), .C(net8943), .Q(bist_adr[9]) );
  DFFQX1 adr_reg_8_ ( .D(N95), .C(net8943), .Q(bist_adr[8]) );
  DFFQX1 adr_reg_10_ ( .D(N97), .C(net8943), .Q(bist_adr[10]) );
  DFFQX1 adr_reg_5_ ( .D(N92), .C(net8943), .Q(bist_adr[5]) );
  DFFQX1 adr_reg_4_ ( .D(N91), .C(net8943), .Q(bist_adr[4]) );
  DFFQX1 adr_reg_3_ ( .D(N90), .C(net8943), .Q(bist_adr[3]) );
  DFFQX1 adr_reg_6_ ( .D(N93), .C(net8943), .Q(bist_adr[6]) );
  DFFQX1 adr_reg_7_ ( .D(N94), .C(net8943), .Q(bist_adr[7]) );
  DFFQX1 adr_reg_2_ ( .D(N89), .C(net8943), .Q(bist_adr[2]) );
  DFFQX1 adr_reg_1_ ( .D(N88), .C(net8943), .Q(bist_adr[1]) );
  DFFQX1 adr_reg_0_ ( .D(N87), .C(net8943), .Q(bist_adr[0]) );
  INVX1 U3 ( .A(1'b1), .Y(bist_xram) );
  NOR21XL U5 ( .B(bist_adr[5]), .A(n91), .Y(n96) );
  NAND21X1 U6 ( .B(n98), .A(n97), .Y(n99) );
  OR2X1 U7 ( .A(n107), .B(n106), .Y(n3) );
  INVXL U8 ( .A(n3), .Y(n4) );
  INVXL U9 ( .A(n3), .Y(n5) );
  BUFXL U10 ( .A(o_bistctl[0]), .Y(bist_en) );
  OAI21BBXL U11 ( .A(n93), .B(n16), .C(n5), .Y(n14) );
  NAND21XL U12 ( .B(n51), .A(o_bistctl[0]), .Y(n101) );
  OAI21BBXL U13 ( .A(n6), .B(o_bistctl[0]), .C(n10), .Y(n100) );
  NAND21XL U14 ( .B(n13), .A(bist_adr[1]), .Y(n93) );
  OAI21BBXL U15 ( .A(n4), .B(n13), .C(n7), .Y(N87) );
  NAND21XL U16 ( .B(bist_adr[9]), .A(n98), .Y(n102) );
  INVX1 U17 ( .A(n12), .Y(n11) );
  INVX1 U18 ( .A(n12), .Y(n10) );
  INVX1 U19 ( .A(srstz), .Y(n12) );
  INVX1 U20 ( .A(n108), .Y(n30) );
  NAND21X1 U21 ( .B(n94), .A(n11), .Y(n75) );
  NAND2X1 U22 ( .A(reg_hit[0]), .B(reg_w), .Y(n108) );
  INVX1 U23 ( .A(n82), .Y(n81) );
  INVX1 U24 ( .A(n86), .Y(n114) );
  AND2X1 U25 ( .A(reg_w), .B(reg_hit[1]), .Y(we_1_) );
  XNOR2XL U26 ( .A(bist_wdat[4]), .B(n128), .Y(n44) );
  INVX1 U27 ( .A(n101), .Y(bist_wr) );
  INVX1 U28 ( .A(n57), .Y(n117) );
  INVX1 U29 ( .A(n79), .Y(n98) );
  INVX1 U30 ( .A(n32), .Y(n31) );
  INVX1 U31 ( .A(n76), .Y(n34) );
  INVX1 U32 ( .A(n19), .Y(n18) );
  INVX1 U33 ( .A(n22), .Y(n21) );
  INVX1 U34 ( .A(n25), .Y(n24) );
  INVX1 U35 ( .A(n28), .Y(n27) );
  NAND21X1 U36 ( .B(n107), .A(n106), .Y(n82) );
  NAND21X1 U37 ( .B(n89), .A(n103), .Y(n84) );
  OAI22X1 U38 ( .A(n103), .B(n86), .C(n114), .D(n84), .Y(bist_wdat[4]) );
  OAI2B11X1 U39 ( .D(N65), .C(n82), .A(n15), .B(n14), .Y(N88) );
  INVX1 U40 ( .A(n75), .Y(n15) );
  NAND2X1 U41 ( .A(n115), .B(n83), .Y(n86) );
  NAND2X1 U42 ( .A(n87), .B(n84), .Y(bist_wdat[0]) );
  NOR2X1 U43 ( .A(n105), .B(n106), .Y(n94) );
  INVX1 U44 ( .A(n85), .Y(n115) );
  AND2X1 U45 ( .A(reg_r), .B(reg_hit[0]), .Y(N21) );
  NAND3X1 U46 ( .A(n105), .B(n11), .C(n107), .Y(N86) );
  XNOR2XL U47 ( .A(n103), .B(n90), .Y(bist_wdat[1]) );
  AOI21X1 U48 ( .B(n86), .C(n115), .A(n89), .Y(n90) );
  XNOR2XL U49 ( .A(n103), .B(n88), .Y(bist_wdat[2]) );
  AOI21X1 U50 ( .B(n86), .C(n83), .A(n89), .Y(n88) );
  OAI221X1 U51 ( .A(n84), .B(n86), .C(n114), .D(n103), .E(n87), .Y(
        bist_wdat[3]) );
  OAI22X1 U52 ( .A(n84), .B(n115), .C(n85), .D(n103), .Y(bist_wdat[5]) );
  XOR2X1 U53 ( .A(bist_wdat[2]), .B(iram_rdat[2]), .Y(n48) );
  XNOR2XL U54 ( .A(n56), .B(n128), .Y(n55) );
  OAI22X1 U55 ( .A(n104), .B(n57), .C(n117), .D(n112), .Y(n56) );
  INVX1 U56 ( .A(iram_rdat[0]), .Y(n129) );
  INVX1 U57 ( .A(iram_rdat[4]), .Y(n128) );
  INVX1 U58 ( .A(iram_rdat[6]), .Y(n126) );
  INVX1 U59 ( .A(iram_rdat[5]), .Y(n127) );
  NOR4XL U60 ( .A(n41), .B(n42), .C(n43), .D(n44), .Y(n39) );
  XNOR2XL U61 ( .A(bist_wdat[0]), .B(n129), .Y(n41) );
  XNOR2XL U62 ( .A(bist_wdat[6]), .B(n126), .Y(n42) );
  XOR2X1 U63 ( .A(bist_wdat[3]), .B(iram_rdat[3]), .Y(n43) );
  NOR4XL U64 ( .A(n45), .B(n46), .C(n47), .D(n48), .Y(n38) );
  XNOR2XL U65 ( .A(bist_wdat[5]), .B(n127), .Y(n45) );
  XOR2X1 U66 ( .A(bist_wdat[1]), .B(iram_rdat[1]), .Y(n47) );
  XNOR2XL U67 ( .A(n103), .B(iram_rdat[7]), .Y(n46) );
  NOR4XL U68 ( .A(n65), .B(n66), .C(n67), .D(n68), .Y(n49) );
  XNOR2XL U69 ( .A(n73), .B(n127), .Y(n65) );
  XNOR2XL U70 ( .A(n104), .B(iram_rdat[7]), .Y(n66) );
  XNOR2XL U71 ( .A(n71), .B(n72), .Y(n67) );
  NOR4XL U72 ( .A(n52), .B(n53), .C(n54), .D(n55), .Y(n50) );
  XNOR2XL U73 ( .A(n63), .B(n129), .Y(n52) );
  XNOR2XL U74 ( .A(n61), .B(n126), .Y(n53) );
  XNOR2XL U75 ( .A(iram_rdat[3]), .B(n58), .Y(n54) );
  NAND3X1 U76 ( .A(n123), .B(n124), .C(n11), .Y(n40) );
  OR2X1 U77 ( .A(n123), .B(n124), .Y(n6) );
  NAND2X1 U78 ( .A(n118), .B(n62), .Y(n57) );
  AOI21X1 U79 ( .B(n57), .C(n118), .A(n64), .Y(n71) );
  INVX1 U80 ( .A(n59), .Y(n112) );
  INVX1 U81 ( .A(n74), .Y(n118) );
  OAI22X1 U82 ( .A(n112), .B(n118), .C(n74), .D(n104), .Y(n73) );
  NAND2X1 U83 ( .A(n60), .B(n112), .Y(n63) );
  NAND3X1 U84 ( .A(bist_adr[9]), .B(bist_adr[10]), .C(n99), .Y(o_bistctl[0])
         );
  NAND21X1 U85 ( .B(bist_adr[1]), .A(n13), .Y(n16) );
  NAND21X1 U86 ( .B(bist_adr[6]), .A(n27), .Y(n32) );
  NAND21X1 U87 ( .B(bist_adr[7]), .A(n31), .Y(n76) );
  NAND21X1 U88 ( .B(bist_adr[8]), .A(n34), .Y(n79) );
  OR2X1 U89 ( .A(bist_adr[2]), .B(n16), .Y(n19) );
  NAND21X1 U90 ( .B(bist_adr[3]), .A(n18), .Y(n22) );
  NAND21X1 U91 ( .B(bist_adr[4]), .A(n21), .Y(n25) );
  NAND21X1 U92 ( .B(bist_adr[5]), .A(n24), .Y(n28) );
  INVX1 U93 ( .A(bist_adr[0]), .Y(n13) );
  NOR43XL U94 ( .B(bist_adr[3]), .C(bist_adr[4]), .D(bist_adr[2]), .A(n93), 
        .Y(n95) );
  NAND4X1 U95 ( .A(bist_adr[8]), .B(bist_adr[7]), .C(n96), .D(n95), .Y(n97) );
  INVX1 U96 ( .A(bist_adr[6]), .Y(n91) );
  NAND42X1 U97 ( .C(o_bistdat[6]), .D(n108), .A(reg_wdat[0]), .B(o_bistdat[7]), 
        .Y(n105) );
  AOI22AXL U98 ( .A(o_bistctl[1]), .B(n108), .D(n108), .C(reg_wdat[1]), .Y(
        n106) );
  AOI21X1 U99 ( .B(N64), .C(n81), .A(n75), .Y(n7) );
  AO21X1 U100 ( .B(N73), .C(n81), .A(n80), .Y(N96) );
  GEN2XL U101 ( .D(bist_adr[9]), .E(n79), .C(n78), .B(n4), .A(n12), .Y(n80) );
  INVX1 U102 ( .A(n102), .Y(n78) );
  AO21X1 U103 ( .B(N72), .C(n81), .A(n77), .Y(N95) );
  GEN2XL U104 ( .D(bist_adr[8]), .E(n76), .C(n98), .B(n5), .A(n75), .Y(n77) );
  AO21X1 U105 ( .B(N71), .C(n81), .A(n33), .Y(N94) );
  GEN2XL U106 ( .D(bist_adr[7]), .E(n32), .C(n34), .B(n4), .A(n75), .Y(n33) );
  AO21X1 U107 ( .B(N70), .C(n81), .A(n29), .Y(N93) );
  GEN2XL U108 ( .D(bist_adr[6]), .E(n28), .C(n31), .B(n5), .A(n75), .Y(n29) );
  AO21X1 U109 ( .B(N69), .C(n81), .A(n26), .Y(N92) );
  GEN2XL U110 ( .D(bist_adr[5]), .E(n25), .C(n27), .B(n4), .A(n75), .Y(n26) );
  AO21X1 U111 ( .B(N68), .C(n81), .A(n23), .Y(N91) );
  GEN2XL U112 ( .D(bist_adr[4]), .E(n22), .C(n24), .B(n5), .A(n75), .Y(n23) );
  AO21X1 U113 ( .B(N67), .C(n81), .A(n20), .Y(N90) );
  GEN2XL U114 ( .D(bist_adr[3]), .E(n19), .C(n21), .B(n4), .A(n75), .Y(n20) );
  AO21X1 U115 ( .B(N66), .C(n81), .A(n17), .Y(N89) );
  GEN2XL U116 ( .D(bist_adr[2]), .E(n16), .C(n18), .B(n5), .A(n75), .Y(n17) );
  INVX1 U117 ( .A(o_bistdat[5]), .Y(n103) );
  NOR2X1 U118 ( .A(n116), .B(o_bistdat[2]), .Y(n85) );
  NOR2X1 U119 ( .A(o_bistdat[3]), .B(o_bistdat[2]), .Y(n89) );
  NAND2X1 U120 ( .A(o_bistdat[2]), .B(n116), .Y(n83) );
  OAI2B11X1 U121 ( .D(N74), .C(n82), .A(n92), .B(srstz), .Y(N97) );
  AOI21X1 U122 ( .B(N63), .C(n4), .A(n94), .Y(n92) );
  NAND2X1 U123 ( .A(n109), .B(n105), .Y(n107) );
  OAI32X1 U124 ( .A(n124), .B(rw_sta[0]), .C(n120), .D(o_bistctl[2]), .E(n51), 
        .Y(n109) );
  INVX1 U125 ( .A(o_bistctl[2]), .Y(n120) );
  NAND2X1 U126 ( .A(o_bistdat[5]), .B(n89), .Y(n87) );
  INVX1 U127 ( .A(o_bistdat[3]), .Y(n116) );
  BUFX3 U128 ( .A(o_bistdat[5]), .Y(bist_wdat[7]) );
  ENOX1 U129 ( .A(n83), .B(n84), .C(n83), .D(o_bistdat[5]), .Y(bist_wdat[6])
         );
  XNOR2XL U130 ( .A(n69), .B(n70), .Y(n68) );
  AOI21X1 U131 ( .B(n57), .C(n62), .A(n64), .Y(n69) );
  XNOR2XL U132 ( .A(o_bistdat[4]), .B(iram_rdat[2]), .Y(n70) );
  XNOR2XL U133 ( .A(o_bistdat[4]), .B(iram_rdat[1]), .Y(n72) );
  OAI31XL U134 ( .A(n125), .B(bistctl_re), .C(n12), .D(n35), .Y(n110) );
  AOI33X1 U135 ( .A(busy_dly), .B(n37), .C(o_bistctl[2]), .D(n36), .E(n10), 
        .F(n122), .Y(n35) );
  AOI211X1 U136 ( .C(n38), .D(n39), .A(n40), .B(bistctl_re), .Y(n37) );
  AOI21X1 U137 ( .B(n49), .C(n50), .A(n51), .Y(n36) );
  MUX2BXL U138 ( .D0(rw_sta[0]), .D1(n40), .S(n100), .Y(n111) );
  NOR2X1 U139 ( .A(n119), .B(o_bistdat[0]), .Y(n74) );
  NOR2X1 U140 ( .A(n64), .B(o_bistdat[4]), .Y(n59) );
  NAND2X1 U141 ( .A(o_bistdat[4]), .B(n64), .Y(n60) );
  NOR2X1 U142 ( .A(o_bistdat[1]), .B(o_bistdat[0]), .Y(n64) );
  OAI32X1 U143 ( .A(n101), .B(n120), .C(n12), .D(n124), .E(n100), .Y(n121) );
  AOI221XL U144 ( .A(o_bistdat[4]), .B(n57), .C(n117), .D(n59), .E(n113), .Y(
        n58) );
  INVX1 U145 ( .A(n60), .Y(n113) );
  ENOX1 U146 ( .A(n62), .B(n112), .C(n62), .D(o_bistdat[4]), .Y(n61) );
  INVX1 U147 ( .A(rw_sta[1]), .Y(n124) );
  NAND2X1 U148 ( .A(o_bistdat[0]), .B(n119), .Y(n62) );
  INVX1 U149 ( .A(o_bistdat[1]), .Y(n119) );
  NAND2X1 U150 ( .A(rw_sta[0]), .B(n124), .Y(n51) );
  INVX1 U151 ( .A(o_bistdat[4]), .Y(n104) );
  INVX1 U152 ( .A(rw_sta[0]), .Y(n123) );
  INVX1 U153 ( .A(bistctl_re), .Y(n122) );
  NOR2X1 U154 ( .A(bistctl_re), .B(n125), .Y(wd_fault) );
  NAND2X1 U155 ( .A(n125), .B(n122), .Y(upd_fault) );
  INVX1 U156 ( .A(r_bistfault), .Y(n125) );
  XNOR2XL U157 ( .A(bist_adr[10]), .B(n102), .Y(N63) );
endmodule


module srambist_a0_DW01_inc_0 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1XL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_srambist_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_6 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net8961;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8961), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net8961), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net8961), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net8961), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net8961), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net8961), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net8961), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net8961), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net8961), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_1 ( clk, arstz, we, wdat, rdat );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we;
  wire   net8979;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8979), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net8979), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net8979), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net8979), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net8979), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net8979), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_0 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module regx_a0 ( regx_r, regx_w, di_drposc, di_imposc, di_rd_det, clk_500k, 
        r_imp_osc, regx_addr, regx_wdat, regx_rdat, regx_hitbst, regx_wrpwm, 
        regx_wrcvc, r_sdischg, r_bistctl, r_bistdat, r_vcomp, r_idacsh, 
        r_cvofsx, r_pwm, regx_wrdac, dac_r_vs, dac_comp, r_dac_en, r_sar_en, 
        r_aopt, r_xtm, r_adummyi, r_bck0, r_bck1, r_bck2, r_i2crout, r_xana, 
        di_xanav, lt_gpi, di_tst, bkpt_pc, bkpt_ena, we_twlb, r_vpp_en, 
        r_vpp0v_en, r_otp_pwdn_en, r_otp_wpls, wd_twlb, r_sap, r_twlb, 
        upd_pwrv, ramacc, sse_idle, bus_idle, r_do_ts, r_dpdo_sel, r_dndo_sel, 
        di_ts, detclk, aswclk, atpg_en, di_aswk, clk, rrstz );
  input [6:0] regx_addr;
  input [7:0] regx_wdat;
  output [7:0] regx_rdat;
  output [1:0] regx_hitbst;
  output [1:0] regx_wrpwm;
  output [3:0] regx_wrcvc;
  input [7:0] r_sdischg;
  input [6:0] r_bistctl;
  input [7:0] r_bistdat;
  input [7:0] r_vcomp;
  input [7:0] r_idacsh;
  input [7:0] r_cvofsx;
  input [15:0] r_pwm;
  output [13:0] regx_wrdac;
  input [79:0] dac_r_vs;
  input [9:0] dac_comp;
  input [9:0] r_dac_en;
  input [9:0] r_sar_en;
  output [7:0] r_aopt;
  output [7:0] r_xtm;
  output [7:0] r_adummyi;
  output [7:0] r_bck0;
  output [7:0] r_bck1;
  output [7:0] r_bck2;
  output [5:0] r_i2crout;
  output [23:0] r_xana;
  input [5:0] di_xanav;
  input [3:0] lt_gpi;
  output [14:0] bkpt_pc;
  output [1:0] wd_twlb;
  output [1:0] r_sap;
  input [1:0] r_twlb;
  output [6:0] r_do_ts;
  output [3:0] r_dpdo_sel;
  output [3:0] r_dndo_sel;
  input [4:0] di_aswk;
  input regx_r, regx_w, di_drposc, di_imposc, di_rd_det, clk_500k, di_tst,
         upd_pwrv, ramacc, sse_idle, bus_idle, di_ts, detclk, aswclk, atpg_en,
         clk, rrstz;
  output r_imp_osc, bkpt_ena, we_twlb, r_vpp_en, r_vpp0v_en, r_otp_pwdn_en,
         r_otp_wpls;
  wire   n129, we_19, we_7, we_6, we_5, we_4, reg1B_3_, reg10_7_, lt_drp,
         i2c_mode_upd, N8, d_we16, lt_reg1C_0, net8997, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n66, n67, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151,
         SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153,
         SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155,
         SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157,
         SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159,
         SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161,
         SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163,
         SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165,
         SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167,
         SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169,
         SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171,
         SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173,
         SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175,
         SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177,
         SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179,
         SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181,
         SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183,
         SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185,
         SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187,
         SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189,
         SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191,
         SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193,
         SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195,
         SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197,
         SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199,
         SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201,
         SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203,
         SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205,
         SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207,
         SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209,
         SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211,
         SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213,
         SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215,
         SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217,
         SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219,
         SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221,
         SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223,
         SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225,
         SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227,
         SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229,
         SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231,
         SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233,
         SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235,
         SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237,
         SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239,
         SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241,
         SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243,
         SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245,
         SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247,
         SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249,
         SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251,
         SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253,
         SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255,
         SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257,
         SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259,
         SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261,
         SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263,
         SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265,
         SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267,
         SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269,
         SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271,
         SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273,
         SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275,
         SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277,
         SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279,
         SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281,
         SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283,
         SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285,
         SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287,
         SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289,
         SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291,
         SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293,
         SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295,
         SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297,
         SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299,
         SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301,
         SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303,
         SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305,
         SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307,
         SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309,
         SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311,
         SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313,
         SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315,
         SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317,
         SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319,
         SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321,
         SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323,
         SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325,
         SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327,
         SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329,
         SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331,
         SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333,
         SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335,
         SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337,
         SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339,
         SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341,
         SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343,
         SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345,
         SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347,
         SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349,
         SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351,
         SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353,
         SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355,
         SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357,
         SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359,
         SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361,
         SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363,
         SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365,
         SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367,
         SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369,
         SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371,
         SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373,
         SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375,
         SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377,
         SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379,
         SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381,
         SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383,
         SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385,
         SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387,
         SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389,
         SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391,
         SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393,
         SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395,
         SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397,
         SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399,
         SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401,
         SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403,
         SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405,
         SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407,
         SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409,
         SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411,
         SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413,
         SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415,
         SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417,
         SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419,
         SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421,
         SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423,
         SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425,
         SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427,
         SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429,
         SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431,
         SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433,
         SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435,
         SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437,
         SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439,
         SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441,
         SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443,
         SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445,
         SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447,
         SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449,
         SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451,
         SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453,
         SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455,
         SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457,
         SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459,
         SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461,
         SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463,
         SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465,
         SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467,
         SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469,
         SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471,
         SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473,
         SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475,
         SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477,
         SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479,
         SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481,
         SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483,
         SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485,
         SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487,
         SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489,
         SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491,
         SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493,
         SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495,
         SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497,
         SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499,
         SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501,
         SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503,
         SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505,
         SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507,
         SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509,
         SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511,
         SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513,
         SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515,
         SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517,
         SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519,
         SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521,
         SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523,
         SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525,
         SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527,
         SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529,
         SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531,
         SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533,
         SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535,
         SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537,
         SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539,
         SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541,
         SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543,
         SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545,
         SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547,
         SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549,
         SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551,
         SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553,
         SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555,
         SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557,
         SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559,
         SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561,
         SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563,
         SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565,
         SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567,
         SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569,
         SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571,
         SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573,
         SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575,
         SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577,
         SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579,
         SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581,
         SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583,
         SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585,
         SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587,
         SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589,
         SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591,
         SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593,
         SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595,
         SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597,
         SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599,
         SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601,
         SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603,
         SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605,
         SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607,
         SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609,
         SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611,
         SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613,
         SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615,
         SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617,
         SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619,
         SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621,
         SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623,
         SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625,
         SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627,
         SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629,
         SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631,
         SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633,
         SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635,
         SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637,
         SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639,
         SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641,
         SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643,
         SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645,
         SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647,
         SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649,
         SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651,
         SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653,
         SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655,
         SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657,
         SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659,
         SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661,
         SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663,
         SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665,
         SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667,
         SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669,
         SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671,
         SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673,
         SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675,
         SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677,
         SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679,
         SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681,
         SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683,
         SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685,
         SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687,
         SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689,
         SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691,
         SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693,
         SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695,
         SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697,
         SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699,
         SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701,
         SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703,
         SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705,
         SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707,
         SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709,
         SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711,
         SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713,
         SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715,
         SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717,
         SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719,
         SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721,
         SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723,
         SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725,
         SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727,
         SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729,
         SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731,
         SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733,
         SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735,
         SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737,
         SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739,
         SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741,
         SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743,
         SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745,
         SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747,
         SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749,
         SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751,
         SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753,
         SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755,
         SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757,
         SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759,
         SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761,
         SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763,
         SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765,
         SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767,
         SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769,
         SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771,
         SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773,
         SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775,
         SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777,
         SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779,
         SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781,
         SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783,
         SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785,
         SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787,
         SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789,
         SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791,
         SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793,
         SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795,
         SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797,
         SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799,
         SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801,
         SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803,
         SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805,
         SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807,
         SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809,
         SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811,
         SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813,
         SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815,
         SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817,
         SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819,
         SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821,
         SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823,
         SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825,
         SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827,
         SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829,
         SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831,
         SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833,
         SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835,
         SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837,
         SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839,
         SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841,
         SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843,
         SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845,
         SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847,
         SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849,
         SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851,
         SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853,
         SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855,
         SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857,
         SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859,
         SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861,
         SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863,
         SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865,
         SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867,
         SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869,
         SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871,
         SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873,
         SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875,
         SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877,
         SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879,
         SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881,
         SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883,
         SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885,
         SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887,
         SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889,
         SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891,
         SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893,
         SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895,
         SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897,
         SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899,
         SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901,
         SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903,
         SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905,
         SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907,
         SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909,
         SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911,
         SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913,
         SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915,
         SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917,
         SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919,
         SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921,
         SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923,
         SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925,
         SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927,
         SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929,
         SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931,
         SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933,
         SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935,
         SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937,
         SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939,
         SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941,
         SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943,
         SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945,
         SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947,
         SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949,
         SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951,
         SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953,
         SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955,
         SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957,
         SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959,
         SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961,
         SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963,
         SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965,
         SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967,
         SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969,
         SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971,
         SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973,
         SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975,
         SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977,
         SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979,
         SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981,
         SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983,
         SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985,
         SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987,
         SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989,
         SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991,
         SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993,
         SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995,
         SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997,
         SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999,
         SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001,
         SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003,
         SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005,
         SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007,
         SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009,
         SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011,
         SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013,
         SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015,
         SYNOPSYS_UNCONNECTED_1016;
  wire   [30:23] we;
  wire   [6:0] d_regx_addr;
  wire   [7:0] reg1F;
  wire   [3:2] reg1E;
  wire   [3:0] reg14;
  wire   [3:0] d_lt_gpi;
  wire   [5:0] lt_reg15_5_0;
  wire   [5:0] i2c_mode_wdat;
  wire   [5:0] d_lt_aswk;
  wire   [5:0] lt_aswk;
  wire   [7:0] wd18;

  glreg_a0_19 u0_reg04 ( .clk(clk), .arstz(n70), .we(we_4), .wdat({n17, n9, 
        n13, n5, n4, n19, n11, wd_twlb[0]}), .rdat(r_bck0) );
  glreg_a0_18 u0_reg05 ( .clk(clk), .arstz(n71), .we(we_5), .wdat({n16, n9, 
        n14, n6, n4, n20, regx_wdat[1], wd_twlb[0]}), .rdat(r_bck1) );
  glreg_a0_17 u0_reg06 ( .clk(clk), .arstz(n72), .we(we_6), .wdat({n17, 
        regx_wdat[6], n13, n5, n3, n20, n11, wd_twlb[0]}), .rdat(r_bck2) );
  glreg_a0_16 u0_reg07 ( .clk(clk), .arstz(n73), .we(we_7), .wdat({n16, n8, 
        n14, n6, n4, regx_wdat[2], n11, wd_twlb[0]}), .rdat(r_adummyi) );
  glreg_WIDTH1_2 u0_reg10 ( .clk(clk), .arstz(n91), .we(1'b1), .wdat(ramacc), 
        .rdat(reg10_7_) );
  glreg_6_00000002 u0_reg12 ( .clk(clk), .arstz(n84), .we(we_twlb), .wdat({n17, 
        n9, n14, n6, n4, n19}), .rdat({r_vpp_en, r_vpp0v_en, r_otp_pwdn_en, 
        r_otp_wpls, r_sap}) );
  glreg_a0_15 u0_reg13 ( .clk(clk), .arstz(n74), .we(we_19), .wdat({n17, n9, 
        n14, n6, n4, n20, n11, wd_twlb[0]}), .rdat({r_dpdo_sel, r_dndo_sel})
         );
  glreg_WIDTH6_1 u0_reg15 ( .clk(clk), .arstz(n86), .we(n21), .wdat({n13, n5, 
        n4, n20, wd_twlb[1], n96}), .rdat(lt_reg15_5_0) );
  glreg_WIDTH6_0 u1_reg15 ( .clk(clk), .arstz(n85), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat({n129, r_i2crout[4:0]}) );
  glreg_a0_14 u0_reg17 ( .clk(clk), .arstz(n75), .we(we[23]), .wdat({n17, 
        regx_wdat[6], n13, n5, n3, n19, regx_wdat[1], n96}), .rdat(r_aopt) );
  glreg_a0_13 u0_tmp18 ( .clk(clk), .arstz(n76), .we(we[24]), .wdat({n16, n8, 
        n13, n5, n4, n19, n11, n96}), .rdat(wd18) );
  glreg_a0_12 u0_reg18 ( .clk(clk), .arstz(n77), .we(we[25]), .wdat(wd18), 
        .rdat(bkpt_pc[7:0]) );
  glreg_a0_11 u0_reg19 ( .clk(clk), .arstz(n78), .we(we[25]), .wdat({n17, n9, 
        n14, n6, n4, n20, n11, n96}), .rdat({bkpt_ena, bkpt_pc[14:8]}) );
  glreg_a0_10 u0_reg1A ( .clk(clk), .arstz(n79), .we(we[26]), .wdat({n17, n9, 
        n13, n5, n4, n20, wd_twlb[1], n96}), .rdat(r_xtm) );
  dbnc_WIDTH2_TIMEOUT2_8 u0_ts_db ( .o_dbc(reg1B_3_), .o_chg(), .i_org(di_ts), 
        .clk(clk), .rstz(n89) );
  glreg_WIDTH7_0 u0_reg1B ( .clk(clk), .arstz(n83), .we(we[27]), .wdat({n17, 
        n9, n14, n6, n20, n11, n96}), .rdat(r_do_ts) );
  glreg_WIDTH1_1 u1_reg1C ( .clk(clk), .arstz(n91), .we(upd_pwrv), .wdat(
        lt_reg1C_0), .rdat(r_xana[0]) );
  glreg_a0_9 u0_reg1C ( .clk(clk), .arstz(n82), .we(we[28]), .wdat({n16, n8, 
        n14, n6, n3, n19, n11, n96}), .rdat({r_xana[7:1], lt_reg1C_0}) );
  glreg_a0_8 u0_reg1D ( .clk(clk), .arstz(n81), .we(we[29]), .wdat({n17, n9, 
        n14, n6, regx_wdat[3], n20, n11, wd_twlb[0]}), .rdat(r_xana[15:8]) );
  glreg_a0_7 u0_reg1E ( .clk(clk), .arstz(n80), .we(we[30]), .wdat({n17, n9, 
        n13, n5, n4, n20, wd_twlb}), .rdat({r_xana[23], r_imp_osc, 
        r_xana[21:20], reg1E, r_xana[17:16]}) );
  dbnc_WIDTH2_TIMEOUT2_7 u0_dosc_db ( .o_dbc(reg14[1]), .o_chg(), .i_org(
        di_imposc), .clk(clk), .rstz(n91) );
  dbnc_WIDTH2_TIMEOUT2_6 u0_iosc_db ( .o_dbc(reg14[2]), .o_chg(), .i_org(
        di_drposc), .clk(clk), .rstz(n91) );
  dbnc_WIDTH2_TIMEOUT2_5 u0_xana_db ( .o_dbc(reg1F[0]), .o_chg(), .i_org(
        di_xanav[0]), .clk(clk), .rstz(n90) );
  dbnc_WIDTH2_TIMEOUT2_4 u1_xana_db ( .o_dbc(reg1F[1]), .o_chg(), .i_org(
        di_xanav[1]), .clk(clk), .rstz(n90) );
  dbnc_WIDTH2_TIMEOUT2_3 u2_xana_db ( .o_dbc(reg1F[2]), .o_chg(), .i_org(
        di_xanav[2]), .clk(clk), .rstz(n88) );
  dbnc_WIDTH2_TIMEOUT2_2 u3_xana_db ( .o_dbc(reg1F[3]), .o_chg(), .i_org(
        di_xanav[3]), .clk(clk), .rstz(n89) );
  dbnc_WIDTH2_TIMEOUT2_1 u4_xana_db ( .o_dbc(reg1F[4]), .o_chg(), .i_org(
        di_xanav[4]), .clk(clk), .rstz(n86) );
  dbnc_WIDTH2_TIMEOUT2_0 u5_xana_db ( .o_dbc(reg1F[5]), .o_chg(), .i_org(
        di_xanav[5]), .clk(clk), .rstz(n84) );
  dbnc_a0_1 u6_xana_db ( .o_dbc(reg1F[6]), .o_chg(), .i_org(di_xanav[0]), 
        .clk(clk_500k), .rstz(n87) );
  dbnc_a0_0 u0_rdet_db ( .o_dbc(reg1F[7]), .o_chg(), .i_org(di_rd_det), .clk(
        clk_500k), .rstz(n88) );
  SNPS_CLOCK_GATE_HIGH_regx_a0 clk_gate_d_lt_gpi_reg ( .CLK(clk), .EN(n94), 
        .ENCLK(net8997), .TE(1'b0) );
  regx_a0_DW_rightsh_0 srl_66 ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        dac_comp[9:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_sar_en[9:8], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_dac_en[9:8], 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_comp[7:0], r_sar_en[7:0], r_dac_en[7:0], dac_r_vs[63:0], 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_r_vs[79:64], reg1F, r_xana[23], r_imp_osc, r_xana[21:20], reg1E, 
        r_xana[17:0], r_do_ts[6:3], reg1B_3_, r_do_ts[2:0], r_xtm, bkpt_ena, 
        bkpt_pc, r_aopt, 1'b0, 1'b0, d_lt_aswk, sse_idle, 1'b0, r_i2crout, 
        d_lt_gpi, reg14, r_dpdo_sel, r_dndo_sel, r_vpp_en, r_vpp0v_en, 
        r_otp_pwdn_en, r_otp_wpls, r_sap, r_twlb, r_bistdat, reg10_7_, 
        r_bistctl, r_sdischg, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_pwm, r_adummyi, 
        r_bck2, r_bck1, r_bck0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_cvofsx, r_idacsh, r_vcomp}), .DATA_TC(1'b0), .SH({d_regx_addr, 1'b0, 
        1'b0, 1'b0}), .B({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, 
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, 
        SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, 
        SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, 
        SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, 
        SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, 
        SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, 
        SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, 
        SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186, 
        SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188, 
        SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190, 
        SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192, 
        SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194, 
        SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196, 
        SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198, 
        SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200, 
        SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202, 
        SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204, 
        SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206, 
        SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208, 
        SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210, 
        SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212, 
        SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214, 
        SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216, 
        SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218, 
        SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220, 
        SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222, 
        SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224, 
        SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226, 
        SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228, 
        SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230, 
        SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232, 
        SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234, 
        SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236, 
        SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238, 
        SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240, 
        SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242, 
        SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244, 
        SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246, 
        SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248, 
        SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250, 
        SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252, 
        SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254, 
        SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256, 
        SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258, 
        SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260, 
        SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262, 
        SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264, 
        SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266, 
        SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268, 
        SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270, 
        SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272, 
        SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274, 
        SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276, 
        SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278, 
        SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280, 
        SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282, 
        SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, 
        SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314, 
        SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316, 
        SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318, 
        SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322, 
        SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324, 
        SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326, 
        SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328, 
        SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330, 
        SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332, 
        SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334, 
        SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, 
        SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380, 
        SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382, 
        SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384, 
        SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386, 
        SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388, 
        SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390, 
        SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392, 
        SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394, 
        SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396, 
        SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398, 
        SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400, 
        SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402, 
        SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404, 
        SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406, 
        SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408, 
        SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410, 
        SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412, 
        SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414, 
        SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416, 
        SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418, 
        SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420, 
        SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422, 
        SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424, 
        SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426, 
        SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428, 
        SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430, 
        SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432, 
        SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434, 
        SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436, 
        SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438, 
        SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440, 
        SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442, 
        SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444, 
        SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446, 
        SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448, 
        SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450, 
        SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452, 
        SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454, 
        SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456, 
        SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458, 
        SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460, 
        SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462, 
        SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464, 
        SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466, 
        SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468, 
        SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470, 
        SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472, 
        SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474, 
        SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476, 
        SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478, 
        SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480, 
        SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482, 
        SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484, 
        SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486, 
        SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488, 
        SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490, 
        SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492, 
        SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494, 
        SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496, 
        SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498, 
        SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500, 
        SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502, 
        SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504, 
        SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506, 
        SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508, 
        SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510, 
        SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512, 
        SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514, 
        SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516, 
        SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518, 
        SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520, 
        SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522, 
        SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524, 
        SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526, 
        SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528, 
        SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530, 
        SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532, 
        SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534, 
        SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536, 
        SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538, 
        SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540, 
        SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542, 
        SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544, 
        SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546, 
        SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548, 
        SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550, 
        SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552, 
        SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554, 
        SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556, 
        SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558, 
        SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560, 
        SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562, 
        SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564, 
        SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566, 
        SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568, 
        SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570, 
        SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572, 
        SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574, 
        SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576, 
        SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578, 
        SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580, 
        SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582, 
        SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584, 
        SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586, 
        SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588, 
        SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590, 
        SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592, 
        SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594, 
        SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596, 
        SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598, 
        SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600, 
        SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602, 
        SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604, 
        SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606, 
        SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608, 
        SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610, 
        SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612, 
        SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614, 
        SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616, 
        SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618, 
        SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620, 
        SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622, 
        SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624, 
        SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626, 
        SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628, 
        SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630, 
        SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632, 
        SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634, 
        SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636, 
        SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638, 
        SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640, 
        SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642, 
        SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644, 
        SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646, 
        SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648, 
        SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650, 
        SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652, 
        SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654, 
        SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656, 
        SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658, 
        SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660, 
        SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662, 
        SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664, 
        SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666, 
        SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668, 
        SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670, 
        SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672, 
        SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674, 
        SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676, 
        SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678, 
        SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680, 
        SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682, 
        SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684, 
        SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686, 
        SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688, 
        SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690, 
        SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692, 
        SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694, 
        SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696, 
        SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698, 
        SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700, 
        SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702, 
        SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704, 
        SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706, 
        SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708, 
        SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710, 
        SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712, 
        SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714, 
        SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716, 
        SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718, 
        SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720, 
        SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722, 
        SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724, 
        SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726, 
        SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728, 
        SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730, 
        SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732, 
        SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734, 
        SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736, 
        SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738, 
        SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740, 
        SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742, 
        SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744, 
        SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746, 
        SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748, 
        SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750, 
        SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752, 
        SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754, 
        SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756, 
        SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758, 
        SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760, 
        SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762, 
        SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764, 
        SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766, 
        SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768, 
        SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770, 
        SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772, 
        SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774, 
        SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776, 
        SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778, 
        SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780, 
        SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782, 
        SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784, 
        SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786, 
        SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788, 
        SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790, 
        SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792, 
        SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794, 
        SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796, 
        SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798, 
        SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800, 
        SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802, 
        SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804, 
        SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806, 
        SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808, 
        SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810, 
        SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812, 
        SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814, 
        SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816, 
        SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818, 
        SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820, 
        SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822, 
        SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824, 
        SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826, 
        SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828, 
        SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830, 
        SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832, 
        SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834, 
        SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836, 
        SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838, 
        SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840, 
        SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842, 
        SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844, 
        SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846, 
        SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848, 
        SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850, 
        SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852, 
        SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854, 
        SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856, 
        SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858, 
        SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860, 
        SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862, 
        SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864, 
        SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866, 
        SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868, 
        SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870, 
        SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872, 
        SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874, 
        SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876, 
        SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878, 
        SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880, 
        SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882, 
        SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884, 
        SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886, 
        SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888, 
        SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890, 
        SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892, 
        SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894, 
        SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896, 
        SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898, 
        SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900, 
        SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902, 
        SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904, 
        SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906, 
        SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908, 
        SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910, 
        SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912, 
        SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914, 
        SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916, 
        SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918, 
        SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920, 
        SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922, 
        SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924, 
        SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926, 
        SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928, 
        SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930, 
        SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932, 
        SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934, 
        SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936, 
        SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938, 
        SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940, 
        SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942, 
        SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944, 
        SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946, 
        SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948, 
        SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950, 
        SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952, 
        SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954, 
        SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956, 
        SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958, 
        SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960, 
        SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962, 
        SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964, 
        SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966, 
        SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968, 
        SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970, 
        SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972, 
        SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974, 
        SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976, 
        SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978, 
        SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980, 
        SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982, 
        SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984, 
        SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986, 
        SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988, 
        SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990, 
        SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992, 
        SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994, 
        SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996, 
        SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998, 
        SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000, 
        SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002, 
        SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004, 
        SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006, 
        SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008, 
        SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010, 
        SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012, 
        SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014, 
        SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016, regx_rdat}) );
  DFFQX1 d_we16_reg ( .D(N8), .C(clk), .Q(d_we16) );
  DFFQX1 d_lt_aswk_reg_2_ ( .D(lt_aswk[2]), .C(clk), .Q(d_lt_aswk[2]) );
  DFFQX1 d_lt_aswk_reg_1_ ( .D(lt_aswk[1]), .C(clk), .Q(d_lt_aswk[1]) );
  DFFQX1 d_lt_drp_reg ( .D(lt_drp), .C(clk), .Q(reg14[0]) );
  DFFQX1 d_di_tst_reg ( .D(di_tst), .C(clk), .Q(reg14[3]) );
  DFFQX1 d_lt_gpi_reg_1_ ( .D(lt_gpi[1]), .C(net8997), .Q(d_lt_gpi[1]) );
  DFFQX1 d_lt_gpi_reg_0_ ( .D(lt_gpi[0]), .C(net8997), .Q(d_lt_gpi[0]) );
  DFFQX1 d_lt_aswk_reg_5_ ( .D(lt_aswk[5]), .C(clk), .Q(d_lt_aswk[5]) );
  DFFQX1 d_lt_aswk_reg_4_ ( .D(lt_aswk[4]), .C(clk), .Q(d_lt_aswk[4]) );
  DFFQX1 d_lt_aswk_reg_3_ ( .D(lt_aswk[3]), .C(clk), .Q(d_lt_aswk[3]) );
  DFFQX1 d_lt_aswk_reg_0_ ( .D(lt_aswk[0]), .C(clk), .Q(d_lt_aswk[0]) );
  DFFQX1 d_lt_gpi_reg_2_ ( .D(lt_gpi[2]), .C(net8997), .Q(d_lt_gpi[2]) );
  DFFQX1 d_regx_addr_reg_4_ ( .D(n56), .C(clk), .Q(d_regx_addr[4]) );
  DFFQX1 d_lt_gpi_reg_3_ ( .D(lt_gpi[3]), .C(net8997), .Q(d_lt_gpi[3]) );
  DFFQX1 d_regx_addr_reg_3_ ( .D(n48), .C(clk), .Q(d_regx_addr[3]) );
  DFFQX1 d_regx_addr_reg_2_ ( .D(n63), .C(clk), .Q(d_regx_addr[2]) );
  DFFQX1 d_regx_addr_reg_1_ ( .D(n62), .C(clk), .Q(d_regx_addr[1]) );
  DFFQX1 d_regx_addr_reg_0_ ( .D(n54), .C(clk), .Q(d_regx_addr[0]) );
  DFFQX1 d_regx_addr_reg_6_ ( .D(n46), .C(clk), .Q(d_regx_addr[6]) );
  DFFQX1 d_regx_addr_reg_5_ ( .D(n45), .C(clk), .Q(d_regx_addr[5]) );
  DFFRQX1 lt_aswk_reg_5_ ( .D(1'b1), .C(aswclk), .XR(n128), .Q(lt_aswk[5]) );
  DFFRQX1 lt_aswk_reg_4_ ( .D(di_aswk[4]), .C(aswclk), .XR(n128), .Q(
        lt_aswk[4]) );
  DFFRQX1 lt_aswk_reg_3_ ( .D(di_aswk[3]), .C(aswclk), .XR(n128), .Q(
        lt_aswk[3]) );
  DFFRQX1 lt_aswk_reg_2_ ( .D(di_aswk[2]), .C(aswclk), .XR(n128), .Q(
        lt_aswk[2]) );
  DFFRQX1 lt_aswk_reg_1_ ( .D(di_aswk[1]), .C(aswclk), .XR(n128), .Q(
        lt_aswk[1]) );
  DFFRQX1 lt_aswk_reg_0_ ( .D(di_aswk[0]), .C(aswclk), .XR(n128), .Q(
        lt_aswk[0]) );
  DFFRQX1 lt_drp_reg ( .D(di_drposc), .C(detclk), .XR(n87), .Q(lt_drp) );
  NOR31XL U3 ( .C(regx_addr[0]), .A(n63), .B(n101), .Y(n41) );
  AND3XL U5 ( .A(n63), .B(n54), .C(n101), .Y(n28) );
  INVX2 U6 ( .A(regx_addr[2]), .Y(n103) );
  AND2X2 U7 ( .A(n112), .B(n66), .Y(regx_wrdac[6]) );
  NOR31X2 U8 ( .C(n101), .A(n54), .B(n103), .Y(n66) );
  NOR21X1 U9 ( .B(regx_addr[2]), .A(n101), .Y(n60) );
  NOR2X2 U10 ( .A(n104), .B(n33), .Y(regx_wrdac[12]) );
  NAND42X2 U11 ( .C(regx_addr[6]), .D(regx_addr[4]), .A(n37), .B(n58), .Y(n111) );
  NAND5X1 U12 ( .A(n117), .B(n118), .C(n116), .D(n58), .E(regx_w), .Y(n33) );
  NAND21X2 U13 ( .B(n36), .A(n23), .Y(n24) );
  AND2X2 U14 ( .A(regx_addr[4]), .B(regx_w), .Y(n23) );
  AND3X4 U15 ( .A(n52), .B(n31), .C(n53), .Y(regx_wrdac[1]) );
  NOR21X2 U16 ( .B(regx_w), .A(n118), .Y(n37) );
  AND3X2 U17 ( .A(n53), .B(n31), .C(n125), .Y(regx_wrdac[0]) );
  AND2X1 U18 ( .A(n61), .B(n112), .Y(regx_wrdac[9]) );
  NOR21X1 U19 ( .B(n54), .A(n100), .Y(n61) );
  NOR3X1 U20 ( .A(n54), .B(n49), .C(n63), .Y(n34) );
  BUFX1 U21 ( .A(n101), .Y(n49) );
  INVX1 U22 ( .A(n60), .Y(n100) );
  AND2X1 U23 ( .A(n41), .B(n112), .Y(regx_wrdac[5]) );
  NOR2X1 U24 ( .A(n100), .B(n54), .Y(n38) );
  NAND21X1 U25 ( .B(n36), .A(n59), .Y(n109) );
  INVX2 U26 ( .A(n104), .Y(n125) );
  AND2X1 U27 ( .A(n112), .B(n34), .Y(regx_wrdac[4]) );
  INVX1 U28 ( .A(n30), .Y(n31) );
  INVX2 U29 ( .A(regx_addr[3]), .Y(n118) );
  BUFX3 U30 ( .A(regx_addr[0]), .Y(n54) );
  AND2XL U31 ( .A(regx_addr[4]), .B(regx_w), .Y(n59) );
  INVX3 U32 ( .A(n111), .Y(n112) );
  INVX1 U33 ( .A(n109), .Y(n115) );
  INVX1 U34 ( .A(regx_wdat[3]), .Y(n2) );
  INVX1 U35 ( .A(n2), .Y(n3) );
  INVX1 U36 ( .A(n2), .Y(n4) );
  INVX1 U37 ( .A(n127), .Y(n5) );
  INVX1 U38 ( .A(n127), .Y(n6) );
  INVX1 U39 ( .A(regx_wdat[6]), .Y(n7) );
  INVX1 U40 ( .A(n7), .Y(n8) );
  INVX1 U41 ( .A(n7), .Y(n9) );
  INVX1 U42 ( .A(regx_wdat[1]), .Y(n10) );
  INVX1 U43 ( .A(n10), .Y(n11) );
  INVX1 U44 ( .A(regx_wdat[5]), .Y(n12) );
  INVX1 U45 ( .A(n12), .Y(n13) );
  INVX1 U46 ( .A(n12), .Y(n14) );
  INVX1 U47 ( .A(regx_wdat[7]), .Y(n15) );
  INVX1 U48 ( .A(n15), .Y(n16) );
  INVX1 U49 ( .A(n15), .Y(n17) );
  INVX1 U50 ( .A(regx_wdat[2]), .Y(n18) );
  INVX1 U51 ( .A(n18), .Y(n19) );
  INVX1 U52 ( .A(n18), .Y(n20) );
  INVXL U53 ( .A(n1047), .Y(n21) );
  INVXL U54 ( .A(n21), .Y(n22) );
  INVXL U55 ( .A(n49), .Y(n62) );
  INVX3 U56 ( .A(n103), .Y(n63) );
  INVX2 U57 ( .A(n119), .Y(n120) );
  INVX3 U58 ( .A(regx_addr[1]), .Y(n101) );
  NOR32X2 U59 ( .B(n101), .C(regx_addr[0]), .A(n63), .Y(n52) );
  NAND21X2 U60 ( .B(regx_addr[6]), .A(n27), .Y(n113) );
  BUFXL U61 ( .A(n34), .Y(n25) );
  BUFXL U62 ( .A(n28), .Y(n26) );
  INVX2 U63 ( .A(regx_addr[4]), .Y(n116) );
  BUFX3 U64 ( .A(regx_addr[5]), .Y(n58) );
  INVXL U65 ( .A(n118), .Y(n27) );
  INVXL U66 ( .A(n104), .Y(n29) );
  INVXL U67 ( .A(n117), .Y(n30) );
  INVX2 U68 ( .A(regx_addr[6]), .Y(n117) );
  INVXL U69 ( .A(regx_addr[2]), .Y(n32) );
  INVXL U70 ( .A(n113), .Y(n114) );
  BUFXL U71 ( .A(n52), .Y(n35) );
  INVXL U72 ( .A(regx_addr[5]), .Y(n36) );
  NOR2X2 U73 ( .A(n24), .B(n48), .Y(n53) );
  AND2X2 U74 ( .A(n112), .B(n38), .Y(regx_wrdac[8]) );
  BUFXL U75 ( .A(n58), .Y(n39) );
  NOR3X1 U76 ( .A(n104), .B(n24), .C(n113), .Y(regx_wrdac[10]) );
  BUFXL U77 ( .A(n61), .Y(n40) );
  AND2XL U78 ( .A(n105), .B(n26), .Y(we[29]) );
  AND2XL U79 ( .A(n121), .B(n26), .Y(we_5) );
  BUFXL U80 ( .A(n38), .Y(n42) );
  INVXL U81 ( .A(n118), .Y(n48) );
  INVXL U82 ( .A(n39), .Y(n43) );
  INVXL U83 ( .A(n43), .Y(n44) );
  BUFXL U84 ( .A(n44), .Y(n45) );
  INVXL U85 ( .A(n31), .Y(n46) );
  INVXL U86 ( .A(n48), .Y(n47) );
  BUFXL U87 ( .A(n66), .Y(n50) );
  INVXL U88 ( .A(n26), .Y(n51) );
  INVXL U89 ( .A(n35), .Y(n110) );
  AND2XL U90 ( .A(n40), .B(n107), .Y(we[23]) );
  NAND32X2 U91 ( .B(regx_addr[0]), .C(regx_addr[1]), .A(n32), .Y(n104) );
  AND3X2 U92 ( .A(n52), .B(n115), .C(n114), .Y(regx_wrdac[11]) );
  BUFXL U93 ( .A(n41), .Y(n55) );
  NAND21XL U94 ( .B(n51), .A(n107), .Y(n1047) );
  INVXL U95 ( .A(n116), .Y(n56) );
  INVX1 U96 ( .A(n56), .Y(n57) );
  AND2XL U97 ( .A(n105), .B(n25), .Y(we[26]) );
  NAND21XL U98 ( .B(n106), .A(n25), .Y(n98) );
  AND2XL U99 ( .A(n121), .B(n34), .Y(regx_wrcvc[2]) );
  AND2XL U100 ( .A(n55), .B(n107), .Y(we_19) );
  AND2XL U101 ( .A(n105), .B(n55), .Y(we[27]) );
  AND2XL U102 ( .A(n40), .B(n123), .Y(regx_wrcvc[3]) );
  AND2XL U103 ( .A(n121), .B(n40), .Y(we_7) );
  NAND5X2 U104 ( .A(n117), .B(n118), .C(n116), .D(n58), .E(regx_w), .Y(n119)
         );
  AND2X2 U105 ( .A(n120), .B(n52), .Y(regx_wrdac[13]) );
  AND2X2 U106 ( .A(n28), .B(n112), .Y(regx_wrdac[7]) );
  INVX1 U107 ( .A(n129), .Y(n64) );
  INVX1 U108 ( .A(n64), .Y(r_i2crout[5]) );
  BUFX3 U109 ( .A(r_imp_osc), .Y(r_xana[22]) );
  AND2XL U110 ( .A(n29), .B(n126), .Y(regx_hitbst[0]) );
  AND2XL U111 ( .A(n121), .B(n29), .Y(regx_wrcvc[0]) );
  AND2XL U112 ( .A(n123), .B(n29), .Y(regx_wrpwm[0]) );
  AND2XL U113 ( .A(n105), .B(n42), .Y(we[30]) );
  AND2XL U114 ( .A(n105), .B(n29), .Y(we[24]) );
  AND2XL U115 ( .A(n121), .B(n42), .Y(we_6) );
  INVX1 U116 ( .A(n92), .Y(n91) );
  INVX1 U117 ( .A(n92), .Y(n88) );
  INVX1 U118 ( .A(n93), .Y(n90) );
  INVX1 U119 ( .A(n92), .Y(n89) );
  INVX1 U120 ( .A(n93), .Y(n80) );
  INVX1 U121 ( .A(n93), .Y(n81) );
  INVX1 U122 ( .A(n92), .Y(n82) );
  INVX1 U123 ( .A(n93), .Y(n79) );
  INVX1 U124 ( .A(n94), .Y(n78) );
  INVX1 U125 ( .A(n94), .Y(n77) );
  INVX1 U126 ( .A(n94), .Y(n76) );
  INVX1 U127 ( .A(n92), .Y(n75) );
  INVX1 U128 ( .A(n93), .Y(n74) );
  INVX1 U129 ( .A(n92), .Y(n73) );
  INVX1 U130 ( .A(n93), .Y(n72) );
  INVX1 U131 ( .A(n93), .Y(n71) );
  INVX1 U132 ( .A(n92), .Y(n70) );
  INVX1 U133 ( .A(n93), .Y(n83) );
  INVX1 U134 ( .A(n93), .Y(n84) );
  INVX1 U135 ( .A(n92), .Y(n87) );
  INVX1 U136 ( .A(n92), .Y(n85) );
  INVX1 U137 ( .A(n93), .Y(n86) );
  INVX1 U138 ( .A(n97), .Y(wd_twlb[0]) );
  INVX1 U139 ( .A(n97), .Y(n96) );
  INVX1 U140 ( .A(rrstz), .Y(n94) );
  INVX1 U141 ( .A(rrstz), .Y(n92) );
  INVX1 U142 ( .A(rrstz), .Y(n93) );
  INVX1 U143 ( .A(n124), .Y(n126) );
  INVX1 U144 ( .A(n106), .Y(n107) );
  AND2XL U145 ( .A(n123), .B(n35), .Y(regx_wrpwm[1]) );
  AND2XL U146 ( .A(n121), .B(n35), .Y(regx_wrcvc[1]) );
  INVX1 U147 ( .A(regx_wdat[0]), .Y(n97) );
  AND2XL U148 ( .A(n112), .B(n125), .Y(regx_wrdac[2]) );
  AND2XL U149 ( .A(n112), .B(n52), .Y(regx_wrdac[3]) );
  NAND32XL U150 ( .B(n57), .C(n67), .A(n47), .Y(n124) );
  INVX1 U151 ( .A(n122), .Y(n123) );
  NAND21X1 U152 ( .B(n124), .A(regx_w), .Y(n106) );
  INVX1 U153 ( .A(n98), .Y(we_twlb) );
  INVX1 U154 ( .A(n102), .Y(we[25]) );
  INVX1 U155 ( .A(n99), .Y(n105) );
  INVX1 U156 ( .A(n108), .Y(n121) );
  NAND5XL U157 ( .A(regx_w), .B(n47), .C(n57), .D(n43), .E(n31), .Y(n108) );
  AND2XL U158 ( .A(n35), .B(n126), .Y(regx_hitbst[1]) );
  AND2X1 U159 ( .A(n105), .B(n50), .Y(we[28]) );
  AND2X1 U160 ( .A(n50), .B(n121), .Y(we_4) );
  OR2XL U161 ( .A(n45), .B(n46), .Y(n67) );
  OAI31XL U162 ( .A(n15), .B(n9), .C(n22), .D(n1048), .Y(i2c_mode_upd) );
  OAI21X1 U163 ( .B(n1049), .C(n1050), .A(bus_idle), .Y(n1048) );
  NAND3X1 U164 ( .A(n1051), .B(n1052), .C(n1053), .Y(n1050) );
  NOR4XL U165 ( .A(n1057), .B(n1058), .C(regx_wdat[3]), .D(n19), .Y(N8) );
  NAND3X1 U166 ( .A(n12), .B(n10), .C(n127), .Y(n1058) );
  NAND5XL U167 ( .A(n16), .B(n1059), .C(n8), .D(n42), .E(n126), .Y(n1057) );
  AND2X1 U168 ( .A(regx_w), .B(wd_twlb[0]), .Y(n1059) );
  INVXL U169 ( .A(regx_wdat[4]), .Y(n127) );
  XNOR2XL U170 ( .A(reg1E[3]), .B(n1046), .Y(r_xana[19]) );
  XNOR2XL U171 ( .A(reg1E[2]), .B(n1046), .Y(r_xana[18]) );
  NAND2X1 U172 ( .A(r_xana[20]), .B(di_drposc), .Y(n1046) );
  BUFX3 U173 ( .A(n11), .Y(wd_twlb[1]) );
  NAND4X1 U174 ( .A(n1054), .B(n1055), .C(n1056), .D(n22), .Y(n1049) );
  XNOR2XL U175 ( .A(r_i2crout[3]), .B(lt_reg15_5_0[3]), .Y(n1054) );
  XNOR2XL U176 ( .A(r_i2crout[4]), .B(lt_reg15_5_0[4]), .Y(n1055) );
  XNOR2XL U177 ( .A(n129), .B(lt_reg15_5_0[5]), .Y(n1056) );
  AO22X1 U178 ( .A(n21), .B(wd_twlb[0]), .C(n22), .D(lt_reg15_5_0[0]), .Y(
        i2c_mode_wdat[0]) );
  AO22X1 U179 ( .A(n21), .B(n20), .C(n1047), .D(lt_reg15_5_0[2]), .Y(
        i2c_mode_wdat[2]) );
  AO22X1 U180 ( .A(n21), .B(n3), .C(n22), .D(lt_reg15_5_0[3]), .Y(
        i2c_mode_wdat[3]) );
  ENOX1 U181 ( .A(n1047), .B(n127), .C(n22), .D(lt_reg15_5_0[4]), .Y(
        i2c_mode_wdat[4]) );
  ENOX1 U182 ( .A(n22), .B(n12), .C(n1047), .D(lt_reg15_5_0[5]), .Y(
        i2c_mode_wdat[5]) );
  ENOX1 U183 ( .A(n1047), .B(n10), .C(n22), .D(lt_reg15_5_0[1]), .Y(
        i2c_mode_wdat[1]) );
  XNOR2XL U184 ( .A(r_i2crout[2]), .B(lt_reg15_5_0[2]), .Y(n1051) );
  XNOR2XL U185 ( .A(r_i2crout[0]), .B(lt_reg15_5_0[0]), .Y(n1052) );
  XNOR2XL U186 ( .A(r_i2crout[1]), .B(lt_reg15_5_0[1]), .Y(n1053) );
  INVX1 U187 ( .A(n1060), .Y(n128) );
  OAI21BX1 U188 ( .C(d_we16), .B(atpg_en), .A(n85), .Y(n1060) );
  NAND21XL U189 ( .B(n110), .A(n105), .Y(n102) );
  NAND32XL U190 ( .B(n56), .C(n67), .A(n37), .Y(n122) );
  NAND32XL U191 ( .B(n67), .C(n47), .A(n23), .Y(n99) );
endmodule


module regx_a0_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680;

  NOR21X1 U2149 ( .B(n3362), .A(n3277), .Y(n3361) );
  MUX2X1 U2150 ( .D0(n3327), .D1(n3328), .S(n3213), .Y(n3210) );
  NOR2X1 U2151 ( .A(n3202), .B(n3277), .Y(n3323) );
  MUX2X1 U2152 ( .D0(A[79]), .D1(A[335]), .S(n3227), .Y(n3202) );
  INVX1 U2153 ( .A(n3228), .Y(n3199) );
  INVX1 U2154 ( .A(n3228), .Y(n3192) );
  NOR21XL U2155 ( .B(n3411), .A(n3274), .Y(n3410) );
  INVX1 U2156 ( .A(n3228), .Y(n3197) );
  NOR21XL U2157 ( .B(n3461), .A(n3279), .Y(n3460) );
  INVX1 U2158 ( .A(n3189), .Y(n3461) );
  INVX1 U2159 ( .A(SH[7]), .Y(n3196) );
  MUX2X1 U2160 ( .D0(n3373), .D1(n3209), .S(n3225), .Y(n3354) );
  MUX2X1 U2161 ( .D0(n3623), .D1(n3207), .S(SH[4]), .Y(n3604) );
  MUX2X1 U2162 ( .D0(n3472), .D1(n3208), .S(n3225), .Y(n3453) );
  NOR21XL U2163 ( .B(n3317), .A(n3278), .Y(n3316) );
  INVX1 U2164 ( .A(SH[6]), .Y(n3201) );
  NAND2X1 U2165 ( .A(A[380]), .B(n3186), .Y(n3187) );
  NAND2X1 U2166 ( .A(A[124]), .B(n3191), .Y(n3188) );
  NAND2X1 U2167 ( .A(n3187), .B(n3188), .Y(n3189) );
  INVX1 U2168 ( .A(n3191), .Y(n3186) );
  INVX1 U2169 ( .A(n3233), .Y(n3191) );
  INVX1 U2170 ( .A(n3197), .Y(n3195) );
  MUX2X1 U2171 ( .D0(n3311), .D1(n3310), .S(n3201), .Y(n3190) );
  NOR32XL U2172 ( .B(n3254), .C(n3280), .A(A[375]), .Y(n3314) );
  NOR21X1 U2173 ( .B(n3510), .A(n3275), .Y(n3509) );
  MUX2IX1 U2174 ( .D0(A[271]), .D1(A[15]), .S(n3192), .Y(n3329) );
  MUX4IX1 U2175 ( .D0(n3314), .D1(n3313), .D2(n3316), .D3(n3315), .S0(n3226), 
        .S1(n3216), .Y(n3193) );
  NAND2X1 U2176 ( .A(n3196), .B(n3203), .Y(n3194) );
  MUX2IX1 U2177 ( .D0(A[127]), .D1(A[383]), .S(n3195), .Y(n3317) );
  MUX2IX1 U2178 ( .D0(n3193), .D1(n3200), .S(n3194), .Y(n3287) );
  NOR2X1 U2179 ( .A(SH[7]), .B(SH[5]), .Y(n3198) );
  MUX2IX1 U2180 ( .D0(A[263]), .D1(A[7]), .S(n3199), .Y(n3330) );
  MUX2IX1 U2181 ( .D0(n3205), .D1(n3312), .S(n3196), .Y(n3200) );
  MUX4X1 U2182 ( .D0(n3324), .D1(n3325), .D2(n3322), .D3(n3323), .S0(n3212), 
        .S1(n3226), .Y(n3311) );
  BUFX3 U2183 ( .A(SH[6]), .Y(n3203) );
  BUFX3 U2184 ( .A(SH[5]), .Y(n3204) );
  NOR4XL U2185 ( .A(n3274), .B(n3234), .C(n3218), .D(A[17]), .Y(n3207) );
  NOR4XL U2186 ( .A(n3274), .B(n3235), .C(n3218), .D(A[20]), .Y(n3208) );
  NOR4XL U2187 ( .A(n3273), .B(n3234), .C(SH[3]), .D(A[22]), .Y(n3209) );
  MUX2IX1 U2188 ( .D0(n3287), .D1(n3190), .S(n3198), .Y(B[7]) );
  MUX4X1 U2189 ( .D0(n3288), .D1(n3289), .D2(n3290), .D3(n3291), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3205) );
  MUX2IX1 U2190 ( .D0(n3577), .D1(n3206), .S(SH[7]), .Y(B[1]) );
  MUX4X1 U2191 ( .D0(n3578), .D1(n3579), .D2(n3580), .D3(n3581), .S0(n3204), 
        .S1(n3203), .Y(n3206) );
  INVX1 U2192 ( .A(n3247), .Y(n3228) );
  INVX1 U2193 ( .A(n3248), .Y(n3227) );
  INVX1 U2194 ( .A(n3280), .Y(n3260) );
  INVX1 U2195 ( .A(n3245), .Y(n3234) );
  INVX1 U2196 ( .A(n3282), .Y(n3268) );
  INVX1 U2197 ( .A(n3281), .Y(n3263) );
  INVX1 U2198 ( .A(n3281), .Y(n3269) );
  INVX1 U2199 ( .A(n3282), .Y(n3278) );
  INVX1 U2200 ( .A(n3282), .Y(n3277) );
  INVX1 U2201 ( .A(n3245), .Y(n3235) );
  INVX1 U2202 ( .A(n3244), .Y(n3236) );
  INVX1 U2203 ( .A(n3242), .Y(n3240) );
  INVX1 U2204 ( .A(n3282), .Y(n3279) );
  INVX1 U2205 ( .A(n3242), .Y(n3241) );
  INVX1 U2206 ( .A(n3280), .Y(n3261) );
  INVX1 U2207 ( .A(n3286), .Y(n3274) );
  INVX1 U2208 ( .A(n3246), .Y(n3232) );
  INVX1 U2209 ( .A(n3247), .Y(n3229) );
  INVX1 U2210 ( .A(n3246), .Y(n3231) );
  INVX1 U2211 ( .A(n3246), .Y(n3233) );
  INVX1 U2212 ( .A(n3247), .Y(n3230) );
  INVX1 U2213 ( .A(n3281), .Y(n3262) );
  INVX1 U2214 ( .A(n3281), .Y(n3271) );
  INVX1 U2215 ( .A(n3281), .Y(n3264) );
  INVX1 U2216 ( .A(n3281), .Y(n3270) );
  INVX1 U2217 ( .A(n3243), .Y(n3239) );
  INVX1 U2218 ( .A(n3243), .Y(n3237) );
  INVX1 U2219 ( .A(n3280), .Y(n3267) );
  INVX1 U2220 ( .A(n3282), .Y(n3266) );
  INVX1 U2221 ( .A(n3282), .Y(n3272) );
  INVX1 U2222 ( .A(n3286), .Y(n3265) );
  INVX1 U2223 ( .A(n3281), .Y(n3273) );
  INVX1 U2224 ( .A(n3282), .Y(n3276) );
  INVX1 U2225 ( .A(n3282), .Y(n3275) );
  INVX1 U2226 ( .A(n3243), .Y(n3238) );
  INVX1 U2227 ( .A(n3256), .Y(n3248) );
  INVX1 U2228 ( .A(n3285), .Y(n3280) );
  INVX1 U2229 ( .A(n3257), .Y(n3247) );
  INVX1 U2230 ( .A(n3257), .Y(n3245) );
  INVX1 U2231 ( .A(n3258), .Y(n3244) );
  INVX1 U2232 ( .A(n3283), .Y(n3282) );
  INVX1 U2233 ( .A(n3258), .Y(n3242) );
  INVX1 U2234 ( .A(n3285), .Y(n3281) );
  INVX1 U2235 ( .A(n3255), .Y(n3250) );
  INVX1 U2236 ( .A(n3257), .Y(n3246) );
  INVX1 U2237 ( .A(n3258), .Y(n3243) );
  INVX1 U2238 ( .A(n3255), .Y(n3249) );
  INVX1 U2239 ( .A(n3255), .Y(n3251) );
  INVX1 U2240 ( .A(n3254), .Y(n3252) );
  INVX1 U2241 ( .A(n3259), .Y(n3257) );
  INVX1 U2242 ( .A(n3286), .Y(n3284) );
  INVX1 U2243 ( .A(n3259), .Y(n3256) );
  INVX1 U2244 ( .A(n3286), .Y(n3283) );
  INVX1 U2245 ( .A(n3259), .Y(n3258) );
  INVX1 U2246 ( .A(n3286), .Y(n3285) );
  INVX1 U2247 ( .A(n3219), .Y(n3212) );
  INVX1 U2248 ( .A(n3226), .Y(n3224) );
  INVX1 U2249 ( .A(n3219), .Y(n3213) );
  INVX1 U2250 ( .A(n3219), .Y(n3216) );
  INVX1 U2251 ( .A(n3219), .Y(n3218) );
  INVX1 U2252 ( .A(n3243), .Y(n3255) );
  INVX1 U2253 ( .A(n3226), .Y(n3225) );
  INVX1 U2254 ( .A(n3226), .Y(n3221) );
  INVX1 U2255 ( .A(n3243), .Y(n3254) );
  INVX1 U2256 ( .A(n3255), .Y(n3253) );
  INVX1 U2257 ( .A(n3226), .Y(n3222) );
  INVX1 U2258 ( .A(n3226), .Y(n3223) );
  INVX1 U2259 ( .A(n3219), .Y(n3217) );
  INVX1 U2260 ( .A(n3219), .Y(n3215) );
  INVX1 U2261 ( .A(n3219), .Y(n3214) );
  MUX2IX1 U2262 ( .D0(n3210), .D1(n3211), .S(n3225), .Y(n3310) );
  OR4X1 U2263 ( .A(n3274), .B(n3234), .C(n3218), .D(A[23]), .Y(n3211) );
  INVX1 U2264 ( .A(SH[8]), .Y(n3259) );
  INVX1 U2265 ( .A(SH[9]), .Y(n3286) );
  INVX1 U2266 ( .A(SH[3]), .Y(n3219) );
  INVX1 U2267 ( .A(n3226), .Y(n3220) );
  INVX1 U2268 ( .A(SH[4]), .Y(n3226) );
  MUX4X1 U2269 ( .D0(n3292), .D1(n3293), .D2(n3294), .D3(n3295), .S0(n3220), 
        .S1(n3216), .Y(n3291) );
  NOR3XL U2270 ( .A(A[255]), .B(n3263), .C(n3236), .Y(n3295) );
  NOR3XL U2271 ( .A(A[239]), .B(n3268), .C(n3235), .Y(n3294) );
  NOR3XL U2272 ( .A(A[247]), .B(n3268), .C(n3241), .Y(n3293) );
  NOR3XL U2273 ( .A(A[231]), .B(n3268), .C(n3241), .Y(n3292) );
  MUX4X1 U2274 ( .D0(n3296), .D1(n3297), .D2(n3298), .D3(n3299), .S0(n3220), 
        .S1(n3218), .Y(n3290) );
  NOR3XL U2275 ( .A(A[223]), .B(n3268), .C(n3241), .Y(n3299) );
  AOI21X1 U2276 ( .B(A[207]), .C(n3248), .A(n3260), .Y(n3298) );
  AOI21X1 U2277 ( .B(A[215]), .C(n3248), .A(n3260), .Y(n3297) );
  AOI21X1 U2278 ( .B(A[199]), .C(n3248), .A(n3260), .Y(n3296) );
  MUX3X1 U2279 ( .D0(n3300), .D1(n3301), .D2(n3302), .S0(n3218), .S1(n3225), 
        .Y(n3289) );
  AOI211X1 U2280 ( .C(n3218), .D(A[191]), .A(n3261), .B(n3234), .Y(n3302) );
  NOR3XL U2281 ( .A(A[175]), .B(n3268), .C(n3241), .Y(n3301) );
  NOR3XL U2282 ( .A(A[167]), .B(n3268), .C(n3241), .Y(n3300) );
  MUX4X1 U2283 ( .D0(n3303), .D1(n3304), .D2(n3305), .D3(n3306), .S0(n3220), 
        .S1(n3216), .Y(n3288) );
  NOR3XL U2284 ( .A(A[159]), .B(n3268), .C(n3241), .Y(n3306) );
  NOR21XL U2285 ( .B(n3307), .A(n3279), .Y(n3305) );
  MUX2IX1 U2286 ( .D0(A[143]), .D1(A[399]), .S(n3227), .Y(n3307) );
  NOR21XL U2287 ( .B(n3308), .A(n3278), .Y(n3304) );
  MUX2IX1 U2288 ( .D0(A[151]), .D1(A[407]), .S(n3227), .Y(n3308) );
  NOR21XL U2289 ( .B(n3309), .A(n3278), .Y(n3303) );
  MUX2IX1 U2290 ( .D0(A[135]), .D1(A[391]), .S(n3227), .Y(n3309) );
  NOR3XL U2291 ( .A(n3250), .B(n3269), .C(A[367]), .Y(n3315) );
  NOR3XL U2292 ( .A(n3253), .B(n3269), .C(A[359]), .Y(n3313) );
  MUX4X1 U2293 ( .D0(n3318), .D1(n3319), .D2(n3320), .D3(n3321), .S0(n3220), 
        .S1(n3216), .Y(n3312) );
  NOR3XL U2294 ( .A(A[63]), .B(n3269), .C(n3241), .Y(n3321) );
  NOR3XL U2295 ( .A(A[47]), .B(n3269), .C(n3240), .Y(n3320) );
  NOR3XL U2296 ( .A(A[55]), .B(n3269), .C(n3240), .Y(n3319) );
  NOR3XL U2297 ( .A(A[39]), .B(n3269), .C(n3240), .Y(n3318) );
  NOR3XL U2298 ( .A(n3243), .B(n3269), .C(A[351]), .Y(n3325) );
  NOR3XL U2299 ( .A(n3243), .B(n3269), .C(A[343]), .Y(n3324) );
  NOR21XL U2300 ( .B(n3326), .A(n3277), .Y(n3322) );
  MUX2IX1 U2301 ( .D0(A[71]), .D1(A[327]), .S(n3228), .Y(n3326) );
  NAND2X1 U2302 ( .A(n3329), .B(n3280), .Y(n3328) );
  NAND2X1 U2303 ( .A(n3330), .B(n3286), .Y(n3327) );
  MUX2IX1 U2304 ( .D0(n3331), .D1(n3332), .S(SH[7]), .Y(B[6]) );
  MUX4X1 U2305 ( .D0(n3333), .D1(n3334), .D2(n3335), .D3(n3336), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3332) );
  MUX4X1 U2306 ( .D0(n3337), .D1(n3338), .D2(n3339), .D3(n3340), .S0(n3220), 
        .S1(n3215), .Y(n3336) );
  NOR3XL U2307 ( .A(A[254]), .B(n3269), .C(n3240), .Y(n3340) );
  NOR3XL U2308 ( .A(A[238]), .B(SH[9]), .C(n3240), .Y(n3339) );
  NOR3XL U2309 ( .A(A[246]), .B(n3285), .C(n3240), .Y(n3338) );
  NOR3XL U2310 ( .A(A[230]), .B(SH[9]), .C(n3240), .Y(n3337) );
  MUX4X1 U2311 ( .D0(n3341), .D1(n3342), .D2(n3343), .D3(n3344), .S0(n3220), 
        .S1(n3214), .Y(n3335) );
  NOR3XL U2312 ( .A(A[222]), .B(SH[9]), .C(n3240), .Y(n3344) );
  AOI21X1 U2313 ( .B(A[206]), .C(n3243), .A(n3260), .Y(n3343) );
  AOI21X1 U2314 ( .B(A[214]), .C(n3243), .A(n3261), .Y(n3342) );
  AOI21X1 U2315 ( .B(A[198]), .C(n3252), .A(n3261), .Y(n3341) );
  MUX2X1 U2316 ( .D0(n3345), .D1(n3346), .S(n3225), .Y(n3334) );
  AOI211X1 U2317 ( .C(n3218), .D(A[190]), .A(n3262), .B(n3234), .Y(n3346) );
  AOI211X1 U2318 ( .C(A[166]), .D(n3219), .A(n3261), .B(n3234), .Y(n3345) );
  MUX4X1 U2319 ( .D0(n3347), .D1(n3348), .D2(n3349), .D3(n3350), .S0(n3221), 
        .S1(n3214), .Y(n3333) );
  NOR3XL U2320 ( .A(A[158]), .B(SH[9]), .C(n3240), .Y(n3350) );
  NOR21XL U2321 ( .B(n3351), .A(n3277), .Y(n3349) );
  MUX2IX1 U2322 ( .D0(A[142]), .D1(A[398]), .S(n3229), .Y(n3351) );
  NOR21XL U2323 ( .B(n3352), .A(n3275), .Y(n3348) );
  MUX2IX1 U2324 ( .D0(A[150]), .D1(A[406]), .S(n3229), .Y(n3352) );
  NOR21XL U2325 ( .B(n3353), .A(n3275), .Y(n3347) );
  MUX2IX1 U2326 ( .D0(A[134]), .D1(A[390]), .S(n3228), .Y(n3353) );
  MUX4X1 U2327 ( .D0(n3354), .D1(n3355), .D2(n3356), .D3(n3357), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3331) );
  MUX4X1 U2328 ( .D0(n3358), .D1(n3359), .D2(n3360), .D3(n3361), .S0(n3221), 
        .S1(n3213), .Y(n3357) );
  MUX2IX1 U2329 ( .D0(A[126]), .D1(A[382]), .S(n3229), .Y(n3362) );
  NOR3XL U2330 ( .A(n3250), .B(SH[9]), .C(A[366]), .Y(n3360) );
  NOR3XL U2331 ( .A(n3253), .B(n3284), .C(A[374]), .Y(n3359) );
  NOR3XL U2332 ( .A(n3253), .B(n3283), .C(A[358]), .Y(n3358) );
  MUX4X1 U2333 ( .D0(n3363), .D1(n3364), .D2(n3365), .D3(n3366), .S0(n3221), 
        .S1(n3213), .Y(n3356) );
  NOR3XL U2334 ( .A(A[62]), .B(SH[9]), .C(n3240), .Y(n3366) );
  NOR3XL U2335 ( .A(A[46]), .B(n3285), .C(n3257), .Y(n3365) );
  NOR3XL U2336 ( .A(A[54]), .B(n3270), .C(n3195), .Y(n3364) );
  NOR3XL U2337 ( .A(A[38]), .B(n3270), .C(n3257), .Y(n3363) );
  MUX4X1 U2338 ( .D0(n3367), .D1(n3368), .D2(n3369), .D3(n3370), .S0(n3212), 
        .S1(n3225), .Y(n3355) );
  NOR3XL U2339 ( .A(n3253), .B(n3270), .C(A[350]), .Y(n3370) );
  NOR3XL U2340 ( .A(n3253), .B(n3270), .C(A[342]), .Y(n3369) );
  NOR21XL U2341 ( .B(n3371), .A(n3275), .Y(n3368) );
  MUX2IX1 U2342 ( .D0(A[78]), .D1(A[334]), .S(n3229), .Y(n3371) );
  NOR21XL U2343 ( .B(n3372), .A(n3276), .Y(n3367) );
  MUX2IX1 U2344 ( .D0(A[70]), .D1(A[326]), .S(n3230), .Y(n3372) );
  MUX2IX1 U2345 ( .D0(n3374), .D1(n3375), .S(n3213), .Y(n3373) );
  NAND2X1 U2346 ( .A(n3376), .B(n3280), .Y(n3375) );
  MUX2IX1 U2347 ( .D0(A[14]), .D1(A[270]), .S(n3229), .Y(n3376) );
  NAND2X1 U2348 ( .A(n3377), .B(n3280), .Y(n3374) );
  MUX2IX1 U2349 ( .D0(A[6]), .D1(A[262]), .S(n3230), .Y(n3377) );
  MUX2IX1 U2350 ( .D0(n3378), .D1(n3379), .S(SH[7]), .Y(B[5]) );
  MUX4X1 U2351 ( .D0(n3380), .D1(n3381), .D2(n3382), .D3(n3383), .S0(SH[5]), 
        .S1(n3203), .Y(n3379) );
  MUX4X1 U2352 ( .D0(n3384), .D1(n3385), .D2(n3386), .D3(n3387), .S0(n3221), 
        .S1(n3213), .Y(n3383) );
  NOR3XL U2353 ( .A(A[253]), .B(n3270), .C(n3257), .Y(n3387) );
  NOR3XL U2354 ( .A(A[237]), .B(n3270), .C(n3256), .Y(n3386) );
  NOR3XL U2355 ( .A(A[245]), .B(n3270), .C(n3257), .Y(n3385) );
  NOR3XL U2356 ( .A(A[229]), .B(n3270), .C(n3257), .Y(n3384) );
  MUX4X1 U2357 ( .D0(n3388), .D1(n3389), .D2(n3390), .D3(n3391), .S0(n3221), 
        .S1(n3214), .Y(n3382) );
  NOR3XL U2358 ( .A(A[221]), .B(n3270), .C(n3195), .Y(n3391) );
  AOI21X1 U2359 ( .B(A[205]), .C(n3251), .A(n3261), .Y(n3390) );
  AOI21X1 U2360 ( .B(A[213]), .C(n3250), .A(n3261), .Y(n3389) );
  AOI21X1 U2361 ( .B(A[197]), .C(n3252), .A(n3261), .Y(n3388) );
  MUX4X1 U2362 ( .D0(n3392), .D1(n3393), .D2(n3394), .D3(n3395), .S0(n3221), 
        .S1(n3214), .Y(n3381) );
  NOR3XL U2363 ( .A(A[189]), .B(n3270), .C(n3257), .Y(n3395) );
  NOR3XL U2364 ( .A(A[173]), .B(n3271), .C(n3257), .Y(n3394) );
  NOR3XL U2365 ( .A(A[181]), .B(n3271), .C(n3239), .Y(n3393) );
  NOR3XL U2366 ( .A(A[165]), .B(n3271), .C(n3239), .Y(n3392) );
  MUX4X1 U2367 ( .D0(n3396), .D1(n3397), .D2(n3398), .D3(n3399), .S0(n3221), 
        .S1(n3214), .Y(n3380) );
  NOR3XL U2368 ( .A(A[157]), .B(n3271), .C(n3239), .Y(n3399) );
  NOR21XL U2369 ( .B(n3400), .A(n3274), .Y(n3398) );
  MUX2IX1 U2370 ( .D0(A[141]), .D1(A[397]), .S(n3230), .Y(n3400) );
  NOR21XL U2371 ( .B(n3401), .A(n3274), .Y(n3397) );
  MUX2IX1 U2372 ( .D0(A[149]), .D1(A[405]), .S(n3231), .Y(n3401) );
  NOR21XL U2373 ( .B(n3402), .A(n3275), .Y(n3396) );
  MUX2IX1 U2374 ( .D0(A[133]), .D1(A[389]), .S(n3231), .Y(n3402) );
  MUX4X1 U2375 ( .D0(n3403), .D1(n3404), .D2(n3405), .D3(n3406), .S0(SH[6]), 
        .S1(n3204), .Y(n3378) );
  MUX4X1 U2376 ( .D0(n3407), .D1(n3408), .D2(n3409), .D3(n3410), .S0(n3222), 
        .S1(n3214), .Y(n3406) );
  MUX2IX1 U2377 ( .D0(A[125]), .D1(A[381]), .S(n3230), .Y(n3411) );
  NOR3XL U2378 ( .A(n3253), .B(n3271), .C(A[365]), .Y(n3409) );
  NOR3XL U2379 ( .A(n3253), .B(n3271), .C(A[373]), .Y(n3408) );
  NOR3XL U2380 ( .A(n3252), .B(n3272), .C(A[357]), .Y(n3407) );
  MUX4X1 U2381 ( .D0(n3412), .D1(n3413), .D2(n3414), .D3(n3415), .S0(n3222), 
        .S1(n3214), .Y(n3405) );
  NOR3XL U2382 ( .A(A[61]), .B(n3271), .C(n3239), .Y(n3415) );
  NOR3XL U2383 ( .A(A[45]), .B(n3272), .C(n3239), .Y(n3414) );
  NOR3XL U2384 ( .A(A[53]), .B(n3272), .C(n3239), .Y(n3413) );
  NOR3XL U2385 ( .A(A[37]), .B(n3271), .C(n3239), .Y(n3412) );
  MUX4X1 U2386 ( .D0(n3416), .D1(n3417), .D2(n3418), .D3(n3419), .S0(n3212), 
        .S1(n3224), .Y(n3404) );
  NOR3XL U2387 ( .A(n3252), .B(n3272), .C(A[349]), .Y(n3419) );
  NOR3XL U2388 ( .A(n3252), .B(n3273), .C(A[341]), .Y(n3418) );
  NOR21XL U2389 ( .B(n3420), .A(n3276), .Y(n3417) );
  MUX2IX1 U2390 ( .D0(A[77]), .D1(A[333]), .S(n3232), .Y(n3420) );
  NOR21XL U2391 ( .B(n3421), .A(n3276), .Y(n3416) );
  MUX2IX1 U2392 ( .D0(A[69]), .D1(A[325]), .S(n3230), .Y(n3421) );
  MUX2X1 U2393 ( .D0(n3422), .D1(n3423), .S(n3225), .Y(n3403) );
  NOR4XL U2394 ( .A(n3274), .B(n3234), .C(n3218), .D(A[21]), .Y(n3423) );
  MUX2IX1 U2395 ( .D0(n3424), .D1(n3425), .S(n3213), .Y(n3422) );
  NAND2X1 U2396 ( .A(n3426), .B(n3281), .Y(n3425) );
  MUX2IX1 U2397 ( .D0(A[13]), .D1(A[269]), .S(n3232), .Y(n3426) );
  NAND2X1 U2398 ( .A(n3427), .B(n3286), .Y(n3424) );
  MUX2IX1 U2399 ( .D0(A[5]), .D1(A[261]), .S(n3231), .Y(n3427) );
  MUX2IX1 U2400 ( .D0(n3428), .D1(n3429), .S(SH[7]), .Y(B[4]) );
  MUX4X1 U2401 ( .D0(n3430), .D1(n3431), .D2(n3432), .D3(n3433), .S0(SH[5]), 
        .S1(n3203), .Y(n3429) );
  MUX4X1 U2402 ( .D0(n3434), .D1(n3435), .D2(n3436), .D3(n3437), .S0(n3220), 
        .S1(n3213), .Y(n3433) );
  NOR3XL U2403 ( .A(A[252]), .B(n3271), .C(n3239), .Y(n3437) );
  NOR3XL U2404 ( .A(A[236]), .B(n3273), .C(n3239), .Y(n3436) );
  NOR3XL U2405 ( .A(A[244]), .B(n3272), .C(n3239), .Y(n3435) );
  NOR3XL U2406 ( .A(A[228]), .B(n3272), .C(n3238), .Y(n3434) );
  MUX4X1 U2407 ( .D0(n3438), .D1(n3439), .D2(n3440), .D3(n3441), .S0(n3222), 
        .S1(n3214), .Y(n3432) );
  NOR3XL U2408 ( .A(A[220]), .B(n3272), .C(n3238), .Y(n3441) );
  AOI21X1 U2409 ( .B(A[204]), .C(n3249), .A(n3260), .Y(n3440) );
  AOI21X1 U2410 ( .B(A[212]), .C(n3250), .A(n3261), .Y(n3439) );
  AOI21X1 U2411 ( .B(A[196]), .C(n3249), .A(n3260), .Y(n3438) );
  MUX4X1 U2412 ( .D0(n3442), .D1(n3443), .D2(n3444), .D3(n3445), .S0(n3221), 
        .S1(n3214), .Y(n3431) );
  NOR3XL U2413 ( .A(A[188]), .B(n3272), .C(n3238), .Y(n3445) );
  NOR3XL U2414 ( .A(A[172]), .B(n3273), .C(n3238), .Y(n3444) );
  NOR3XL U2415 ( .A(A[180]), .B(n3273), .C(n3238), .Y(n3443) );
  NOR3XL U2416 ( .A(A[164]), .B(n3272), .C(n3238), .Y(n3442) );
  MUX4X1 U2417 ( .D0(n3446), .D1(n3447), .D2(n3448), .D3(n3449), .S0(n3222), 
        .S1(n3215), .Y(n3430) );
  NOR3XL U2418 ( .A(A[156]), .B(n3273), .C(n3238), .Y(n3449) );
  NOR21XL U2419 ( .B(n3450), .A(n3278), .Y(n3448) );
  MUX2IX1 U2420 ( .D0(A[140]), .D1(A[396]), .S(n3233), .Y(n3450) );
  NOR21XL U2421 ( .B(n3451), .A(n3279), .Y(n3447) );
  MUX2IX1 U2422 ( .D0(A[148]), .D1(A[404]), .S(n3231), .Y(n3451) );
  NOR21XL U2423 ( .B(n3452), .A(n3279), .Y(n3446) );
  MUX2IX1 U2424 ( .D0(A[132]), .D1(A[388]), .S(n3233), .Y(n3452) );
  MUX4X1 U2425 ( .D0(n3453), .D1(n3454), .D2(n3455), .D3(n3456), .S0(SH[6]), 
        .S1(n3204), .Y(n3428) );
  MUX4X1 U2426 ( .D0(n3457), .D1(n3458), .D2(n3459), .D3(n3460), .S0(n3222), 
        .S1(n3215), .Y(n3456) );
  NOR3XL U2427 ( .A(n3252), .B(n3273), .C(A[364]), .Y(n3459) );
  NOR3XL U2428 ( .A(n3249), .B(n3272), .C(A[372]), .Y(n3458) );
  NOR3XL U2429 ( .A(n3252), .B(n3273), .C(A[356]), .Y(n3457) );
  MUX4X1 U2430 ( .D0(n3462), .D1(n3463), .D2(n3464), .D3(n3465), .S0(n3222), 
        .S1(n3215), .Y(n3455) );
  NOR3XL U2431 ( .A(A[60]), .B(n3265), .C(n3238), .Y(n3465) );
  NOR3XL U2432 ( .A(A[44]), .B(n3262), .C(n3238), .Y(n3464) );
  NOR3XL U2433 ( .A(A[52]), .B(n3262), .C(n3238), .Y(n3463) );
  NOR3XL U2434 ( .A(A[36]), .B(n3262), .C(n3237), .Y(n3462) );
  MUX4X1 U2435 ( .D0(n3466), .D1(n3467), .D2(n3468), .D3(n3469), .S0(n3212), 
        .S1(n3224), .Y(n3454) );
  NOR3XL U2436 ( .A(n3252), .B(n3262), .C(A[348]), .Y(n3469) );
  NOR3XL U2437 ( .A(n3252), .B(n3262), .C(A[340]), .Y(n3468) );
  NOR21XL U2438 ( .B(n3470), .A(n3279), .Y(n3467) );
  MUX2IX1 U2439 ( .D0(A[76]), .D1(A[332]), .S(n3233), .Y(n3470) );
  NOR21XL U2440 ( .B(n3471), .A(n3278), .Y(n3466) );
  MUX2IX1 U2441 ( .D0(A[68]), .D1(A[324]), .S(n3233), .Y(n3471) );
  MUX2IX1 U2442 ( .D0(n3473), .D1(n3474), .S(n3213), .Y(n3472) );
  NAND2X1 U2443 ( .A(n3475), .B(n3281), .Y(n3474) );
  MUX2IX1 U2444 ( .D0(A[12]), .D1(A[268]), .S(n3233), .Y(n3475) );
  NAND2X1 U2445 ( .A(n3476), .B(n3280), .Y(n3473) );
  MUX2IX1 U2446 ( .D0(A[4]), .D1(A[260]), .S(n3233), .Y(n3476) );
  MUX2IX1 U2447 ( .D0(n3477), .D1(n3478), .S(SH[7]), .Y(B[3]) );
  MUX4X1 U2448 ( .D0(n3479), .D1(n3480), .D2(n3481), .D3(n3482), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3478) );
  MUX4X1 U2449 ( .D0(n3483), .D1(n3484), .D2(n3485), .D3(n3486), .S0(n3223), 
        .S1(n3215), .Y(n3482) );
  NOR3XL U2450 ( .A(A[251]), .B(n3264), .C(n3237), .Y(n3486) );
  NOR3XL U2451 ( .A(A[235]), .B(n3262), .C(n3237), .Y(n3485) );
  NOR3XL U2452 ( .A(A[243]), .B(n3262), .C(n3237), .Y(n3484) );
  NOR3XL U2453 ( .A(A[227]), .B(n3263), .C(n3237), .Y(n3483) );
  MUX4X1 U2454 ( .D0(n3487), .D1(n3488), .D2(n3489), .D3(n3490), .S0(n3223), 
        .S1(n3215), .Y(n3481) );
  NOR3XL U2455 ( .A(A[219]), .B(n3262), .C(n3237), .Y(n3490) );
  AOI21X1 U2456 ( .B(A[203]), .C(n3249), .A(n3261), .Y(n3489) );
  AOI21X1 U2457 ( .B(A[211]), .C(n3249), .A(n3260), .Y(n3488) );
  AOI21X1 U2458 ( .B(A[195]), .C(n3249), .A(n3260), .Y(n3487) );
  MUX4X1 U2459 ( .D0(n3491), .D1(n3492), .D2(n3493), .D3(n3494), .S0(n3222), 
        .S1(n3214), .Y(n3480) );
  NOR3XL U2460 ( .A(A[187]), .B(n3263), .C(n3237), .Y(n3494) );
  NOR3XL U2461 ( .A(A[171]), .B(n3264), .C(n3237), .Y(n3493) );
  NOR3XL U2462 ( .A(A[179]), .B(n3263), .C(n3237), .Y(n3492) );
  NOR3XL U2463 ( .A(A[163]), .B(n3262), .C(n3237), .Y(n3491) );
  MUX4X1 U2464 ( .D0(n3495), .D1(n3496), .D2(n3497), .D3(n3498), .S0(n3223), 
        .S1(n3215), .Y(n3479) );
  NOR3XL U2465 ( .A(A[155]), .B(n3264), .C(n3255), .Y(n3498) );
  NOR21XL U2466 ( .B(n3499), .A(n3276), .Y(n3497) );
  MUX2IX1 U2467 ( .D0(A[139]), .D1(A[395]), .S(n3232), .Y(n3499) );
  NOR21XL U2468 ( .B(n3500), .A(n3275), .Y(n3496) );
  MUX2IX1 U2469 ( .D0(A[147]), .D1(A[403]), .S(n3230), .Y(n3500) );
  NOR21XL U2470 ( .B(n3501), .A(n3277), .Y(n3495) );
  MUX2IX1 U2471 ( .D0(A[131]), .D1(A[387]), .S(n3232), .Y(n3501) );
  MUX4X1 U2472 ( .D0(n3502), .D1(n3503), .D2(n3504), .D3(n3505), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3477) );
  MUX4X1 U2473 ( .D0(n3506), .D1(n3507), .D2(n3508), .D3(n3509), .S0(n3223), 
        .S1(n3215), .Y(n3505) );
  MUX2IX1 U2474 ( .D0(A[123]), .D1(A[379]), .S(n3231), .Y(n3510) );
  NOR3XL U2475 ( .A(n3250), .B(n3263), .C(A[363]), .Y(n3508) );
  NOR3XL U2476 ( .A(n3251), .B(n3263), .C(A[371]), .Y(n3507) );
  NOR3XL U2477 ( .A(n3249), .B(n3263), .C(A[355]), .Y(n3506) );
  MUX4X1 U2478 ( .D0(n3511), .D1(n3512), .D2(n3513), .D3(n3514), .S0(n3223), 
        .S1(n3215), .Y(n3504) );
  NOR3XL U2479 ( .A(A[59]), .B(n3263), .C(n3241), .Y(n3514) );
  NOR3XL U2480 ( .A(A[43]), .B(n3265), .C(n3258), .Y(n3513) );
  NOR3XL U2481 ( .A(A[51]), .B(n3264), .C(n3255), .Y(n3512) );
  NOR3XL U2482 ( .A(A[35]), .B(n3263), .C(n3254), .Y(n3511) );
  MUX4X1 U2483 ( .D0(n3515), .D1(n3516), .D2(n3517), .D3(n3518), .S0(n3212), 
        .S1(n3224), .Y(n3503) );
  NOR3XL U2484 ( .A(n3249), .B(n3263), .C(A[347]), .Y(n3518) );
  NOR3XL U2485 ( .A(n3251), .B(n3264), .C(A[339]), .Y(n3517) );
  NOR21XL U2486 ( .B(n3519), .A(n3279), .Y(n3516) );
  MUX2IX1 U2487 ( .D0(A[75]), .D1(A[331]), .S(n3230), .Y(n3519) );
  NOR21XL U2488 ( .B(n3520), .A(n3275), .Y(n3515) );
  MUX2IX1 U2489 ( .D0(A[67]), .D1(A[323]), .S(n3229), .Y(n3520) );
  MUX2X1 U2490 ( .D0(n3521), .D1(n3522), .S(n3225), .Y(n3502) );
  NOR4XL U2491 ( .A(n3273), .B(n3234), .C(SH[3]), .D(A[19]), .Y(n3522) );
  MUX2IX1 U2492 ( .D0(n3523), .D1(n3524), .S(n3213), .Y(n3521) );
  NAND2X1 U2493 ( .A(n3525), .B(n3282), .Y(n3524) );
  MUX2IX1 U2494 ( .D0(A[11]), .D1(A[267]), .S(n3228), .Y(n3525) );
  NAND2X1 U2495 ( .A(n3526), .B(n3281), .Y(n3523) );
  MUX2IX1 U2496 ( .D0(A[3]), .D1(A[259]), .S(n3227), .Y(n3526) );
  MUX2IX1 U2497 ( .D0(n3527), .D1(n3528), .S(SH[7]), .Y(B[2]) );
  MUX4X1 U2498 ( .D0(n3529), .D1(n3530), .D2(n3531), .D3(n3532), .S0(n3204), 
        .S1(n3203), .Y(n3528) );
  MUX4X1 U2499 ( .D0(n3533), .D1(n3534), .D2(n3535), .D3(n3536), .S0(n3223), 
        .S1(n3216), .Y(n3532) );
  NOR3XL U2500 ( .A(A[250]), .B(n3265), .C(n3258), .Y(n3536) );
  NOR3XL U2501 ( .A(A[234]), .B(n3264), .C(n3258), .Y(n3535) );
  NOR3XL U2502 ( .A(A[242]), .B(n3264), .C(n3258), .Y(n3534) );
  NOR3XL U2503 ( .A(A[226]), .B(n3264), .C(n3258), .Y(n3533) );
  MUX4X1 U2504 ( .D0(n3537), .D1(n3538), .D2(n3539), .D3(n3540), .S0(n3223), 
        .S1(n3216), .Y(n3531) );
  NOR3XL U2505 ( .A(A[218]), .B(n3264), .C(n3258), .Y(n3540) );
  AOI21X1 U2506 ( .B(A[202]), .C(n3252), .A(n3260), .Y(n3539) );
  AOI21X1 U2507 ( .B(A[210]), .C(n3249), .A(n3261), .Y(n3538) );
  AOI21X1 U2508 ( .B(A[194]), .C(n3243), .A(n3260), .Y(n3537) );
  MUX4X1 U2509 ( .D0(n3541), .D1(n3542), .D2(n3543), .D3(n3544), .S0(n3222), 
        .S1(n3216), .Y(n3530) );
  NOR3XL U2510 ( .A(A[186]), .B(n3264), .C(n3236), .Y(n3544) );
  NOR3XL U2511 ( .A(A[170]), .B(n3265), .C(n3195), .Y(n3543) );
  NOR3XL U2512 ( .A(A[178]), .B(n3265), .C(n3235), .Y(n3542) );
  NOR3XL U2513 ( .A(A[162]), .B(n3265), .C(n3235), .Y(n3541) );
  MUX4X1 U2514 ( .D0(n3545), .D1(n3546), .D2(n3547), .D3(n3548), .S0(n3223), 
        .S1(n3216), .Y(n3529) );
  NOR3XL U2515 ( .A(A[154]), .B(n3265), .C(n3235), .Y(n3548) );
  NOR21XL U2516 ( .B(n3549), .A(n3274), .Y(n3547) );
  MUX2IX1 U2517 ( .D0(A[138]), .D1(A[394]), .S(n3227), .Y(n3549) );
  NOR21XL U2518 ( .B(n3550), .A(n3276), .Y(n3546) );
  MUX2IX1 U2519 ( .D0(A[146]), .D1(A[402]), .S(n3229), .Y(n3550) );
  NOR21XL U2520 ( .B(n3551), .A(n3274), .Y(n3545) );
  MUX2IX1 U2521 ( .D0(A[130]), .D1(A[386]), .S(n3229), .Y(n3551) );
  MUX4X1 U2522 ( .D0(n3552), .D1(n3553), .D2(n3554), .D3(n3555), .S0(n3203), 
        .S1(n3204), .Y(n3527) );
  MUX4X1 U2523 ( .D0(n3556), .D1(n3557), .D2(n3558), .D3(n3559), .S0(n3221), 
        .S1(n3215), .Y(n3555) );
  NOR21XL U2524 ( .B(n3560), .A(n3277), .Y(n3559) );
  MUX2IX1 U2525 ( .D0(A[122]), .D1(A[378]), .S(n3230), .Y(n3560) );
  NOR3XL U2526 ( .A(n3250), .B(n3265), .C(A[362]), .Y(n3558) );
  NOR3XL U2527 ( .A(n3253), .B(n3265), .C(A[370]), .Y(n3557) );
  NOR3XL U2528 ( .A(n3251), .B(n3265), .C(A[354]), .Y(n3556) );
  MUX4X1 U2529 ( .D0(n3561), .D1(n3562), .D2(n3563), .D3(n3564), .S0(n3224), 
        .S1(n3216), .Y(n3554) );
  NOR3XL U2530 ( .A(A[58]), .B(n3266), .C(n3235), .Y(n3564) );
  NOR3XL U2531 ( .A(A[42]), .B(n3266), .C(n3235), .Y(n3563) );
  NOR3XL U2532 ( .A(A[50]), .B(n3266), .C(n3235), .Y(n3562) );
  NOR3XL U2533 ( .A(A[34]), .B(n3266), .C(n3235), .Y(n3561) );
  MUX4X1 U2534 ( .D0(n3565), .D1(n3566), .D2(n3567), .D3(n3568), .S0(n3212), 
        .S1(SH[4]), .Y(n3553) );
  NOR3XL U2535 ( .A(n3251), .B(n3266), .C(A[346]), .Y(n3568) );
  NOR3XL U2536 ( .A(n3253), .B(n3266), .C(A[338]), .Y(n3567) );
  NOR21XL U2537 ( .B(n3569), .A(n3276), .Y(n3566) );
  MUX2IX1 U2538 ( .D0(A[74]), .D1(A[330]), .S(n3232), .Y(n3569) );
  NOR21XL U2539 ( .B(n3570), .A(n3275), .Y(n3565) );
  MUX2IX1 U2540 ( .D0(A[66]), .D1(A[322]), .S(n3231), .Y(n3570) );
  MUX2X1 U2541 ( .D0(n3571), .D1(n3572), .S(SH[4]), .Y(n3552) );
  NOR4XL U2542 ( .A(n3273), .B(n3234), .C(n3218), .D(A[18]), .Y(n3572) );
  MUX2IX1 U2543 ( .D0(n3573), .D1(n3574), .S(n3212), .Y(n3571) );
  NAND2X1 U2544 ( .A(n3575), .B(n3282), .Y(n3574) );
  MUX2IX1 U2545 ( .D0(A[10]), .D1(A[266]), .S(n3233), .Y(n3575) );
  NAND2X1 U2546 ( .A(n3576), .B(n3286), .Y(n3573) );
  MUX2IX1 U2547 ( .D0(A[2]), .D1(A[258]), .S(n3232), .Y(n3576) );
  MUX4X1 U2548 ( .D0(n3582), .D1(n3583), .D2(n3584), .D3(n3585), .S0(n3224), 
        .S1(n3217), .Y(n3581) );
  NOR3XL U2549 ( .A(A[249]), .B(n3266), .C(n3235), .Y(n3585) );
  NOR3XL U2550 ( .A(A[233]), .B(n3271), .C(n3195), .Y(n3584) );
  NOR3XL U2551 ( .A(A[241]), .B(n3266), .C(n3195), .Y(n3583) );
  NOR3XL U2552 ( .A(A[225]), .B(n3266), .C(n3195), .Y(n3582) );
  MUX4X1 U2553 ( .D0(n3586), .D1(n3587), .D2(n3588), .D3(n3589), .S0(n3224), 
        .S1(n3216), .Y(n3580) );
  NOR3XL U2554 ( .A(A[217]), .B(n3266), .C(n3195), .Y(n3589) );
  NOR21XL U2555 ( .B(n3590), .A(n3275), .Y(n3588) );
  MUX2IX1 U2556 ( .D0(A[201]), .D1(A[457]), .S(n3233), .Y(n3590) );
  NOR21XL U2557 ( .B(n3591), .A(n3276), .Y(n3587) );
  MUX2IX1 U2558 ( .D0(A[209]), .D1(A[465]), .S(n3232), .Y(n3591) );
  NOR21XL U2559 ( .B(n3592), .A(n3275), .Y(n3586) );
  MUX2IX1 U2560 ( .D0(A[193]), .D1(A[449]), .S(n3233), .Y(n3592) );
  MUX4X1 U2561 ( .D0(n3593), .D1(n3594), .D2(n3595), .D3(n3596), .S0(n3222), 
        .S1(n3217), .Y(n3579) );
  NOR3XL U2562 ( .A(A[185]), .B(n3267), .C(n3241), .Y(n3596) );
  NOR3XL U2563 ( .A(A[169]), .B(n3267), .C(n3195), .Y(n3595) );
  NOR3XL U2564 ( .A(A[177]), .B(n3267), .C(n3241), .Y(n3594) );
  NOR3XL U2565 ( .A(A[161]), .B(n3267), .C(n3258), .Y(n3593) );
  MUX4X1 U2566 ( .D0(n3597), .D1(n3598), .D2(n3599), .D3(n3600), .S0(n3224), 
        .S1(n3217), .Y(n3578) );
  NOR3XL U2567 ( .A(A[153]), .B(n3267), .C(n3195), .Y(n3600) );
  NOR21XL U2568 ( .B(n3601), .A(n3276), .Y(n3599) );
  MUX2IX1 U2569 ( .D0(A[137]), .D1(A[393]), .S(n3232), .Y(n3601) );
  NOR21XL U2570 ( .B(n3602), .A(n3276), .Y(n3598) );
  MUX2IX1 U2571 ( .D0(A[145]), .D1(A[401]), .S(n3231), .Y(n3602) );
  NOR21XL U2572 ( .B(n3603), .A(n3277), .Y(n3597) );
  MUX2IX1 U2573 ( .D0(A[129]), .D1(A[385]), .S(n3232), .Y(n3603) );
  MUX4X1 U2574 ( .D0(n3604), .D1(n3605), .D2(n3606), .D3(n3607), .S0(n3203), 
        .S1(n3204), .Y(n3577) );
  MUX4X1 U2575 ( .D0(n3608), .D1(n3609), .D2(n3610), .D3(n3611), .S0(n3224), 
        .S1(n3217), .Y(n3607) );
  NOR21XL U2576 ( .B(n3612), .A(n3276), .Y(n3611) );
  MUX2IX1 U2577 ( .D0(A[121]), .D1(A[377]), .S(n3232), .Y(n3612) );
  NOR3XL U2578 ( .A(n3251), .B(n3267), .C(A[361]), .Y(n3610) );
  NOR3XL U2579 ( .A(n3251), .B(n3267), .C(A[369]), .Y(n3609) );
  NOR3XL U2580 ( .A(n3251), .B(n3267), .C(A[353]), .Y(n3608) );
  MUX4X1 U2581 ( .D0(n3613), .D1(n3614), .D2(n3615), .D3(n3616), .S0(n3224), 
        .S1(n3217), .Y(n3606) );
  NOR3XL U2582 ( .A(A[57]), .B(n3267), .C(n3255), .Y(n3616) );
  NOR3XL U2583 ( .A(A[41]), .B(n3267), .C(n3254), .Y(n3615) );
  NOR3XL U2584 ( .A(A[49]), .B(n3283), .C(n3255), .Y(n3614) );
  NOR3XL U2585 ( .A(A[33]), .B(SH[9]), .C(n3254), .Y(n3613) );
  MUX4X1 U2586 ( .D0(n3617), .D1(n3618), .D2(n3619), .D3(n3620), .S0(n3212), 
        .S1(n3225), .Y(n3605) );
  NOR3XL U2587 ( .A(n3250), .B(n3285), .C(A[345]), .Y(n3620) );
  NOR3XL U2588 ( .A(n3251), .B(SH[9]), .C(A[337]), .Y(n3619) );
  NOR21XL U2589 ( .B(n3621), .A(n3277), .Y(n3618) );
  MUX2IX1 U2590 ( .D0(A[73]), .D1(A[329]), .S(n3231), .Y(n3621) );
  NOR21XL U2591 ( .B(n3622), .A(n3278), .Y(n3617) );
  MUX2IX1 U2592 ( .D0(A[65]), .D1(A[321]), .S(n3231), .Y(n3622) );
  MUX2IX1 U2593 ( .D0(n3624), .D1(n3625), .S(n3212), .Y(n3623) );
  NAND2X1 U2594 ( .A(n3626), .B(n3286), .Y(n3625) );
  MUX2IX1 U2595 ( .D0(A[9]), .D1(A[265]), .S(n3229), .Y(n3626) );
  NAND2X1 U2596 ( .A(n3627), .B(n3280), .Y(n3624) );
  MUX2IX1 U2597 ( .D0(A[1]), .D1(A[257]), .S(n3231), .Y(n3627) );
  MUX2IX1 U2598 ( .D0(n3628), .D1(n3629), .S(SH[7]), .Y(B[0]) );
  MUX4X1 U2599 ( .D0(n3630), .D1(n3631), .D2(n3632), .D3(n3633), .S0(SH[5]), 
        .S1(n3203), .Y(n3629) );
  MUX4X1 U2600 ( .D0(n3634), .D1(n3635), .D2(n3636), .D3(n3637), .S0(n3223), 
        .S1(n3217), .Y(n3633) );
  NOR3XL U2601 ( .A(A[248]), .B(n3284), .C(n3254), .Y(n3637) );
  NOR3XL U2602 ( .A(A[232]), .B(n3284), .C(n3254), .Y(n3636) );
  NOR3XL U2603 ( .A(A[240]), .B(n3284), .C(n3254), .Y(n3635) );
  NOR3XL U2604 ( .A(A[224]), .B(n3285), .C(n3255), .Y(n3634) );
  MUX4X1 U2605 ( .D0(n3638), .D1(n3639), .D2(n3640), .D3(n3641), .S0(n3223), 
        .S1(n3217), .Y(n3632) );
  NOR3XL U2606 ( .A(A[216]), .B(n3285), .C(n3255), .Y(n3641) );
  NOR21XL U2607 ( .B(n3642), .A(n3277), .Y(n3640) );
  MUX2IX1 U2608 ( .D0(A[200]), .D1(A[456]), .S(n3230), .Y(n3642) );
  NOR21XL U2609 ( .B(n3643), .A(n3277), .Y(n3639) );
  MUX2IX1 U2610 ( .D0(A[208]), .D1(A[464]), .S(n3230), .Y(n3643) );
  NOR21XL U2611 ( .B(n3644), .A(n3278), .Y(n3638) );
  MUX2IX1 U2612 ( .D0(A[192]), .D1(A[448]), .S(n3229), .Y(n3644) );
  MUX4X1 U2613 ( .D0(n3645), .D1(n3646), .D2(n3647), .D3(n3648), .S0(n3222), 
        .S1(n3217), .Y(n3631) );
  NOR3XL U2614 ( .A(A[184]), .B(n3284), .C(n3254), .Y(n3648) );
  NOR3XL U2615 ( .A(A[168]), .B(n3283), .C(n3236), .Y(n3647) );
  NOR3XL U2616 ( .A(A[176]), .B(n3279), .C(n3236), .Y(n3646) );
  NOR3XL U2617 ( .A(A[160]), .B(n3284), .C(n3236), .Y(n3645) );
  MUX4X1 U2618 ( .D0(n3649), .D1(n3650), .D2(n3651), .D3(n3652), .S0(n3221), 
        .S1(n3217), .Y(n3630) );
  NOR3XL U2619 ( .A(A[152]), .B(n3284), .C(n3236), .Y(n3652) );
  NOR21XL U2620 ( .B(n3653), .A(n3278), .Y(n3651) );
  MUX2IX1 U2621 ( .D0(A[136]), .D1(A[392]), .S(n3228), .Y(n3653) );
  NOR21XL U2622 ( .B(n3654), .A(n3278), .Y(n3650) );
  MUX2IX1 U2623 ( .D0(A[144]), .D1(A[400]), .S(n3228), .Y(n3654) );
  NOR21XL U2624 ( .B(n3655), .A(n3278), .Y(n3649) );
  MUX2IX1 U2625 ( .D0(A[128]), .D1(A[384]), .S(n3228), .Y(n3655) );
  MUX4X1 U2626 ( .D0(n3656), .D1(n3657), .D2(n3658), .D3(n3659), .S0(SH[6]), 
        .S1(n3204), .Y(n3628) );
  MUX4X1 U2627 ( .D0(n3660), .D1(n3661), .D2(n3662), .D3(n3663), .S0(n3220), 
        .S1(n3217), .Y(n3659) );
  NOR21XL U2628 ( .B(n3664), .A(n3279), .Y(n3663) );
  MUX2IX1 U2629 ( .D0(A[120]), .D1(A[376]), .S(n3228), .Y(n3664) );
  NOR3XL U2630 ( .A(n3250), .B(n3285), .C(A[360]), .Y(n3662) );
  NOR3XL U2631 ( .A(n3250), .B(n3284), .C(A[368]), .Y(n3661) );
  NOR3XL U2632 ( .A(n3251), .B(n3283), .C(A[352]), .Y(n3660) );
  MUX4X1 U2633 ( .D0(n3665), .D1(n3666), .D2(n3667), .D3(n3668), .S0(n3220), 
        .S1(n3218), .Y(n3658) );
  NOR3XL U2634 ( .A(A[56]), .B(n3284), .C(n3236), .Y(n3668) );
  NOR3XL U2635 ( .A(A[40]), .B(n3283), .C(n3236), .Y(n3667) );
  NOR3XL U2636 ( .A(A[48]), .B(n3283), .C(n3236), .Y(n3666) );
  NOR3XL U2637 ( .A(A[32]), .B(n3268), .C(n3236), .Y(n3665) );
  MUX4X1 U2638 ( .D0(n3669), .D1(n3670), .D2(n3671), .D3(n3672), .S0(n3212), 
        .S1(n3224), .Y(n3657) );
  NOR3XL U2639 ( .A(n3249), .B(n3268), .C(A[344]), .Y(n3672) );
  NOR3XL U2640 ( .A(n3250), .B(n3268), .C(A[336]), .Y(n3671) );
  NOR21XL U2641 ( .B(n3673), .A(n3279), .Y(n3670) );
  MUX2IX1 U2642 ( .D0(A[72]), .D1(A[328]), .S(n3227), .Y(n3673) );
  NOR21XL U2643 ( .B(n3674), .A(n3279), .Y(n3669) );
  MUX2IX1 U2644 ( .D0(A[64]), .D1(A[320]), .S(n3227), .Y(n3674) );
  MUX2X1 U2645 ( .D0(n3675), .D1(n3676), .S(n3225), .Y(n3656) );
  NOR4XL U2646 ( .A(n3274), .B(n3234), .C(SH[3]), .D(A[16]), .Y(n3676) );
  MUX2IX1 U2647 ( .D0(n3677), .D1(n3678), .S(n3213), .Y(n3675) );
  NAND2X1 U2648 ( .A(n3679), .B(n3280), .Y(n3678) );
  MUX2IX1 U2649 ( .D0(A[8]), .D1(A[264]), .S(n3227), .Y(n3679) );
  NAND2X1 U2650 ( .A(n3680), .B(n3286), .Y(n3677) );
  MUX2IX1 U2651 ( .D0(A[0]), .D1(A[256]), .S(n3227), .Y(n3680) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regx_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_0 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N16, N17, N18, N19, N20, net9015, n5, n6, n7, n8, n9, n10,
         n11, n12, n1, n2, n3, n4;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9015), .TE(1'b0) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N20), .C(net9015), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N19), .C(net9015), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N18), .C(net9015), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N17), .C(net9015), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n12), .C(net9015), .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n1) );
  NOR2X1 U4 ( .A(n6), .B(n5), .Y(n8) );
  NOR2X1 U5 ( .A(n3), .B(n7), .Y(n5) );
  OAI22X1 U6 ( .A(n1), .B(n3), .C(n7), .D(n1), .Y(N20) );
  NOR2X1 U7 ( .A(n10), .B(n1), .Y(N18) );
  XNOR2XL U8 ( .A(n4), .B(n2), .Y(n10) );
  GEN2XL U9 ( .D(n8), .E(n4), .C(N17), .B(db_cnt[2]), .A(n9), .Y(N19) );
  NOR4XL U10 ( .A(db_cnt[2]), .B(n2), .C(n4), .D(n1), .Y(n9) );
  NAND3X1 U11 ( .A(db_cnt[1]), .B(db_cnt[0]), .C(db_cnt[2]), .Y(n7) );
  NOR2X1 U12 ( .A(n1), .B(db_cnt[0]), .Y(N17) );
  XNOR2XL U13 ( .A(o_dbc), .B(d_org_0_), .Y(n6) );
  AO22AXL U14 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR21XL U15 ( .B(n5), .A(n6), .Y(o_chg) );
  INVX1 U16 ( .A(db_cnt[3]), .Y(n3) );
  INVX1 U17 ( .A(db_cnt[0]), .Y(n2) );
  INVX1 U18 ( .A(db_cnt[1]), .Y(n4) );
  NAND3X1 U19 ( .A(n6), .B(n2), .C(n11), .Y(N16) );
  NOR3XL U20 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_1 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N16, N17, N18, N19, N20, net9033, n5, n6, n7, n8, n9, n10,
         n11, n12, n1, n2, n3, n4;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9033), .TE(1'b0) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N20), .C(net9033), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N19), .C(net9033), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N18), .C(net9033), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N17), .C(net9033), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n12), .C(net9033), .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n1) );
  NOR2X1 U4 ( .A(n6), .B(n5), .Y(n8) );
  NOR2X1 U5 ( .A(n3), .B(n7), .Y(n5) );
  OAI22X1 U6 ( .A(n1), .B(n3), .C(n7), .D(n1), .Y(N20) );
  NOR2X1 U7 ( .A(n10), .B(n1), .Y(N18) );
  XNOR2XL U8 ( .A(n4), .B(n2), .Y(n10) );
  GEN2XL U9 ( .D(n8), .E(n4), .C(N17), .B(db_cnt[2]), .A(n9), .Y(N19) );
  NOR4XL U10 ( .A(db_cnt[2]), .B(n2), .C(n4), .D(n1), .Y(n9) );
  NAND3X1 U11 ( .A(db_cnt[1]), .B(db_cnt[0]), .C(db_cnt[2]), .Y(n7) );
  NOR2X1 U12 ( .A(n1), .B(db_cnt[0]), .Y(N17) );
  XNOR2XL U13 ( .A(o_dbc), .B(d_org_0_), .Y(n6) );
  AO22AXL U14 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR21XL U15 ( .B(n5), .A(n6), .Y(o_chg) );
  INVX1 U16 ( .A(db_cnt[3]), .Y(n3) );
  INVX1 U17 ( .A(db_cnt[0]), .Y(n2) );
  INVX1 U18 ( .A(db_cnt[1]), .Y(n4) );
  NAND3X1 U19 ( .A(n6), .B(n2), .C(n11), .Y(N16) );
  NOR3XL U20 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_0 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_1 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_2 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_3 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_4 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_5 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_6 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_7 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module glreg_a0_7 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9051;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_7 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9051), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9051), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9051), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9051), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9051), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9051), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9051), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9051), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9051), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_8 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9069;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_8 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9069), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9069), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9069), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9069), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9069), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9069), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9069), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9069), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9069), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_9 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9087;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_9 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9087), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9087), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9087), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9087), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9087), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9087), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9087), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9087), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9087), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_1 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH7_0 ( clk, arstz, we, wdat, rdat );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we;
  wire   net9105;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9105), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9105), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9105), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9105), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9105), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9105), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9105), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9105), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_8 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module glreg_a0_10 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9123;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_10 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9123), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9123), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9123), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9123), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9123), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9123), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9123), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9123), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9123), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_11 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9141;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_11 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9141), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9141), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9141), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9141), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9141), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9141), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9141), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9141), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9141), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_12 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9159;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_12 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9159), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9159), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9159), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9159), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9159), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9159), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9159), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9159), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9159), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_13 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9177;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_13 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9177), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9177), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9177), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9177), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9177), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9177), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9177), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9177), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9177), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_14 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9195;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_14 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9195), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9195), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9195), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9195), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9195), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9195), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9195), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9195), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9195), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_0 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net9213;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9213), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9213), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9213), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9213), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9213), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9213), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9213), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_1 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net9231;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9231), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9231), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9231), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9231), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9231), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9231), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9231), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_15 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9249;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_15 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9249), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9249), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9249), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9249), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9249), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9249), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9249), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9249), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9249), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_6_00000002 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net9267;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9267), .TE(1'b0) );
  DFFSQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9267), .XS(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9267), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9267), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9267), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9267), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9267), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_2 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_a0_16 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9285;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_16 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9285), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9285), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9285), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9285), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9285), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9285), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9285), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9285), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9285), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_17 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9303;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_17 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9303), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9303), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9303), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9303), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9303), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9303), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9303), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9303), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9303), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_18 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9321;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_18 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9321), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9321), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9321), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9321), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9321), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9321), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9321), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9321), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9321), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_19 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9339;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_19 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9339), .TE(1'b0) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9339), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9339), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9339), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9339), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9339), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9339), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9339), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9339), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module cvctl_a0 ( r_cvcwr, wdat, r_sdischg, r_vcomp, r_idacsh, r_cvofsx, 
        r_cvofs, sdischg_duty, r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, 
        r_fw_pwrv, r_dac0, r_dac3, clk_100k, clk, srstz );
  input [5:0] r_cvcwr;
  input [7:0] wdat;
  output [7:0] r_sdischg;
  output [7:0] r_vcomp;
  output [7:0] r_idacsh;
  output [7:0] r_cvofsx;
  output [15:0] r_cvofs;
  input [11:0] r_fw_pwrv;
  output [10:0] r_dac0;
  output [5:0] r_dac3;
  input r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, clk_100k, clk, srstz;
  output sdischg_duty;
  wire   clk_5k, N29, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N46,
         N47, N84, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N106, N107, N108, N109, N115, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N129, N130, net9357, n81, N83, N82, N81, N80, N79,
         N78, N77, N76, N75, N74, N73, N72, N68, N67, N66, N65, N64, N63, N62,
         N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48,
         sub_62_carry_2_, sub_62_carry_3_, sub_62_carry_4_, sub_62_carry_5_,
         n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;
  wire   [4:0] div20_cnt;
  wire   [10:1] cv_code;
  wire   [4:0] sdischg_cnt;
  wire   [4:2] add_81_carry;
  wire   [4:2] add_41_carry;
  wire   [7:1] add_3_root_sub_0_root_add_46_3_carry;

  glreg_a0_25 u0_v_comp ( .clk(clk), .arstz(n8), .we(r_cvcwr[3]), .wdat(wdat), 
        .rdat(r_vcomp) );
  glreg_a0_24 u0_idac_shift ( .clk(clk), .arstz(n7), .we(r_cvcwr[4]), .wdat(
        wdat), .rdat(r_idacsh) );
  glreg_a0_23 u0_cv_ofsx ( .clk(clk), .arstz(n6), .we(r_cvcwr[5]), .wdat(wdat), 
        .rdat(r_cvofsx) );
  glreg_a0_22 u0_cvofs01 ( .clk(clk), .arstz(n5), .we(r_cvcwr[0]), .wdat(wdat), 
        .rdat(r_cvofs[7:0]) );
  glreg_a0_21 u0_cvofs23 ( .clk(clk), .arstz(n4), .we(r_cvcwr[1]), .wdat(wdat), 
        .rdat(r_cvofs[15:8]) );
  glreg_a0_20 u0_sdischg ( .clk(clk), .arstz(n2), .we(r_cvcwr[2]), .wdat(wdat), 
        .rdat(r_sdischg) );
  SNPS_CLOCK_GATE_HIGH_cvctl_a0 clk_gate_sdischg_cnt_reg ( .CLK(clk_100k), 
        .EN(N115), .ENCLK(net9357), .TE(1'b0) );
  cvctl_a0_DW01_add_0 add_62 ( .A({N99, N98, N97, N96, N95, N94}), .B({1'b0, 
        1'b0, N109, N108, N107, N106}), .CI(1'b0), .SUM(r_dac3), .CO() );
  cvctl_a0_DW01_sub_1 sub_2_root_sub_0_root_add_46_3 ( .A(r_fw_pwrv), .B({1'b0, 
        1'b0, 1'b0, 1'b0, r_idacsh}), .CI(1'b0), .DIFF({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .CO() );
  cvctl_a0_DW01_add_2 add_1_root_sub_0_root_add_46_3 ( .A({r_cvofsx[7], 
        r_cvofsx[7], r_cvofsx[7], r_cvofsx[7], r_cvofsx}), .B({1'b0, 1'b0, 
        1'b0, N68, N67, N66, N65, N64, N63, N62, N61, N60}), .CI(1'b0), .SUM({
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}), .CO() );
  cvctl_a0_DW01_add_1 add_0_root_sub_0_root_add_46_3 ( .A({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .B({N83, N82, N81, N80, N79, 
        N78, N77, N76, N75, N74, N73, N72}), .CI(1'b0), .SUM({N84, cv_code, 
        r_dac0[0]}), .CO() );
  HAD1X1 add_81_U1_1_1 ( .A(sdischg_cnt[1]), .B(sdischg_cnt[0]), .CO(
        add_81_carry[2]), .SO(N121) );
  HAD1X1 add_81_U1_1_2 ( .A(sdischg_cnt[2]), .B(add_81_carry[2]), .CO(
        add_81_carry[3]), .SO(N122) );
  HAD1X1 add_81_U1_1_3 ( .A(sdischg_cnt[3]), .B(add_81_carry[3]), .CO(
        add_81_carry[4]), .SO(N123) );
  HAD1X1 add_41_U1_1_1 ( .A(div20_cnt[1]), .B(div20_cnt[0]), .CO(
        add_41_carry[2]), .SO(N34) );
  HAD1X1 add_41_U1_1_2 ( .A(div20_cnt[2]), .B(add_41_carry[2]), .CO(
        add_41_carry[3]), .SO(N35) );
  HAD1X1 add_41_U1_1_3 ( .A(div20_cnt[3]), .B(add_41_carry[3]), .CO(
        add_41_carry[4]), .SO(N36) );
  FAD1X1 add_3_root_sub_0_root_add_46_3_U1_1 ( .A(N47), .B(r_vcomp[1]), .CI(
        add_3_root_sub_0_root_add_46_3_carry[1]), .CO(
        add_3_root_sub_0_root_add_46_3_carry[2]), .SO(N61) );
  DFFRQX1 sdischg_cnt_reg_4_ ( .D(N130), .C(net9357), .XR(n6), .Q(
        sdischg_cnt[4]) );
  DFFRQX1 sdischg_cnt_reg_0_ ( .D(N126), .C(net9357), .XR(srstz), .Q(
        sdischg_cnt[0]) );
  DFFRQX1 div20_cnt_reg_1_ ( .D(N39), .C(clk_100k), .XR(n5), .Q(div20_cnt[1])
         );
  DFFRQX1 div20_cnt_reg_3_ ( .D(N41), .C(clk_100k), .XR(n4), .Q(div20_cnt[3])
         );
  DFFRQX1 div20_cnt_reg_0_ ( .D(N38), .C(clk_100k), .XR(n8), .Q(div20_cnt[0])
         );
  DFFRQX1 div20_cnt_reg_2_ ( .D(N40), .C(clk_100k), .XR(n2), .Q(div20_cnt[2])
         );
  DFFRQX1 div20_cnt_reg_4_ ( .D(N42), .C(clk_100k), .XR(n8), .Q(div20_cnt[4])
         );
  DFFRQX1 sdischg_cnt_reg_2_ ( .D(N128), .C(net9357), .XR(n4), .Q(
        sdischg_cnt[2]) );
  DFFRQX1 sdischg_cnt_reg_3_ ( .D(N129), .C(net9357), .XR(n6), .Q(
        sdischg_cnt[3]) );
  DFFRQX1 sdischg_cnt_reg_1_ ( .D(N127), .C(net9357), .XR(srstz), .Q(
        sdischg_cnt[1]) );
  DFFRQX1 sdischg_reg ( .D(n81), .C(net9357), .XR(n7), .Q(sdischg_duty) );
  DFFRQX1 clk_5k_reg ( .D(N29), .C(clk_100k), .XR(n5), .Q(clk_5k) );
  INVX1 U3 ( .A(n37), .Y(n1) );
  INVX1 U4 ( .A(n9), .Y(n8) );
  INVX1 U5 ( .A(n9), .Y(n4) );
  INVX1 U6 ( .A(n9), .Y(n5) );
  INVX1 U7 ( .A(n9), .Y(n6) );
  INVX1 U8 ( .A(n9), .Y(n7) );
  INVX1 U9 ( .A(n9), .Y(n2) );
  INVX1 U10 ( .A(srstz), .Y(n9) );
  INVX1 U12 ( .A(r_sdischg[3]), .Y(n18) );
  INVX1 U13 ( .A(sdischg_cnt[1]), .Y(n16) );
  INVX1 U14 ( .A(r_sdischg[2]), .Y(n17) );
  INVX1 U15 ( .A(r_sdischg[4]), .Y(n19) );
  AND2X1 U16 ( .A(r_vcomp[7]), .B(add_3_root_sub_0_root_add_46_3_carry[7]), 
        .Y(N68) );
  XOR2X1 U17 ( .A(add_3_root_sub_0_root_add_46_3_carry[7]), .B(r_vcomp[7]), 
        .Y(N67) );
  XOR2X1 U18 ( .A(cv_code[6]), .B(sub_62_carry_5_), .Y(N93) );
  AND2X1 U19 ( .A(cv_code[5]), .B(sub_62_carry_4_), .Y(sub_62_carry_5_) );
  XOR2X1 U20 ( .A(sub_62_carry_4_), .B(cv_code[5]), .Y(N92) );
  AND2X1 U21 ( .A(cv_code[4]), .B(sub_62_carry_3_), .Y(sub_62_carry_4_) );
  XOR2X1 U22 ( .A(sub_62_carry_3_), .B(cv_code[4]), .Y(N91) );
  AND2X1 U23 ( .A(cv_code[3]), .B(sub_62_carry_2_), .Y(sub_62_carry_3_) );
  XOR2X1 U24 ( .A(sub_62_carry_2_), .B(cv_code[3]), .Y(N90) );
  AND2X1 U25 ( .A(cv_code[2]), .B(cv_code[1]), .Y(sub_62_carry_2_) );
  XOR2X1 U26 ( .A(cv_code[1]), .B(cv_code[2]), .Y(N89) );
  AND2X1 U27 ( .A(r_vcomp[6]), .B(add_3_root_sub_0_root_add_46_3_carry[6]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[7]) );
  XOR2X1 U28 ( .A(add_3_root_sub_0_root_add_46_3_carry[6]), .B(r_vcomp[6]), 
        .Y(N66) );
  AND2X1 U29 ( .A(r_vcomp[5]), .B(add_3_root_sub_0_root_add_46_3_carry[5]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[6]) );
  XOR2X1 U30 ( .A(add_3_root_sub_0_root_add_46_3_carry[5]), .B(r_vcomp[5]), 
        .Y(N65) );
  AND2X1 U31 ( .A(r_vcomp[4]), .B(add_3_root_sub_0_root_add_46_3_carry[4]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[5]) );
  XOR2X1 U32 ( .A(add_3_root_sub_0_root_add_46_3_carry[4]), .B(r_vcomp[4]), 
        .Y(N64) );
  AND2X1 U33 ( .A(r_vcomp[3]), .B(add_3_root_sub_0_root_add_46_3_carry[3]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[4]) );
  XOR2X1 U34 ( .A(add_3_root_sub_0_root_add_46_3_carry[3]), .B(r_vcomp[3]), 
        .Y(N63) );
  AND2X1 U35 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[3]) );
  XOR2X1 U36 ( .A(add_3_root_sub_0_root_add_46_3_carry[2]), .B(r_vcomp[2]), 
        .Y(N62) );
  AND2X1 U37 ( .A(r_vcomp[0]), .B(N46), .Y(
        add_3_root_sub_0_root_add_46_3_carry[1]) );
  XOR2X1 U38 ( .A(N46), .B(r_vcomp[0]), .Y(N60) );
  INVX1 U39 ( .A(cv_code[1]), .Y(N88) );
  INVX1 U40 ( .A(div20_cnt[0]), .Y(N33) );
  XOR2X1 U41 ( .A(add_41_carry[4]), .B(div20_cnt[4]), .Y(N37) );
  INVX1 U42 ( .A(sdischg_cnt[0]), .Y(N120) );
  XOR2X1 U43 ( .A(add_81_carry[4]), .B(sdischg_cnt[4]), .Y(N124) );
  AND2X1 U44 ( .A(sdischg_cnt[3]), .B(n18), .Y(n11) );
  OAI32X1 U45 ( .A(n17), .B(sdischg_cnt[2]), .C(n11), .D(sdischg_cnt[3]), .E(
        n18), .Y(n12) );
  AOI22BXL U46 ( .B(r_sdischg[1]), .A(sdischg_cnt[1]), .D(r_sdischg[0]), .C(
        sdischg_cnt[0]), .Y(n10) );
  AOI211X1 U47 ( .C(r_sdischg[1]), .D(n16), .A(n12), .B(n10), .Y(n15) );
  AOI21X1 U48 ( .B(sdischg_cnt[2]), .C(n17), .A(n11), .Y(n13) );
  ENOX1 U49 ( .A(n13), .B(n12), .C(n19), .D(sdischg_cnt[4]), .Y(n14) );
  OAI22X1 U50 ( .A(sdischg_cnt[4]), .B(n19), .C(n15), .D(n14), .Y(N125) );
  OR2X1 U51 ( .A(cv_code[8]), .B(N84), .Y(r_dac0[8]) );
  OR2X1 U52 ( .A(cv_code[7]), .B(n1), .Y(r_dac0[7]) );
  OR2X1 U53 ( .A(cv_code[6]), .B(N84), .Y(r_dac0[6]) );
  OR2X1 U54 ( .A(cv_code[5]), .B(n1), .Y(r_dac0[5]) );
  OR2X1 U55 ( .A(cv_code[4]), .B(n1), .Y(r_dac0[4]) );
  OR2X1 U56 ( .A(cv_code[3]), .B(n1), .Y(r_dac0[3]) );
  OR2X1 U57 ( .A(cv_code[2]), .B(n1), .Y(r_dac0[2]) );
  OR2X1 U58 ( .A(cv_code[1]), .B(n1), .Y(r_dac0[1]) );
  MUX2X1 U59 ( .D0(N125), .D1(sdischg_duty), .S(n20), .Y(n81) );
  AND2X1 U60 ( .A(N93), .B(N84), .Y(N99) );
  AND2X1 U61 ( .A(N92), .B(N84), .Y(N98) );
  AND2X1 U62 ( .A(N91), .B(N84), .Y(N97) );
  AND2X1 U63 ( .A(N90), .B(N84), .Y(N96) );
  AND2X1 U64 ( .A(N89), .B(N84), .Y(N95) );
  AND2X1 U65 ( .A(N88), .B(N84), .Y(N94) );
  NOR32XL U66 ( .B(r_hlsb_en), .C(clk_5k), .A(r_hlsb_sel), .Y(N47) );
  NOR32XL U67 ( .B(r_hlsb_sel), .C(clk_5k), .A(n21), .Y(N46) );
  NOR21XL U68 ( .B(N37), .A(n22), .Y(N42) );
  NOR21XL U69 ( .B(N36), .A(n22), .Y(N41) );
  NOR21XL U70 ( .B(N35), .A(n22), .Y(N40) );
  NOR21XL U71 ( .B(N34), .A(n22), .Y(N39) );
  NOR21XL U72 ( .B(N33), .A(n22), .Y(N38) );
  OAI221X1 U73 ( .A(n23), .B(n24), .C(n25), .D(n26), .E(r_hlsb_en), .Y(n22) );
  AOI221XL U74 ( .A(div20_cnt[3]), .B(n24), .C(div20_cnt[1]), .D(div20_cnt[0]), 
        .E(div20_cnt[2]), .Y(n25) );
  INVX1 U75 ( .A(r_hlsb_freq), .Y(n24) );
  AOI21BX1 U76 ( .C(n26), .B(n27), .A(div20_cnt[4]), .Y(n23) );
  MUX2IX1 U77 ( .D0(div20_cnt[4]), .D1(div20_cnt[3]), .S(r_hlsb_freq), .Y(n26)
         );
  AOI31X1 U78 ( .A(n28), .B(n29), .C(n30), .D(n21), .Y(N29) );
  INVX1 U79 ( .A(r_hlsb_en), .Y(n21) );
  OAI31XL U80 ( .A(n31), .B(r_hlsb_freq), .C(div20_cnt[2]), .D(div20_cnt[3]), 
        .Y(n30) );
  AO21X1 U81 ( .B(div20_cnt[0]), .C(r_hlsb_duty), .A(div20_cnt[1]), .Y(n31) );
  INVX1 U82 ( .A(div20_cnt[4]), .Y(n29) );
  OAI211X1 U83 ( .C(r_hlsb_duty), .D(n27), .A(r_hlsb_freq), .B(div20_cnt[2]), 
        .Y(n28) );
  OR2X1 U84 ( .A(div20_cnt[0]), .B(div20_cnt[1]), .Y(n27) );
  NOR21XL U85 ( .B(N124), .A(n20), .Y(N130) );
  NOR21XL U86 ( .B(N123), .A(n20), .Y(N129) );
  NOR21XL U87 ( .B(N122), .A(n20), .Y(N128) );
  NOR21XL U88 ( .B(N121), .A(n20), .Y(N127) );
  NOR21XL U89 ( .B(N120), .A(n20), .Y(N126) );
  NAND42X1 U90 ( .C(sdischg_cnt[1]), .D(sdischg_cnt[0]), .A(n20), .B(n32), .Y(
        N115) );
  NOR3XL U91 ( .A(sdischg_cnt[2]), .B(sdischg_cnt[4]), .C(sdischg_cnt[3]), .Y(
        n32) );
  NOR2X1 U92 ( .A(r_sdischg[6]), .B(r_sdischg[5]), .Y(n20) );
  AO2222XL U93 ( .A(r_cvofs[7]), .B(n33), .C(r_cvofs[15]), .D(n34), .E(
        r_cvofs[14]), .F(n35), .G(r_cvofs[6]), .H(n36), .Y(N109) );
  AO2222XL U94 ( .A(r_cvofs[2]), .B(n33), .C(r_cvofs[10]), .D(n34), .E(
        r_cvofs[13]), .F(n35), .G(r_cvofs[5]), .H(n36), .Y(N108) );
  AO2222XL U95 ( .A(r_cvofs[1]), .B(n33), .C(r_cvofs[9]), .D(n34), .E(
        r_cvofs[12]), .F(n35), .G(r_cvofs[4]), .H(n36), .Y(N107) );
  AO2222XL U96 ( .A(r_cvofs[0]), .B(n33), .C(r_cvofs[8]), .D(n34), .E(
        r_cvofs[11]), .F(n35), .G(r_cvofs[3]), .H(n36), .Y(N106) );
  NOR2X1 U97 ( .A(n33), .B(r_dac0[10]), .Y(n36) );
  OAI21BBX1 U98 ( .A(cv_code[10]), .B(cv_code[9]), .C(n37), .Y(n35) );
  NOR2X1 U99 ( .A(n38), .B(r_dac0[9]), .Y(n34) );
  NAND21X1 U100 ( .B(cv_code[9]), .A(n37), .Y(r_dac0[9]) );
  INVX1 U101 ( .A(N84), .Y(n37) );
  NOR2X1 U102 ( .A(r_dac0[10]), .B(cv_code[9]), .Y(n33) );
  INVX1 U103 ( .A(n38), .Y(r_dac0[10]) );
  NOR2X1 U104 ( .A(cv_code[10]), .B(N84), .Y(n38) );
endmodule


module cvctl_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module cvctl_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  XOR2X1 U2 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  XOR2X1 U3 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  AND2X1 U4 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U5 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U6 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  AND2X1 U7 ( .A(carry[10]), .B(A[10]), .Y(carry[11]) );
endmodule


module cvctl_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [10:1] carry;

  FAD1X1 U2_7 ( .A(A[7]), .B(n3), .CI(carry[7]), .CO(carry[8]), .SO(DIFF[7])
         );
  FAD1X1 U2_6 ( .A(A[6]), .B(n4), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n5), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n6), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n7), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n8), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n9), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  NOR2X1 U1 ( .A(A[10]), .B(carry[10]), .Y(n1) );
  XOR2X1 U2 ( .A(n1), .B(A[11]), .Y(DIFF[11]) );
  XNOR2XL U3 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2XL U4 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2XL U5 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  INVX1 U6 ( .A(B[7]), .Y(n3) );
  INVX1 U7 ( .A(B[2]), .Y(n8) );
  INVX1 U8 ( .A(B[3]), .Y(n7) );
  INVX1 U9 ( .A(B[4]), .Y(n6) );
  INVX1 U10 ( .A(B[5]), .Y(n5) );
  INVX1 U11 ( .A(B[6]), .Y(n4) );
  INVX1 U12 ( .A(B[1]), .Y(n9) );
  NAND21X1 U13 ( .B(n10), .A(n2), .Y(carry[1]) );
  INVX1 U14 ( .A(A[0]), .Y(n2) );
  OR2X1 U15 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  XNOR2XL U16 ( .A(n10), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U17 ( .A(B[0]), .Y(n10) );
  OR2X1 U18 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
endmodule


module cvctl_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [5:0] A;
  input [5:0] B;
  output [5:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [5:1] carry;

  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  INVX1 U1 ( .A(A[4]), .Y(n1) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  XOR2X1 U3 ( .A(carry[4]), .B(A[4]), .Y(SUM[4]) );
  XOR2X1 U4 ( .A(A[5]), .B(carry[5]), .Y(SUM[5]) );
  NOR21XL U5 ( .B(carry[4]), .A(n1), .Y(carry[5]) );
  XOR2X1 U6 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  NOR21XL U7 ( .B(A[0]), .A(n2), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_cvctl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_20 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9375;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_20 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9375), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9375), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9375), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9375), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9375), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9375), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9375), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9375), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9375), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_21 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9393;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_21 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9393), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9393), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9393), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9393), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9393), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9393), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9393), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9393), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9393), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_22 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9411;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_22 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9411), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9411), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9411), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9411), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9411), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9411), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9411), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9411), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9411), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_23 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9429;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_23 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9429), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9429), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9429), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9429), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9429), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9429), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9429), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9429), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9429), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_24 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9447;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_24 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9447), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9447), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9447), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9447), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9447), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9447), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9447), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9447), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9447), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_25 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9465;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_25 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9465), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9465), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9465), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9465), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9465), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9465), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9465), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9465), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9465), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcp_a0 ( dp_comp, dm_comp, id_comp, intr, tx_en, tx_dat, r_dat, r_sta, 
        r_ctl, r_msk, r_crc, r_acc, r_dpdmsta, r_wdat, r_wr, r_re, clk, srstz, 
        r_tui );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  output [7:0] r_crc;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input [7:0] r_wdat;
  input [6:0] r_wr;
  output [7:0] r_tui;
  input dp_comp, dm_comp, id_comp, r_re, clk, srstz;
  output intr, tx_en, tx_dat;
  wire   r_dm, r_dmchg, r_acc_int, r_wr_last, r_wr_other, n1, n2, n3;

  dpdmacc_a0 u0_dpdmacc ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(
        id_comp), .r_re_0(r_re), .r_wr_1(r_wr[6]), .r_wdat(r_wdat), .r_acc(
        r_acc), .r_dpdmsta(r_dpdmsta), .r_dm(r_dm), .r_dmchg(r_dmchg), .r_int(
        r_acc_int), .clk(clk), .rstz(srstz) );
  fcpegn_a0 u0_fcpegn ( .intr(intr), .tx_en(tx_en), .tx_dat(tx_dat), .r_dat(
        r_dat), .r_sta(r_sta), .r_ctl(r_ctl), .r_msk(r_msk), .r_wr(r_wr[4:0]), 
        .r_wdat(r_wdat), .ff_idn(r_dm), .ff_chg(n1), .r_acc_int(r_acc_int), 
        .clk(clk), .srstz(n2), .r_tui(r_tui) );
  fcpcrc_a0 u0_fcpcrc ( .tx_crc(r_crc), .crc_din(r_wdat), .crc_en(r_ctl[2]), 
        .crc_shfi(r_wr_other), .crc_shfl(r_wr_last), .clk(clk), .srstz(n2) );
  BUFX3 U1 ( .A(r_dmchg), .Y(n1) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(srstz), .Y(n3) );
  AND2X1 U4 ( .A(r_wr[5]), .B(r_ctl[3]), .Y(r_wr_last) );
  NOR21XL U5 ( .B(r_wr[5]), .A(r_ctl[3]), .Y(r_wr_other) );
endmodule


module fcpcrc_a0 ( tx_crc, crc_din, crc_en, crc_shfi, crc_shfl, clk, srstz );
  output [7:0] tx_crc;
  input [7:0] crc_din;
  input crc_en, crc_shfi, crc_shfl, clk, srstz;
  wire   N81, N82, N83, N84, N85, N86, N87, N88, N89, net9483, n5, n6, n8, n15,
         n22, n24, n1, n2, n3, n4, n7, n9, n10, n11, n12, n13, n14, n16, n17,
         n18, n19, n20, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48;

  SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 clk_gate_crc8_r_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net9483), .TE(1'b0) );
  DFFRQX1 crc8_r_reg_7_ ( .D(N89), .C(net9483), .XR(srstz), .Q(tx_crc[7]) );
  DFFRQX1 crc8_r_reg_6_ ( .D(N88), .C(net9483), .XR(srstz), .Q(tx_crc[6]) );
  DFFRQX1 crc8_r_reg_4_ ( .D(N86), .C(net9483), .XR(srstz), .Q(tx_crc[4]) );
  DFFRQX1 crc8_r_reg_5_ ( .D(N87), .C(net9483), .XR(srstz), .Q(tx_crc[5]) );
  DFFRQX1 crc8_r_reg_3_ ( .D(N85), .C(net9483), .XR(srstz), .Q(tx_crc[3]) );
  DFFRQX1 crc8_r_reg_2_ ( .D(N84), .C(net9483), .XR(srstz), .Q(tx_crc[2]) );
  DFFRQX1 crc8_r_reg_1_ ( .D(N83), .C(net9483), .XR(srstz), .Q(tx_crc[1]) );
  DFFRQX1 crc8_r_reg_0_ ( .D(N82), .C(net9483), .XR(srstz), .Q(tx_crc[0]) );
  XOR3X1 U3 ( .A(tx_crc[5]), .B(n34), .C(n12), .Y(n30) );
  XNOR2XL U4 ( .A(n15), .B(n24), .Y(n8) );
  INVX1 U5 ( .A(n29), .Y(n36) );
  INVX1 U6 ( .A(n15), .Y(n39) );
  XOR3X1 U7 ( .A(n4), .B(n44), .C(n28), .Y(n29) );
  XOR2X1 U8 ( .A(n26), .B(n4), .Y(n15) );
  XOR2X1 U9 ( .A(n37), .B(n36), .Y(n43) );
  XNOR2XL U10 ( .A(n22), .B(n5), .Y(n24) );
  XNOR3X1 U11 ( .A(n8), .B(n44), .C(n47), .Y(n1) );
  INVX1 U12 ( .A(n5), .Y(n20) );
  XOR3X1 U13 ( .A(crc_din[4]), .B(n34), .C(n33), .Y(n22) );
  INVX1 U14 ( .A(n37), .Y(n32) );
  XOR3X1 U15 ( .A(n16), .B(n18), .C(n2), .Y(n5) );
  XNOR2XL U16 ( .A(n10), .B(crc_din[7]), .Y(n2) );
  XOR3X1 U17 ( .A(n44), .B(n31), .C(n3), .Y(n37) );
  XNOR2XL U18 ( .A(n41), .B(n24), .Y(n3) );
  OAI22X1 U19 ( .A(n27), .B(n48), .C(n6), .D(n26), .Y(N85) );
  XOR2X1 U20 ( .A(n39), .B(n1), .Y(n27) );
  XNOR2XL U21 ( .A(n41), .B(n20), .Y(n4) );
  OAI22X1 U22 ( .A(n42), .B(n48), .C(n6), .D(n41), .Y(N88) );
  XOR3X1 U23 ( .A(n40), .B(n39), .C(n38), .Y(n42) );
  INVX1 U24 ( .A(n41), .Y(n40) );
  INVX1 U25 ( .A(n43), .Y(n38) );
  OAI22X1 U26 ( .A(n21), .B(n48), .C(n6), .D(n5), .Y(N89) );
  XOR3X1 U27 ( .A(n8), .B(n20), .C(n36), .Y(n21) );
  OAI22X1 U28 ( .A(n46), .B(n48), .C(n6), .D(n45), .Y(N87) );
  XOR3X1 U29 ( .A(n44), .B(n1), .C(n43), .Y(n46) );
  OAI22X1 U30 ( .A(n35), .B(n48), .C(n6), .D(n22), .Y(N86) );
  XOR3X1 U31 ( .A(n24), .B(n1), .C(n32), .Y(n35) );
  OAI22X1 U32 ( .A(n32), .B(n48), .C(n6), .D(n31), .Y(N83) );
  OAI22X1 U33 ( .A(n29), .B(n48), .C(n6), .D(n28), .Y(N84) );
  OAI22X1 U34 ( .A(n1), .B(n48), .C(n6), .D(n47), .Y(N82) );
  INVX1 U35 ( .A(n45), .Y(n44) );
  XOR2X1 U36 ( .A(n30), .B(crc_din[1]), .Y(n31) );
  XOR3X1 U37 ( .A(crc_din[3]), .B(n23), .C(n25), .Y(n26) );
  XOR2X1 U38 ( .A(n19), .B(crc_din[2]), .Y(n28) );
  XOR2X1 U39 ( .A(n25), .B(crc_din[0]), .Y(n47) );
  XOR2X1 U40 ( .A(n11), .B(n23), .Y(n16) );
  XOR2X1 U41 ( .A(n25), .B(n17), .Y(n33) );
  INVX1 U42 ( .A(n13), .Y(n23) );
  INVX1 U43 ( .A(n30), .Y(n17) );
  INVX1 U44 ( .A(n11), .Y(n34) );
  INVX1 U45 ( .A(n19), .Y(n18) );
  XOR3X1 U46 ( .A(n18), .B(n17), .C(n14), .Y(n41) );
  XOR3X1 U47 ( .A(tx_crc[6]), .B(crc_din[6]), .C(n13), .Y(n14) );
  NAND21X1 U48 ( .B(crc_shfl), .A(crc_en), .Y(n6) );
  NAND2X1 U49 ( .A(crc_en), .B(crc_shfl), .Y(n48) );
  OR2X1 U50 ( .A(crc_shfi), .B(n6), .Y(N81) );
  XNOR3X1 U51 ( .A(n7), .B(n18), .C(n33), .Y(n45) );
  XNOR2XL U52 ( .A(tx_crc[5]), .B(crc_din[5]), .Y(n7) );
  XOR3X1 U53 ( .A(tx_crc[5]), .B(tx_crc[0]), .C(n16), .Y(n25) );
  XOR2X1 U54 ( .A(n9), .B(tx_crc[3]), .Y(n13) );
  XOR2X1 U55 ( .A(n10), .B(tx_crc[4]), .Y(n11) );
  XOR2X1 U56 ( .A(n10), .B(tx_crc[6]), .Y(n9) );
  INVX1 U57 ( .A(tx_crc[7]), .Y(n10) );
  XNOR2XL U58 ( .A(tx_crc[6]), .B(tx_crc[1]), .Y(n12) );
  XOR3X1 U59 ( .A(tx_crc[2]), .B(tx_crc[5]), .C(n9), .Y(n19) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcpegn_a0 ( intr, tx_en, tx_dat, r_dat, r_sta, r_ctl, r_msk, r_wr, 
        r_wdat, ff_idn, ff_chg, r_acc_int, clk, srstz, r_tui );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  input [4:0] r_wr;
  input [7:0] r_wdat;
  output [7:0] r_tui;
  input ff_idn, ff_chg, r_acc_int, clk, srstz;
  output intr, tx_en, tx_dat;
  wire   N22, upd_dbuf_en, N85, N87, N88, N95, N96, N97, N98, N99, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N186, N187, N188, N189, N190, N192, adp_tx_ui_7_, adp_tx_ui_6_,
         adp_tx_ui_5_, tui_upd, N205, N219, N221, N222, N223, N224, N225, N226,
         N227, N228, N260, N261, N324, N326, N328, N331, N336, N337, N338,
         N348, N349, N356, N362, N363, N418, N419, N444, rx_trans_8_chg, N1005,
         N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015,
         N1016, N1043, net9505, net9509, net9512, net9513, net9514, net9515,
         net9516, net9517, net9520, net9523, net9528, net9533, net9538, n26,
         n27, n28, n29, n30, n31, n32, n516, n517, n525, n526, N1259, N1258,
         N1257, N1256, N1255, N1254, N1253, N1252, N168, N167, N166, N165,
         N164, N163, N162, N161, N160, N159, N116, N115, N114, N113, N112,
         N111, N110, N109, N108, N107, gt_647_B_3_, add_423_carry_5_,
         sub_423_carry_5_, add_264_A_0_, add_282_carry_7_, mult_274_2_n7,
         mult_274_2_n6, mult_274_2_n5, mult_274_2_n4, mult_274_2_n3,
         mult_274_2_n2, mult_274_n7, mult_274_n6, mult_274_n5, mult_274_n4,
         mult_274_n3, mult_274_n2, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;
  wire   [6:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;
  wire   [7:0] upd_dbuf;
  wire   [10:0] rxtx_buf;
  wire   [3:0] us_cnt;
  wire   [6:4] rx_ui_1_2;
  wire   [6:0] rx_ui_3_8;
  wire   [7:0] rx_ui_5_8;
  wire   [5:0] catch_sync;
  wire   [7:0] ui_intv_cnt;
  wire   [6:2] symb_cnt;
  wire   [15:3] catch_ping;
  wire   [12:5] ui_by_ping;
  wire   [6:0] adp_tx_1_4;
  wire   [7:0] tui_wdat;
  wire   [11:0] trans_buf;
  wire   [1:0] new_rx_sync_cnt;
  wire   [3:0] fcp_state;
  wire   [11:1] add_277_carry;
  wire   [6:1] add_264_carry;
  wire   [5:1] add_263_carry;
  wire   [14:6] add_274_2_carry;
  wire   [15:6] add_274_carry;

  glreg_8_00000000 u0_fcpctl ( .clk(clk), .arstz(n51), .we(r_wr[0]), .wdat({
        n45, n43, r_wdat[5:0]}), .rdat({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, r_ctl[4:0]}) );
  glsta_a0_0 u0_fcpsta ( .clk(clk), .arstz(n50), .rst0(1'b0), .set2({r_acc_int, 
        setsta[6:3], n525, n517, setsta[0]}), .clr1(clrsta), .rdat(r_sta), 
        .irq(r_irq) );
  glreg_a0_4 u0_fcpmsk ( .clk(clk), .arstz(n49), .we(r_wr[2]), .wdat({n45, n43, 
        r_wdat[5:0]}), .rdat(r_msk) );
  glreg_a0_3 u0_fcpdat ( .clk(clk), .arstz(n48), .we(upd_dbuf_en), .wdat(
        upd_dbuf), .rdat(r_dat) );
  glreg_a0_2 u0_fcptui ( .clk(clk), .arstz(n47), .we(tui_upd), .wdat(tui_wdat), 
        .rdat(r_tui) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 clk_gate_catch_sync_reg ( .CLK(clk), .EN(
        n526), .ENCLK(net9505), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 clk_gate_ui_intv_cnt_reg ( .CLK(clk), .EN(
        N205), .ENCLK(net9523), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 clk_gate_rxtx_buf_reg ( .CLK(clk), .EN(N22), 
        .ENCLK(net9528), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 clk_gate_fcp_state_reg ( .CLK(clk), .EN(
        N1005), .ENCLK(net9533), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 clk_gate_symb_cnt_reg ( .CLK(clk), .EN(
        N1043), .ENCLK(net9538), .TE(1'b0) );
  fcpegn_a0_DW01_inc_0 r611 ( .A({symb_cnt[6:4], n18, symb_cnt[2], n13, n21}), 
        .SUM({n26, n27, n28, n29, n30, n31, n32}) );
  fcpegn_a0_DW01_inc_1 add_283_round ( .A({1'b0, adp_tx_ui_7_, adp_tx_ui_6_, 
        adp_tx_ui_5_, r_tui[4:1]}), .SUM({adp_tx_1_4, SYNOPSYS_UNCONNECTED_4})
         );
  fcpegn_a0_DW01_inc_2 add_316_aco ( .A({N1259, N1258, N1257, N1256, N1255, 
        N1254, N1253, N1252}), .SUM({N228, N227, N226, N225, N224, N223, N222, 
        N221}) );
  FAD1X1 add_264_U1_1 ( .A(N324), .B(n12), .CI(add_264_carry[1]), .CO(
        add_264_carry[2]), .SO(rx_ui_5_8[1]) );
  FAD1X1 add_264_U1_2 ( .A(n5), .B(rx_ui_1_2[4]), .CI(add_264_carry[2]), .CO(
        add_264_carry[3]), .SO(rx_ui_5_8[2]) );
  FAD1X1 add_264_U1_3 ( .A(n12), .B(gt_647_B_3_), .CI(add_264_carry[3]), .CO(
        add_264_carry[4]), .SO(rx_ui_5_8[3]) );
  FAD1X1 add_264_U1_4 ( .A(n355), .B(rx_ui_1_2[6]), .CI(add_264_carry[4]), 
        .CO(add_264_carry[5]), .SO(rx_ui_5_8[4]) );
  FAD1X1 add_263_U1_1 ( .A(n5), .B(n11), .CI(add_263_carry[1]), .CO(
        add_263_carry[2]), .SO(rx_ui_3_8[1]) );
  FAD1X1 add_263_U1_2 ( .A(n11), .B(rx_ui_1_2[4]), .CI(add_263_carry[2]), .CO(
        add_263_carry[3]), .SO(rx_ui_3_8[2]) );
  FAD1X1 add_263_U1_3 ( .A(rx_ui_1_2[4]), .B(gt_647_B_3_), .CI(
        add_263_carry[3]), .CO(add_263_carry[4]), .SO(rx_ui_3_8[3]) );
  FAD1X1 add_263_U1_4 ( .A(gt_647_B_3_), .B(rx_ui_1_2[6]), .CI(
        add_263_carry[4]), .CO(add_263_carry[5]), .SO(rx_ui_3_8[4]) );
  FAD1X1 add_274_2_U1_6 ( .A(N160), .B(ui_intv_cnt[6]), .CI(add_274_2_carry[6]), .CO(add_274_2_carry[7]), .SO(N172) );
  FAD1X1 add_274_2_U1_7 ( .A(N161), .B(ui_intv_cnt[7]), .CI(add_274_2_carry[7]), .CO(add_274_2_carry[8]), .SO(N173) );
  HAD1X1 mult_274_2_U8 ( .A(symb_cnt[2]), .B(N159), .CO(mult_274_2_n7), .SO(
        N161) );
  FAD1X1 mult_274_2_U7 ( .A(symb_cnt[3]), .B(N160), .CI(mult_274_2_n7), .CO(
        mult_274_2_n6), .SO(N162) );
  FAD1X1 mult_274_2_U6 ( .A(symb_cnt[4]), .B(symb_cnt[2]), .CI(mult_274_2_n6), 
        .CO(mult_274_2_n5), .SO(N163) );
  FAD1X1 mult_274_2_U5 ( .A(symb_cnt[5]), .B(symb_cnt[3]), .CI(mult_274_2_n5), 
        .CO(mult_274_2_n4), .SO(N164) );
  FAD1X1 mult_274_2_U4 ( .A(symb_cnt[6]), .B(symb_cnt[4]), .CI(mult_274_2_n4), 
        .CO(mult_274_2_n3), .SO(N165) );
  HAD1X1 mult_274_2_U3 ( .A(mult_274_2_n3), .B(symb_cnt[5]), .CO(mult_274_2_n2), .SO(N166) );
  HAD1X1 mult_274_2_U2 ( .A(mult_274_2_n2), .B(symb_cnt[6]), .CO(N168), .SO(
        N167) );
  FAD1X1 add_274_U1_6 ( .A(N107), .B(ui_intv_cnt[6]), .CI(add_274_carry[6]), 
        .CO(add_274_carry[7]), .SO(N144) );
  FAD1X1 add_274_U1_7 ( .A(N108), .B(ui_intv_cnt[7]), .CI(add_274_carry[7]), 
        .CO(add_274_carry[8]), .SO(N145) );
  HAD1X1 mult_274_U29 ( .A(N95), .B(n206), .CO(mult_274_n7), .SO(N108) );
  FAD1X1 mult_274_U28 ( .A(N96), .B(N107), .CI(mult_274_n7), .CO(mult_274_n6), 
        .SO(N109) );
  FAD1X1 mult_274_U27 ( .A(N97), .B(N95), .CI(mult_274_n6), .CO(mult_274_n5), 
        .SO(N110) );
  FAD1X1 mult_274_U26 ( .A(N98), .B(N96), .CI(mult_274_n5), .CO(mult_274_n4), 
        .SO(N111) );
  FAD1X1 mult_274_U25 ( .A(N99), .B(N97), .CI(mult_274_n4), .CO(mult_274_n3), 
        .SO(N112) );
  FAD1X1 mult_274_U24 ( .A(N116), .B(N98), .CI(mult_274_n3), .CO(mult_274_n2), 
        .SO(N113) );
  FAD1X1 mult_274_U23 ( .A(N116), .B(N99), .CI(mult_274_n2), .CO(N115), .SO(
        N114) );
  DFFRQX1 rxtx_buf_reg_8_ ( .D(trans_buf[8]), .C(net9528), .XR(n52), .Q(
        rxtx_buf[8]) );
  DFFRQX1 rxtx_buf_reg_9_ ( .D(trans_buf[9]), .C(net9528), .XR(n52), .Q(
        rxtx_buf[9]) );
  DFFRQX1 rxtx_buf_reg_10_ ( .D(trans_buf[10]), .C(net9528), .XR(n52), .Q(
        rxtx_buf[10]) );
  DFFRQX1 rxtx_buf_reg_7_ ( .D(trans_buf[7]), .C(net9528), .XR(n52), .Q(
        rxtx_buf[7]) );
  DFFRQX1 rx_byte_pchk_reg ( .D(N356), .C(clk), .XR(n55), .Q(setsta[5]) );
  DFFRQX1 rxtx_buf_reg_1_ ( .D(trans_buf[1]), .C(net9528), .XR(n54), .Q(
        rxtx_buf[1]) );
  DFFRQX1 rxtx_buf_reg_2_ ( .D(trans_buf[2]), .C(net9528), .XR(n52), .Q(
        rxtx_buf[2]) );
  DFFRQX1 rxtx_buf_reg_3_ ( .D(trans_buf[3]), .C(net9528), .XR(n53), .Q(
        rxtx_buf[3]) );
  DFFRQX1 rxtx_buf_reg_5_ ( .D(trans_buf[5]), .C(net9528), .XR(n52), .Q(
        rxtx_buf[5]) );
  DFFRQX1 rxtx_buf_reg_4_ ( .D(trans_buf[4]), .C(net9528), .XR(n52), .Q(
        rxtx_buf[4]) );
  DFFRQX1 rxtx_buf_reg_6_ ( .D(trans_buf[6]), .C(net9528), .XR(n52), .Q(
        rxtx_buf[6]) );
  DFFRQX1 new_rx_sync_cnt_reg_0_ ( .D(N348), .C(clk), .XR(n47), .Q(
        new_rx_sync_cnt[0]) );
  DFFRQX1 new_rx_sync_cnt_reg_1_ ( .D(N349), .C(clk), .XR(n49), .Q(
        new_rx_sync_cnt[1]) );
  DFFRQX1 rxtx_buf_reg_0_ ( .D(trans_buf[0]), .C(net9528), .XR(n53), .Q(
        rxtx_buf[0]) );
  DFFQX1 rx_trans_8_chg_reg ( .D(n516), .C(clk), .Q(rx_trans_8_chg) );
  DFFSQX1 catch_sync_reg_5_ ( .D(n9), .C(net9505), .XS(n51), .Q(catch_sync[5])
         );
  DFFSQX1 catch_sync_reg_3_ ( .D(n17), .C(net9505), .XS(n51), .Q(catch_sync[3]) );
  DFFRQX1 catch_sync_reg_4_ ( .D(n20), .C(net9505), .XR(n53), .Q(catch_sync[4]) );
  DFFRQX1 us_cnt_reg_1_ ( .D(n506), .C(clk), .XR(n48), .Q(us_cnt[1]) );
  DFFRQX1 us_cnt_reg_0_ ( .D(N85), .C(clk), .XR(n52), .Q(us_cnt[0]) );
  DFFRQX1 us_cnt_reg_2_ ( .D(N87), .C(clk), .XR(n50), .Q(us_cnt[2]) );
  DFFRQX1 us_cnt_reg_3_ ( .D(N88), .C(clk), .XR(srstz), .Q(us_cnt[3]) );
  DFFRQX1 catch_sync_reg_1_ ( .D(n16), .C(net9505), .XR(n53), .Q(catch_sync[1]) );
  DFFRQX1 catch_sync_reg_0_ ( .D(ui_intv_cnt[0]), .C(net9505), .XR(n53), .Q(
        catch_sync[0]) );
  DFFRQX1 catch_sync_reg_2_ ( .D(ui_intv_cnt[2]), .C(net9505), .XR(n53), .Q(
        catch_sync[2]) );
  DFFRQX1 sync_length_reg_1_ ( .D(N261), .C(net9523), .XR(n54), .Q(N363) );
  DFFRQX1 ui_intv_cnt_reg_0_ ( .D(net9520), .C(net9523), .XR(n53), .Q(
        ui_intv_cnt[0]) );
  DFFRQX1 ui_intv_cnt_reg_1_ ( .D(net9517), .C(net9523), .XR(n53), .Q(
        ui_intv_cnt[1]) );
  DFFRQX1 sync_length_reg_0_ ( .D(N260), .C(net9523), .XR(n54), .Q(N362) );
  DFFRQX1 ui_intv_cnt_reg_6_ ( .D(net9512), .C(net9523), .XR(n54), .Q(
        ui_intv_cnt[6]) );
  DFFRQX1 ui_intv_cnt_reg_4_ ( .D(net9514), .C(net9523), .XR(n54), .Q(N142) );
  DFFRQX1 symb_cnt_reg_6_ ( .D(N1016), .C(net9538), .XR(n54), .Q(symb_cnt[6])
         );
  DFFRQX1 ui_intv_cnt_reg_7_ ( .D(net9509), .C(net9523), .XR(n54), .Q(
        ui_intv_cnt[7]) );
  DFFRQX1 ui_intv_cnt_reg_2_ ( .D(net9516), .C(net9523), .XR(n53), .Q(
        ui_intv_cnt[2]) );
  DFFRQX1 symb_cnt_reg_4_ ( .D(N1014), .C(net9538), .XR(n55), .Q(symb_cnt[4])
         );
  DFFRQX1 ui_intv_cnt_reg_5_ ( .D(net9513), .C(net9523), .XR(n54), .Q(
        ui_intv_cnt[5]) );
  DFFRQX1 symb_cnt_reg_5_ ( .D(N1015), .C(net9538), .XR(n55), .Q(symb_cnt[5])
         );
  DFFRQX1 ui_intv_cnt_reg_3_ ( .D(net9515), .C(net9523), .XR(n53), .Q(N141) );
  DFFRQX1 symb_cnt_reg_2_ ( .D(N1012), .C(net9538), .XR(n55), .Q(symb_cnt[2])
         );
  DFFRQX1 symb_cnt_reg_3_ ( .D(N1013), .C(net9538), .XR(n55), .Q(symb_cnt[3])
         );
  DFFRQX1 symb_cnt_reg_1_ ( .D(N1011), .C(net9538), .XR(n55), .Q(N160) );
  DFFRQX1 symb_cnt_reg_0_ ( .D(N1010), .C(net9538), .XR(n55), .Q(N159) );
  DFFSQX1 tx_dbuf_keep_empty_reg ( .D(N444), .C(clk), .XS(n52), .Q(r_ctl[7])
         );
  DFFRQX1 rxtx_buf_reg_11_ ( .D(trans_buf[11]), .C(net9528), .XR(n54), .Q(
        tx_dat) );
  DFFRQX1 fcp_state_reg_2_ ( .D(N1008), .C(net9533), .XR(n55), .Q(fcp_state[2]) );
  DFFRQX1 fcp_state_reg_3_ ( .D(N1009), .C(net9533), .XR(n54), .Q(fcp_state[3]) );
  DFFRQX1 fcp_state_reg_1_ ( .D(N1007), .C(net9533), .XR(n55), .Q(fcp_state[1]) );
  DFFRQX1 fcp_state_reg_0_ ( .D(N1006), .C(net9533), .XR(n55), .Q(fcp_state[0]) );
  OA21X1 U3 ( .B(n155), .C(n154), .A(n153), .Y(n1) );
  NOR2X1 U4 ( .A(sub_423_carry_5_), .B(rx_ui_1_2[6]), .Y(n2) );
  INVX1 U5 ( .A(n325), .Y(n3) );
  INVX1 U6 ( .A(n207), .Y(n4) );
  INVX1 U7 ( .A(n445), .Y(n5) );
  INVX1 U8 ( .A(n180), .Y(n6) );
  INVX1 U9 ( .A(n441), .Y(n7) );
  INVX1 U10 ( .A(n365), .Y(n8) );
  BUFX3 U11 ( .A(ui_intv_cnt[5]), .Y(n9) );
  INVX1 U12 ( .A(r_ctl[0]), .Y(n10) );
  MUX2IX1 U13 ( .D0(catch_sync[2]), .D1(r_tui[4]), .S(n252), .Y(N326) );
  INVX1 U14 ( .A(N326), .Y(n11) );
  INVX1 U15 ( .A(N326), .Y(n12) );
  INVX1 U16 ( .A(n208), .Y(n13) );
  INVX1 U17 ( .A(n323), .Y(n35) );
  INVX1 U18 ( .A(n35), .Y(n14) );
  NAND2X1 U19 ( .A(n188), .B(n139), .Y(n15) );
  INVX1 U20 ( .A(n247), .Y(n16) );
  INVX1 U21 ( .A(n241), .Y(n17) );
  INVX1 U22 ( .A(n210), .Y(n18) );
  BUFX3 U23 ( .A(n168), .Y(n19) );
  INVX1 U24 ( .A(n324), .Y(n20) );
  INVX1 U25 ( .A(n206), .Y(n21) );
  INVX1 U26 ( .A(n56), .Y(n51) );
  INVX1 U27 ( .A(n56), .Y(n52) );
  INVX1 U28 ( .A(n56), .Y(n53) );
  INVX1 U29 ( .A(n56), .Y(n54) );
  INVX1 U30 ( .A(n56), .Y(n55) );
  INVX1 U31 ( .A(n56), .Y(n50) );
  INVX1 U32 ( .A(n56), .Y(n48) );
  INVX1 U33 ( .A(n56), .Y(n49) );
  INVX1 U34 ( .A(n56), .Y(n47) );
  INVX1 U35 ( .A(srstz), .Y(n56) );
  INVX1 U36 ( .A(n46), .Y(n45) );
  INVX1 U37 ( .A(n44), .Y(n43) );
  INVX1 U38 ( .A(r_wdat[7]), .Y(n46) );
  INVX1 U39 ( .A(r_wdat[0]), .Y(n36) );
  INVX1 U40 ( .A(r_wdat[1]), .Y(n37) );
  INVX1 U41 ( .A(r_wdat[6]), .Y(n44) );
  INVX1 U42 ( .A(r_wdat[5]), .Y(n41) );
  INVX1 U43 ( .A(r_wdat[4]), .Y(n40) );
  INVX1 U44 ( .A(r_wdat[3]), .Y(n39) );
  INVX1 U45 ( .A(r_wdat[2]), .Y(n38) );
  INVX1 U46 ( .A(n96), .Y(n84) );
  NAND21X1 U47 ( .B(ui_by_ping[5]), .A(n253), .Y(n257) );
  INVX1 U48 ( .A(n292), .Y(n204) );
  BUFX3 U49 ( .A(tx_en), .Y(r_ctl[6]) );
  INVX1 U50 ( .A(n175), .Y(n177) );
  NAND21X1 U51 ( .B(n178), .A(n84), .Y(tx_en) );
  NAND21X1 U52 ( .B(n134), .A(n132), .Y(n96) );
  INVX1 U53 ( .A(n152), .Y(n134) );
  NAND2X1 U54 ( .A(n168), .B(n167), .Y(n292) );
  INVX1 U55 ( .A(n290), .Y(n203) );
  INVX1 U56 ( .A(n157), .Y(n198) );
  NAND21X1 U57 ( .B(n191), .A(n195), .Y(n157) );
  INVX1 U58 ( .A(n192), .Y(n190) );
  INVX1 U59 ( .A(n193), .Y(n194) );
  NAND21X1 U60 ( .B(n192), .A(n191), .Y(n193) );
  XOR2X1 U61 ( .A(sub_423_carry_5_), .B(rx_ui_1_2[6]), .Y(n22) );
  NAND21X1 U62 ( .B(n180), .A(n169), .Y(n175) );
  NAND32X1 U63 ( .B(n423), .C(n84), .A(n83), .Y(n153) );
  INVX1 U64 ( .A(n169), .Y(n176) );
  NAND21X1 U65 ( .B(n367), .A(n242), .Y(n308) );
  NAND21X1 U66 ( .B(n483), .A(n179), .Y(n102) );
  INVX1 U67 ( .A(n221), .Y(n229) );
  NAND21X1 U68 ( .B(n132), .A(n488), .Y(n111) );
  NAND2X1 U69 ( .A(n67), .B(n134), .Y(n120) );
  NAND21X1 U70 ( .B(n123), .A(n103), .Y(n116) );
  INVX1 U71 ( .A(n80), .Y(n114) );
  NAND21X1 U72 ( .B(n125), .A(n124), .Y(n80) );
  INVX1 U74 ( .A(n242), .Y(n131) );
  INVX1 U75 ( .A(n148), .Y(n150) );
  INVX1 U76 ( .A(n63), .Y(n123) );
  NAND21X1 U77 ( .B(n131), .A(n62), .Y(n63) );
  INVX1 U78 ( .A(n189), .Y(n191) );
  OAI211X1 U79 ( .C(n418), .D(n179), .A(n368), .B(n178), .Y(N1043) );
  INVX1 U80 ( .A(n185), .Y(n526) );
  NAND32X1 U81 ( .B(n181), .C(n76), .A(n75), .Y(n152) );
  NAND21X1 U82 ( .B(n62), .A(n149), .Y(n178) );
  INVX1 U83 ( .A(n133), .Y(n62) );
  NOR2X1 U84 ( .A(n75), .B(n181), .Y(n23) );
  NAND21X1 U85 ( .B(n75), .A(n59), .Y(n132) );
  NAND21X1 U86 ( .B(n164), .A(r_wr[3]), .Y(n168) );
  OAI33XL U87 ( .A(tx_en), .B(n209), .C(n292), .D(n290), .E(n143), .F(n142), 
        .Y(trans_buf[0]) );
  INVX1 U88 ( .A(n295), .Y(n143) );
  INVX1 U89 ( .A(n296), .Y(n142) );
  INVX1 U90 ( .A(n286), .Y(n289) );
  INVX1 U91 ( .A(n288), .Y(n293) );
  NAND42X1 U92 ( .C(n10), .D(n204), .A(n141), .B(n140), .Y(n290) );
  NAND21X1 U93 ( .B(n364), .A(n15), .Y(n141) );
  NAND21X1 U94 ( .B(n25), .A(n19), .Y(n140) );
  NAND43X1 U95 ( .B(n114), .C(n113), .D(n112), .A(n111), .Y(N1006) );
  INVX1 U96 ( .A(n102), .Y(n113) );
  GEN3XL U97 ( .F(n123), .G(n213), .E(n110), .D(n122), .C(n121), .B(n214), .A(
        n109), .Y(n112) );
  INVX1 U98 ( .A(n103), .Y(n110) );
  INVX1 U99 ( .A(n121), .Y(n69) );
  OAI211X1 U100 ( .C(n274), .D(tx_en), .A(n1), .B(n19), .Y(n192) );
  OA22X1 U101 ( .A(n364), .B(n19), .C(n167), .D(n25), .Y(n366) );
  AO21X1 U102 ( .B(N225), .C(n195), .A(n194), .Y(net9514) );
  AO21X1 U103 ( .B(N227), .C(n195), .A(n194), .Y(net9512) );
  NAND32X1 U104 ( .B(n184), .C(n192), .A(n189), .Y(N205) );
  INVX1 U105 ( .A(n313), .Y(n184) );
  INVX1 U106 ( .A(n156), .Y(n195) );
  NAND21X1 U107 ( .B(n313), .A(n190), .Y(n156) );
  OAI31XL U108 ( .A(n275), .B(n274), .C(n169), .D(n256), .Y(tui_upd) );
  OAI2B11X1 U109 ( .D(N221), .C(n313), .A(n190), .B(n189), .Y(net9520) );
  INVX1 U110 ( .A(n280), .Y(n201) );
  INVX1 U111 ( .A(n287), .Y(n200) );
  NAND2X1 U112 ( .A(n188), .B(n139), .Y(n167) );
  NAND21X1 U113 ( .B(n138), .A(n137), .Y(n188) );
  AOI31X1 U114 ( .A(n179), .B(n136), .C(n24), .D(n135), .Y(n137) );
  AND3X1 U115 ( .A(n369), .B(n370), .C(n148), .Y(n138) );
  AND4X1 U116 ( .A(n373), .B(n374), .C(n134), .D(n151), .Y(n135) );
  GEN2XL U117 ( .D(n249), .E(n324), .C(n248), .B(n325), .A(n326), .Y(n323) );
  AOI33X1 U118 ( .A(n433), .B(n332), .C(n96), .D(n426), .E(n425), .F(n180), 
        .Y(n97) );
  OAI221X1 U119 ( .A(n274), .B(n164), .C(n345), .D(n310), .E(n163), .Y(n343)
         );
  NAND32X1 U120 ( .B(n212), .C(n162), .A(N331), .Y(n163) );
  AO21X1 U121 ( .B(n310), .C(n185), .A(n346), .Y(n162) );
  INVX1 U122 ( .A(n389), .Y(gt_647_B_3_) );
  NAND2X1 U123 ( .A(n374), .B(n210), .Y(n368) );
  INVX1 U124 ( .A(n311), .Y(n213) );
  INVX1 U125 ( .A(n442), .Y(rx_ui_1_2[4]) );
  INVX1 U126 ( .A(n371), .Y(n136) );
  INVX1 U127 ( .A(n164), .Y(n159) );
  INVX1 U128 ( .A(n166), .Y(n196) );
  OAI211X1 U129 ( .C(n331), .D(n446), .A(n169), .B(n165), .Y(n166) );
  INVX1 U130 ( .A(n343), .Y(n165) );
  INVX1 U131 ( .A(n173), .Y(n180) );
  INVX1 U132 ( .A(n441), .Y(rx_ui_1_2[6]) );
  OAI22X1 U133 ( .A(n175), .B(n170), .C(n389), .D(n173), .Y(n388) );
  INVX1 U134 ( .A(adp_tx_ui_6_), .Y(n170) );
  NAND21X1 U135 ( .B(n158), .A(n316), .Y(n315) );
  INVX1 U136 ( .A(n484), .Y(n211) );
  NAND32X1 U137 ( .B(n75), .C(n77), .A(n76), .Y(n169) );
  NAND21X1 U138 ( .B(n370), .A(n213), .Y(n67) );
  NAND21X1 U139 ( .B(n425), .A(n180), .Y(n367) );
  NAND2X1 U140 ( .A(n132), .B(n133), .Y(n148) );
  INVX1 U141 ( .A(n331), .Y(n212) );
  INVX1 U142 ( .A(n332), .Y(n83) );
  INVX1 U143 ( .A(n149), .Y(n179) );
  INVX1 U144 ( .A(n61), .Y(n517) );
  OAI221X1 U145 ( .A(n178), .B(n83), .C(n213), .D(n96), .E(n60), .Y(n61) );
  AND3X1 U146 ( .A(n331), .B(n206), .C(tx_en), .Y(n60) );
  AOI221XL U147 ( .A(adp_tx_ui_5_), .B(n177), .C(rx_ui_1_2[4]), .D(n180), .E(
        n176), .Y(n398) );
  OAI211X1 U148 ( .C(n486), .D(n133), .A(n111), .B(n66), .Y(n129) );
  NAND43X1 U149 ( .B(n6), .C(n344), .D(n209), .A(n345), .Y(n66) );
  OA22X1 U150 ( .A(n152), .B(n72), .C(n371), .D(n132), .Y(n74) );
  INVX1 U151 ( .A(n370), .Y(n72) );
  OA21X1 U152 ( .B(n427), .C(n186), .A(n95), .Y(n98) );
  AOI32X1 U153 ( .A(n422), .B(n161), .C(n94), .D(n93), .E(n92), .Y(n95) );
  OAI22AX1 U154 ( .D(n427), .C(n186), .A(n211), .B(n158), .Y(n93) );
  INVX1 U155 ( .A(n88), .Y(n158) );
  OAI31XL U156 ( .A(n164), .B(n108), .C(n107), .D(n106), .Y(n109) );
  INVX1 U157 ( .A(n128), .Y(n106) );
  INVX1 U158 ( .A(n490), .Y(n107) );
  NAND21X1 U159 ( .B(n173), .A(ff_chg), .Y(n310) );
  NAND32X1 U160 ( .B(n77), .C(n76), .A(n75), .Y(n186) );
  NAND21X1 U161 ( .B(n274), .A(n161), .Y(n185) );
  INVX1 U162 ( .A(n422), .Y(n81) );
  INVX1 U163 ( .A(n94), .Y(n125) );
  OR3XL U164 ( .A(n209), .B(n173), .C(n275), .Y(n189) );
  OR3XL U165 ( .A(n424), .B(n149), .C(n368), .Y(n103) );
  INVX1 U166 ( .A(n424), .Y(n73) );
  INVX1 U167 ( .A(n92), .Y(n82) );
  INVX1 U168 ( .A(n160), .Y(n197) );
  NAND21X1 U169 ( .B(n159), .A(n313), .Y(n160) );
  INVX1 U170 ( .A(n79), .Y(n124) );
  NAND21X1 U171 ( .B(n209), .A(n161), .Y(n79) );
  NAND21X1 U172 ( .B(fcp_state[2]), .A(n23), .Y(n133) );
  NAND21X1 U173 ( .B(fcp_state[0]), .A(fcp_state[3]), .Y(n181) );
  NAND21X1 U174 ( .B(fcp_state[1]), .A(n59), .Y(n149) );
  INVX1 U175 ( .A(fcp_state[1]), .Y(n75) );
  INVX1 U176 ( .A(n58), .Y(n59) );
  NAND32X1 U177 ( .B(n65), .C(n57), .A(n76), .Y(n58) );
  INVX1 U178 ( .A(fcp_state[3]), .Y(n57) );
  INVX1 U179 ( .A(fcp_state[2]), .Y(n76) );
  INVX1 U180 ( .A(fcp_state[0]), .Y(n65) );
  OAI22AX1 U181 ( .D(r_dat[7]), .C(n15), .A(n168), .B(n46), .Y(n280) );
  OAI22AX1 U182 ( .D(r_dat[0]), .C(n167), .A(n168), .B(n36), .Y(n288) );
  OAI22AX1 U183 ( .D(r_dat[2]), .C(n167), .A(n168), .B(n38), .Y(n286) );
  OAI22AX1 U184 ( .D(r_dat[1]), .C(n167), .A(n168), .B(n37), .Y(n287) );
  OAI22X1 U185 ( .A(n15), .B(n144), .C(n41), .D(n168), .Y(n278) );
  INVX1 U186 ( .A(r_dat[5]), .Y(n144) );
  OAI22X1 U187 ( .A(n167), .B(n145), .C(n40), .D(n168), .Y(n281) );
  INVX1 U188 ( .A(r_dat[4]), .Y(n145) );
  OAI22X1 U189 ( .A(n15), .B(n146), .C(n44), .D(n168), .Y(n283) );
  INVX1 U190 ( .A(r_dat[6]), .Y(n146) );
  OAI22X1 U191 ( .A(n15), .B(n147), .C(n39), .D(n168), .Y(n284) );
  INVX1 U192 ( .A(r_dat[3]), .Y(n147) );
  OAI32X1 U193 ( .A(n490), .B(n19), .C(n108), .D(r_ctl[7]), .E(n64), .Y(n121)
         );
  OA22X1 U194 ( .A(n152), .B(n67), .C(n488), .D(n132), .Y(n64) );
  NAND32X1 U195 ( .B(n129), .C(n128), .A(n127), .Y(N1007) );
  AOI22X1 U196 ( .A(n485), .B(n126), .C(n125), .D(n124), .Y(n127) );
  GEN2XL U197 ( .D(n483), .E(n179), .C(n123), .B(n122), .A(n121), .Y(n126) );
  OAI211X1 U198 ( .C(r_ctl[7]), .D(n71), .A(n102), .B(n70), .Y(N1009) );
  INVX1 U199 ( .A(n116), .Y(n71) );
  AND3X1 U200 ( .A(n69), .B(n68), .C(n120), .Y(n70) );
  INVX1 U201 ( .A(n129), .Y(n68) );
  OAI211X1 U202 ( .C(n209), .D(n186), .A(n120), .B(n119), .Y(N1008) );
  AOI31X1 U203 ( .A(r_ctl[0]), .B(r_ctl[1]), .C(n118), .D(n117), .Y(n119) );
  AO21X1 U204 ( .B(n139), .C(n116), .A(n121), .Y(n118) );
  NAND43X1 U205 ( .B(n313), .C(n6), .D(n131), .A(n243), .Y(n231) );
  AOI21BBXL U206 ( .B(r_ctl[7]), .C(n517), .A(r_wr[3]), .Y(N444) );
  NAND21X1 U207 ( .B(symb_cnt[5]), .A(n205), .Y(n307) );
  NAND21X1 U208 ( .B(n100), .A(n99), .Y(n420) );
  GEN2XL U209 ( .D(n423), .E(n96), .C(n91), .B(n311), .A(n117), .Y(n100) );
  OA21X1 U210 ( .B(n209), .C(n98), .A(n97), .Y(n99) );
  OAI31XL U211 ( .A(n133), .B(symb_cnt[2]), .C(n215), .D(n149), .Y(n91) );
  OAI211X1 U212 ( .C(n311), .D(n87), .A(n86), .B(n85), .Y(n419) );
  AOI32X1 U213 ( .A(n82), .B(ff_idn), .C(n93), .D(n114), .E(n81), .Y(n86) );
  OA222X1 U214 ( .A(n18), .B(n133), .C(n74), .D(n433), .E(n149), .F(n73), .Y(
        n87) );
  OA21X1 U215 ( .B(n421), .C(n367), .A(n153), .Y(n85) );
  OAI31XL U216 ( .A(n133), .B(n18), .C(n213), .D(n101), .Y(n130) );
  INVX1 U217 ( .A(n420), .Y(n101) );
  AO22X1 U218 ( .A(symb_cnt[6]), .B(n130), .C(n26), .D(n419), .Y(N1016) );
  AO22X1 U219 ( .A(n130), .B(symb_cnt[5]), .C(n27), .D(n419), .Y(N1015) );
  AO22X1 U220 ( .A(n130), .B(symb_cnt[4]), .C(n28), .D(n419), .Y(N1014) );
  AO22X1 U221 ( .A(n130), .B(symb_cnt[2]), .C(n30), .D(n419), .Y(N1012) );
  AO22X1 U222 ( .A(n130), .B(n13), .C(n31), .D(n419), .Y(N1011) );
  AO22X1 U223 ( .A(n130), .B(n21), .C(n32), .D(n419), .Y(N1010) );
  INVX1 U224 ( .A(N159), .Y(n206) );
  INVX1 U225 ( .A(symb_cnt[4]), .Y(n205) );
  OAI21AX1 U226 ( .B(n404), .C(n405), .A(n406), .Y(n24) );
  NAND42X1 U227 ( .C(us_cnt[2]), .D(n159), .A(us_cnt[3]), .B(n328), .Y(n313)
         );
  NAND32X1 U228 ( .B(fcp_state[2]), .C(n77), .A(n75), .Y(n164) );
  INVX1 U229 ( .A(n372), .Y(n151) );
  NAND21X1 U230 ( .B(fcp_state[3]), .A(n65), .Y(n77) );
  INVX1 U231 ( .A(ui_intv_cnt[5]), .Y(n249) );
  INVX1 U232 ( .A(symb_cnt[3]), .Y(n210) );
  INVX1 U233 ( .A(symb_cnt[2]), .Y(n207) );
  INVX1 U234 ( .A(n115), .Y(n139) );
  NAND21X1 U235 ( .B(r_ctl[7]), .A(n213), .Y(n115) );
  INVX1 U236 ( .A(r_tui[5]), .Y(adp_tx_ui_5_) );
  AOI221XL U237 ( .A(adp_tx_ui_7_), .B(n177), .C(rx_ui_1_2[6]), .D(n180), .E(
        n176), .Y(n390) );
  NAND43X1 U238 ( .B(fcp_state[2]), .C(fcp_state[3]), .D(n65), .A(fcp_state[1]), .Y(n173) );
  INVX1 U239 ( .A(n224), .Y(n230) );
  OA21X1 U240 ( .B(n173), .C(r_tui[7]), .A(n175), .Y(n387) );
  INVX1 U241 ( .A(N160), .Y(n208) );
  OA22X1 U242 ( .A(n175), .B(n172), .C(n173), .D(n445), .Y(n395) );
  INVX1 U243 ( .A(r_tui[3]), .Y(n172) );
  OAI22X1 U244 ( .A(n175), .B(n171), .C(n314), .D(n173), .Y(n394) );
  INVX1 U245 ( .A(r_tui[2]), .Y(n171) );
  AND3X1 U246 ( .A(r_ctl[7]), .B(n213), .C(n188), .Y(setsta[0]) );
  OA222X1 U247 ( .A(n152), .B(n151), .C(n150), .D(n369), .E(n149), .F(n24), 
        .Y(n155) );
  GEN2XL U248 ( .D(n8), .E(n399), .C(N363), .B(n400), .A(n311), .Y(n154) );
  AOI22BXL U249 ( .B(n175), .A(r_tui[4]), .D(n173), .C(n12), .Y(n391) );
  OAI22X1 U250 ( .A(n175), .B(n174), .C(n397), .D(n173), .Y(n396) );
  INVX1 U251 ( .A(r_tui[1]), .Y(n174) );
  NAND41X1 U252 ( .D(n313), .A(n326), .B(ui_intv_cnt[6]), .C(N142), .Y(n92) );
  AO21X1 U253 ( .B(n23), .C(fcp_state[2]), .A(n176), .Y(n88) );
  NAND21X1 U254 ( .B(n105), .A(n104), .Y(n128) );
  AO21X1 U255 ( .B(n345), .C(n446), .A(n173), .Y(n104) );
  AND4X1 U256 ( .A(n21), .B(n331), .C(n161), .D(n209), .Y(n105) );
  INVX1 U257 ( .A(n90), .Y(n117) );
  NAND21X1 U258 ( .B(n89), .A(ff_idn), .Y(n90) );
  AOI32X1 U259 ( .A(n446), .B(n345), .C(n180), .D(n88), .E(n211), .Y(n89) );
  OR3XL U260 ( .A(n21), .B(n208), .C(n417), .Y(n94) );
  INVX1 U261 ( .A(ff_idn), .Y(n209) );
  XOR2X1 U262 ( .A(r_dat[7]), .B(n209), .Y(n25) );
  INVX1 U263 ( .A(n78), .Y(n161) );
  NAND43X1 U264 ( .B(fcp_state[1]), .C(fcp_state[3]), .D(fcp_state[2]), .A(
        fcp_state[0]), .Y(n78) );
  NOR32XL U265 ( .B(symb_cnt[6]), .C(n187), .A(n306), .Y(setsta[6]) );
  INVX1 U266 ( .A(n186), .Y(n187) );
  NAND5XL U267 ( .A(fcp_state[1]), .B(ff_idn), .C(n183), .D(n484), .E(n182), 
        .Y(N1005) );
  AOI221XL U268 ( .A(n316), .B(ff_chg), .C(fcp_state[2]), .D(n181), .E(n180), 
        .Y(n182) );
  INVX1 U269 ( .A(tx_en), .Y(n183) );
  INVX1 U270 ( .A(n310), .Y(n199) );
  INVX1 U271 ( .A(r_ctl[0]), .Y(n279) );
  INVX1 U272 ( .A(r_ctl[4]), .Y(n108) );
  INVX1 U273 ( .A(r_ctl[7]), .Y(n122) );
  INVX1 U274 ( .A(r_ctl[1]), .Y(n214) );
  INVX1 U275 ( .A(rxtx_buf[0]), .Y(n202) );
  BUFX3 U276 ( .A(ff_idn), .Y(r_ctl[5]) );
  AND2X1 U277 ( .A(catch_ping[15]), .B(add_277_carry[11]), .Y(ui_by_ping[12])
         );
  XOR2X1 U278 ( .A(add_277_carry[11]), .B(catch_ping[15]), .Y(ui_by_ping[11])
         );
  AND2X1 U279 ( .A(add_277_carry[10]), .B(catch_ping[14]), .Y(
        add_277_carry[11]) );
  XOR2X1 U280 ( .A(add_277_carry[10]), .B(catch_ping[14]), .Y(ui_by_ping[10])
         );
  AND2X1 U281 ( .A(add_277_carry[9]), .B(catch_ping[13]), .Y(add_277_carry[10]) );
  XOR2X1 U282 ( .A(add_277_carry[9]), .B(catch_ping[13]), .Y(ui_by_ping[9]) );
  AND2X1 U283 ( .A(add_277_carry[8]), .B(catch_ping[12]), .Y(add_277_carry[9])
         );
  XOR2X1 U284 ( .A(add_277_carry[8]), .B(catch_ping[12]), .Y(ui_by_ping[8]) );
  AND2X1 U285 ( .A(add_277_carry[7]), .B(catch_ping[11]), .Y(add_277_carry[8])
         );
  XOR2X1 U286 ( .A(add_277_carry[7]), .B(catch_ping[11]), .Y(ui_by_ping[7]) );
  AND2X1 U287 ( .A(N168), .B(add_274_2_carry[14]), .Y(N181) );
  XOR2X1 U288 ( .A(add_274_2_carry[14]), .B(N168), .Y(N180) );
  AND2X1 U289 ( .A(N167), .B(add_274_2_carry[13]), .Y(add_274_2_carry[14]) );
  XOR2X1 U290 ( .A(add_274_2_carry[13]), .B(N167), .Y(N179) );
  AND2X1 U291 ( .A(N166), .B(add_274_2_carry[12]), .Y(add_274_2_carry[13]) );
  XOR2X1 U292 ( .A(add_274_2_carry[12]), .B(N166), .Y(N178) );
  AND2X1 U293 ( .A(N165), .B(add_274_2_carry[11]), .Y(add_274_2_carry[12]) );
  XOR2X1 U294 ( .A(add_274_2_carry[11]), .B(N165), .Y(N177) );
  XOR2X1 U295 ( .A(N116), .B(add_274_carry[15]), .Y(N153) );
  AND2X1 U296 ( .A(N115), .B(add_274_carry[14]), .Y(add_274_carry[15]) );
  XOR2X1 U297 ( .A(add_274_carry[14]), .B(N115), .Y(N152) );
  AND2X1 U298 ( .A(N114), .B(add_274_carry[13]), .Y(add_274_carry[14]) );
  XOR2X1 U299 ( .A(add_274_carry[13]), .B(N114), .Y(N151) );
  AND2X1 U300 ( .A(N113), .B(add_274_carry[12]), .Y(add_274_carry[13]) );
  XOR2X1 U301 ( .A(add_274_carry[12]), .B(N113), .Y(N150) );
  AND2X1 U302 ( .A(N112), .B(add_274_carry[11]), .Y(add_274_carry[12]) );
  XOR2X1 U303 ( .A(add_274_carry[11]), .B(N112), .Y(N149) );
  XNOR2XL U304 ( .A(ui_by_ping[6]), .B(ui_by_ping[5]), .Y(N192) );
  AND2X1 U305 ( .A(add_277_carry[6]), .B(catch_ping[10]), .Y(add_277_carry[7])
         );
  XOR2X1 U306 ( .A(add_277_carry[6]), .B(catch_ping[10]), .Y(ui_by_ping[6]) );
  AND2X1 U307 ( .A(add_277_carry[5]), .B(catch_ping[9]), .Y(add_277_carry[6])
         );
  XOR2X1 U308 ( .A(add_277_carry[5]), .B(catch_ping[9]), .Y(ui_by_ping[5]) );
  AND2X1 U309 ( .A(catch_ping[8]), .B(add_277_carry[4]), .Y(add_277_carry[5])
         );
  XOR2X1 U310 ( .A(add_277_carry[4]), .B(catch_ping[8]), .Y(N190) );
  AND2X1 U311 ( .A(catch_ping[7]), .B(add_277_carry[3]), .Y(add_277_carry[4])
         );
  XOR2X1 U312 ( .A(add_277_carry[3]), .B(catch_ping[7]), .Y(N189) );
  AND2X1 U313 ( .A(catch_ping[6]), .B(add_277_carry[2]), .Y(add_277_carry[3])
         );
  XOR2X1 U314 ( .A(add_277_carry[2]), .B(catch_ping[6]), .Y(N188) );
  AND2X1 U315 ( .A(catch_ping[5]), .B(add_277_carry[1]), .Y(add_277_carry[2])
         );
  XOR2X1 U316 ( .A(add_277_carry[1]), .B(catch_ping[5]), .Y(N187) );
  AND2X1 U317 ( .A(catch_ping[3]), .B(catch_ping[4]), .Y(add_277_carry[1]) );
  XOR2X1 U318 ( .A(catch_ping[4]), .B(catch_ping[3]), .Y(N186) );
  AND2X1 U319 ( .A(N164), .B(add_274_2_carry[10]), .Y(add_274_2_carry[11]) );
  XOR2X1 U320 ( .A(add_274_2_carry[10]), .B(N164), .Y(N176) );
  AND2X1 U321 ( .A(N163), .B(add_274_2_carry[9]), .Y(add_274_2_carry[10]) );
  XOR2X1 U322 ( .A(add_274_2_carry[9]), .B(N163), .Y(N175) );
  AND2X1 U323 ( .A(N162), .B(add_274_2_carry[8]), .Y(add_274_2_carry[9]) );
  XOR2X1 U324 ( .A(add_274_2_carry[8]), .B(N162), .Y(N174) );
  AND2X1 U325 ( .A(ui_intv_cnt[5]), .B(N159), .Y(add_274_2_carry[6]) );
  XOR2X1 U326 ( .A(N159), .B(ui_intv_cnt[5]), .Y(N171) );
  AND2X1 U327 ( .A(N111), .B(add_274_carry[10]), .Y(add_274_carry[11]) );
  XOR2X1 U328 ( .A(add_274_carry[10]), .B(N111), .Y(N148) );
  AND2X1 U329 ( .A(N110), .B(add_274_carry[9]), .Y(add_274_carry[10]) );
  XOR2X1 U330 ( .A(add_274_carry[9]), .B(N110), .Y(N147) );
  AND2X1 U331 ( .A(N109), .B(add_274_carry[8]), .Y(add_274_carry[9]) );
  XOR2X1 U332 ( .A(add_274_carry[8]), .B(N109), .Y(N146) );
  AND2X1 U333 ( .A(ui_intv_cnt[5]), .B(n206), .Y(add_274_carry[6]) );
  XOR2X1 U334 ( .A(n206), .B(ui_intv_cnt[5]), .Y(N143) );
  AND2X1 U335 ( .A(n7), .B(add_264_carry[6]), .Y(rx_ui_5_8[7]) );
  XOR2X1 U336 ( .A(add_264_carry[6]), .B(n7), .Y(rx_ui_5_8[6]) );
  AND2X1 U337 ( .A(add_264_carry[5]), .B(gt_647_B_3_), .Y(add_264_carry[6]) );
  XOR2X1 U338 ( .A(add_264_carry[5]), .B(gt_647_B_3_), .Y(rx_ui_5_8[5]) );
  AND2X1 U339 ( .A(add_264_A_0_), .B(n5), .Y(add_264_carry[1]) );
  XOR2X1 U340 ( .A(add_264_A_0_), .B(n5), .Y(rx_ui_5_8[0]) );
  OR2X1 U341 ( .A(rx_ui_1_2[4]), .B(gt_647_B_3_), .Y(sub_423_carry_5_) );
  XNOR2XL U342 ( .A(n355), .B(gt_647_B_3_), .Y(N328) );
  AND2X1 U343 ( .A(rx_ui_1_2[6]), .B(add_423_carry_5_), .Y(N338) );
  XOR2X1 U344 ( .A(add_423_carry_5_), .B(rx_ui_1_2[6]), .Y(N337) );
  AND2X1 U345 ( .A(gt_647_B_3_), .B(rx_ui_1_2[4]), .Y(add_423_carry_5_) );
  XOR2X1 U346 ( .A(rx_ui_1_2[4]), .B(gt_647_B_3_), .Y(N336) );
  AND2X1 U347 ( .A(rx_ui_1_2[6]), .B(add_263_carry[5]), .Y(rx_ui_3_8[6]) );
  XOR2X1 U348 ( .A(add_263_carry[5]), .B(rx_ui_1_2[6]), .Y(rx_ui_3_8[5]) );
  AND2X1 U349 ( .A(N324), .B(n5), .Y(add_263_carry[1]) );
  XOR2X1 U350 ( .A(N324), .B(n5), .Y(rx_ui_3_8[0]) );
  AND2X1 U351 ( .A(N363), .B(N362), .Y(N419) );
  XOR2X1 U352 ( .A(N362), .B(N363), .Y(N418) );
  XNOR2XL U353 ( .A(r_tui[6]), .B(add_282_carry_7_), .Y(adp_tx_ui_7_) );
  AND2X1 U354 ( .A(r_tui[5]), .B(r_tui[6]), .Y(add_282_carry_7_) );
  XOR2X1 U355 ( .A(r_tui[5]), .B(r_tui[6]), .Y(adp_tx_ui_6_) );
  AND2X1 U356 ( .A(ui_intv_cnt[0]), .B(N219), .Y(N1252) );
  AND2X1 U357 ( .A(n16), .B(N219), .Y(N1253) );
  AND2X1 U358 ( .A(ui_intv_cnt[2]), .B(N219), .Y(N1254) );
  AND2X1 U359 ( .A(n17), .B(N219), .Y(N1255) );
  AND2X1 U360 ( .A(n20), .B(N219), .Y(N1256) );
  AND2X1 U361 ( .A(n9), .B(N219), .Y(N1257) );
  AND2X1 U362 ( .A(ui_intv_cnt[6]), .B(N219), .Y(N1258) );
  AND2X1 U363 ( .A(N219), .B(ui_intv_cnt[7]), .Y(N1259) );
  OR2X1 U364 ( .A(N160), .B(N159), .Y(n215) );
  OAI21BBX1 U365 ( .A(N159), .B(N160), .C(n215), .Y(N107) );
  OR2X1 U366 ( .A(n215), .B(n4), .Y(n216) );
  OAI21BBX1 U367 ( .A(n215), .B(symb_cnt[2]), .C(n216), .Y(N95) );
  OR2X1 U368 ( .A(n216), .B(symb_cnt[3]), .Y(n217) );
  OAI21BBX1 U369 ( .A(n216), .B(symb_cnt[3]), .C(n217), .Y(N96) );
  OR2X1 U370 ( .A(n217), .B(symb_cnt[4]), .Y(n218) );
  OAI21BBX1 U371 ( .A(n217), .B(symb_cnt[4]), .C(n218), .Y(N97) );
  XNOR2XL U372 ( .A(n218), .B(symb_cnt[5]), .Y(N98) );
  OR2X1 U373 ( .A(symb_cnt[5]), .B(n218), .Y(n219) );
  NOR3XL U374 ( .A(symb_cnt[5]), .B(symb_cnt[6]), .C(n218), .Y(N116) );
  AO21X1 U375 ( .B(n219), .C(symb_cnt[6]), .A(N116), .Y(N99) );
  NOR2X1 U376 ( .A(n22), .B(n9), .Y(n224) );
  AOI32X1 U377 ( .A(n230), .B(N336), .C(n20), .D(n9), .E(n22), .Y(n228) );
  AND2X1 U378 ( .A(n442), .B(n241), .Y(n223) );
  OAI32X1 U379 ( .A(n357), .B(n12), .C(n223), .D(n442), .E(n241), .Y(n221) );
  AOI22BXL U380 ( .B(ui_intv_cnt[1]), .A(n5), .D(ui_intv_cnt[0]), .C(N324), 
        .Y(n220) );
  AOI211X1 U381 ( .C(ui_intv_cnt[1]), .D(n445), .A(n221), .B(n220), .Y(n222)
         );
  GEN2XL U382 ( .D(n12), .E(n357), .C(n223), .B(n229), .A(n222), .Y(n225) );
  AOI211X1 U383 ( .C(N328), .D(n324), .A(n225), .B(n224), .Y(n226) );
  NOR3XL U384 ( .A(n226), .B(ui_intv_cnt[7]), .C(ui_intv_cnt[6]), .Y(n227) );
  AOI21X1 U385 ( .B(n228), .C(n227), .A(n2), .Y(N331) );
  OAI21X1 U386 ( .B(n231), .C(n232), .A(n233), .Y(upd_dbuf_en) );
  NAND4X1 U387 ( .A(n234), .B(n235), .C(n236), .D(n237), .Y(n232) );
  XNOR2XL U388 ( .A(ui_intv_cnt[2]), .B(rx_ui_5_8[2]), .Y(n237) );
  NOR2X1 U389 ( .A(n238), .B(n239), .Y(n236) );
  XNOR2XL U390 ( .A(rx_ui_5_8[0]), .B(n240), .Y(n239) );
  XNOR2XL U391 ( .A(rx_ui_5_8[3]), .B(n241), .Y(n238) );
  XNOR2XL U392 ( .A(n20), .B(rx_ui_5_8[4]), .Y(n235) );
  XNOR2XL U393 ( .A(ui_intv_cnt[7]), .B(rx_ui_5_8[7]), .Y(n234) );
  NOR3XL U394 ( .A(n244), .B(n245), .C(n246), .Y(n243) );
  XNOR2XL U395 ( .A(rx_ui_5_8[1]), .B(n247), .Y(n246) );
  XNOR2XL U396 ( .A(rx_ui_5_8[6]), .B(n248), .Y(n245) );
  XNOR2XL U397 ( .A(rx_ui_5_8[5]), .B(n249), .Y(n244) );
  MUX2X1 U398 ( .D0(n45), .D1(rxtx_buf[7]), .S(n233), .Y(upd_dbuf[7]) );
  MUX2X1 U399 ( .D0(n43), .D1(rxtx_buf[6]), .S(n233), .Y(upd_dbuf[6]) );
  MUX2X1 U400 ( .D0(r_wdat[5]), .D1(rxtx_buf[5]), .S(n233), .Y(upd_dbuf[5]) );
  MUX2X1 U401 ( .D0(r_wdat[4]), .D1(rxtx_buf[4]), .S(n233), .Y(upd_dbuf[4]) );
  MUX2X1 U402 ( .D0(r_wdat[3]), .D1(rxtx_buf[3]), .S(n233), .Y(upd_dbuf[3]) );
  INVX1 U403 ( .A(r_wr[3]), .Y(n233) );
  MUX2IX1 U404 ( .D0(n250), .D1(n38), .S(r_wr[3]), .Y(upd_dbuf[2]) );
  MUX2IX1 U405 ( .D0(n251), .D1(n37), .S(r_wr[3]), .Y(upd_dbuf[1]) );
  MUX2IX1 U406 ( .D0(n202), .D1(n36), .S(r_wr[3]), .Y(upd_dbuf[0]) );
  MUX2IX1 U407 ( .D0(n252), .D1(n46), .S(r_wr[4]), .Y(tui_wdat[7]) );
  OAI21BBX1 U408 ( .A(N192), .B(n253), .C(n254), .Y(tui_wdat[6]) );
  MUX2IX1 U409 ( .D0(n255), .D1(n43), .S(r_wr[4]), .Y(n254) );
  OAI211X1 U410 ( .C(n41), .D(n256), .A(n257), .B(n258), .Y(tui_wdat[5]) );
  OAI211X1 U411 ( .C(n40), .D(n256), .A(n259), .B(n258), .Y(tui_wdat[4]) );
  NAND2X1 U412 ( .A(N190), .B(n253), .Y(n259) );
  OAI211X1 U413 ( .C(n39), .D(n256), .A(n260), .B(n258), .Y(tui_wdat[3]) );
  NAND2X1 U414 ( .A(N189), .B(n253), .Y(n260) );
  OAI2B11X1 U415 ( .D(n253), .C(n261), .A(n258), .B(n262), .Y(tui_wdat[2]) );
  MUX2IX1 U416 ( .D0(n255), .D1(r_wdat[2]), .S(r_wr[4]), .Y(n262) );
  NAND2X1 U417 ( .A(n263), .B(n256), .Y(n258) );
  INVX1 U418 ( .A(N188), .Y(n261) );
  ENOX1 U419 ( .A(n37), .B(n256), .C(N187), .D(n253), .Y(tui_wdat[1]) );
  ENOX1 U420 ( .A(n36), .B(n256), .C(N186), .D(n253), .Y(tui_wdat[0]) );
  NOR3XL U421 ( .A(n255), .B(r_wr[4]), .C(n263), .Y(n253) );
  NAND43X1 U422 ( .B(ui_by_ping[8]), .C(ui_by_ping[9]), .D(ui_by_ping[12]), 
        .A(n264), .Y(n263) );
  AOI211X1 U423 ( .C(n265), .D(n266), .A(ui_by_ping[11]), .B(ui_by_ping[10]), 
        .Y(n264) );
  OAI21BX1 U424 ( .C(N190), .B(n267), .A(n268), .Y(n266) );
  OAI21BX1 U425 ( .C(N189), .B(n269), .A(n268), .Y(n265) );
  NAND21X1 U426 ( .B(n267), .A(ui_by_ping[5]), .Y(n268) );
  NAND2X1 U427 ( .A(ui_by_ping[7]), .B(ui_by_ping[6]), .Y(n267) );
  OAI21X1 U428 ( .B(N186), .C(N187), .A(N188), .Y(n269) );
  AND2X1 U429 ( .A(n270), .B(n271), .Y(n255) );
  NOR4XL U430 ( .A(ui_by_ping[9]), .B(ui_by_ping[8]), .C(ui_by_ping[7]), .D(
        ui_by_ping[12]), .Y(n271) );
  AOI211X1 U431 ( .C(n272), .D(ui_by_ping[6]), .A(ui_by_ping[11]), .B(
        ui_by_ping[10]), .Y(n270) );
  INVX1 U432 ( .A(n273), .Y(n272) );
  OAI31XL U433 ( .A(N189), .B(N190), .C(N188), .D(ui_by_ping[5]), .Y(n273) );
  INVX1 U434 ( .A(r_wr[4]), .Y(n256) );
  NAND2X1 U435 ( .A(n276), .B(n277), .Y(trans_buf[9]) );
  AOI22X1 U436 ( .A(n278), .B(n279), .C(rxtx_buf[8]), .D(n204), .Y(n276) );
  AO2222XL U437 ( .A(n204), .B(rxtx_buf[7]), .C(n203), .D(n280), .E(n281), .F(
        n279), .G(n282), .H(n283), .Y(trans_buf[8]) );
  AO2222XL U438 ( .A(n204), .B(rxtx_buf[6]), .C(n203), .D(n283), .E(n284), .F(
        n279), .G(n285), .H(n278), .Y(trans_buf[7]) );
  AO2222XL U439 ( .A(n204), .B(rxtx_buf[5]), .C(n203), .D(n278), .E(n286), .F(
        n279), .G(n285), .H(n281), .Y(trans_buf[6]) );
  AO2222XL U440 ( .A(n204), .B(rxtx_buf[4]), .C(n287), .D(n279), .E(n203), .F(
        n281), .G(n285), .H(n284), .Y(trans_buf[5]) );
  AO2222XL U441 ( .A(n204), .B(rxtx_buf[3]), .C(n288), .D(n279), .E(n203), .F(
        n284), .G(n285), .H(n286), .Y(trans_buf[4]) );
  OAI222XL U442 ( .A(n289), .B(n290), .C(n200), .D(n291), .E(n250), .F(n292), 
        .Y(trans_buf[3]) );
  INVX1 U443 ( .A(rxtx_buf[2]), .Y(n250) );
  OAI222XL U444 ( .A(n200), .B(n290), .C(n293), .D(n291), .E(n251), .F(n292), 
        .Y(trans_buf[2]) );
  INVX1 U445 ( .A(rxtx_buf[1]), .Y(n251) );
  OAI21X1 U446 ( .B(n202), .C(n292), .A(n294), .Y(trans_buf[1]) );
  AOI32X1 U447 ( .A(n282), .B(n295), .C(n296), .D(n203), .E(n288), .Y(n294) );
  NAND2X1 U448 ( .A(n297), .B(n277), .Y(trans_buf[11]) );
  MUX2IX1 U449 ( .D0(n285), .D1(n203), .S(n201), .Y(n277) );
  AOI22X1 U450 ( .A(n280), .B(n279), .C(rxtx_buf[10]), .D(n204), .Y(n297) );
  NAND2X1 U451 ( .A(n298), .B(n299), .Y(trans_buf[10]) );
  MUX2IX1 U452 ( .D0(n203), .D1(n282), .S(n201), .Y(n299) );
  INVX1 U453 ( .A(n291), .Y(n282) );
  NAND2X1 U454 ( .A(n285), .B(n292), .Y(n291) );
  NOR2X1 U455 ( .A(n279), .B(n203), .Y(n285) );
  AOI22X1 U456 ( .A(n283), .B(n279), .C(rxtx_buf[9]), .D(n204), .Y(n298) );
  XNOR2XL U457 ( .A(n300), .B(n301), .Y(n296) );
  XNOR2XL U458 ( .A(n302), .B(n303), .Y(n301) );
  XNOR2XL U459 ( .A(n286), .B(n280), .Y(n303) );
  XNOR2XL U460 ( .A(n287), .B(n288), .Y(n302) );
  XNOR2XL U461 ( .A(n304), .B(n305), .Y(n300) );
  XNOR2XL U462 ( .A(n283), .B(n278), .Y(n305) );
  XNOR2XL U463 ( .A(n284), .B(n281), .Y(n304) );
  NAND3X1 U464 ( .A(ff_chg), .B(n307), .C(ff_idn), .Y(n306) );
  INVX1 U465 ( .A(n308), .Y(setsta[4]) );
  NOR32XL U466 ( .B(new_rx_sync_cnt[1]), .C(n309), .A(n310), .Y(setsta[3]) );
  AOI21BBXL U467 ( .B(us_cnt[1]), .C(us_cnt[0]), .A(n312), .Y(n506) );
  AND2X1 U468 ( .A(N222), .B(n198), .Y(net9517) );
  AND2X1 U469 ( .A(N223), .B(n198), .Y(net9516) );
  AND2X1 U470 ( .A(N224), .B(n198), .Y(net9515) );
  AND2X1 U471 ( .A(N226), .B(n198), .Y(net9513) );
  AND2X1 U472 ( .A(N228), .B(n198), .Y(net9509) );
  INVX1 U473 ( .A(n314), .Y(N324) );
  NOR4XL U474 ( .A(n211), .B(n315), .C(n274), .D(n209), .Y(n525) );
  MUX2IX1 U475 ( .D0(n317), .D1(ff_chg), .S(rx_trans_8_chg), .Y(n516) );
  NAND2X1 U476 ( .A(n199), .B(n242), .Y(n317) );
  NAND4X1 U477 ( .A(n318), .B(n319), .C(n320), .D(n321), .Y(intr) );
  AOI22X1 U478 ( .A(r_msk[0]), .B(r_irq[0]), .C(r_msk[1]), .D(r_irq[1]), .Y(
        n321) );
  AOI22X1 U479 ( .A(r_msk[2]), .B(r_irq[2]), .C(r_msk[3]), .D(r_irq[3]), .Y(
        n320) );
  AOI22X1 U480 ( .A(r_msk[4]), .B(r_irq[4]), .C(r_msk[5]), .D(r_irq[5]), .Y(
        n319) );
  AOI22X1 U481 ( .A(r_msk[6]), .B(r_irq[6]), .C(r_msk[7]), .D(r_irq[7]), .Y(
        n318) );
  NOR2X1 U482 ( .A(n46), .B(n322), .Y(clrsta[7]) );
  NOR2X1 U483 ( .A(n44), .B(n322), .Y(clrsta[6]) );
  NOR2X1 U484 ( .A(n41), .B(n322), .Y(clrsta[5]) );
  NOR2X1 U485 ( .A(n40), .B(n322), .Y(clrsta[4]) );
  NOR2X1 U486 ( .A(n39), .B(n322), .Y(clrsta[3]) );
  NOR2X1 U487 ( .A(n38), .B(n322), .Y(clrsta[2]) );
  NOR2X1 U488 ( .A(n37), .B(n322), .Y(clrsta[1]) );
  NOR2X1 U489 ( .A(n36), .B(n322), .Y(clrsta[0]) );
  INVX1 U490 ( .A(r_wr[1]), .Y(n322) );
  MUX2X1 U491 ( .D0(N147), .D1(N175), .S(n14), .Y(catch_ping[9]) );
  MUX2X1 U492 ( .D0(N146), .D1(N174), .S(n14), .Y(catch_ping[8]) );
  MUX2X1 U493 ( .D0(N145), .D1(N173), .S(n14), .Y(catch_ping[7]) );
  MUX2X1 U494 ( .D0(N144), .D1(N172), .S(n14), .Y(catch_ping[6]) );
  MUX2X1 U495 ( .D0(N143), .D1(N171), .S(n323), .Y(catch_ping[5]) );
  MUX2X1 U496 ( .D0(N142), .D1(N142), .S(n323), .Y(catch_ping[4]) );
  MUX2X1 U497 ( .D0(N141), .D1(N141), .S(n323), .Y(catch_ping[3]) );
  MUX2X1 U498 ( .D0(N153), .D1(N181), .S(n14), .Y(catch_ping[15]) );
  MUX2X1 U499 ( .D0(N152), .D1(N180), .S(n14), .Y(catch_ping[14]) );
  MUX2X1 U500 ( .D0(N151), .D1(N179), .S(n14), .Y(catch_ping[13]) );
  MUX2X1 U501 ( .D0(N150), .D1(N178), .S(n14), .Y(catch_ping[12]) );
  MUX2X1 U502 ( .D0(N149), .D1(N177), .S(n14), .Y(catch_ping[11]) );
  MUX2X1 U503 ( .D0(N148), .D1(N176), .S(n14), .Y(catch_ping[10]) );
  MUX2IX1 U504 ( .D0(n327), .D1(n312), .S(us_cnt[3]), .Y(N88) );
  NAND3X1 U505 ( .A(n197), .B(n328), .C(us_cnt[2]), .Y(n327) );
  MUX2IX1 U506 ( .D0(n329), .D1(n312), .S(us_cnt[2]), .Y(N87) );
  NAND2X1 U507 ( .A(n197), .B(n330), .Y(n312) );
  NAND2X1 U508 ( .A(n197), .B(n328), .Y(n329) );
  NOR21XL U509 ( .B(n197), .A(us_cnt[0]), .Y(N85) );
  NOR2X1 U510 ( .A(n308), .B(n333), .Y(N356) );
  XNOR2XL U511 ( .A(rxtx_buf[7]), .B(n334), .Y(n333) );
  XNOR2XL U512 ( .A(n335), .B(n336), .Y(n334) );
  XNOR2XL U513 ( .A(n337), .B(n338), .Y(n336) );
  XNOR2XL U514 ( .A(rxtx_buf[6]), .B(rxtx_buf[5]), .Y(n338) );
  XNOR2XL U515 ( .A(rxtx_buf[4]), .B(rxtx_buf[3]), .Y(n337) );
  XNOR2XL U516 ( .A(n339), .B(n340), .Y(n335) );
  XNOR2XL U517 ( .A(rxtx_buf[2]), .B(rxtx_buf[1]), .Y(n340) );
  XNOR2XL U518 ( .A(rxtx_buf[0]), .B(ff_idn), .Y(n339) );
  MUX2IX1 U519 ( .D0(n341), .D1(n342), .S(new_rx_sync_cnt[1]), .Y(N349) );
  AOI21X1 U520 ( .B(n343), .C(n309), .A(n196), .Y(n342) );
  NAND2X1 U521 ( .A(new_rx_sync_cnt[0]), .B(n343), .Y(n341) );
  MUX2X1 U522 ( .D0(n196), .D1(n343), .S(n309), .Y(N348) );
  INVX1 U523 ( .A(new_rx_sync_cnt[0]), .Y(n309) );
  OAI2B11X1 U524 ( .D(n347), .C(n348), .A(n325), .B(n349), .Y(n346) );
  AOI32X1 U525 ( .A(n350), .B(n347), .C(n351), .D(ui_intv_cnt[6]), .E(n352), 
        .Y(n349) );
  INVX1 U526 ( .A(N338), .Y(n352) );
  AOI22AXL U527 ( .A(N336), .B(n324), .D(n353), .C(n354), .Y(n351) );
  NAND2X1 U528 ( .A(n17), .B(n355), .Y(n354) );
  OAI31XL U529 ( .A(n356), .B(n12), .C(n357), .D(n358), .Y(n353) );
  INVX1 U530 ( .A(n359), .Y(n358) );
  AOI211X1 U531 ( .C(n12), .D(n357), .A(n360), .B(n356), .Y(n359) );
  AOI22AXL U532 ( .A(n361), .B(ui_intv_cnt[0]), .D(n5), .C(ui_intv_cnt[1]), 
        .Y(n360) );
  AOI21X1 U533 ( .B(n5), .C(n247), .A(N324), .Y(n361) );
  NOR2X1 U534 ( .A(n355), .B(N141), .Y(n356) );
  INVX1 U535 ( .A(n442), .Y(n355) );
  AOI32X1 U536 ( .A(n350), .B(N328), .C(N142), .D(ui_intv_cnt[5]), .E(n362), 
        .Y(n348) );
  INVX1 U537 ( .A(N337), .Y(n362) );
  NAND2X1 U538 ( .A(N337), .B(n249), .Y(n350) );
  NAND2X1 U539 ( .A(N338), .B(n248), .Y(n347) );
  OAI21X1 U540 ( .B(n363), .C(n292), .A(n290), .Y(N261) );
  OAI22X1 U541 ( .A(n365), .B(n292), .C(n366), .D(n279), .Y(N260) );
  XNOR2XL U542 ( .A(n45), .B(ff_idn), .Y(n364) );
  OAI211X1 U543 ( .C(n367), .D(n368), .A(n204), .B(n1), .Y(N22) );
  AOI211X1 U544 ( .C(n8), .D(n21), .A(n375), .B(n376), .Y(n373) );
  INVX1 U545 ( .A(n377), .Y(n369) );
  NAND4X1 U546 ( .A(n378), .B(n379), .C(n380), .D(n381), .Y(N219) );
  NOR4XL U547 ( .A(n382), .B(n383), .C(n384), .D(n385), .Y(n381) );
  XNOR2XL U548 ( .A(ui_intv_cnt[0]), .B(n386), .Y(n385) );
  NAND21X1 U549 ( .B(n387), .A(r_tui[0]), .Y(n386) );
  XNOR2XL U550 ( .A(n388), .B(n248), .Y(n384) );
  XNOR2XL U551 ( .A(ui_intv_cnt[7]), .B(n390), .Y(n383) );
  XNOR2XL U552 ( .A(N142), .B(n391), .Y(n382) );
  NOR2X1 U553 ( .A(n392), .B(n393), .Y(n380) );
  XNOR2XL U554 ( .A(n394), .B(n357), .Y(n393) );
  XNOR2XL U555 ( .A(N141), .B(n395), .Y(n392) );
  XNOR2XL U556 ( .A(ui_intv_cnt[1]), .B(n396), .Y(n379) );
  XNOR2XL U557 ( .A(n398), .B(n249), .Y(n378) );
  OAI31XL U558 ( .A(n401), .B(n402), .C(n403), .D(n368), .Y(n377) );
  AOI21X1 U559 ( .B(N362), .C(n399), .A(N363), .Y(n403) );
  AOI21X1 U560 ( .B(n8), .C(n206), .A(n208), .Y(n402) );
  AOI21X1 U561 ( .B(n407), .C(symb_cnt[2]), .A(symb_cnt[3]), .Y(n405) );
  AOI211X1 U562 ( .C(n408), .D(n409), .A(n410), .B(n411), .Y(n404) );
  OAI22X1 U563 ( .A(n407), .B(n207), .C(n407), .D(n208), .Y(n410) );
  NAND2X1 U564 ( .A(n365), .B(n206), .Y(n409) );
  OAI2B11X1 U565 ( .D(N419), .C(n401), .A(n412), .B(n368), .Y(n372) );
  NAND42X1 U566 ( .C(n413), .D(n414), .A(n415), .B(n416), .Y(n412) );
  NOR2X1 U567 ( .A(n376), .B(n375), .Y(n416) );
  NOR2X1 U568 ( .A(n208), .B(N418), .Y(n375) );
  NOR2X1 U569 ( .A(n207), .B(N419), .Y(n376) );
  OAI21X1 U570 ( .B(N159), .C(n8), .A(N160), .Y(n415) );
  AOI21X1 U571 ( .B(n206), .C(n365), .A(N418), .Y(n413) );
  OAI31XL U572 ( .A(n417), .B(n21), .C(n365), .D(n212), .Y(n400) );
  INVX1 U573 ( .A(N362), .Y(n365) );
  AOI21X1 U574 ( .B(symb_cnt[3]), .C(n13), .A(n316), .Y(n275) );
  AO22X1 U575 ( .A(n18), .B(n420), .C(n29), .D(n419), .Y(N1013) );
  INVX1 U576 ( .A(n426), .Y(n421) );
  NOR43XL U577 ( .B(n247), .C(n357), .D(n428), .A(ui_intv_cnt[0]), .Y(n326) );
  NOR3XL U578 ( .A(N141), .B(n3), .C(ui_intv_cnt[5]), .Y(n428) );
  NAND4X1 U579 ( .A(N142), .B(ui_intv_cnt[2]), .C(n429), .D(n430), .Y(n422) );
  NOR4XL U580 ( .A(ui_intv_cnt[7]), .B(ui_intv_cnt[6]), .C(ui_intv_cnt[1]), 
        .D(ui_intv_cnt[0]), .Y(n430) );
  NOR2X1 U581 ( .A(n313), .B(n431), .Y(n429) );
  XNOR2XL U582 ( .A(ui_intv_cnt[5]), .B(n241), .Y(n431) );
  NAND3X1 U583 ( .A(symb_cnt[6]), .B(n432), .C(symb_cnt[5]), .Y(n427) );
  NAND3X1 U584 ( .A(n210), .B(n205), .C(n207), .Y(n432) );
  NAND4X1 U585 ( .A(n434), .B(n435), .C(n436), .D(n437), .Y(n425) );
  NOR4XL U586 ( .A(n313), .B(n438), .C(n439), .D(n440), .Y(n437) );
  XNOR2XL U587 ( .A(ui_intv_cnt[6]), .B(n441), .Y(n440) );
  XNOR2XL U588 ( .A(N142), .B(n442), .Y(n439) );
  XNOR2XL U589 ( .A(add_264_A_0_), .B(n240), .Y(n438) );
  INVX1 U590 ( .A(n397), .Y(add_264_A_0_) );
  NAND2X1 U591 ( .A(r_tui[1]), .B(n252), .Y(n397) );
  NOR3XL U592 ( .A(n443), .B(ui_intv_cnt[7]), .C(n444), .Y(n436) );
  XNOR2XL U593 ( .A(ui_intv_cnt[1]), .B(n314), .Y(n444) );
  MUX2IX1 U594 ( .D0(r_tui[2]), .D1(catch_sync[0]), .S(r_tui[7]), .Y(n314) );
  XNOR2XL U595 ( .A(gt_647_B_3_), .B(n249), .Y(n443) );
  XNOR2XL U596 ( .A(ui_intv_cnt[2]), .B(n5), .Y(n435) );
  XNOR2XL U597 ( .A(n17), .B(n12), .Y(n434) );
  OAI32X1 U598 ( .A(n345), .B(new_rx_sync_cnt[1]), .C(new_rx_sync_cnt[0]), .D(
        n446), .E(n447), .Y(n426) );
  NOR43XL U599 ( .B(rx_trans_8_chg), .C(n448), .D(ff_chg), .A(n449), .Y(n447)
         );
  OAI31XL U600 ( .A(n450), .B(ui_intv_cnt[6]), .C(ui_intv_cnt[5]), .D(n368), 
        .Y(n449) );
  OAI21X1 U601 ( .B(rx_ui_1_2[6]), .C(n324), .A(n451), .Y(n450) );
  OAI22X1 U602 ( .A(N142), .B(n441), .C(n452), .D(n453), .Y(n451) );
  AOI211X1 U603 ( .C(n12), .D(n454), .A(n455), .B(n456), .Y(n453) );
  AOI21BBXL U604 ( .B(n454), .C(n12), .A(ui_intv_cnt[1]), .Y(n456) );
  OAI22X1 U605 ( .A(ui_intv_cnt[2]), .B(n442), .C(N141), .D(n389), .Y(n455) );
  NAND2X1 U606 ( .A(ui_intv_cnt[0]), .B(n445), .Y(n454) );
  MUX2IX1 U607 ( .D0(r_tui[3]), .D1(catch_sync[1]), .S(r_tui[7]), .Y(n445) );
  INVX1 U608 ( .A(r_tui[7]), .Y(n252) );
  MAJ3X1 U609 ( .A(n389), .B(n457), .C(N141), .Y(n452) );
  NOR2X1 U610 ( .A(rx_ui_1_2[4]), .B(n357), .Y(n457) );
  MUX2IX1 U611 ( .D0(adp_tx_ui_5_), .D1(catch_sync[3]), .S(r_tui[7]), .Y(n442)
         );
  MUX2IX1 U612 ( .D0(adp_tx_ui_6_), .D1(catch_sync[4]), .S(r_tui[7]), .Y(n389)
         );
  MUX2IX1 U613 ( .D0(adp_tx_ui_7_), .D1(catch_sync[5]), .S(r_tui[7]), .Y(n441)
         );
  OAI21X1 U614 ( .B(n458), .C(n459), .A(n460), .Y(n448) );
  OAI211X1 U615 ( .C(rx_ui_3_8[5]), .D(n249), .A(n461), .B(n462), .Y(n460) );
  AOI22AXL U616 ( .A(n463), .B(n464), .D(rx_ui_3_8[4]), .C(N142), .Y(n462) );
  NAND3X1 U617 ( .A(n465), .B(n466), .C(n467), .Y(n464) );
  AOI22AXL U618 ( .A(n468), .B(n469), .D(rx_ui_3_8[2]), .C(ui_intv_cnt[2]), 
        .Y(n467) );
  OAI21X1 U619 ( .B(n468), .C(n469), .A(ui_intv_cnt[1]), .Y(n465) );
  INVX1 U620 ( .A(rx_ui_3_8[1]), .Y(n469) );
  NAND2X1 U621 ( .A(rx_ui_3_8[0]), .B(n240), .Y(n468) );
  AOI32X1 U622 ( .A(n466), .B(n357), .C(rx_ui_3_8[2]), .D(rx_ui_3_8[3]), .E(
        n241), .Y(n463) );
  INVX1 U623 ( .A(ui_intv_cnt[2]), .Y(n357) );
  OR2X1 U624 ( .A(rx_ui_3_8[3]), .B(n241), .Y(n466) );
  INVX1 U625 ( .A(n459), .Y(n461) );
  OAI21X1 U626 ( .B(rx_ui_3_8[6]), .C(n248), .A(n325), .Y(n459) );
  AOI221XL U627 ( .A(rx_ui_3_8[5]), .B(n249), .C(rx_ui_3_8[6]), .D(n248), .E(
        n470), .Y(n458) );
  INVX1 U628 ( .A(n471), .Y(n470) );
  OAI211X1 U629 ( .C(n249), .D(rx_ui_3_8[5]), .A(rx_ui_3_8[4]), .B(n324), .Y(
        n471) );
  NAND4X1 U630 ( .A(n472), .B(n473), .C(n474), .D(n475), .Y(n332) );
  NOR4XL U631 ( .A(n476), .B(n477), .C(n478), .D(n479), .Y(n475) );
  XNOR2XL U632 ( .A(adp_tx_1_4[6]), .B(n248), .Y(n479) );
  XNOR2XL U633 ( .A(adp_tx_1_4[5]), .B(n249), .Y(n478) );
  XNOR2XL U634 ( .A(adp_tx_1_4[4]), .B(n324), .Y(n477) );
  XNOR2XL U635 ( .A(adp_tx_1_4[3]), .B(n241), .Y(n476) );
  INVX1 U636 ( .A(N141), .Y(n241) );
  NOR3XL U637 ( .A(n480), .B(ui_intv_cnt[7]), .C(n313), .Y(n474) );
  XNOR2XL U638 ( .A(adp_tx_1_4[0]), .B(n240), .Y(n480) );
  XNOR2XL U639 ( .A(ui_intv_cnt[1]), .B(adp_tx_1_4[1]), .Y(n473) );
  XNOR2XL U640 ( .A(ui_intv_cnt[2]), .B(adp_tx_1_4[2]), .Y(n472) );
  INVX1 U641 ( .A(n433), .Y(n423) );
  OAI21X1 U642 ( .B(n363), .C(n212), .A(n481), .Y(n433) );
  OAI21X1 U643 ( .B(n8), .C(n206), .A(n482), .Y(n481) );
  OAI21X1 U644 ( .B(n363), .C(n417), .A(n212), .Y(n482) );
  INVX1 U645 ( .A(N363), .Y(n363) );
  OAI21X1 U646 ( .B(r_ctl[0]), .C(n214), .A(n295), .Y(n485) );
  NAND2X1 U647 ( .A(r_ctl[0]), .B(n214), .Y(n295) );
  INVX1 U648 ( .A(n344), .Y(n446) );
  NOR3XL U649 ( .A(n311), .B(n487), .C(n418), .Y(n486) );
  NAND4X1 U650 ( .A(n21), .B(n489), .C(symb_cnt[3]), .D(n208), .Y(n345) );
  NOR3XL U651 ( .A(n368), .B(n311), .C(n424), .Y(n483) );
  GEN2XL U652 ( .D(N362), .E(n208), .C(n491), .B(n489), .A(n344), .Y(n370) );
  NAND2X1 U653 ( .A(n368), .B(n418), .Y(n344) );
  OA21X1 U654 ( .B(n492), .C(N362), .A(N363), .Y(n491) );
  NAND2X1 U655 ( .A(n213), .B(n371), .Y(n488) );
  GEN3XL U656 ( .F(N362), .G(N159), .E(N160), .D(n493), .C(symb_cnt[2]), .B(
        symb_cnt[3]), .A(n406), .Y(n371) );
  OAI21BBX1 U657 ( .A(symb_cnt[3]), .B(n407), .C(n374), .Y(n406) );
  NOR2X1 U658 ( .A(n408), .B(N362), .Y(n407) );
  INVX1 U659 ( .A(n494), .Y(n408) );
  NAND2X1 U660 ( .A(n494), .B(n492), .Y(n493) );
  XNOR2XL U661 ( .A(N363), .B(N362), .Y(n494) );
  NAND2X1 U662 ( .A(n411), .B(symb_cnt[2]), .Y(n424) );
  INVX1 U663 ( .A(n492), .Y(n411) );
  NAND2X1 U664 ( .A(N159), .B(N160), .Y(n492) );
  NAND4X1 U665 ( .A(n495), .B(n496), .C(n497), .D(n498), .Y(n311) );
  NOR4XL U666 ( .A(n499), .B(n500), .C(n501), .D(n502), .Y(n498) );
  XNOR2XL U667 ( .A(n325), .B(adp_tx_ui_7_), .Y(n502) );
  INVX1 U668 ( .A(ui_intv_cnt[7]), .Y(n325) );
  XNOR2XL U669 ( .A(n248), .B(adp_tx_ui_6_), .Y(n501) );
  INVX1 U670 ( .A(ui_intv_cnt[6]), .Y(n248) );
  XNOR2XL U671 ( .A(n249), .B(adp_tx_ui_5_), .Y(n500) );
  XNOR2XL U672 ( .A(n324), .B(r_tui[4]), .Y(n499) );
  INVX1 U673 ( .A(N142), .Y(n324) );
  NOR3XL U674 ( .A(n503), .B(n313), .C(n504), .Y(n497) );
  XNOR2XL U675 ( .A(r_tui[1]), .B(n247), .Y(n504) );
  INVX1 U676 ( .A(ui_intv_cnt[1]), .Y(n247) );
  INVX1 U677 ( .A(n330), .Y(n328) );
  NAND2X1 U678 ( .A(us_cnt[1]), .B(us_cnt[0]), .Y(n330) );
  XNOR2XL U679 ( .A(n240), .B(r_tui[0]), .Y(n503) );
  INVX1 U680 ( .A(ui_intv_cnt[0]), .Y(n240) );
  XNOR2XL U681 ( .A(ui_intv_cnt[2]), .B(r_tui[2]), .Y(n496) );
  XNOR2XL U682 ( .A(N141), .B(r_tui[3]), .Y(n495) );
  NOR2X1 U683 ( .A(n418), .B(n210), .Y(n242) );
  NAND2X1 U684 ( .A(n489), .B(n399), .Y(n418) );
  INVX1 U685 ( .A(n401), .Y(n489) );
  NAND2X1 U686 ( .A(n374), .B(n207), .Y(n401) );
  NOR3XL U687 ( .A(n274), .B(n21), .C(n212), .Y(n490) );
  NOR2X1 U688 ( .A(n417), .B(N160), .Y(n331) );
  INVX1 U689 ( .A(ff_chg), .Y(n274) );
  NAND2X1 U690 ( .A(n487), .B(n207), .Y(n417) );
  INVX1 U691 ( .A(n368), .Y(n487) );
  OAI21X1 U692 ( .B(n210), .C(n207), .A(n374), .Y(n316) );
  OAI31XL U693 ( .A(n505), .B(symb_cnt[6]), .C(symb_cnt[5]), .D(n414), .Y(n484) );
  INVX1 U694 ( .A(n374), .Y(n414) );
  NOR2X1 U695 ( .A(n307), .B(symb_cnt[6]), .Y(n374) );
  OAI21X1 U696 ( .B(n399), .C(n207), .A(n210), .Y(n505) );
  NOR2X1 U697 ( .A(N160), .B(N159), .Y(n399) );
endmodule


module fcpegn_a0_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module fcpegn_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(SUM[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
endmodule


module fcpegn_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_2 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9555;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9555), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9555), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9555), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9555), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9555), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9555), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9555), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9555), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9555), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_3 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9573;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9573), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9573), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9573), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9573), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9573), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9573), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9573), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9573), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9573), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_4 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9591;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9591), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9591), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9591), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9591), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9591), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9591), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9591), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9591), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9591), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_0 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_0 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[4]), .Y(n2) );
  INVX1 U4 ( .A(set2[2]), .Y(n7) );
  INVX1 U5 ( .A(set2[1]), .Y(n1) );
  NAND3X1 U6 ( .A(n6), .B(n4), .C(n16), .Y(n21) );
  INVX1 U7 ( .A(set2[0]), .Y(n3) );
  INVX1 U8 ( .A(set2[3]), .Y(n5) );
  NAND4X1 U9 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U10 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U11 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U12 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U13 ( .C(n3), .D(n15), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U14 ( .A(rdat[0]), .Y(n15) );
  AOI211X1 U15 ( .C(n1), .D(n14), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U16 ( .A(rdat[1]), .Y(n14) );
  AOI211X1 U17 ( .C(n7), .D(n13), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U18 ( .A(rdat[2]), .Y(n13) );
  AOI211X1 U19 ( .C(n5), .D(n12), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U20 ( .A(rdat[3]), .Y(n12) );
  AOI211X1 U21 ( .C(n2), .D(n11), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U22 ( .A(rdat[4]), .Y(n11) );
  AOI211X1 U23 ( .C(n16), .D(n10), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U24 ( .A(rdat[5]), .Y(n10) );
  AOI211X1 U25 ( .C(n6), .D(n9), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U26 ( .A(rdat[6]), .Y(n9) );
  AOI211X1 U27 ( .C(n4), .D(n8), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U28 ( .A(rdat[7]), .Y(n8) );
  NOR2X1 U29 ( .A(rdat[6]), .B(n6), .Y(irq[6]) );
  NOR2X1 U30 ( .A(rdat[7]), .B(n4), .Y(irq[7]) );
  INVX1 U31 ( .A(set2[7]), .Y(n4) );
  NOR2X1 U32 ( .A(rdat[0]), .B(n3), .Y(irq[0]) );
  NOR2X1 U33 ( .A(rdat[1]), .B(n1), .Y(irq[1]) );
  NOR2X1 U34 ( .A(rdat[2]), .B(n7), .Y(irq[2]) );
  NOR2X1 U35 ( .A(rdat[4]), .B(n2), .Y(irq[4]) );
  NOR2X1 U36 ( .A(rdat[3]), .B(n5), .Y(irq[3]) );
  INVX1 U37 ( .A(set2[6]), .Y(n6) );
  NOR2X1 U38 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
  INVX1 U39 ( .A(set2[5]), .Y(n16) );
endmodule


module glreg_WIDTH8_0 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9609;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9609), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9609), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9609), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9609), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9609), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9609), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9609), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9609), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9609), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000000 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9627;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9627), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9627), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9627), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9627), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9627), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9627), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9627), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9627), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9627), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dpdmacc_a0 ( dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, r_wdat, r_acc, 
        r_dpdmsta, r_dm, r_dmchg, r_int, clk, rstz );
  input [7:0] r_wdat;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, clk, rstz;
  output r_dm, r_dmchg, r_int;
  wire   dp_chg, dp_rise, dm_fall, dp_active_acc, dp_inacti_acc, dm_active_acc,
         dm_inacti_acc, upd00, N12, N15, N16, N17, N18, N19, N22, N23, N24,
         N25, n21, n22, n23, n24, n25, n26, N34, N35, n1, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [7:0] wd00;

  ff_sync_2 u0_dpsync ( .i_org(dp_comp), .o_dbc(r_dpdmsta[6]), .o_chg(dp_chg), 
        .clk(clk), .rstz(n4) );
  ff_sync_1 u0_dmsync ( .i_org(dm_comp), .o_dbc(r_dm), .o_chg(r_dmchg), .clk(
        clk), .rstz(n4) );
  ff_sync_0 u0_idsync ( .i_org(id_comp), .o_dbc(r_dpdmsta[5]), .o_chg(), .clk(
        clk), .rstz(n5) );
  filter150us_a0_1 u0_dpfltr ( .active_hit(dp_active_acc), .inacti_hit(
        dp_inacti_acc), .start_edge(dp_rise), .any_edge(dp_chg), .clk(clk), 
        .rstz(n5) );
  filter150us_a0_0 u0_dmfltr ( .active_hit(dm_active_acc), .inacti_hit(
        dm_inacti_acc), .start_edge(dm_fall), .any_edge(r_dmchg), .clk(clk), 
        .rstz(n5) );
  glreg_a0_5 u0_accmltr ( .clk(clk), .arstz(n3), .we(upd00), .wdat(wd00), 
        .rdat(r_acc) );
  glreg_WIDTH5_0 u0_dpdmsta ( .clk(clk), .arstz(n4), .we(r_wr_1), .wdat(
        r_wdat[4:0]), .rdat(r_dpdmsta[4:0]) );
  INVX1 U3 ( .A(r_re_0), .Y(n1) );
  INVX1 U4 ( .A(n6), .Y(n4) );
  INVX1 U5 ( .A(n6), .Y(n3) );
  INVX1 U6 ( .A(n6), .Y(n5) );
  INVX1 U7 ( .A(rstz), .Y(n6) );
  NAND2X1 U8 ( .A(n23), .B(n1), .Y(upd00) );
  INVX1 U9 ( .A(r_re_0), .Y(n9) );
  NOR2X1 U10 ( .A(n7), .B(n11), .Y(n23) );
  NOR21XL U11 ( .B(r_dmchg), .A(n8), .Y(dm_fall) );
  INVX1 U12 ( .A(n22), .Y(n11) );
  INVX1 U13 ( .A(n21), .Y(n7) );
  OAI21X1 U14 ( .B(n23), .C(n9), .A(n24), .Y(r_int) );
  AOI33X1 U15 ( .A(n7), .B(n13), .C(n25), .D(n11), .E(n14), .F(n26), .Y(n24)
         );
  INVX1 U16 ( .A(r_acc[0]), .Y(n14) );
  ENOX1 U17 ( .A(n22), .B(n9), .C(N22), .D(n9), .Y(wd00[0]) );
  XOR2X1 U18 ( .A(N34), .B(r_acc[0]), .Y(N22) );
  ENOX1 U19 ( .A(n21), .B(n1), .C(N15), .D(n9), .Y(wd00[4]) );
  XOR2X1 U20 ( .A(N35), .B(r_acc[4]), .Y(N15) );
  AND2X1 U21 ( .A(N23), .B(n9), .Y(wd00[1]) );
  XNOR2XL U22 ( .A(r_acc[1]), .B(n20), .Y(N23) );
  AND2X1 U23 ( .A(N24), .B(n9), .Y(wd00[2]) );
  XOR2X1 U24 ( .A(n19), .B(r_acc[2]), .Y(N24) );
  NOR21XL U25 ( .B(r_acc[1]), .A(n20), .Y(n19) );
  AND2X1 U26 ( .A(N25), .B(n9), .Y(wd00[3]) );
  XNOR2XL U27 ( .A(r_acc[3]), .B(n18), .Y(N25) );
  NAND4X1 U28 ( .A(r_acc[2]), .B(r_acc[1]), .C(N34), .D(r_acc[0]), .Y(n18) );
  AND2X1 U29 ( .A(N16), .B(n9), .Y(wd00[5]) );
  XNOR2XL U30 ( .A(r_acc[5]), .B(n17), .Y(N16) );
  AND2X1 U31 ( .A(N17), .B(n9), .Y(wd00[6]) );
  XOR2X1 U32 ( .A(n16), .B(r_acc[6]), .Y(N17) );
  NOR21XL U33 ( .B(r_acc[5]), .A(n17), .Y(n16) );
  AND2X1 U34 ( .A(N18), .B(n9), .Y(wd00[7]) );
  XNOR2XL U35 ( .A(r_acc[7]), .B(n15), .Y(N18) );
  NAND4X1 U36 ( .A(r_acc[6]), .B(r_acc[5]), .C(N35), .D(r_acc[4]), .Y(n15) );
  AOI32X1 U37 ( .A(n10), .B(n8), .C(dm_active_acc), .D(r_dpdmsta[1]), .E(
        dm_inacti_acc), .Y(n21) );
  INVX1 U38 ( .A(r_dpdmsta[1]), .Y(n10) );
  AOI32X1 U39 ( .A(dp_active_acc), .B(n12), .C(r_dpdmsta[6]), .D(r_dpdmsta[0]), 
        .E(dp_inacti_acc), .Y(n22) );
  INVX1 U40 ( .A(r_dpdmsta[0]), .Y(n12) );
  NOR21XL U41 ( .B(dp_chg), .A(r_dpdmsta[6]), .Y(dp_rise) );
  INVX1 U42 ( .A(r_dm), .Y(n8) );
  AND2X1 U43 ( .A(N19), .B(n11), .Y(N34) );
  NAND4X1 U44 ( .A(r_acc[3]), .B(r_acc[2]), .C(r_acc[1]), .D(r_acc[0]), .Y(N19) );
  AND2X1 U45 ( .A(N12), .B(n7), .Y(N35) );
  NAND4X1 U46 ( .A(r_acc[7]), .B(r_acc[6]), .C(r_acc[5]), .D(r_acc[4]), .Y(N12) );
  NAND2X1 U47 ( .A(N34), .B(r_acc[0]), .Y(n20) );
  NAND2X1 U48 ( .A(N35), .B(r_acc[4]), .Y(n17) );
  NOR3XL U49 ( .A(r_acc[1]), .B(r_acc[3]), .C(r_acc[2]), .Y(n26) );
  NOR3XL U50 ( .A(r_acc[5]), .B(r_acc[7]), .C(r_acc[6]), .Y(n25) );
  INVX1 U51 ( .A(r_acc[4]), .Y(n13) );
  BUFX3 U52 ( .A(r_dm), .Y(r_dpdmsta[7]) );
endmodule


module glreg_WIDTH5_0 ( clk, arstz, we, wdat, rdat );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we;
  wire   net9645;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9645), .TE(1'b0) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9645), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9645), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9645), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9645), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9645), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_5 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9663;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9663), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9663), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9663), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9663), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9663), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9663), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9663), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9663), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9663), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_0 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz );
  input start_edge, any_edge, clk, rstz;
  output active_hit, inacti_hit;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, net9681, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [11:0] dbcnt;

  SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9681), .TE(1'b0) );
  filter150us_a0_0_DW01_inc_0 add_76 ( .A(dbcnt), .SUM({N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12}) );
  DFFRQX1 dbcnt_reg_11_ ( .D(N36), .C(net9681), .XR(n2), .Q(dbcnt[11]) );
  DFFRQX1 dbcnt_reg_1_ ( .D(N26), .C(net9681), .XR(rstz), .Q(dbcnt[1]) );
  DFFRQX1 dbcnt_reg_9_ ( .D(N34), .C(net9681), .XR(n2), .Q(dbcnt[9]) );
  DFFRQX1 dbcnt_reg_2_ ( .D(N27), .C(net9681), .XR(rstz), .Q(dbcnt[2]) );
  DFFRQX1 dbcnt_reg_8_ ( .D(N33), .C(net9681), .XR(n2), .Q(dbcnt[8]) );
  DFFRQX1 dbcnt_reg_10_ ( .D(N35), .C(net9681), .XR(n2), .Q(dbcnt[10]) );
  DFFRQX1 dbcnt_reg_0_ ( .D(N25), .C(net9681), .XR(n2), .Q(dbcnt[0]) );
  DFFRQX1 dbcnt_reg_6_ ( .D(N31), .C(net9681), .XR(n2), .Q(dbcnt[6]) );
  DFFRQX1 dbcnt_reg_5_ ( .D(N30), .C(net9681), .XR(n2), .Q(dbcnt[5]) );
  DFFRQX1 dbcnt_reg_7_ ( .D(N32), .C(net9681), .XR(n2), .Q(dbcnt[7]) );
  DFFRQX1 dbcnt_reg_3_ ( .D(N28), .C(net9681), .XR(n2), .Q(dbcnt[3]) );
  DFFRQX1 dbcnt_reg_4_ ( .D(N29), .C(net9681), .XR(n2), .Q(dbcnt[4]) );
  BUFX3 U3 ( .A(n11), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  NOR3XL U6 ( .A(n13), .B(any_edge), .C(n14), .Y(n11) );
  AOI211X1 U7 ( .C(n4), .D(n5), .A(n6), .B(start_edge), .Y(inacti_hit) );
  INVX1 U8 ( .A(any_edge), .Y(n6) );
  AO21X1 U9 ( .B(n7), .C(n8), .A(n9), .Y(n5) );
  NOR4XL U10 ( .A(dbcnt[11]), .B(n10), .C(n9), .D(n7), .Y(active_hit) );
  NAND3X1 U11 ( .A(dbcnt[1]), .B(dbcnt[0]), .C(dbcnt[2]), .Y(n7) );
  AND2X1 U12 ( .A(N23), .B(n1), .Y(N36) );
  AND2X1 U13 ( .A(N22), .B(n1), .Y(N35) );
  AND2X1 U14 ( .A(N21), .B(n1), .Y(N34) );
  AND2X1 U15 ( .A(N20), .B(n1), .Y(N33) );
  AND2X1 U16 ( .A(N19), .B(n11), .Y(N32) );
  AND2X1 U17 ( .A(N18), .B(n11), .Y(N31) );
  AND2X1 U18 ( .A(N17), .B(n11), .Y(N30) );
  AND2X1 U19 ( .A(N16), .B(n11), .Y(N29) );
  AND2X1 U20 ( .A(N15), .B(n11), .Y(N28) );
  AND2X1 U21 ( .A(N14), .B(n11), .Y(N27) );
  AND2X1 U22 ( .A(N13), .B(n11), .Y(N26) );
  OAI21BBX1 U23 ( .A(N12), .B(n11), .C(n12), .Y(N25) );
  OAI21X1 U24 ( .B(n13), .C(n14), .A(any_edge), .Y(n12) );
  OR2X1 U25 ( .A(n11), .B(any_edge), .Y(N24) );
  OAI21X1 U26 ( .B(n8), .C(n9), .A(n4), .Y(n14) );
  INVX1 U27 ( .A(dbcnt[11]), .Y(n4) );
  NAND3X1 U28 ( .A(dbcnt[8]), .B(dbcnt[10]), .C(dbcnt[9]), .Y(n9) );
  NOR42XL U29 ( .C(n8), .D(n15), .A(dbcnt[0]), .B(dbcnt[10]), .Y(n13) );
  NOR4XL U30 ( .A(dbcnt[9]), .B(dbcnt[8]), .C(dbcnt[2]), .D(dbcnt[1]), .Y(n15)
         );
  INVX1 U31 ( .A(n10), .Y(n8) );
  NAND32X1 U32 ( .B(dbcnt[4]), .C(dbcnt[3]), .A(n16), .Y(n10) );
  NOR3XL U33 ( .A(dbcnt[5]), .B(dbcnt[7]), .C(dbcnt[6]), .Y(n16) );
endmodule


module filter150us_a0_0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_1 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz );
  input start_edge, any_edge, clk, rstz;
  output active_hit, inacti_hit;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, net9699, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [11:0] dbcnt;

  SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9699), .TE(1'b0) );
  filter150us_a0_1_DW01_inc_0 add_76 ( .A(dbcnt), .SUM({N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12}) );
  DFFRQX1 dbcnt_reg_4_ ( .D(N29), .C(net9699), .XR(n2), .Q(dbcnt[4]) );
  DFFRQX1 dbcnt_reg_11_ ( .D(N36), .C(net9699), .XR(n2), .Q(dbcnt[11]) );
  DFFRQX1 dbcnt_reg_1_ ( .D(N26), .C(net9699), .XR(rstz), .Q(dbcnt[1]) );
  DFFRQX1 dbcnt_reg_9_ ( .D(N34), .C(net9699), .XR(n2), .Q(dbcnt[9]) );
  DFFRQX1 dbcnt_reg_2_ ( .D(N27), .C(net9699), .XR(rstz), .Q(dbcnt[2]) );
  DFFRQX1 dbcnt_reg_8_ ( .D(N33), .C(net9699), .XR(n2), .Q(dbcnt[8]) );
  DFFRQX1 dbcnt_reg_10_ ( .D(N35), .C(net9699), .XR(n2), .Q(dbcnt[10]) );
  DFFRQX1 dbcnt_reg_0_ ( .D(N25), .C(net9699), .XR(n2), .Q(dbcnt[0]) );
  DFFRQX1 dbcnt_reg_6_ ( .D(N31), .C(net9699), .XR(n2), .Q(dbcnt[6]) );
  DFFRQX1 dbcnt_reg_5_ ( .D(N30), .C(net9699), .XR(n2), .Q(dbcnt[5]) );
  DFFRQX1 dbcnt_reg_7_ ( .D(N32), .C(net9699), .XR(n2), .Q(dbcnt[7]) );
  DFFRQX1 dbcnt_reg_3_ ( .D(N28), .C(net9699), .XR(n2), .Q(dbcnt[3]) );
  BUFX3 U3 ( .A(n11), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  NOR3XL U6 ( .A(n13), .B(any_edge), .C(n14), .Y(n11) );
  AOI211X1 U7 ( .C(n4), .D(n5), .A(n6), .B(start_edge), .Y(inacti_hit) );
  INVX1 U8 ( .A(any_edge), .Y(n6) );
  AO21X1 U9 ( .B(n7), .C(n8), .A(n9), .Y(n5) );
  NOR4XL U10 ( .A(dbcnt[11]), .B(n10), .C(n9), .D(n7), .Y(active_hit) );
  NAND3X1 U11 ( .A(dbcnt[1]), .B(dbcnt[0]), .C(dbcnt[2]), .Y(n7) );
  AND2X1 U12 ( .A(N23), .B(n1), .Y(N36) );
  AND2X1 U13 ( .A(N22), .B(n1), .Y(N35) );
  AND2X1 U14 ( .A(N21), .B(n1), .Y(N34) );
  AND2X1 U15 ( .A(N20), .B(n1), .Y(N33) );
  AND2X1 U16 ( .A(N19), .B(n11), .Y(N32) );
  AND2X1 U17 ( .A(N18), .B(n11), .Y(N31) );
  AND2X1 U18 ( .A(N17), .B(n11), .Y(N30) );
  AND2X1 U19 ( .A(N16), .B(n11), .Y(N29) );
  AND2X1 U20 ( .A(N15), .B(n11), .Y(N28) );
  AND2X1 U21 ( .A(N14), .B(n11), .Y(N27) );
  AND2X1 U22 ( .A(N13), .B(n11), .Y(N26) );
  OAI21BBX1 U23 ( .A(N12), .B(n11), .C(n12), .Y(N25) );
  OAI21X1 U24 ( .B(n13), .C(n14), .A(any_edge), .Y(n12) );
  OR2X1 U25 ( .A(n11), .B(any_edge), .Y(N24) );
  OAI21X1 U26 ( .B(n8), .C(n9), .A(n4), .Y(n14) );
  INVX1 U27 ( .A(dbcnt[11]), .Y(n4) );
  NAND3X1 U28 ( .A(dbcnt[8]), .B(dbcnt[10]), .C(dbcnt[9]), .Y(n9) );
  NOR42XL U29 ( .C(n8), .D(n15), .A(dbcnt[0]), .B(dbcnt[10]), .Y(n13) );
  NOR4XL U30 ( .A(dbcnt[9]), .B(dbcnt[8]), .C(dbcnt[2]), .D(dbcnt[1]), .Y(n15)
         );
  INVX1 U31 ( .A(n10), .Y(n8) );
  NAND32X1 U32 ( .B(dbcnt[4]), .C(dbcnt[3]), .A(n16), .Y(n10) );
  NOR3XL U33 ( .A(dbcnt[5]), .B(dbcnt[7]), .C(dbcnt[6]), .Y(n16) );
endmodule


module filter150us_a0_1_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ff_sync_0 ( i_org, o_dbc, o_chg, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_;

  DFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .C(clk), .XR(rstz), .Q(o_dbc) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_1 ( i_org, o_dbc, o_chg, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   n3, d_org_0_, n1;

  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .C(clk), .XR(rstz), .Q(n3) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(o_dbc) );
  XOR2X1 U5 ( .A(n3), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_2 ( i_org, o_dbc, o_chg, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_;

  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .C(clk), .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module dacmux_a0 ( clk, srstz, i_comp, r_comp_opt, r_wdat, r_adofs, r_isofs, 
        r_wr, dacv_wr, o_dacv, o_shrst, o_hold, o_dac1, o_daci_sel, o_dat, 
        r_dac_en, r_sar_en, o_dactl, o_cmpsta, x_daclsb, o_intr, o_smpl );
  input [2:0] r_comp_opt;
  input [7:0] r_wdat;
  output [7:0] r_adofs;
  output [7:0] r_isofs;
  input [10:0] r_wr;
  input [17:0] dacv_wr;
  output [143:0] o_dacv;
  output [9:0] o_dac1;
  output [17:0] o_daci_sel;
  output [17:0] o_dat;
  output [17:0] r_dac_en;
  output [17:0] r_sar_en;
  output [7:0] o_dactl;
  output [7:0] o_cmpsta;
  output [5:0] x_daclsb;
  output [4:0] o_smpl;
  input clk, srstz, i_comp;
  output o_shrst, o_hold, o_intr;
  wire   n566, n567, n568, n569, n570, n571, n572, n573, dacyc_done, updcmp,
         semi_start, auto_start, auto_sar, sacyc_done, sar_ini, sar_nxt,
         ps_sample, sampl_begn, sampl_done, ps_md4ch, updlsb, N859, tochg,
         N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1250,
         N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1261, N1262,
         N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1272, N1273, N1274,
         N1275, N1276, N1277, N1278, N1279, N1280, N1283, N1284, N1285, N1286,
         N1287, N1288, N1289, N1290, N1291, N1294, N1295, N1296, N1297, N1298,
         N1299, N1300, N1301, N1302, N1305, N1306, N1307, N1308, N1309, N1310,
         N1311, N1312, N1313, N1316, N1317, N1318, N1319, N1320, N1321, N1322,
         N1323, N1324, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334,
         N1335, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346,
         N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1360,
         N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1371, N1372,
         N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1382, N1383, N1384,
         N1385, N1386, N1387, N1388, N1389, N1390, N1393, N1394, N1395, N1396,
         N1397, N1398, N1399, N1400, N1401, N1404, N1405, N1406, N1407, N1408,
         N1409, N1410, N1411, N1412, N1415, N1416, N1417, N1418, N1419, N1420,
         N1421, N1422, N1423, N1426, N1427, N1428, N1429, N1430, N1431, N1432,
         N1433, N1434, n63, n99, n101, n148, n149, n150, n152, n159, n160,
         n199, n200, n201, n202, n203, n263, n264, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, net145949, net156831, net162211,
         net162210, net167900, net168001, net169004, net169040, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n86, n87, n88, n90, n91, n92, n94, n95, n96, n97, n98,
         n100, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n151, n153, n154, n155, n156, n157, n158, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565;
  wire   [1:0] syn_comp;
  wire   [4:0] cs_ptr;
  wire   [17:0] datcmp;
  wire   [4:0] ps_ptr;
  wire   [9:0] r_dac1v;
  wire   [9:0] r_rpt_v;
  wire   [17:0] app_dacis;
  wire   [17:0] pos_dacis;
  wire   [5:0] wdlsb;
  wire   [17:0] upd;
  wire   [7:0] wda;
  wire   [143:0] r_dacvs;
  wire   [7:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;

  glreg_00000012 u0_compi ( .clk(clk), .arstz(n198), .we(updcmp), .wdat(datcmp), .rdat(o_dat) );
  dac2sar_a0 u0_dac2sar ( .r_dac_t(o_dactl[3:2]), .r_dacyc(o_dactl[7]), 
        .r_sar10(n63), .sar_ini(sar_ini), .sar_nxt(sar_nxt), .semi_nxt(n99), 
        .auto_sar(auto_sar), .busy(o_dactl[0]), .stop(net145949), .sync_i(
        syn_comp[1]), .ps_sample(ps_sample), .sampl_begn(sampl_begn), 
        .sampl_done(sampl_done), .sh_rst(o_shrst), .dacyc_done(dacyc_done), 
        .sacyc_done(sacyc_done), .dac_v(r_dac1v), .rpt_v(r_rpt_v), .clk(clk), 
        .srstz(n198) );
  shmux_00000005_00000012_00000012 u0_shmux ( .ps_md4ch(ps_md4ch), 
        .r_comp_swtch(r_comp_opt[2]), .r_semi(n101), .r_loop(o_dactl[1]), 
        .r_dac_en({r_dac_en[17:4], n100, r_dac_en[2:0]}), .wr_dacv(dacv_wr), 
        .busy(o_dactl[0]), .sh_hold(o_hold), .stop(net145949), .semi_start(
        semi_start), .auto_start(auto_start), .mxcyc_done(n111), .sampl_begn(
        sampl_begn), .sampl_done(sampl_done), .app_dacis(app_dacis), 
        .pos_dacis(pos_dacis), .cs_ptr(cs_ptr), .ps_ptr(ps_ptr), .clk(clk), 
        .srstz(n198) );
  glreg_WIDTH7_1 u0_dactl ( .clk(clk), .arstz(n197), .we(net169040), .wdat({
        r_wdat[7:6], n27, net156831, r_wdat[3], n21, n24}), .rdat(o_dactl[7:1]) );
  glreg_a0_49 u0_dacen ( .clk(clk), .arstz(n172), .we(r_wr[1]), .wdat({
        r_wdat[7:6], n27, net167900, r_wdat[3], n21, n24, n32}), .rdat({
        r_dac_en[7:4], n573, r_dac_en[2:0]}) );
  glreg_a0_48 u0_saren ( .clk(clk), .arstz(n173), .we(r_wr[2]), .wdat({
        r_wdat[7:6], n27, net156831, r_wdat[3], n21, n23, n32}), .rdat(
        r_sar_en[7:0]) );
  glreg_WIDTH6_2 u0_daclsb ( .clk(clk), .arstz(n198), .we(updlsb), .wdat(wdlsb), .rdat(x_daclsb) );
  glreg_a0_47 dacvs_0__u0 ( .clk(clk), .arstz(n174), .we(upd[0]), .wdat({n43, 
        n45, n46, n70, n48, n52, n56, n62}), .rdat(r_dacvs[7:0]) );
  glreg_a0_46 dacvs_1__u0 ( .clk(clk), .arstz(n185), .we(upd[1]), .wdat({n43, 
        n45, n47, n71, n49, n53, n57, n64}), .rdat(r_dacvs[15:8]) );
  glreg_a0_45 dacvs_2__u0 ( .clk(clk), .arstz(n175), .we(upd[2]), .wdat({n43, 
        n45, n47, n71, n49, n53, n57, n64}), .rdat(r_dacvs[23:16]) );
  glreg_a0_44 dacvs_3__u0 ( .clk(clk), .arstz(n176), .we(upd[3]), .wdat({
        wda[7:6], n46, n71, n48, n52, n56, n62}), .rdat(r_dacvs[31:24]) );
  glreg_a0_43 dacvs_4__u0 ( .clk(clk), .arstz(n177), .we(upd[4]), .wdat({n43, 
        n45, n47, n70, n49, n53, n57, n64}), .rdat(r_dacvs[39:32]) );
  glreg_a0_42 dacvs_5__u0 ( .clk(clk), .arstz(n178), .we(upd[5]), .wdat({
        wda[7:6], n47, n71, n49, n53, n56, n62}), .rdat(r_dacvs[47:40]) );
  glreg_a0_41 dacvs_6__u0 ( .clk(clk), .arstz(n179), .we(upd[6]), .wdat({
        wda[7:6], n47, n71, n48, n52, n57, n64}), .rdat(r_dacvs[55:48]) );
  glreg_a0_40 dacvs_7__u0 ( .clk(clk), .arstz(n180), .we(upd[7]), .wdat({
        wda[7:6], n47, n70, n48, n52, n57, n64}), .rdat(r_dacvs[63:56]) );
  glreg_a0_39 dacvs_8__u0 ( .clk(clk), .arstz(n181), .we(upd[8]), .wdat({
        wda[7:6], n47, n70, n49, n53, n57, n64}), .rdat(r_dacvs[71:64]) );
  glreg_a0_38 dacvs_9__u0 ( .clk(clk), .arstz(n182), .we(upd[9]), .wdat({
        wda[7:6], n47, n71, n49, n53, n57, n64}), .rdat(r_dacvs[79:72]) );
  glreg_a0_37 dacvs_10__u0 ( .clk(clk), .arstz(n183), .we(upd[10]), .wdat({
        wda[7:6], n46, n70, n48, n52, n57, n64}), .rdat(r_dacvs[87:80]) );
  glreg_a0_36 dacvs_11__u0 ( .clk(clk), .arstz(n184), .we(upd[11]), .wdat({
        wda[7:6], n47, n70, n48, n52, n56, n62}), .rdat(r_dacvs[95:88]) );
  glreg_a0_35 dacvs_12__u0 ( .clk(clk), .arstz(n186), .we(upd[12]), .wdat({
        wda[7:6], n46, n71, n48, n52, n56, n62}), .rdat(r_dacvs[103:96]) );
  glreg_a0_34 dacvs_13__u0 ( .clk(clk), .arstz(n187), .we(upd[13]), .wdat({n43, 
        n45, n46, n71, n49, n53, n57, n64}), .rdat(r_dacvs[111:104]) );
  glreg_a0_33 dacvs_14__u0 ( .clk(clk), .arstz(n188), .we(upd[14]), .wdat({n43, 
        n45, n46, n70, n48, n52, n56, n62}), .rdat(r_dacvs[119:112]) );
  glreg_a0_32 dacvs_15__u0 ( .clk(clk), .arstz(n189), .we(upd[15]), .wdat({n43, 
        n45, n46, n70, n48, n52, n56, n62}), .rdat(r_dacvs[127:120]) );
  glreg_a0_31 dacvs_16__u0 ( .clk(clk), .arstz(n190), .we(upd[16]), .wdat({n43, 
        n45, n46, n71, n49, n53, n56, n62}), .rdat(r_dacvs[135:128]) );
  glreg_a0_30 dacvs_17__u0 ( .clk(clk), .arstz(n191), .we(upd[17]), .wdat({n43, 
        n45, n46, n70, n49, n53, n56, n62}), .rdat(r_dacvs[143:136]) );
  glsta_a0_1 u0_cmpsta ( .clk(clk), .arstz(n192), .rst0(1'b0), .set2(setsta), 
        .clr1(clrsta), .rdat(o_cmpsta), .irq(r_irq) );
  glreg_a0_29 u0_adofs ( .clk(clk), .arstz(n193), .we(r_wr[5]), .wdat({
        r_wdat[7:6], n26, net167900, r_wdat[3], n21, n24, n31}), .rdat({n566, 
        n567, r_adofs[5], n568, n569, n570, n571, n572}) );
  glreg_a0_28 u0_isofs ( .clk(clk), .arstz(n194), .we(r_wr[6]), .wdat({
        r_wdat[7:6], n27, net156831, r_wdat[3], n21, n24, n32}), .rdat(r_isofs) );
  glreg_a0_27 u1_dacen ( .clk(clk), .arstz(n195), .we(r_wr[7]), .wdat({
        r_wdat[7:6], n27, net167900, r_wdat[3], n21, n24, n31}), .rdat(
        r_dac_en[15:8]) );
  glreg_a0_26 u1_saren ( .clk(clk), .arstz(n196), .we(r_wr[8]), .wdat({
        r_wdat[7:6], n27, net156831, r_wdat[3], n21, n24, n32}), .rdat(
        r_sar_en[15:8]) );
  glreg_WIDTH2_1 u2_dacen ( .clk(clk), .arstz(n186), .we(r_wr[9]), .wdat({n24, 
        n32}), .rdat(r_dac_en[17:16]) );
  glreg_WIDTH2_0 u2_saren ( .clk(clk), .arstz(n197), .we(r_wr[10]), .wdat({n24, 
        n31}), .rdat(r_sar_en[17:16]) );
  dacmux_a0_DW01_add_0 add_235_I18 ( .A({1'b0, r_dacvs[143:136]}), .B({n166, 
        n166, r_adofs[6:5], n95, n75, n91, n87, n40}), .CI(1'b0), .SUM({N1434, 
        N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426}), .CO() );
  dacmux_a0_DW01_add_1 add_235_I17 ( .A({1'b0, r_dacvs[135:128]}), .B({n166, 
        n166, n567, n97, n94, n74, n90, n86, r_adofs[0]}), .CI(1'b0), .SUM({
        N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415}), .CO()
         );
  dacmux_a0_DW01_add_2 add_235_I16 ( .A({1'b0, r_dacvs[127:120]}), .B({n166, 
        n166, r_adofs[6], n97, r_adofs[4:1], n40}), .CI(1'b0), .SUM({N1412, 
        N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404}), .CO() );
  dacmux_a0_DW01_add_3 add_235_I15 ( .A({1'b0, r_dacvs[119:112]}), .B({n166, 
        n166, r_adofs[6:5], n95, n75, n91, n87, n38}), .CI(1'b0), .SUM({N1401, 
        N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393}), .CO() );
  dacmux_a0_DW01_add_4 add_235_I14 ( .A({1'b0, r_dacvs[111:104]}), .B({n166, 
        n166, n567, r_adofs[5], n95, n75, n91, n87, n38}), .CI(1'b0), .SUM({
        N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382}), .CO()
         );
  dacmux_a0_DW01_add_5 add_235_I13 ( .A({1'b0, r_dacvs[103:96]}), .B({n167, 
        n167, n567, n97, n94, n74, n90, n86, n38}), .CI(1'b0), .SUM({N1379, 
        N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371}), .CO() );
  dacmux_a0_DW01_add_6 add_235_I12 ( .A({1'b0, r_dacvs[95:88]}), .B({n167, 
        n167, n567, r_adofs[5:1], n38}), .CI(1'b0), .SUM({N1368, N1367, N1366, 
        N1365, N1364, N1363, N1362, N1361, N1360}), .CO() );
  dacmux_a0_DW01_add_7 add_235_I11 ( .A({1'b0, r_dacvs[87:80]}), .B({n167, 
        n167, r_adofs[6:0]}), .CI(1'b0), .SUM({N1357, N1356, N1355, N1354, 
        N1353, N1352, N1351, N1350, N1349}), .CO() );
  dacmux_a0_DW01_add_8 add_235_I10 ( .A({1'b0, r_dacvs[79:72]}), .B({n167, 
        n167, n567, n97, n92, n72, n88, n84, r_adofs[0]}), .CI(1'b0), .SUM({
        N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338}), .CO()
         );
  dacmux_a0_DW01_add_9 add_235_I9 ( .A({1'b0, r_dacvs[71:64]}), .B({n167, n168, 
        n567, n97, n92, n72, n88, n84, n40}), .CI(1'b0), .SUM({N1335, N1334, 
        N1333, N1332, N1331, N1330, N1329, N1328, N1327}), .CO() );
  dacmux_a0_DW01_add_10 add_235_I8 ( .A({1'b0, r_dacvs[63:56]}), .B({n168, 
        n168, n567, r_adofs[5:1], n40}), .CI(1'b0), .SUM({N1324, N1323, N1322, 
        N1321, N1320, N1319, N1318, N1317, N1316}), .CO() );
  dacmux_a0_DW01_add_11 add_235_I7 ( .A({1'b0, r_dacvs[55:48]}), .B({n168, 
        n168, n567, n97, n94, n74, n90, n86, n38}), .CI(1'b0), .SUM({N1313, 
        N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305}), .CO() );
  dacmux_a0_DW01_add_12 add_235_I6 ( .A({1'b0, r_dacvs[47:40]}), .B({n168, 
        n168, r_adofs[6], n97, n95, n75, n91, n87, n38}), .CI(1'b0), .SUM({
        N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294}), .CO()
         );
  dacmux_a0_DW01_add_13 add_235_I5 ( .A({1'b0, r_dacvs[39:32]}), .B({n168, 
        n168, r_adofs[6], n97, n94, n74, n90, n86, n38}), .CI(1'b0), .SUM({
        N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283}), .CO()
         );
  dacmux_a0_DW01_add_14 add_235_I4 ( .A({1'b0, r_dacvs[31:24]}), .B({n168, 
        n169, r_adofs[6:5], n95, n75, n91, n87, r_adofs[0]}), .CI(1'b0), .SUM(
        {N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272}), 
        .CO() );
  dacmux_a0_DW01_add_15 add_235_I3 ( .A({1'b0, r_dacvs[23:16]}), .B({
        r_isofs[7], r_isofs}), .CI(1'b0), .SUM({N1269, N1268, N1267, N1266, 
        N1265, N1264, N1263, N1262, N1261}), .CO() );
  dacmux_a0_DW01_add_16 add_235_I2 ( .A({1'b0, r_dacvs[15:8]}), .B({n169, n169, 
        r_adofs[6], n97, n94, n74, n90, n86, n38}), .CI(1'b0), .SUM({N1258, 
        N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250}), .CO() );
  dacmux_a0_DW01_add_17 add_235 ( .A({1'b0, r_dacvs[7:0]}), .B({n169, n167, 
        n567, r_adofs[5:0]}), .CI(1'b0), .SUM({N1247, N1246, N1245, N1244, 
        N1243, N1242, N1241, N1240, N1239}), .CO() );
  DFFQX1 syn_comp_reg_1_ ( .D(syn_comp[0]), .C(clk), .Q(syn_comp[1]) );
  DFFQX1 syn_comp_reg_0_ ( .D(i_comp), .C(clk), .Q(syn_comp[0]) );
  INVX1 U3 ( .A(N1434), .Y(n533) );
  AO21X1 U4 ( .B(N1407), .C(n41), .A(n526), .Y(o_dacv[123]) );
  INVX1 U5 ( .A(n404), .Y(n407) );
  AO21X1 U6 ( .B(n445), .C(n428), .A(n427), .Y(n432) );
  INVX2 U7 ( .A(n414), .Y(n417) );
  MUX2IX4 U8 ( .D0(n112), .D1(n104), .S(pos_dacis[14]), .Y(n460) );
  AND4X2 U9 ( .A(n469), .B(n474), .C(n456), .D(n459), .Y(n104) );
  NAND21X2 U10 ( .B(n19), .A(n436), .Y(n453) );
  INVXL U11 ( .A(n406), .Y(n395) );
  INVXL U12 ( .A(N1390), .Y(n521) );
  INVXL U13 ( .A(r_wdat[4]), .Y(net162211) );
  MUX2BXL U14 ( .D0(n399), .D1(n398), .S(pos_dacis[3]), .Y(n414) );
  MUX2X1 U15 ( .D0(n395), .D1(n394), .S(pos_dacis[2]), .Y(n399) );
  BUFX3 U16 ( .A(n571), .Y(r_adofs[1]) );
  BUFX3 U17 ( .A(n570), .Y(n88) );
  BUFX3 U18 ( .A(n570), .Y(r_adofs[2]) );
  BUFX3 U19 ( .A(n569), .Y(n72) );
  BUFX3 U20 ( .A(n568), .Y(n92) );
  BUFX3 U21 ( .A(n568), .Y(r_adofs[4]) );
  INVX1 U22 ( .A(pos_dacis[0]), .Y(n401) );
  BUFX3 U23 ( .A(n571), .Y(n84) );
  INVX1 U42 ( .A(n486), .Y(n487) );
  INVX1 U43 ( .A(n507), .Y(n508) );
  INVX1 U44 ( .A(N1346), .Y(n509) );
  AO21X1 U45 ( .B(n409), .C(n408), .A(n407), .Y(n437) );
  MUX2X1 U46 ( .D0(n278), .D1(n277), .S(ps_ptr[3]), .Y(n279) );
  AO21X1 U47 ( .B(r_dac_en[16]), .C(ps_ptr[4]), .A(n383), .Y(n392) );
  AO21X1 U48 ( .B(n464), .C(n463), .A(n468), .Y(n472) );
  INVX1 U49 ( .A(r_wr[0]), .Y(n33) );
  BUFX3 U50 ( .A(n569), .Y(r_adofs[3]) );
  AO21X1 U51 ( .B(N1408), .C(n41), .A(n526), .Y(o_dacv[124]) );
  OA22X1 U52 ( .A(n434), .B(n440), .C(pos_dacis[10]), .D(n433), .Y(n19) );
  INVX1 U53 ( .A(r_adofs[5]), .Y(n96) );
  INVX1 U54 ( .A(n566), .Y(n171) );
  NAND21X1 U55 ( .B(n31), .A(r_wr[0]), .Y(net169004) );
  INVX1 U56 ( .A(n36), .Y(net169040) );
  INVX1 U57 ( .A(r_wdat[2]), .Y(n20) );
  INVX1 U58 ( .A(n20), .Y(n21) );
  INVX1 U59 ( .A(r_wdat[1]), .Y(n22) );
  INVX1 U60 ( .A(n22), .Y(n23) );
  INVX1 U61 ( .A(n22), .Y(n24) );
  INVX1 U62 ( .A(r_wdat[5]), .Y(n25) );
  INVX1 U63 ( .A(n25), .Y(n26) );
  INVX1 U64 ( .A(n25), .Y(n27) );
  INVX1 U65 ( .A(n567), .Y(n28) );
  INVX1 U66 ( .A(n28), .Y(r_adofs[6]) );
  INVXL U67 ( .A(r_wdat[0]), .Y(n30) );
  INVXL U68 ( .A(n30), .Y(n31) );
  INVXL U69 ( .A(n30), .Y(n32) );
  XNOR2X1 U70 ( .A(pos_dacis[0]), .B(pos_dacis[1]), .Y(n406) );
  INVXL U71 ( .A(N1401), .Y(n524) );
  NAND32XL U72 ( .B(n446), .C(n429), .A(n432), .Y(n433) );
  INVX1 U73 ( .A(N1412), .Y(n527) );
  INVXL U74 ( .A(N1379), .Y(n518) );
  BUFX3 U75 ( .A(n527), .Y(n41) );
  INVX3 U76 ( .A(n525), .Y(n526) );
  AO21X4 U77 ( .B(n431), .C(n430), .A(n452), .Y(n436) );
  NAND3X1 U78 ( .A(n460), .B(n459), .C(n458), .Y(n114) );
  OAI211X1 U79 ( .C(n420), .D(n447), .A(n419), .B(n418), .Y(n421) );
  MUX2AX2 U80 ( .D0(n105), .D1(n415), .S(pos_dacis[6]), .Y(n420) );
  BUFX6 U81 ( .A(n572), .Y(n40) );
  BUFX6 U82 ( .A(n572), .Y(n38) );
  MUX2IX2 U83 ( .D0(net162210), .D1(net162211), .S(n34), .Y(ps_sample) );
  NAND21X1 U84 ( .B(n33), .A(n37), .Y(n36) );
  NOR21X2 U85 ( .B(r_wr[0]), .A(n35), .Y(n34) );
  NAND2X1 U86 ( .A(n32), .B(o_dactl[0]), .Y(n37) );
  AND2X2 U87 ( .A(r_wdat[0]), .B(o_dactl[0]), .Y(n35) );
  BUFX6 U88 ( .A(n572), .Y(r_adofs[0]) );
  INVX3 U89 ( .A(n519), .Y(n520) );
  NAND21X1 U90 ( .B(r_adofs[7]), .A(N1346), .Y(n507) );
  BUFXL U91 ( .A(net162211), .Y(net168001) );
  INVXL U92 ( .A(dacv_wr[13]), .Y(n247) );
  INVXL U93 ( .A(net168001), .Y(net167900) );
  INVXL U94 ( .A(net169004), .Y(net145949) );
  INVXL U95 ( .A(dacv_wr[12]), .Y(n248) );
  INVX1 U96 ( .A(wda[7]), .Y(n42) );
  INVX1 U97 ( .A(n42), .Y(n43) );
  INVX1 U98 ( .A(wda[6]), .Y(n44) );
  INVX1 U99 ( .A(n44), .Y(n45) );
  BUFX3 U100 ( .A(n220), .Y(wda[5]) );
  INVX1 U101 ( .A(wda[5]), .Y(n46) );
  INVX1 U102 ( .A(wda[5]), .Y(n47) );
  BUFX3 U103 ( .A(n218), .Y(wda[3]) );
  INVX1 U104 ( .A(wda[3]), .Y(n48) );
  INVX1 U105 ( .A(wda[3]), .Y(n49) );
  NAND2X1 U106 ( .A(n378), .B(n199), .Y(n298) );
  INVX1 U107 ( .A(n298), .Y(n50) );
  INVX1 U108 ( .A(n298), .Y(n51) );
  BUFX3 U109 ( .A(n217), .Y(wda[2]) );
  INVX1 U110 ( .A(wda[2]), .Y(n52) );
  INVX1 U111 ( .A(wda[2]), .Y(n53) );
  NAND2X1 U112 ( .A(n378), .B(n375), .Y(n294) );
  INVX1 U113 ( .A(n294), .Y(n54) );
  INVX1 U114 ( .A(n294), .Y(n55) );
  BUFX3 U115 ( .A(n216), .Y(wda[1]) );
  INVX1 U116 ( .A(wda[1]), .Y(n56) );
  INVX1 U117 ( .A(wda[1]), .Y(n57) );
  NAND2X1 U118 ( .A(n374), .B(n199), .Y(n296) );
  INVX1 U119 ( .A(n296), .Y(n58) );
  INVX1 U120 ( .A(n296), .Y(n59) );
  NAND2X1 U121 ( .A(n377), .B(n375), .Y(n291) );
  INVX1 U122 ( .A(n291), .Y(n60) );
  INVX1 U123 ( .A(n291), .Y(n61) );
  BUFX3 U124 ( .A(n215), .Y(wda[0]) );
  INVX1 U125 ( .A(wda[0]), .Y(n62) );
  INVX1 U126 ( .A(wda[0]), .Y(n64) );
  INVX1 U127 ( .A(n379), .Y(n65) );
  NAND2X1 U128 ( .A(n377), .B(n199), .Y(n297) );
  INVX1 U129 ( .A(n297), .Y(n66) );
  INVX1 U130 ( .A(n297), .Y(n67) );
  NAND2X1 U131 ( .A(n375), .B(n376), .Y(n292) );
  INVX1 U132 ( .A(n292), .Y(n68) );
  INVX1 U133 ( .A(n292), .Y(n69) );
  BUFX3 U134 ( .A(n219), .Y(wda[4]) );
  INVX1 U135 ( .A(wda[4]), .Y(n70) );
  INVX1 U136 ( .A(wda[4]), .Y(n71) );
  BUFX1 U137 ( .A(n569), .Y(n74) );
  BUFX1 U138 ( .A(n569), .Y(n75) );
  NAND2X1 U139 ( .A(n376), .B(n199), .Y(n295) );
  INVX1 U140 ( .A(n295), .Y(n76) );
  INVX1 U141 ( .A(n295), .Y(n77) );
  NAND2X1 U142 ( .A(n374), .B(n375), .Y(n293) );
  INVX1 U143 ( .A(n293), .Y(n78) );
  INVX1 U144 ( .A(n293), .Y(n79) );
  BUFX3 U145 ( .A(n299), .Y(n80) );
  NOR2X1 U146 ( .A(o_dactl[0]), .B(semi_start), .Y(n267) );
  INVX1 U147 ( .A(n267), .Y(n81) );
  INVX1 U148 ( .A(n267), .Y(n82) );
  INVX1 U149 ( .A(r_comp_opt[0]), .Y(n147) );
  INVX1 U150 ( .A(n147), .Y(n83) );
  BUFX1 U151 ( .A(n571), .Y(n86) );
  BUFX1 U152 ( .A(n571), .Y(n87) );
  BUFX1 U153 ( .A(n570), .Y(n90) );
  BUFX1 U154 ( .A(n570), .Y(n91) );
  BUFX1 U155 ( .A(n568), .Y(n94) );
  BUFX1 U156 ( .A(n568), .Y(n95) );
  INVX1 U157 ( .A(n96), .Y(n97) );
  INVX1 U158 ( .A(n573), .Y(n98) );
  INVX1 U159 ( .A(n98), .Y(n100) );
  INVX1 U160 ( .A(n98), .Y(r_dac_en[3]) );
  NAND21X1 U161 ( .B(ps_ptr[2]), .A(n275), .Y(n272) );
  NAND21XL U162 ( .B(ps_ptr[2]), .A(ps_ptr[1]), .Y(n271) );
  NAND21XL U163 ( .B(ps_ptr[1]), .A(ps_ptr[2]), .Y(n274) );
  AO21XL U164 ( .B(N1240), .C(n482), .A(n481), .Y(o_dacv[1]) );
  AO21XL U165 ( .B(N1295), .C(n497), .A(n496), .Y(o_dacv[41]) );
  AO21XL U166 ( .B(N1306), .C(n500), .A(n499), .Y(o_dacv[49]) );
  AO21XL U167 ( .B(N1318), .C(n503), .A(n502), .Y(o_dacv[58]) );
  INVXL U168 ( .A(N1269), .Y(n488) );
  OAI22AX1 U169 ( .D(n453), .C(n442), .A(n435), .B(n473), .Y(n441) );
  INVX1 U170 ( .A(n413), .Y(n419) );
  NAND21XL U171 ( .B(n452), .A(n451), .Y(n456) );
  AO21XL U172 ( .B(n466), .C(n470), .A(n108), .Y(o_smpl[0]) );
  NAND21XL U173 ( .B(n479), .A(n478), .Y(o_smpl[4]) );
  INVX1 U174 ( .A(o_dactl[4]), .Y(net162210) );
  AO21XL U175 ( .B(N1317), .C(n503), .A(n502), .Y(o_dacv[57]) );
  OAI21BBXL U176 ( .A(ps_ptr[4]), .B(r_dac_en[17]), .C(n103), .Y(n391) );
  MUX2IX1 U177 ( .D0(n390), .D1(n389), .S(ps_ptr[3]), .Y(n103) );
  OAI22XL U178 ( .A(n427), .B(n426), .C(n425), .D(n424), .Y(n438) );
  OAI21BXL U179 ( .C(n472), .B(pos_dacis[17]), .A(n471), .Y(o_smpl[2]) );
  INVXL U180 ( .A(n438), .Y(n439) );
  INVXL U181 ( .A(n455), .Y(n466) );
  OAI211XL U182 ( .C(n460), .D(n454), .A(n459), .B(n458), .Y(n455) );
  AOI21XL U183 ( .B(n417), .C(n409), .A(n407), .Y(n105) );
  NAND3XL U184 ( .A(n110), .B(n418), .C(n448), .Y(n113) );
  INVX1 U185 ( .A(n399), .Y(n396) );
  NAND21X1 U186 ( .B(pos_dacis[0]), .A(n406), .Y(n397) );
  AND3X1 U187 ( .A(n226), .B(n225), .C(n106), .Y(n233) );
  AOI22XL U188 ( .A(r_sar_en[8]), .B(dacv_wr[8]), .C(r_sar_en[9]), .D(
        dacv_wr[9]), .Y(n106) );
  AND4X1 U189 ( .A(n229), .B(n228), .C(n227), .D(n107), .Y(n230) );
  AOI22X1 U190 ( .A(dacv_wr[0]), .B(r_sar_en[0]), .C(dacv_wr[1]), .D(
        r_sar_en[1]), .Y(n107) );
  AOI22XL U191 ( .A(r_dacvs[35]), .B(n58), .C(r_dacvs[51]), .D(n66), .Y(n337)
         );
  AOI22XL U192 ( .A(r_dacvs[43]), .B(n58), .C(r_dacvs[59]), .D(n66), .Y(n341)
         );
  INVX1 U193 ( .A(dacv_wr[4]), .Y(n257) );
  INVX1 U194 ( .A(dacv_wr[2]), .Y(n261) );
  INVX1 U195 ( .A(dacv_wr[3]), .Y(n259) );
  INVX1 U196 ( .A(n204), .Y(n198) );
  INVX1 U197 ( .A(n155), .Y(n146) );
  INVX1 U198 ( .A(n155), .Y(n145) );
  INVX1 U199 ( .A(r_wr[4]), .Y(n536) );
  INVX1 U200 ( .A(n204), .Y(n192) );
  INVX1 U201 ( .A(n204), .Y(n191) );
  INVX1 U202 ( .A(n205), .Y(n190) );
  INVX1 U203 ( .A(n206), .Y(n189) );
  INVX1 U204 ( .A(n206), .Y(n188) );
  INVX1 U205 ( .A(n205), .Y(n187) );
  INVX1 U206 ( .A(n204), .Y(n186) );
  INVX1 U207 ( .A(n205), .Y(n184) );
  INVX1 U208 ( .A(n205), .Y(n183) );
  INVX1 U209 ( .A(n206), .Y(n182) );
  INVX1 U210 ( .A(n204), .Y(n181) );
  INVX1 U211 ( .A(n205), .Y(n180) );
  INVX1 U212 ( .A(n206), .Y(n179) );
  INVX1 U213 ( .A(n205), .Y(n178) );
  INVX1 U214 ( .A(n205), .Y(n177) );
  INVX1 U215 ( .A(n206), .Y(n176) );
  INVX1 U216 ( .A(n206), .Y(n175) );
  INVX1 U217 ( .A(n206), .Y(n185) );
  INVX1 U218 ( .A(n206), .Y(n174) );
  INVX1 U219 ( .A(n205), .Y(n196) );
  INVX1 U220 ( .A(n205), .Y(n195) );
  INVX1 U221 ( .A(n205), .Y(n194) );
  INVX1 U222 ( .A(n204), .Y(n193) );
  INVX1 U223 ( .A(n206), .Y(n173) );
  INVX1 U224 ( .A(n204), .Y(n197) );
  INVX1 U225 ( .A(srstz), .Y(n204) );
  INVX1 U226 ( .A(r_wr[3]), .Y(n537) );
  NOR2X1 U227 ( .A(n156), .B(n158), .Y(n378) );
  NAND2X1 U228 ( .A(n154), .B(n156), .Y(n564) );
  NAND21X1 U229 ( .B(n156), .A(n154), .Y(n262) );
  NAND21X1 U230 ( .B(n154), .A(n156), .Y(n260) );
  NAND21X1 U231 ( .B(n265), .A(n256), .Y(n544) );
  NAND21X1 U232 ( .B(n262), .A(n256), .Y(n557) );
  NAND21X1 U233 ( .B(n265), .A(n253), .Y(n545) );
  NAND21X1 U234 ( .B(n262), .A(n253), .Y(n558) );
  NAND21X1 U235 ( .B(n265), .A(n243), .Y(n543) );
  NAND21X1 U236 ( .B(n262), .A(n243), .Y(n555) );
  NAND21X1 U237 ( .B(n260), .A(n256), .Y(n549) );
  NAND21X1 U238 ( .B(n258), .A(n256), .Y(n553) );
  NAND21X1 U239 ( .B(n260), .A(n253), .Y(n546) );
  NAND21X1 U240 ( .B(n258), .A(n253), .Y(n550) );
  OR2X1 U241 ( .A(n266), .B(n265), .Y(n541) );
  OR2X1 U242 ( .A(n266), .B(n262), .Y(n556) );
  OR2X1 U243 ( .A(n266), .B(n260), .Y(n548) );
  OR2X1 U244 ( .A(n266), .B(n258), .Y(n552) );
  INVX1 U245 ( .A(n206), .Y(n172) );
  INVX1 U246 ( .A(srstz), .Y(n206) );
  INVX1 U247 ( .A(srstz), .Y(n205) );
  INVX1 U248 ( .A(n276), .Y(n385) );
  NAND21X1 U249 ( .B(n275), .A(ps_ptr[2]), .Y(n276) );
  INVX1 U250 ( .A(n272), .Y(n388) );
  INVX1 U251 ( .A(n273), .Y(n384) );
  NAND21X1 U252 ( .B(ps_ptr[4]), .A(n388), .Y(n273) );
  NAND21X1 U253 ( .B(n393), .A(n270), .Y(semi_start) );
  INVX1 U254 ( .A(n270), .Y(n99) );
  INVX1 U255 ( .A(n155), .Y(n154) );
  AND2X1 U256 ( .A(net167900), .B(r_wr[4]), .Y(clrsta[4]) );
  NOR2X1 U257 ( .A(n535), .B(n536), .Y(clrsta[6]) );
  NOR2X1 U258 ( .A(n534), .B(n536), .Y(clrsta[7]) );
  NOR2X1 U259 ( .A(n65), .B(n154), .Y(n285) );
  INVX1 U260 ( .A(n142), .Y(n144) );
  INVX1 U261 ( .A(n157), .Y(n156) );
  INVX1 U262 ( .A(n161), .Y(n158) );
  NOR2X1 U263 ( .A(n161), .B(n156), .Y(n374) );
  NOR2X1 U264 ( .A(n157), .B(n158), .Y(n376) );
  NOR2X1 U265 ( .A(n157), .B(n161), .Y(n377) );
  NOR2X1 U266 ( .A(n565), .B(n561), .Y(setsta[4]) );
  NOR2X1 U267 ( .A(n565), .B(n562), .Y(setsta[5]) );
  NOR2X1 U268 ( .A(n565), .B(n563), .Y(setsta[6]) );
  NOR2X1 U269 ( .A(n565), .B(n564), .Y(setsta[7]) );
  INVX1 U270 ( .A(n538), .Y(n151) );
  INVX1 U271 ( .A(n538), .Y(n153) );
  INVX1 U272 ( .A(n142), .Y(n143) );
  NAND2X1 U273 ( .A(n156), .B(n155), .Y(n563) );
  NAND2X1 U274 ( .A(n154), .B(n157), .Y(n562) );
  NAND21X1 U275 ( .B(n154), .A(n157), .Y(n265) );
  NAND21X1 U276 ( .B(n157), .A(n154), .Y(n258) );
  NAND32X1 U277 ( .B(n162), .C(n158), .A(n142), .Y(n266) );
  NAND21X1 U278 ( .B(n265), .A(n109), .Y(n542) );
  NAND21X1 U279 ( .B(n262), .A(n109), .Y(n554) );
  NAND21X1 U280 ( .B(n260), .A(n109), .Y(n547) );
  NAND21X1 U281 ( .B(n258), .A(n109), .Y(n551) );
  INVX1 U282 ( .A(n255), .Y(n256) );
  NAND32X1 U283 ( .B(n162), .C(n161), .A(n142), .Y(n255) );
  INVX1 U284 ( .A(n249), .Y(n253) );
  NAND32X1 U285 ( .B(n158), .C(n142), .A(n163), .Y(n249) );
  INVX1 U286 ( .A(n241), .Y(n243) );
  NAND32X1 U287 ( .B(n158), .C(n163), .A(n142), .Y(n241) );
  NAND21X1 U288 ( .B(r_adofs[7]), .A(N1412), .Y(n525) );
  INVX1 U289 ( .A(N1423), .Y(n530) );
  INVX1 U290 ( .A(N1368), .Y(n515) );
  INVX1 U291 ( .A(N1357), .Y(n512) );
  INVX1 U292 ( .A(N1335), .Y(n506) );
  INVX1 U293 ( .A(n531), .Y(n532) );
  NAND21X1 U294 ( .B(r_adofs[7]), .A(N1434), .Y(n531) );
  INVX1 U295 ( .A(n528), .Y(n529) );
  NAND21X1 U296 ( .B(r_adofs[7]), .A(N1423), .Y(n528) );
  INVX1 U297 ( .A(n513), .Y(n514) );
  NAND21X1 U298 ( .B(r_adofs[7]), .A(N1368), .Y(n513) );
  INVX1 U299 ( .A(n510), .Y(n511) );
  NAND21X1 U300 ( .B(r_adofs[7]), .A(N1357), .Y(n510) );
  INVX1 U301 ( .A(n522), .Y(n523) );
  NAND21X1 U302 ( .B(r_adofs[7]), .A(N1401), .Y(n522) );
  INVX1 U303 ( .A(n516), .Y(n517) );
  NAND21X1 U304 ( .B(r_adofs[7]), .A(N1379), .Y(n516) );
  NAND21X1 U305 ( .B(n566), .A(N1390), .Y(n519) );
  INVX1 U306 ( .A(n504), .Y(n505) );
  NAND21X1 U307 ( .B(r_adofs[7]), .A(N1335), .Y(n504) );
  INVX1 U308 ( .A(n483), .Y(n484) );
  NAND21X1 U309 ( .B(n169), .A(N1258), .Y(n483) );
  INVX1 U310 ( .A(n489), .Y(n490) );
  NAND21X1 U311 ( .B(n169), .A(N1280), .Y(n489) );
  INVX1 U312 ( .A(n480), .Y(n481) );
  NAND21X1 U313 ( .B(n169), .A(N1247), .Y(n480) );
  INVX1 U314 ( .A(n422), .Y(n425) );
  NAND21X1 U315 ( .B(n446), .A(n428), .Y(n422) );
  AND2X1 U316 ( .A(n472), .B(n465), .Y(n108) );
  INVX1 U317 ( .A(n492), .Y(n493) );
  NAND21X1 U318 ( .B(n169), .A(N1291), .Y(n492) );
  INVX1 U319 ( .A(N1258), .Y(n485) );
  INVX1 U320 ( .A(N1280), .Y(n491) );
  INVX1 U321 ( .A(N1247), .Y(n482) );
  INVX1 U322 ( .A(N1291), .Y(n494) );
  INVX1 U323 ( .A(N1313), .Y(n500) );
  INVX1 U324 ( .A(N1324), .Y(n503) );
  INVX1 U325 ( .A(n498), .Y(n499) );
  NAND21X1 U326 ( .B(n169), .A(N1313), .Y(n498) );
  INVX1 U327 ( .A(n501), .Y(n502) );
  NAND21X1 U328 ( .B(n566), .A(N1324), .Y(n501) );
  INVX1 U329 ( .A(n495), .Y(n496) );
  NAND21X1 U330 ( .B(n169), .A(N1302), .Y(n495) );
  INVX1 U331 ( .A(N1302), .Y(n497) );
  INVX1 U332 ( .A(n269), .Y(auto_start) );
  INVX1 U333 ( .A(n271), .Y(n387) );
  INVX1 U334 ( .A(n274), .Y(n386) );
  INVX1 U335 ( .A(ps_ptr[1]), .Y(n275) );
  INVX1 U336 ( .A(n239), .Y(n393) );
  INVX1 U337 ( .A(r_wdat[3]), .Y(n238) );
  NAND6XL U338 ( .A(n27), .B(r_wdat[3]), .C(n21), .D(n240), .E(n30), .F(n535), 
        .Y(n270) );
  OAI22X1 U339 ( .A(n244), .B(n81), .C(n543), .D(n148), .Y(upd[16]) );
  INVXL U340 ( .A(dacv_wr[16]), .Y(n244) );
  OAI22X1 U341 ( .A(n245), .B(n81), .C(n551), .D(n148), .Y(upd[15]) );
  OAI22X1 U342 ( .A(n246), .B(n81), .C(n547), .D(n148), .Y(upd[14]) );
  OAI22X1 U343 ( .A(n247), .B(n81), .C(n554), .D(n148), .Y(upd[13]) );
  OAI22X1 U344 ( .A(n248), .B(n81), .C(n542), .D(n148), .Y(upd[12]) );
  OAI22X1 U345 ( .A(n250), .B(n81), .C(n550), .D(n153), .Y(upd[11]) );
  INVXL U346 ( .A(dacv_wr[11]), .Y(n250) );
  OAI22X1 U347 ( .A(n251), .B(n81), .C(n546), .D(n153), .Y(upd[10]) );
  OAI22X1 U348 ( .A(n252), .B(n81), .C(n558), .D(n153), .Y(upd[9]) );
  INVXL U349 ( .A(dacv_wr[9]), .Y(n252) );
  OAI22X1 U350 ( .A(n254), .B(n81), .C(n545), .D(n153), .Y(upd[8]) );
  INVXL U351 ( .A(dacv_wr[8]), .Y(n254) );
  OAI22AX1 U352 ( .D(dacv_wr[7]), .C(n82), .A(n553), .B(n153), .Y(upd[7]) );
  OAI22AX1 U353 ( .D(dacv_wr[6]), .C(n82), .A(n549), .B(n153), .Y(upd[6]) );
  OAI22AX1 U354 ( .D(dacv_wr[5]), .C(n82), .A(n557), .B(n153), .Y(upd[5]) );
  OAI22X1 U355 ( .A(n257), .B(n82), .C(n544), .D(n153), .Y(upd[4]) );
  OAI22X1 U356 ( .A(n259), .B(n82), .C(n552), .D(n153), .Y(upd[3]) );
  OAI22AX1 U357 ( .D(dacv_wr[1]), .C(n82), .A(n556), .B(n153), .Y(upd[1]) );
  OAI22X1 U358 ( .A(n242), .B(n82), .C(n555), .D(n151), .Y(upd[17]) );
  INVXL U359 ( .A(dacv_wr[17]), .Y(n242) );
  OAI22X1 U360 ( .A(n261), .B(n82), .C(n548), .D(n151), .Y(upd[2]) );
  OAI22AX1 U361 ( .D(dacv_wr[0]), .C(n82), .A(n541), .B(n151), .Y(upd[0]) );
  INVX1 U362 ( .A(cs_ptr[2]), .Y(n161) );
  INVX1 U363 ( .A(cs_ptr[0]), .Y(n155) );
  INVX1 U364 ( .A(cs_ptr[1]), .Y(n157) );
  INVX1 U365 ( .A(r_wdat[6]), .Y(n535) );
  INVX1 U366 ( .A(r_wdat[7]), .Y(n534) );
  AND2X1 U367 ( .A(n27), .B(r_wr[4]), .Y(clrsta[5]) );
  AND2X1 U368 ( .A(n24), .B(r_wr[4]), .Y(clrsta[1]) );
  AND2X1 U369 ( .A(n21), .B(r_wr[4]), .Y(clrsta[2]) );
  AND2X1 U370 ( .A(r_wdat[3]), .B(r_wr[4]), .Y(clrsta[3]) );
  INVX1 U371 ( .A(n163), .Y(n162) );
  INVX1 U372 ( .A(cs_ptr[4]), .Y(n163) );
  NOR2X1 U373 ( .A(cs_ptr[3]), .B(n162), .Y(n199) );
  AND2X1 U374 ( .A(n154), .B(n379), .Y(n283) );
  INVX1 U375 ( .A(n379), .Y(n539) );
  INVX1 U376 ( .A(cs_ptr[3]), .Y(n142) );
  NOR21XL U377 ( .B(cs_ptr[3]), .A(n162), .Y(n375) );
  NOR32XL U378 ( .B(n378), .C(n162), .A(cs_ptr[3]), .Y(n299) );
  INVX1 U379 ( .A(dacyc_done), .Y(n540) );
  OR3XL U380 ( .A(n560), .B(cs_ptr[3]), .C(n162), .Y(n565) );
  NOR2X1 U381 ( .A(n561), .B(n559), .Y(setsta[0]) );
  NOR2X1 U382 ( .A(n563), .B(n559), .Y(setsta[2]) );
  NOR2X1 U383 ( .A(n562), .B(n559), .Y(setsta[1]) );
  NOR2X1 U384 ( .A(n564), .B(n559), .Y(setsta[3]) );
  INVX1 U385 ( .A(n538), .Y(n148) );
  NAND21X1 U386 ( .B(cs_ptr[0]), .A(n157), .Y(n561) );
  NOR31X1 U387 ( .C(cs_ptr[2]), .A(n142), .B(cs_ptr[4]), .Y(n109) );
  AO21X1 U388 ( .B(N1283), .C(n494), .A(n493), .Y(o_dacv[32]) );
  AO21X1 U389 ( .B(N1262), .C(n488), .A(n487), .Y(o_dacv[17]) );
  AO21X1 U390 ( .B(N1263), .C(n488), .A(n487), .Y(o_dacv[18]) );
  AO21XL U391 ( .B(N1241), .C(n482), .A(n481), .Y(o_dacv[2]) );
  AO21X1 U392 ( .B(N1367), .C(n515), .A(n514), .Y(o_dacv[95]) );
  AO21X1 U393 ( .B(N1356), .C(n512), .A(n511), .Y(o_dacv[87]) );
  AO21X1 U394 ( .B(N1400), .C(n524), .A(n523), .Y(o_dacv[119]) );
  AO21X1 U395 ( .B(N1378), .C(n518), .A(n517), .Y(o_dacv[103]) );
  AO21X1 U396 ( .B(N1389), .C(n521), .A(n520), .Y(o_dacv[111]) );
  OR3XL U397 ( .A(n457), .B(n456), .C(n467), .Y(n464) );
  INVX1 U398 ( .A(n450), .Y(n431) );
  INVX1 U399 ( .A(n421), .Y(n428) );
  NAND32X1 U400 ( .B(n468), .C(n467), .A(n471), .Y(n477) );
  AO21X1 U401 ( .B(N1239), .C(n482), .A(n481), .Y(o_dacv[0]) );
  AO21XL U402 ( .B(N1361), .C(n515), .A(n514), .Y(o_dacv[89]) );
  AO21XL U403 ( .B(N1350), .C(n512), .A(n511), .Y(o_dacv[81]) );
  AO21XL U404 ( .B(N1394), .C(n524), .A(n523), .Y(o_dacv[113]) );
  AO21XL U405 ( .B(N1372), .C(n518), .A(n517), .Y(o_dacv[97]) );
  AO21XL U406 ( .B(N1383), .C(n521), .A(n520), .Y(o_dacv[105]) );
  AO21XL U407 ( .B(N1364), .C(n515), .A(n514), .Y(o_dacv[92]) );
  AO21XL U408 ( .B(N1366), .C(n515), .A(n514), .Y(o_dacv[94]) );
  AO21XL U409 ( .B(N1353), .C(n512), .A(n511), .Y(o_dacv[84]) );
  AO21XL U410 ( .B(N1355), .C(n512), .A(n511), .Y(o_dacv[86]) );
  AO21XL U411 ( .B(N1397), .C(n524), .A(n523), .Y(o_dacv[116]) );
  AO21XL U412 ( .B(N1399), .C(n524), .A(n523), .Y(o_dacv[118]) );
  AO21XL U413 ( .B(N1377), .C(n518), .A(n517), .Y(o_dacv[102]) );
  AO21XL U414 ( .B(N1375), .C(n518), .A(n517), .Y(o_dacv[100]) );
  AO21XL U415 ( .B(N1388), .C(n521), .A(n520), .Y(o_dacv[110]) );
  AO21XL U416 ( .B(N1386), .C(n521), .A(n520), .Y(o_dacv[108]) );
  AO21XL U417 ( .B(N1365), .C(n515), .A(n514), .Y(o_dacv[93]) );
  AO21XL U418 ( .B(N1354), .C(n512), .A(n511), .Y(o_dacv[85]) );
  AO21XL U419 ( .B(N1398), .C(n524), .A(n523), .Y(o_dacv[117]) );
  AO21XL U420 ( .B(N1376), .C(n518), .A(n517), .Y(o_dacv[101]) );
  AO21XL U421 ( .B(N1363), .C(n515), .A(n514), .Y(o_dacv[91]) );
  AO21XL U422 ( .B(N1352), .C(n512), .A(n511), .Y(o_dacv[83]) );
  AO21XL U423 ( .B(N1387), .C(n521), .A(n520), .Y(o_dacv[109]) );
  AO21XL U424 ( .B(N1396), .C(n524), .A(n523), .Y(o_dacv[115]) );
  AO21XL U425 ( .B(N1374), .C(n518), .A(n517), .Y(o_dacv[99]) );
  AO21XL U426 ( .B(N1385), .C(n521), .A(n520), .Y(o_dacv[107]) );
  AO21XL U427 ( .B(N1360), .C(n515), .A(n514), .Y(o_dacv[88]) );
  AO21XL U428 ( .B(N1349), .C(n512), .A(n511), .Y(o_dacv[80]) );
  AO21XL U429 ( .B(N1362), .C(n515), .A(n514), .Y(o_dacv[90]) );
  AO21XL U430 ( .B(N1393), .C(n524), .A(n523), .Y(o_dacv[112]) );
  AO21XL U431 ( .B(N1371), .C(n518), .A(n517), .Y(o_dacv[96]) );
  AO21XL U432 ( .B(N1382), .C(n521), .A(n520), .Y(o_dacv[104]) );
  INVX1 U433 ( .A(n430), .Y(n446) );
  AND2X1 U434 ( .A(n437), .B(n419), .Y(n110) );
  INVX1 U435 ( .A(n461), .Y(n465) );
  NAND21X1 U436 ( .B(n478), .A(n466), .Y(n461) );
  INVX1 U437 ( .A(n397), .Y(n394) );
  NAND21X1 U438 ( .B(n409), .A(n403), .Y(n404) );
  OAI211X1 U439 ( .C(n412), .D(n410), .A(n417), .B(n411), .Y(n403) );
  NAND21X1 U440 ( .B(n450), .A(n449), .Y(n451) );
  NAND21X1 U441 ( .B(n448), .A(n447), .Y(n449) );
  AO21XL U442 ( .B(N1284), .C(n494), .A(n493), .Y(o_dacv[33]) );
  AO21XL U443 ( .B(N1351), .C(n512), .A(n511), .Y(o_dacv[82]) );
  AO21XL U444 ( .B(N1395), .C(n524), .A(n523), .Y(o_dacv[114]) );
  AO21XL U445 ( .B(N1373), .C(n518), .A(n517), .Y(o_dacv[98]) );
  AO21XL U446 ( .B(N1384), .C(n521), .A(n520), .Y(o_dacv[106]) );
  OAI211XL U447 ( .C(n417), .D(n412), .A(n411), .B(n410), .Y(n413) );
  NAND32XL U448 ( .B(n417), .C(n416), .A(n418), .Y(n448) );
  AO21XL U449 ( .B(N1285), .C(n494), .A(n493), .Y(o_dacv[34]) );
  AO21XL U450 ( .B(N1296), .C(n497), .A(n496), .Y(o_dacv[42]) );
  INVX1 U451 ( .A(n171), .Y(n166) );
  INVX1 U452 ( .A(n171), .Y(n167) );
  INVX1 U453 ( .A(n171), .Y(n168) );
  INVX1 U454 ( .A(n171), .Y(r_adofs[7]) );
  INVX1 U455 ( .A(n416), .Y(n409) );
  INVX1 U456 ( .A(n171), .Y(n169) );
  INVX1 U457 ( .A(n429), .Y(n445) );
  OR2X1 U458 ( .A(n429), .B(n440), .Y(n450) );
  INVX1 U459 ( .A(n457), .Y(n442) );
  NOR32XL U460 ( .B(n237), .C(n236), .A(n235), .Y(n240) );
  NOR32XL U461 ( .B(n234), .C(n233), .A(n232), .Y(n235) );
  NOR32XL U462 ( .B(n101), .C(r_wdat[7]), .A(o_dactl[0]), .Y(n236) );
  NOR21XL U463 ( .B(n22), .A(net167900), .Y(n237) );
  AO21XL U464 ( .B(N1264), .C(n488), .A(n487), .Y(o_dacv[19]) );
  AO21XL U465 ( .B(N1242), .C(n482), .A(n481), .Y(o_dacv[3]) );
  INVX1 U466 ( .A(n479), .Y(n470) );
  AO21XL U467 ( .B(N1298), .C(n497), .A(n496), .Y(o_dacv[44]) );
  INVX1 U468 ( .A(n149), .Y(n63) );
  AO21XL U469 ( .B(N1299), .C(n497), .A(n496), .Y(o_dacv[45]) );
  AO21XL U470 ( .B(N1297), .C(n497), .A(n496), .Y(o_dacv[43]) );
  AO21XL U471 ( .B(N1286), .C(n494), .A(n493), .Y(o_dacv[35]) );
  AO21XL U472 ( .B(N1319), .C(n503), .A(n502), .Y(o_dacv[59]) );
  AO21XL U473 ( .B(N1290), .C(n494), .A(n493), .Y(o_dacv[39]) );
  AO21XL U474 ( .B(N1267), .C(n488), .A(n487), .Y(o_dacv[22]) );
  AO21XL U475 ( .B(N1245), .C(n482), .A(n481), .Y(o_dacv[6]) );
  AO21XL U476 ( .B(N1244), .C(n482), .A(n481), .Y(o_dacv[5]) );
  AO21XL U477 ( .B(N1243), .C(n482), .A(n481), .Y(o_dacv[4]) );
  AO21XL U478 ( .B(N1288), .C(n494), .A(n493), .Y(o_dacv[37]) );
  AO21XL U479 ( .B(N1287), .C(n494), .A(n493), .Y(o_dacv[36]) );
  NAND2X1 U480 ( .A(o_dactl[0]), .B(n120), .Y(n379) );
  AO21XL U481 ( .B(N1266), .C(n488), .A(n487), .Y(o_dacv[21]) );
  AO21XL U482 ( .B(N1265), .C(n488), .A(n487), .Y(o_dacv[20]) );
  AO21XL U483 ( .B(N1246), .C(n482), .A(n481), .Y(o_dacv[7]) );
  AO21XL U484 ( .B(N1289), .C(n494), .A(n493), .Y(o_dacv[38]) );
  AO21XL U485 ( .B(N1301), .C(n497), .A(n496), .Y(o_dacv[47]) );
  AO21XL U486 ( .B(N1322), .C(n503), .A(n502), .Y(o_dacv[62]) );
  AO21XL U487 ( .B(N1300), .C(n497), .A(n496), .Y(o_dacv[46]) );
  OAI21X1 U488 ( .B(n151), .C(n149), .A(n537), .Y(updlsb) );
  AO21XL U489 ( .B(N1268), .C(n488), .A(n487), .Y(o_dacv[23]) );
  INVX1 U490 ( .A(n159), .Y(n101) );
  MUX2AXL U491 ( .D0(n540), .D1(sacyc_done), .S(auto_sar), .Y(n111) );
  INVX1 U492 ( .A(n268), .Y(auto_sar) );
  NAND21X1 U493 ( .B(n101), .A(n120), .Y(n268) );
  NAND42X1 U494 ( .C(cs_ptr[3]), .D(n162), .A(tochg), .B(n560), .Y(n559) );
  NAND2X1 U495 ( .A(n263), .B(n264), .Y(o_intr) );
  NOR4XL U496 ( .A(r_irq[7]), .B(r_irq[6]), .C(r_irq[5]), .D(r_irq[4]), .Y(
        n264) );
  NOR4XL U497 ( .A(r_irq[3]), .B(r_irq[2]), .C(r_irq[1]), .D(r_irq[0]), .Y(
        n263) );
  NAND2X1 U498 ( .A(n158), .B(tochg), .Y(n560) );
  AO21X1 U499 ( .B(n101), .C(dacyc_done), .A(sacyc_done), .Y(n538) );
  NOR2X1 U500 ( .A(n150), .B(n540), .Y(updcmp) );
  XNOR2XL U501 ( .A(n120), .B(n125), .Y(n150) );
  AOI21X1 U502 ( .B(n159), .C(n160), .A(n540), .Y(sar_nxt) );
  NAND2X1 U503 ( .A(n125), .B(n120), .Y(n160) );
  AO21X1 U504 ( .B(N1250), .C(n485), .A(n484), .Y(o_dacv[8]) );
  AO21X1 U505 ( .B(N1272), .C(n491), .A(n490), .Y(o_dacv[24]) );
  AO21XL U506 ( .B(N1273), .C(n491), .A(n490), .Y(o_dacv[25]) );
  AO21X1 U507 ( .B(N1411), .C(n527), .A(n526), .Y(o_dacv[127]) );
  AO21X1 U508 ( .B(N1305), .C(n500), .A(n499), .Y(o_dacv[48]) );
  AO21X1 U509 ( .B(N1345), .C(n509), .A(n508), .Y(o_dacv[79]) );
  AO21X1 U510 ( .B(N1294), .C(n497), .A(n496), .Y(o_dacv[40]) );
  AO21X1 U511 ( .B(N1433), .C(n533), .A(n532), .Y(o_dacv[143]) );
  AO21XL U512 ( .B(N1307), .C(n500), .A(n499), .Y(o_dacv[50]) );
  AO21XL U513 ( .B(N1274), .C(n491), .A(n490), .Y(o_dacv[26]) );
  AO21X1 U514 ( .B(N1334), .C(n506), .A(n505), .Y(o_dacv[71]) );
  AO21XL U515 ( .B(N1251), .C(n485), .A(n484), .Y(o_dacv[9]) );
  AO21XL U516 ( .B(N1252), .C(n485), .A(n484), .Y(o_dacv[10]) );
  AO21X1 U517 ( .B(N1422), .C(n530), .A(n529), .Y(o_dacv[135]) );
  AO21XL U518 ( .B(N1344), .C(n509), .A(n508), .Y(o_dacv[78]) );
  AO21XL U519 ( .B(N1410), .C(n41), .A(n526), .Y(o_dacv[126]) );
  AO21XL U520 ( .B(N1341), .C(n509), .A(n508), .Y(o_dacv[75]) );
  NAND21X1 U521 ( .B(n108), .A(pos_dacis[17]), .Y(n471) );
  AOI21XL U522 ( .B(n442), .C(n436), .A(n441), .Y(n112) );
  NAND32XL U523 ( .B(pos_dacis[2]), .C(n406), .A(n405), .Y(n408) );
  AO21XL U524 ( .B(N1340), .C(n509), .A(n508), .Y(o_dacv[74]) );
  NAND21X1 U525 ( .B(n397), .A(n396), .Y(n398) );
  NAND32XL U526 ( .B(pos_dacis[6]), .C(n437), .A(n447), .Y(n444) );
  NAND21X1 U527 ( .B(n440), .A(n439), .Y(n443) );
  MUX2X2 U528 ( .D0(n420), .D1(n113), .S(pos_dacis[7]), .Y(n430) );
  MUX2IX1 U529 ( .D0(n460), .D1(n114), .S(pos_dacis[15]), .Y(n478) );
  AO21XL U530 ( .B(n470), .C(n469), .A(n477), .Y(o_smpl[1]) );
  INVX1 U531 ( .A(pos_dacis[9]), .Y(n426) );
  NAND21XL U532 ( .B(n414), .A(n110), .Y(n415) );
  OAI21BBX1 U533 ( .A(pos_dacis[11]), .B(pos_dacis[10]), .C(n115), .Y(n452) );
  OAI21X1 U534 ( .B(n440), .C(n438), .A(n433), .Y(n115) );
  AO21XL U535 ( .B(N1427), .C(n533), .A(n532), .Y(o_dacv[137]) );
  AO21XL U536 ( .B(N1416), .C(n530), .A(n529), .Y(o_dacv[129]) );
  AO21XL U537 ( .B(N1339), .C(n509), .A(n508), .Y(o_dacv[73]) );
  AO21XL U538 ( .B(N1405), .C(n41), .A(n526), .Y(o_dacv[121]) );
  AO21XL U539 ( .B(N1432), .C(n533), .A(n532), .Y(o_dacv[142]) );
  AO21XL U540 ( .B(N1430), .C(n533), .A(n532), .Y(o_dacv[140]) );
  AO21XL U541 ( .B(N1421), .C(n530), .A(n529), .Y(o_dacv[134]) );
  AO21XL U542 ( .B(N1419), .C(n530), .A(n529), .Y(o_dacv[132]) );
  AO21XL U543 ( .B(N1431), .C(n533), .A(n532), .Y(o_dacv[141]) );
  AO21XL U544 ( .B(N1420), .C(n530), .A(n529), .Y(o_dacv[133]) );
  AO21XL U545 ( .B(N1429), .C(n533), .A(n532), .Y(o_dacv[139]) );
  AO21XL U546 ( .B(N1418), .C(n530), .A(n529), .Y(o_dacv[131]) );
  AO21XL U547 ( .B(N1426), .C(n533), .A(n532), .Y(o_dacv[136]) );
  AO21XL U548 ( .B(N1415), .C(n530), .A(n529), .Y(o_dacv[128]) );
  AO21XL U549 ( .B(N1428), .C(n533), .A(n532), .Y(o_dacv[138]) );
  AO21XL U550 ( .B(N1417), .C(n530), .A(n529), .Y(o_dacv[130]) );
  AO21XL U551 ( .B(N1342), .C(n509), .A(n508), .Y(o_dacv[76]) );
  AO21XL U552 ( .B(N1343), .C(n509), .A(n508), .Y(o_dacv[77]) );
  AO21XL U553 ( .B(N1409), .C(n41), .A(n526), .Y(o_dacv[125]) );
  AO21XL U554 ( .B(N1333), .C(n506), .A(n505), .Y(o_dacv[70]) );
  AO21XL U555 ( .B(N1332), .C(n506), .A(n505), .Y(o_dacv[69]) );
  AO21XL U556 ( .B(N1338), .C(n509), .A(n508), .Y(o_dacv[72]) );
  AO21XL U557 ( .B(N1330), .C(n506), .A(n505), .Y(o_dacv[67]) );
  AO21XL U558 ( .B(N1404), .C(n41), .A(n526), .Y(o_dacv[120]) );
  AO21XL U559 ( .B(N1406), .C(n41), .A(n526), .Y(o_dacv[122]) );
  OAI22XL U560 ( .A(pos_dacis[12]), .B(n453), .C(n19), .D(n457), .Y(n459) );
  INVX1 U561 ( .A(n462), .Y(n468) );
  NAND21X1 U562 ( .B(n465), .A(pos_dacis[16]), .Y(n462) );
  INVX1 U563 ( .A(pos_dacis[15]), .Y(n454) );
  INVX1 U564 ( .A(n423), .Y(n427) );
  NAND21X1 U565 ( .B(pos_dacis[8]), .A(n425), .Y(n423) );
  AO21XL U566 ( .B(N1329), .C(n506), .A(n505), .Y(o_dacv[66]) );
  INVX1 U567 ( .A(n402), .Y(n411) );
  OAI211XL U568 ( .C(n406), .D(n405), .A(n401), .B(n400), .Y(n402) );
  INVXL U569 ( .A(pos_dacis[2]), .Y(n400) );
  NAND21XL U570 ( .B(n477), .A(n476), .Y(o_smpl[3]) );
  NAND21X1 U571 ( .B(n479), .A(n475), .Y(n476) );
  NAND21X1 U572 ( .B(n474), .A(n473), .Y(n475) );
  AO21X1 U573 ( .B(N1316), .C(n503), .A(n502), .Y(o_dacv[56]) );
  AO21XL U574 ( .B(N1328), .C(n506), .A(n505), .Y(o_dacv[65]) );
  AO21XL U575 ( .B(N1331), .C(n506), .A(n505), .Y(o_dacv[68]) );
  AO21XL U576 ( .B(N1327), .C(n506), .A(n505), .Y(o_dacv[64]) );
  INVXL U577 ( .A(n432), .Y(n434) );
  AO21X1 U578 ( .B(N1261), .C(n488), .A(n487), .Y(o_dacv[16]) );
  NAND21X1 U579 ( .B(r_isofs[7]), .A(N1269), .Y(n486) );
  INVX1 U580 ( .A(pos_dacis[3]), .Y(n405) );
  OAI21AX1 U581 ( .B(n116), .C(n117), .A(n393), .Y(sar_ini) );
  OAI21X1 U582 ( .B(auto_start), .C(n111), .A(n380), .Y(n116) );
  MUX2IX1 U583 ( .D0(n392), .D1(n391), .S(ps_ptr[0]), .Y(n117) );
  NAND21X1 U584 ( .B(pos_dacis[4]), .A(n412), .Y(n416) );
  AO2222XL U585 ( .A(n387), .B(r_sar_en[2]), .C(n384), .D(r_sar_en[0]), .E(
        n386), .F(r_sar_en[4]), .G(n385), .H(r_sar_en[6]), .Y(n278) );
  AO2222XL U586 ( .A(n388), .B(r_sar_en[8]), .C(n387), .D(r_sar_en[10]), .E(
        n386), .F(r_sar_en[12]), .G(n385), .H(r_sar_en[14]), .Y(n277) );
  MUX2IX1 U587 ( .D0(n118), .D1(n119), .S(ps_ptr[0]), .Y(n380) );
  AOI21XL U588 ( .B(ps_ptr[4]), .C(r_sar_en[16]), .A(n279), .Y(n118) );
  AOI21XL U589 ( .B(ps_ptr[4]), .C(r_sar_en[17]), .A(n282), .Y(n119) );
  MUX2X1 U590 ( .D0(n281), .D1(n280), .S(ps_ptr[3]), .Y(n282) );
  AO2222XL U591 ( .A(n388), .B(r_sar_en[9]), .C(n387), .D(r_sar_en[11]), .E(
        n386), .F(r_sar_en[13]), .G(n385), .H(r_sar_en[15]), .Y(n280) );
  AO2222XL U592 ( .A(n387), .B(r_sar_en[3]), .C(n384), .D(r_sar_en[1]), .E(
        n386), .F(r_sar_en[5]), .G(n385), .H(r_sar_en[7]), .Y(n281) );
  MUX2X1 U593 ( .D0(n382), .D1(n381), .S(ps_ptr[3]), .Y(n383) );
  AO2222XL U594 ( .A(r_dac_en[8]), .B(n388), .C(r_dac_en[10]), .D(n387), .E(
        r_dac_en[12]), .F(n386), .G(r_dac_en[14]), .H(n385), .Y(n381) );
  AO2222XL U595 ( .A(r_dac_en[2]), .B(n387), .C(r_dac_en[0]), .D(n384), .E(
        r_dac_en[4]), .F(n386), .G(r_dac_en[6]), .H(n385), .Y(n382) );
  NAND32XL U596 ( .B(pos_dacis[12]), .C(n450), .A(n446), .Y(n474) );
  AO2222XL U597 ( .A(r_dac_en[9]), .B(n388), .C(r_dac_en[11]), .D(n387), .E(
        r_dac_en[13]), .F(n386), .G(r_dac_en[15]), .H(n385), .Y(n389) );
  AO2222XL U598 ( .A(r_dac_en[3]), .B(n387), .C(r_dac_en[1]), .D(n384), .E(
        r_dac_en[5]), .F(n386), .G(r_dac_en[7]), .H(n385), .Y(n390) );
  INVX1 U599 ( .A(pos_dacis[5]), .Y(n412) );
  INVX1 U600 ( .A(pos_dacis[4]), .Y(n410) );
  INVX1 U601 ( .A(pos_dacis[6]), .Y(n418) );
  INVX1 U602 ( .A(pos_dacis[7]), .Y(n447) );
  NAND21X1 U603 ( .B(pos_dacis[9]), .A(n424), .Y(n429) );
  INVX1 U604 ( .A(pos_dacis[8]), .Y(n424) );
  OR2X1 U605 ( .A(pos_dacis[11]), .B(pos_dacis[10]), .Y(n440) );
  NAND21X1 U606 ( .B(pos_dacis[13]), .A(n435), .Y(n457) );
  INVX1 U607 ( .A(pos_dacis[12]), .Y(n435) );
  INVX1 U608 ( .A(pos_dacis[13]), .Y(n473) );
  NOR43XL U609 ( .B(n224), .C(n223), .D(n222), .A(n221), .Y(n234) );
  NAND21X1 U610 ( .B(n248), .A(r_sar_en[12]), .Y(n223) );
  NAND21X1 U611 ( .B(n247), .A(r_sar_en[13]), .Y(n224) );
  NAND21X1 U612 ( .B(n246), .A(r_sar_en[14]), .Y(n222) );
  NAND2XL U613 ( .A(r_sar_en[11]), .B(dacv_wr[11]), .Y(n225) );
  NOR21XL U614 ( .B(app_dacis[11]), .A(n83), .Y(o_daci_sel[11]) );
  NOR21XL U615 ( .B(app_dacis[5]), .A(n83), .Y(o_daci_sel[5]) );
  NOR21XL U616 ( .B(app_dacis[2]), .A(n83), .Y(o_daci_sel[2]) );
  NOR21XL U617 ( .B(app_dacis[12]), .A(n83), .Y(o_daci_sel[12]) );
  NOR21XL U618 ( .B(app_dacis[14]), .A(n83), .Y(o_daci_sel[14]) );
  NOR21XL U619 ( .B(app_dacis[4]), .A(n83), .Y(o_daci_sel[4]) );
  NOR21XL U620 ( .B(app_dacis[6]), .A(n83), .Y(o_daci_sel[6]) );
  NOR21XL U621 ( .B(app_dacis[7]), .A(n83), .Y(o_daci_sel[7]) );
  NOR21XL U622 ( .B(app_dacis[16]), .A(n83), .Y(o_daci_sel[16]) );
  NOR21XL U623 ( .B(app_dacis[1]), .A(n83), .Y(o_daci_sel[1]) );
  NOR21XL U624 ( .B(app_dacis[3]), .A(r_comp_opt[0]), .Y(o_daci_sel[3]) );
  NOR21XL U625 ( .B(app_dacis[13]), .A(r_comp_opt[0]), .Y(o_daci_sel[13]) );
  NOR21XL U626 ( .B(app_dacis[15]), .A(r_comp_opt[0]), .Y(o_daci_sel[15]) );
  NOR21XL U627 ( .B(app_dacis[9]), .A(r_comp_opt[0]), .Y(o_daci_sel[9]) );
  NOR21XL U628 ( .B(app_dacis[8]), .A(r_comp_opt[0]), .Y(o_daci_sel[8]) );
  NOR21XL U629 ( .B(app_dacis[0]), .A(r_comp_opt[0]), .Y(o_daci_sel[0]) );
  NOR21XL U630 ( .B(app_dacis[17]), .A(r_comp_opt[0]), .Y(o_daci_sel[17]) );
  NAND21X1 U631 ( .B(n231), .A(n230), .Y(n232) );
  AO2222XL U632 ( .A(dacv_wr[7]), .B(r_sar_en[7]), .C(dacv_wr[6]), .D(
        r_sar_en[6]), .E(dacv_wr[17]), .F(r_sar_en[17]), .G(dacv_wr[5]), .H(
        r_sar_en[5]), .Y(n231) );
  NOR21XL U633 ( .B(app_dacis[10]), .A(r_comp_opt[0]), .Y(o_daci_sel[10]) );
  INVX1 U634 ( .A(pos_dacis[14]), .Y(n458) );
  NAND21X1 U635 ( .B(pos_dacis[15]), .A(n458), .Y(n467) );
  AO21XL U636 ( .B(N1275), .C(n491), .A(n490), .Y(o_dacv[27]) );
  NAND21X1 U637 ( .B(pos_dacis[17]), .A(n463), .Y(n479) );
  AO21XL U638 ( .B(N1308), .C(n500), .A(n499), .Y(o_dacv[51]) );
  AO21XL U639 ( .B(N1253), .C(n485), .A(n484), .Y(o_dacv[11]) );
  NAND21X1 U640 ( .B(n259), .A(r_sar_en[3]), .Y(n229) );
  NAND21X1 U641 ( .B(n257), .A(r_sar_en[4]), .Y(n228) );
  NAND21X1 U642 ( .B(n261), .A(r_sar_en[2]), .Y(n227) );
  INVX1 U643 ( .A(pos_dacis[16]), .Y(n463) );
  AO21XL U644 ( .B(N1254), .C(n485), .A(n484), .Y(o_dacv[12]) );
  AO21XL U645 ( .B(N1276), .C(n491), .A(n490), .Y(o_dacv[28]) );
  MUX2XL U646 ( .D0(n27), .D1(o_dactl[5]), .S(n36), .Y(ps_md4ch) );
  AO21XL U647 ( .B(N1310), .C(n500), .A(n499), .Y(o_dacv[53]) );
  AO21XL U648 ( .B(N1309), .C(n500), .A(n499), .Y(o_dacv[52]) );
  AO21XL U649 ( .B(N1321), .C(n503), .A(n502), .Y(o_dacv[61]) );
  AO21XL U650 ( .B(N1320), .C(n503), .A(n502), .Y(o_dacv[60]) );
  NAND4X1 U651 ( .A(o_dactl[6]), .B(n199), .C(n200), .D(n201), .Y(n149) );
  NOR2X1 U652 ( .A(n202), .B(n203), .Y(n201) );
  XNOR2XL U653 ( .A(x_daclsb[3]), .B(n154), .Y(n200) );
  XNOR2XL U654 ( .A(n161), .B(x_daclsb[5]), .Y(n202) );
  XNOR2XL U655 ( .A(n157), .B(x_daclsb[4]), .Y(n203) );
  AO21XL U656 ( .B(N1255), .C(n485), .A(n484), .Y(o_dacv[13]) );
  AO21XL U657 ( .B(N1277), .C(n491), .A(n490), .Y(o_dacv[29]) );
  MUX2AXL U658 ( .D0(r_rpt_v[6]), .D1(net168001), .S(n151), .Y(n219) );
  AO21XL U659 ( .B(N1257), .C(n485), .A(n484), .Y(o_dacv[15]) );
  AO21XL U660 ( .B(N1278), .C(n491), .A(n490), .Y(o_dacv[30]) );
  AO21XL U661 ( .B(N1279), .C(n491), .A(n490), .Y(o_dacv[31]) );
  ENOX1 U662 ( .A(n535), .B(n538), .C(r_rpt_v[8]), .D(n538), .Y(wda[6]) );
  ENOX1 U663 ( .A(n538), .B(n534), .C(r_rpt_v[9]), .D(n538), .Y(wda[7]) );
  AO21XL U664 ( .B(N1312), .C(n500), .A(n499), .Y(o_dacv[55]) );
  AO21XL U665 ( .B(N1311), .C(n500), .A(n499), .Y(o_dacv[54]) );
  AO21XL U666 ( .B(N1323), .C(n503), .A(n502), .Y(o_dacv[63]) );
  MUX2AXL U667 ( .D0(r_rpt_v[7]), .D1(n25), .S(n151), .Y(n220) );
  MUX2AXL U668 ( .D0(r_rpt_v[2]), .D1(n30), .S(n151), .Y(n215) );
  MUX2AXL U669 ( .D0(r_rpt_v[4]), .D1(n20), .S(n151), .Y(n217) );
  MUX2AXL U670 ( .D0(r_rpt_v[5]), .D1(n238), .S(n151), .Y(n218) );
  AO21XL U671 ( .B(N1256), .C(n485), .A(n484), .Y(o_dacv[14]) );
  MUX2X1 U672 ( .D0(n21), .D1(x_daclsb[2]), .S(n537), .Y(wdlsb[2]) );
  MUX2X1 U673 ( .D0(net167900), .D1(x_daclsb[3]), .S(n537), .Y(wdlsb[3]) );
  MUX2X1 U674 ( .D0(n26), .D1(x_daclsb[4]), .S(n537), .Y(wdlsb[4]) );
  MUX2X1 U675 ( .D0(n23), .D1(r_rpt_v[1]), .S(n537), .Y(wdlsb[1]) );
  MUX2AXL U676 ( .D0(r_rpt_v[3]), .D1(n22), .S(n151), .Y(n216) );
  ENOX1 U677 ( .A(n535), .B(n537), .C(n537), .D(x_daclsb[5]), .Y(wdlsb[5]) );
  MUX4X1 U678 ( .D0(r_sar_en[2]), .D1(r_sar_en[3]), .D2(r_sar_en[10]), .D3(
        r_sar_en[11]), .S0(n146), .S1(n144), .Y(n133) );
  MUX4X1 U679 ( .D0(r_sar_en[4]), .D1(r_sar_en[5]), .D2(r_sar_en[12]), .D3(
        r_sar_en[13]), .S0(n146), .S1(n144), .Y(n134) );
  MUX4X1 U680 ( .D0(r_sar_en[0]), .D1(r_sar_en[1]), .D2(r_sar_en[8]), .D3(
        r_sar_en[9]), .S0(n146), .S1(n144), .Y(n135) );
  MUX4X1 U681 ( .D0(r_sar_en[6]), .D1(r_sar_en[7]), .D2(r_sar_en[14]), .D3(
        r_sar_en[15]), .S0(n146), .S1(n144), .Y(n132) );
  AO222X1 U682 ( .A(n283), .B(n344), .C(n285), .D(n345), .E(r_dac1v[4]), .F(
        n539), .Y(o_dac1[4]) );
  NAND4X1 U683 ( .A(n350), .B(n351), .C(n352), .D(n353), .Y(n344) );
  NAND4X1 U684 ( .A(n346), .B(n347), .C(n348), .D(n349), .Y(n345) );
  AOI22XL U685 ( .A(r_dacvs[10]), .B(n51), .C(r_dacvs[138]), .D(n299), .Y(n350) );
  AO222X1 U686 ( .A(n283), .B(n324), .C(n285), .D(n325), .E(r_dac1v[6]), .F(
        n539), .Y(o_dac1[6]) );
  NAND4X1 U687 ( .A(n330), .B(n331), .C(n332), .D(n333), .Y(n324) );
  NAND4X1 U688 ( .A(n326), .B(n327), .C(n328), .D(n329), .Y(n325) );
  AOI22XL U689 ( .A(r_dacvs[12]), .B(n51), .C(r_dacvs[140]), .D(n80), .Y(n330)
         );
  AO222X1 U690 ( .A(n283), .B(n304), .C(n285), .D(n305), .E(r_dac1v[8]), .F(
        n539), .Y(o_dac1[8]) );
  NAND4X1 U691 ( .A(n310), .B(n311), .C(n312), .D(n313), .Y(n304) );
  NAND4X1 U692 ( .A(n306), .B(n307), .C(n308), .D(n309), .Y(n305) );
  AOI22XL U693 ( .A(r_dacvs[14]), .B(n51), .C(r_dacvs[142]), .D(n80), .Y(n310)
         );
  AO222X1 U694 ( .A(n283), .B(n364), .C(n285), .D(n365), .E(r_dac1v[2]), .F(
        n539), .Y(o_dac1[2]) );
  NAND4X1 U695 ( .A(n370), .B(n371), .C(n372), .D(n373), .Y(n364) );
  NAND4X1 U696 ( .A(n366), .B(n367), .C(n368), .D(n369), .Y(n365) );
  AOI22XL U697 ( .A(r_dacvs[8]), .B(n51), .C(r_dacvs[136]), .D(n80), .Y(n370)
         );
  AO222X1 U698 ( .A(n283), .B(n354), .C(n285), .D(n355), .E(r_dac1v[3]), .F(
        n539), .Y(o_dac1[3]) );
  NAND4X1 U699 ( .A(n360), .B(n361), .C(n362), .D(n363), .Y(n354) );
  NAND4X1 U700 ( .A(n356), .B(n357), .C(n358), .D(n359), .Y(n355) );
  AOI22XL U701 ( .A(r_dacvs[9]), .B(n51), .C(r_dacvs[137]), .D(n80), .Y(n360)
         );
  AO222X1 U702 ( .A(n283), .B(n314), .C(n285), .D(n315), .E(r_dac1v[7]), .F(
        n539), .Y(o_dac1[7]) );
  NAND4X1 U703 ( .A(n320), .B(n321), .C(n322), .D(n323), .Y(n314) );
  NAND4X1 U704 ( .A(n316), .B(n317), .C(n318), .D(n319), .Y(n315) );
  AOI22XL U705 ( .A(r_dacvs[13]), .B(n51), .C(r_dacvs[141]), .D(n80), .Y(n320)
         );
  AO222X1 U706 ( .A(n283), .B(n284), .C(n285), .D(n286), .E(r_dac1v[9]), .F(
        n539), .Y(o_dac1[9]) );
  NAND4X1 U707 ( .A(n300), .B(n301), .C(n302), .D(n303), .Y(n284) );
  NAND4X1 U708 ( .A(n287), .B(n288), .C(n289), .D(n290), .Y(n286) );
  AOI22X1 U709 ( .A(r_dacvs[15]), .B(n51), .C(r_dacvs[143]), .D(n80), .Y(n300)
         );
  AO222X1 U710 ( .A(n283), .B(n334), .C(n285), .D(n335), .E(r_dac1v[5]), .F(
        n539), .Y(o_dac1[5]) );
  NAND4X1 U711 ( .A(n340), .B(n341), .C(n342), .D(n343), .Y(n334) );
  NAND4X1 U712 ( .A(n336), .B(n337), .C(n338), .D(n339), .Y(n335) );
  AOI22XL U713 ( .A(r_dacvs[11]), .B(n51), .C(r_dacvs[139]), .D(n299), .Y(n340) );
  MUX2BXL U714 ( .D0(n121), .D1(n122), .S(n162), .Y(n120) );
  MUX4X1 U715 ( .D0(n135), .D1(n133), .D2(n134), .D3(n132), .S0(n156), .S1(
        n158), .Y(n121) );
  MUX2IX1 U716 ( .D0(r_sar_en[16]), .D1(r_sar_en[17]), .S(n145), .Y(n122) );
  AO22X1 U717 ( .A(r_dac1v[0]), .B(n539), .C(x_daclsb[0]), .D(n379), .Y(
        o_dac1[0]) );
  AO22X1 U718 ( .A(r_dac1v[1]), .B(n539), .C(x_daclsb[1]), .D(n379), .Y(
        o_dac1[1]) );
  AOI222XL U719 ( .A(r_dacvs[112]), .B(n60), .C(r_dacvs[80]), .D(n68), .E(
        r_dacvs[96]), .F(n78), .Y(n369) );
  AOI222XL U720 ( .A(r_dacvs[120]), .B(n61), .C(r_dacvs[88]), .D(n69), .E(
        r_dacvs[104]), .F(n79), .Y(n373) );
  AOI222XL U721 ( .A(r_dacvs[113]), .B(n60), .C(r_dacvs[81]), .D(n68), .E(
        r_dacvs[97]), .F(n78), .Y(n359) );
  AOI222XL U722 ( .A(r_dacvs[121]), .B(n61), .C(r_dacvs[89]), .D(n69), .E(
        r_dacvs[105]), .F(n79), .Y(n363) );
  AOI222XL U723 ( .A(r_dacvs[114]), .B(n60), .C(r_dacvs[82]), .D(n68), .E(
        r_dacvs[98]), .F(n78), .Y(n349) );
  AOI222XL U724 ( .A(r_dacvs[122]), .B(n61), .C(r_dacvs[90]), .D(n69), .E(
        r_dacvs[106]), .F(n79), .Y(n353) );
  AOI222XL U725 ( .A(r_dacvs[115]), .B(n60), .C(r_dacvs[83]), .D(n68), .E(
        r_dacvs[99]), .F(n78), .Y(n339) );
  AOI222XL U726 ( .A(r_dacvs[123]), .B(n61), .C(r_dacvs[91]), .D(n69), .E(
        r_dacvs[107]), .F(n79), .Y(n343) );
  AOI222XL U727 ( .A(r_dacvs[116]), .B(n60), .C(r_dacvs[84]), .D(n68), .E(
        r_dacvs[100]), .F(n78), .Y(n329) );
  AOI222XL U728 ( .A(r_dacvs[124]), .B(n61), .C(r_dacvs[92]), .D(n69), .E(
        r_dacvs[108]), .F(n79), .Y(n333) );
  AOI222XL U729 ( .A(r_dacvs[117]), .B(n61), .C(r_dacvs[85]), .D(n69), .E(
        r_dacvs[101]), .F(n79), .Y(n319) );
  AOI222XL U730 ( .A(r_dacvs[125]), .B(n61), .C(r_dacvs[93]), .D(n69), .E(
        r_dacvs[109]), .F(n79), .Y(n323) );
  AOI222XL U731 ( .A(r_dacvs[118]), .B(n60), .C(r_dacvs[86]), .D(n68), .E(
        r_dacvs[102]), .F(n78), .Y(n309) );
  AOI222XL U732 ( .A(r_dacvs[126]), .B(n61), .C(r_dacvs[94]), .D(n69), .E(
        r_dacvs[110]), .F(n79), .Y(n313) );
  AOI222XL U733 ( .A(r_dacvs[119]), .B(n61), .C(r_dacvs[87]), .D(n69), .E(
        r_dacvs[103]), .F(n79), .Y(n290) );
  AOI222XL U734 ( .A(r_dacvs[127]), .B(n61), .C(r_dacvs[95]), .D(n69), .E(
        r_dacvs[111]), .F(n79), .Y(n303) );
  AOI22XL U735 ( .A(r_dacvs[64]), .B(n54), .C(r_dacvs[16]), .D(n76), .Y(n368)
         );
  AOI22XL U736 ( .A(r_dacvs[65]), .B(n54), .C(r_dacvs[17]), .D(n76), .Y(n358)
         );
  AOI22XL U737 ( .A(r_dacvs[66]), .B(n54), .C(r_dacvs[18]), .D(n76), .Y(n348)
         );
  AOI22XL U738 ( .A(r_dacvs[67]), .B(n54), .C(r_dacvs[19]), .D(n76), .Y(n338)
         );
  AOI22XL U739 ( .A(r_dacvs[68]), .B(n54), .C(r_dacvs[20]), .D(n76), .Y(n328)
         );
  AOI22XL U740 ( .A(r_dacvs[69]), .B(n55), .C(r_dacvs[21]), .D(n77), .Y(n318)
         );
  AOI22XL U741 ( .A(r_dacvs[70]), .B(n54), .C(r_dacvs[22]), .D(n76), .Y(n308)
         );
  AOI22X1 U742 ( .A(r_dacvs[71]), .B(n55), .C(r_dacvs[23]), .D(n77), .Y(n289)
         );
  AOI22XL U743 ( .A(r_dacvs[32]), .B(n58), .C(r_dacvs[48]), .D(n66), .Y(n367)
         );
  AOI22XL U744 ( .A(r_dacvs[33]), .B(n58), .C(r_dacvs[49]), .D(n66), .Y(n357)
         );
  AOI22XL U745 ( .A(r_dacvs[34]), .B(n58), .C(r_dacvs[50]), .D(n66), .Y(n347)
         );
  AOI22X1 U746 ( .A(r_dacvs[36]), .B(n59), .C(r_dacvs[52]), .D(n67), .Y(n327)
         );
  AOI22X1 U747 ( .A(r_dacvs[37]), .B(n59), .C(r_dacvs[53]), .D(n67), .Y(n317)
         );
  AOI22X1 U748 ( .A(r_dacvs[38]), .B(n59), .C(r_dacvs[54]), .D(n67), .Y(n307)
         );
  AOI22X1 U749 ( .A(r_dacvs[39]), .B(n59), .C(r_dacvs[55]), .D(n67), .Y(n288)
         );
  AOI22XL U750 ( .A(r_dacvs[72]), .B(n55), .C(r_dacvs[24]), .D(n77), .Y(n372)
         );
  AOI22XL U751 ( .A(r_dacvs[73]), .B(n55), .C(r_dacvs[25]), .D(n77), .Y(n362)
         );
  AOI22XL U752 ( .A(r_dacvs[74]), .B(n55), .C(r_dacvs[26]), .D(n77), .Y(n352)
         );
  AOI22XL U753 ( .A(r_dacvs[75]), .B(n55), .C(r_dacvs[27]), .D(n77), .Y(n342)
         );
  AOI22XL U754 ( .A(r_dacvs[76]), .B(n55), .C(r_dacvs[28]), .D(n77), .Y(n332)
         );
  AOI22XL U755 ( .A(r_dacvs[77]), .B(n55), .C(r_dacvs[29]), .D(n77), .Y(n322)
         );
  AOI22XL U756 ( .A(r_dacvs[78]), .B(n55), .C(r_dacvs[30]), .D(n77), .Y(n312)
         );
  AOI22X1 U757 ( .A(r_dacvs[79]), .B(n55), .C(r_dacvs[31]), .D(n77), .Y(n302)
         );
  AOI22XL U758 ( .A(r_dacvs[40]), .B(n59), .C(r_dacvs[56]), .D(n67), .Y(n371)
         );
  AOI22XL U759 ( .A(r_dacvs[41]), .B(n59), .C(r_dacvs[57]), .D(n67), .Y(n361)
         );
  AOI22XL U760 ( .A(r_dacvs[42]), .B(n58), .C(r_dacvs[58]), .D(n66), .Y(n351)
         );
  AOI22X1 U761 ( .A(r_dacvs[44]), .B(n59), .C(r_dacvs[60]), .D(n67), .Y(n331)
         );
  AOI22X1 U762 ( .A(r_dacvs[45]), .B(n59), .C(r_dacvs[61]), .D(n67), .Y(n321)
         );
  AOI22X1 U763 ( .A(r_dacvs[46]), .B(n59), .C(r_dacvs[62]), .D(n67), .Y(n311)
         );
  AOI22X1 U764 ( .A(r_dacvs[47]), .B(n59), .C(r_dacvs[63]), .D(n67), .Y(n301)
         );
  AOI22XL U765 ( .A(r_dacvs[0]), .B(n50), .C(r_dacvs[128]), .D(n299), .Y(n366)
         );
  AOI22XL U766 ( .A(r_dacvs[1]), .B(n50), .C(r_dacvs[129]), .D(n299), .Y(n356)
         );
  AOI22XL U767 ( .A(r_dacvs[2]), .B(n50), .C(r_dacvs[130]), .D(n299), .Y(n346)
         );
  AOI22XL U768 ( .A(r_dacvs[3]), .B(n50), .C(r_dacvs[131]), .D(n299), .Y(n336)
         );
  AOI22XL U769 ( .A(r_dacvs[4]), .B(n50), .C(r_dacvs[132]), .D(n299), .Y(n326)
         );
  AOI22XL U770 ( .A(r_dacvs[5]), .B(n51), .C(r_dacvs[133]), .D(n299), .Y(n316)
         );
  AOI22XL U771 ( .A(r_dacvs[6]), .B(n50), .C(r_dacvs[134]), .D(n299), .Y(n306)
         );
  AOI22X1 U772 ( .A(r_dacvs[7]), .B(n51), .C(r_dacvs[135]), .D(n80), .Y(n287)
         );
  NAND42X1 U773 ( .C(r_dac_en[2]), .D(n214), .A(n213), .B(n212), .Y(n159) );
  NAND21X1 U774 ( .B(r_dac_en[4]), .A(n98), .Y(n214) );
  NOR32XL U775 ( .B(n124), .C(n123), .A(n207), .Y(n213) );
  NOR43XL U776 ( .B(n211), .C(n210), .D(n209), .A(n208), .Y(n212) );
  OR4X1 U777 ( .A(r_dac_en[1]), .B(r_dac_en[0]), .C(r_dac_en[13]), .D(
        r_dac_en[14]), .Y(n208) );
  OR2X1 U778 ( .A(r_dac_en[6]), .B(r_dac_en[5]), .Y(n207) );
  INVX1 U779 ( .A(r_dac_en[11]), .Y(n211) );
  INVX1 U780 ( .A(r_dac_en[10]), .Y(n209) );
  INVX1 U781 ( .A(r_dac_en[12]), .Y(n210) );
  NOR3XL U782 ( .A(r_dac_en[15]), .B(r_dac_en[16]), .C(r_dac_en[17]), .Y(n123)
         );
  NOR3XL U783 ( .A(r_dac_en[7]), .B(r_dac_en[8]), .C(r_dac_en[9]), .Y(n124) );
  MUX4X1 U784 ( .D0(n140), .D1(n138), .D2(n139), .D3(n137), .S0(n156), .S1(
        n158), .Y(n141) );
  MUX4X1 U785 ( .D0(o_dat[4]), .D1(o_dat[5]), .D2(o_dat[12]), .D3(o_dat[13]), 
        .S0(n145), .S1(n144), .Y(n139) );
  MUX4X1 U786 ( .D0(o_dat[6]), .D1(o_dat[7]), .D2(o_dat[14]), .D3(o_dat[15]), 
        .S0(n146), .S1(n144), .Y(n137) );
  MUX4X1 U787 ( .D0(o_dat[2]), .D1(o_dat[3]), .D2(o_dat[10]), .D3(o_dat[11]), 
        .S0(n145), .S1(n144), .Y(n138) );
  MUX4X1 U788 ( .D0(o_dat[0]), .D1(o_dat[1]), .D2(o_dat[8]), .D3(o_dat[9]), 
        .S0(n146), .S1(n144), .Y(n140) );
  NOR42XL U789 ( .C(o_dactl[1]), .D(dacyc_done), .A(n120), .B(n152), .Y(tochg)
         );
  XNOR2XL U790 ( .A(syn_comp[1]), .B(N859), .Y(n152) );
  MUX2X1 U791 ( .D0(n141), .D1(n136), .S(n162), .Y(N859) );
  MUX2X1 U792 ( .D0(o_dat[16]), .D1(o_dat[17]), .S(n145), .Y(n136) );
  MUX4X1 U793 ( .D0(r_dac_en[2]), .D1(r_dac_en[3]), .D2(r_dac_en[10]), .D3(
        r_dac_en[11]), .S0(n146), .S1(n143), .Y(n129) );
  MUX4X1 U794 ( .D0(r_dac_en[4]), .D1(r_dac_en[5]), .D2(r_dac_en[12]), .D3(
        r_dac_en[13]), .S0(n146), .S1(n144), .Y(n130) );
  MUX4X1 U795 ( .D0(r_dac_en[0]), .D1(r_dac_en[1]), .D2(r_dac_en[8]), .D3(
        r_dac_en[9]), .S0(n146), .S1(n144), .Y(n131) );
  MUX4X1 U796 ( .D0(r_dac_en[6]), .D1(r_dac_en[7]), .D2(r_dac_en[14]), .D3(
        r_dac_en[15]), .S0(n146), .S1(n143), .Y(n128) );
  MUX2BXL U797 ( .D0(n126), .D1(n127), .S(n162), .Y(n125) );
  MUX4X1 U798 ( .D0(n131), .D1(n129), .D2(n130), .D3(n128), .S0(n156), .S1(
        n158), .Y(n126) );
  MUX2IX1 U799 ( .D0(r_dac_en[16]), .D1(r_dac_en[17]), .S(n145), .Y(n127) );
  ENOX1 U800 ( .A(n548), .B(n165), .C(o_dat[2]), .D(n548), .Y(datcmp[2]) );
  ENOX1 U801 ( .A(n552), .B(n165), .C(o_dat[3]), .D(n552), .Y(datcmp[3]) );
  ENOX1 U802 ( .A(n544), .B(n165), .C(o_dat[4]), .D(n544), .Y(datcmp[4]) );
  ENOX1 U803 ( .A(n557), .B(n165), .C(o_dat[5]), .D(n557), .Y(datcmp[5]) );
  ENOX1 U804 ( .A(n549), .B(n165), .C(o_dat[6]), .D(n549), .Y(datcmp[6]) );
  ENOX1 U805 ( .A(n553), .B(n165), .C(o_dat[7]), .D(n553), .Y(datcmp[7]) );
  ENOX1 U806 ( .A(n545), .B(n165), .C(o_dat[8]), .D(n545), .Y(datcmp[8]) );
  ENOX1 U807 ( .A(n558), .B(n165), .C(o_dat[9]), .D(n558), .Y(datcmp[9]) );
  ENOX1 U808 ( .A(n541), .B(n164), .C(o_dat[0]), .D(n541), .Y(datcmp[0]) );
  ENOX1 U809 ( .A(n556), .B(n164), .C(o_dat[1]), .D(n556), .Y(datcmp[1]) );
  ENOX1 U810 ( .A(n546), .B(n164), .C(o_dat[10]), .D(n546), .Y(datcmp[10]) );
  ENOX1 U811 ( .A(n550), .B(n164), .C(o_dat[11]), .D(n550), .Y(datcmp[11]) );
  ENOX1 U812 ( .A(n542), .B(n164), .C(o_dat[12]), .D(n542), .Y(datcmp[12]) );
  ENOX1 U813 ( .A(n554), .B(n164), .C(o_dat[13]), .D(n554), .Y(datcmp[13]) );
  ENOX1 U814 ( .A(n547), .B(n164), .C(o_dat[14]), .D(n547), .Y(datcmp[14]) );
  ENOX1 U815 ( .A(n551), .B(n164), .C(o_dat[15]), .D(n551), .Y(datcmp[15]) );
  ENOX1 U816 ( .A(n543), .B(n164), .C(o_dat[16]), .D(n543), .Y(datcmp[16]) );
  ENOX1 U817 ( .A(n555), .B(n164), .C(o_dat[17]), .D(n555), .Y(datcmp[17]) );
  INVX1 U818 ( .A(syn_comp[1]), .Y(n164) );
  INVX1 U819 ( .A(syn_comp[1]), .Y(n165) );
  BUFXL U820 ( .A(net167900), .Y(net156831) );
  INVXL U821 ( .A(dacv_wr[14]), .Y(n246) );
  INVXL U822 ( .A(dacv_wr[15]), .Y(n245) );
  AO22XL U823 ( .A(dacv_wr[16]), .B(r_sar_en[16]), .C(dacv_wr[15]), .D(
        r_sar_en[15]), .Y(n221) );
  INVXL U824 ( .A(dacv_wr[10]), .Y(n251) );
  NAND2XL U825 ( .A(r_sar_en[10]), .B(dacv_wr[10]), .Y(n226) );
  MUX2XL U826 ( .D0(n32), .D1(r_rpt_v[0]), .S(n537), .Y(wdlsb[0]) );
  AND2XL U827 ( .A(n32), .B(r_wr[4]), .Y(clrsta[0]) );
  NAND6XL U828 ( .A(r_wdat[6]), .B(n32), .C(n240), .D(n20), .E(n238), .F(n25), 
        .Y(n239) );
  NAND32XL U829 ( .B(n101), .C(net145949), .A(net169040), .Y(n269) );
  GEN2X1 U830 ( .D(n445), .E(n444), .C(n443), .B(n442), .A(n441), .Y(n469) );
endmodule


module dacmux_a0_DW01_add_17 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1XL U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_16 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1XL U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_15 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_14 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1XL U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_13 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1XL U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_12 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2XL U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_11 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2XL U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_10 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2XL U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_9 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2XL U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  INVX8 U1 ( .A(n1), .Y(carry[1]) );
  XOR2X4 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(n1) );
  XOR2XL U4 ( .A(A[1]), .B(B[1]), .Y(n2) );
  XOR2XL U5 ( .A(n2), .B(carry[1]), .Y(SUM[1]) );
  NAND2XL U6 ( .A(A[1]), .B(B[1]), .Y(n3) );
  NAND2XL U7 ( .A(A[1]), .B(carry[1]), .Y(n4) );
  NAND2XL U8 ( .A(B[1]), .B(carry[1]), .Y(n5) );
  NAND3X1 U9 ( .A(n3), .B(n4), .C(n5), .Y(carry[2]) );
  XOR2X1 U10 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_6 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  INVX1 U1 ( .A(B[8]), .Y(n1) );
  XNOR2X1 U2 ( .A(n1), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_5 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  INVX1 U1 ( .A(B[8]), .Y(n1) );
  XNOR2X1 U2 ( .A(n1), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  XOR3X1 U1 ( .A(carry[3]), .B(B[3]), .C(A[3]), .Y(SUM[3]) );
  NAND2X1 U2 ( .A(carry[3]), .B(B[3]), .Y(n1) );
  NAND2XL U3 ( .A(carry[3]), .B(A[3]), .Y(n2) );
  NAND2X1 U4 ( .A(B[3]), .B(A[3]), .Y(n3) );
  NAND3X1 U5 ( .A(n3), .B(n2), .C(n1), .Y(carry[4]) );
  XOR2X1 U6 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  NAND3X1 U1 ( .A(n10), .B(n9), .C(n8), .Y(carry[5]) );
  NAND3X1 U2 ( .A(n1), .B(n2), .C(n3), .Y(carry[2]) );
  XOR2X1 U3 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  NAND3X1 U4 ( .A(n5), .B(n6), .C(n7), .Y(carry[3]) );
  XOR3XL U5 ( .A(A[1]), .B(B[1]), .C(carry[1]), .Y(SUM[1]) );
  NAND2X1 U6 ( .A(A[1]), .B(B[1]), .Y(n1) );
  NAND2XL U7 ( .A(A[1]), .B(carry[1]), .Y(n2) );
  NAND2XL U8 ( .A(B[1]), .B(carry[1]), .Y(n3) );
  XOR2XL U9 ( .A(A[2]), .B(B[2]), .Y(n4) );
  XOR2XL U10 ( .A(n4), .B(carry[2]), .Y(SUM[2]) );
  NAND2XL U11 ( .A(A[2]), .B(B[2]), .Y(n5) );
  NAND2X1 U12 ( .A(A[2]), .B(carry[2]), .Y(n6) );
  NAND2X1 U13 ( .A(B[2]), .B(carry[2]), .Y(n7) );
  XOR3X1 U14 ( .A(carry[4]), .B(B[4]), .C(A[4]), .Y(SUM[4]) );
  NAND2X1 U15 ( .A(carry[4]), .B(B[4]), .Y(n8) );
  NAND2XL U16 ( .A(carry[4]), .B(A[4]), .Y(n9) );
  NAND2X1 U17 ( .A(B[4]), .B(A[4]), .Y(n10) );
endmodule


module dacmux_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  FAD1X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(1'b0), .CO(carry[1]), .SO(SUM[0]) );
  INVX1 U1 ( .A(B[8]), .Y(n1) );
  XNOR2X1 U2 ( .A(n1), .B(carry[8]), .Y(SUM[8]) );
endmodule


module glreg_WIDTH2_0 ( clk, arstz, we, wdat, rdat );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we;
  wire   n1, n4, n5;

  DFFRQX1 mem_reg_0_ ( .D(n5), .C(clk), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(n4), .C(clk), .XR(arstz), .Q(rdat[1]) );
  INVXL U2 ( .A(we), .Y(n1) );
  AO22XL U3 ( .A(wdat[1]), .B(we), .C(rdat[1]), .D(n1), .Y(n4) );
  AO22XL U4 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(n1), .Y(n5) );
endmodule


module glreg_WIDTH2_1 ( clk, arstz, we, wdat, rdat );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we;
  wire   n10, n11, n1, n5, n7, n8, n9;

  DFFRQX1 mem_reg_0_ ( .D(n9), .C(clk), .XR(arstz), .Q(n11) );
  DFFRQX1 mem_reg_1_ ( .D(n8), .C(clk), .XR(arstz), .Q(n10) );
  INVXL U2 ( .A(n10), .Y(n1) );
  INVXL U3 ( .A(n1), .Y(rdat[1]) );
  INVXL U4 ( .A(n11), .Y(n5) );
  INVXL U5 ( .A(n5), .Y(rdat[0]) );
  INVXL U6 ( .A(we), .Y(n7) );
  AO22XL U7 ( .A(wdat[1]), .B(we), .C(n10), .D(n7), .Y(n8) );
  AO22XL U8 ( .A(we), .B(wdat[0]), .C(n11), .D(n7), .Y(n9) );
endmodule


module glreg_a0_26 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9717;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_26 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9717), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9717), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9717), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9717), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9717), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9717), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9717), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9717), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9717), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_27 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9735;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_27 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9735), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9735), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9735), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9735), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9735), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9735), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9735), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9735), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9735), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_28 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9753;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_28 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9753), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9753), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9753), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9753), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9753), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9753), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9753), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9753), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9753), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_29 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9771;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_29 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9771), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9771), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9771), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9771), .XR(arstz), .Q(rdat[6]) );
  DFFRQXX2 mem_reg_0_ ( .D(wdat[0]), .C(net9771), .XR(arstz), .Q(rdat[0]), 
        .XQ() );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9771), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9771), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9771), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9771), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_1 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22;
  wire   [7:0] wd_r;

  glreg_WIDTH8_1 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  INVX1 U2 ( .A(set2[4]), .Y(n14) );
  INVX1 U3 ( .A(set2[5]), .Y(n9) );
  NAND31X1 U4 ( .C(set2[5]), .A(n8), .B(n7), .Y(n1) );
  NOR8XL U5 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .E(clr1[7]), 
        .F(clr1[6]), .G(clr1[5]), .H(clr1[4]), .Y(n4) );
  INVX1 U6 ( .A(set2[6]), .Y(n8) );
  INVX1 U7 ( .A(set2[7]), .Y(n7) );
  INVX1 U8 ( .A(set2[0]), .Y(n10) );
  INVX1 U9 ( .A(set2[2]), .Y(n12) );
  INVX1 U10 ( .A(set2[1]), .Y(n11) );
  INVX1 U11 ( .A(set2[3]), .Y(n13) );
  NAND42X1 U12 ( .C(n6), .D(n5), .A(n4), .B(n3), .Y(upd_r) );
  NOR32XL U13 ( .B(n14), .C(n2), .A(n1), .Y(n3) );
  NAND21X1 U14 ( .B(set2[3]), .A(n12), .Y(n6) );
  NAND21X1 U15 ( .B(set2[1]), .A(n10), .Y(n5) );
  AOI211X1 U16 ( .C(n14), .D(n18), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U17 ( .A(rdat[4]), .Y(n18) );
  AOI211X1 U18 ( .C(n8), .D(n16), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U19 ( .A(rdat[6]), .Y(n16) );
  AOI211X1 U20 ( .C(n7), .D(n15), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U21 ( .A(rdat[7]), .Y(n15) );
  AOI211X1 U22 ( .C(n10), .D(n22), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U23 ( .A(rdat[0]), .Y(n22) );
  AOI211X1 U24 ( .C(n11), .D(n21), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U25 ( .A(rdat[1]), .Y(n21) );
  AOI211X1 U26 ( .C(n12), .D(n20), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U27 ( .A(rdat[2]), .Y(n20) );
  AOI211X1 U28 ( .C(n13), .D(n19), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U29 ( .A(rdat[3]), .Y(n19) );
  AOI211X1 U30 ( .C(n9), .D(n17), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U31 ( .A(rdat[5]), .Y(n17) );
  NOR2X1 U32 ( .A(rdat[1]), .B(n11), .Y(irq[1]) );
  NOR2X1 U33 ( .A(rdat[5]), .B(n9), .Y(irq[5]) );
  NOR2X1 U34 ( .A(rdat[0]), .B(n10), .Y(irq[0]) );
  NOR2X1 U35 ( .A(rdat[4]), .B(n14), .Y(irq[4]) );
  NOR2X1 U36 ( .A(rdat[2]), .B(n12), .Y(irq[2]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n8), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[3]), .B(n13), .Y(irq[3]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n7), .Y(irq[7]) );
  INVX1 U40 ( .A(rst0), .Y(n2) );
endmodule


module glreg_WIDTH8_1 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9789;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9789), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9789), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9789), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9789), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9789), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9789), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9789), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9789), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9789), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_30 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9807;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_30 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9807), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9807), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9807), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9807), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9807), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9807), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9807), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9807), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9807), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_31 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9825;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_31 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9825), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9825), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9825), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9825), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9825), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9825), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9825), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9825), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9825), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_32 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9843;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_32 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9843), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9843), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9843), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9843), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9843), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9843), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9843), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9843), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9843), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_33 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9861;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_33 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9861), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9861), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9861), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9861), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9861), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9861), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9861), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9861), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9861), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_34 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9879;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_34 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9879), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9879), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9879), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9879), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9879), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9879), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9879), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9879), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9879), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_35 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9897;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_35 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9897), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9897), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9897), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9897), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9897), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9897), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9897), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9897), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9897), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_36 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9915;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_36 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9915), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9915), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9915), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9915), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9915), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9915), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9915), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9915), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9915), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_37 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9933;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_37 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9933), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9933), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9933), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9933), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9933), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9933), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9933), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9933), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9933), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_38 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9951;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_38 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9951), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9951), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9951), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9951), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9951), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9951), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9951), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9951), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9951), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_39 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9969;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_39 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9969), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9969), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9969), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9969), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9969), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9969), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9969), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9969), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9969), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_40 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9987;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_40 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9987), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9987), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9987), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9987), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9987), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9987), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9987), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9987), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9987), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_41 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10005;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_41 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10005), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10005), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10005), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10005), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10005), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10005), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10005), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10005), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10005), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_42 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10023;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_42 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10023), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10023), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10023), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10023), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10023), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10023), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10023), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10023), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10023), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_43 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10041;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_43 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10041), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10041), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10041), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10041), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10041), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10041), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10041), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10041), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10041), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_44 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10059;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_44 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10059), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10059), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10059), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10059), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10059), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10059), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10059), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10059), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10059), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_45 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10077;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_45 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10077), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10077), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10077), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10077), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10077), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10077), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10077), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10077), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10077), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_46 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10095;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_46 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10095), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10095), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10095), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10095), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10095), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10095), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10095), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10095), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10095), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_47 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10113;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_47 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10113), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10113), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10113), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10113), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10113), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10113), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10113), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10113), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10113), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_2 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net10131;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10131), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10131), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10131), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10131), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10131), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10131), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10131), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_48 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10149;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_48 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10149), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10149), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10149), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10149), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10149), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10149), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10149), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10149), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10149), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_49 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10167;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_49 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10167), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10167), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10167), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10167), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10167), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10167), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10167), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10167), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10167), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH7_1 ( clk, arstz, we, wdat, rdat );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we;
  wire   net10185;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10185), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10185), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10185), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10185), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10185), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10185), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10185), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10185), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module shmux_00000005_00000012_00000012 ( ps_md4ch, r_comp_swtch, r_semi, 
        r_loop, r_dac_en, wr_dacv, busy, sh_hold, stop, semi_start, auto_start, 
        mxcyc_done, sampl_begn, sampl_done, app_dacis, pos_dacis, cs_ptr, 
        ps_ptr, clk, srstz );
  input [17:0] r_dac_en;
  input [17:0] wr_dacv;
  output [17:0] app_dacis;
  output [17:0] pos_dacis;
  output [4:0] cs_ptr;
  output [4:0] ps_ptr;
  input ps_md4ch, r_comp_swtch, r_semi, r_loop, stop, semi_start, auto_start,
         mxcyc_done, sampl_begn, sampl_done, clk, srstz;
  output busy, sh_hold;
  wire   cs_mux_5_, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958,
         N959, N960, N961, N962, N963, N964, N965, N966, N967, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N994, N995, N996, N997, N998,
         N999, N1136, N1137, N1139, N1140, N1145, N1146, N1147, N1148, N1149,
         N1177, N1178, N1179, N1181, N1185, N1186, N1187, N1219, N1220, N1221,
         N1222, N1227, N1228, N1229, N1230, N1231, N1262, N1263, N1268, N1269,
         N1270, N1271, N1303, N1304, N1309, N1310, N1311, N1312, N1313, N1343,
         N1344, N1345, N1350, N1351, N1352, N1354, N1384, N1385, N1386, N1391,
         N1392, N1393, N1394, N1395, N1425, N1426, N1427, N1433, N1436, N1466,
         N1467, N1468, N1469, N1473, N1474, N1477, N1514, N1515, N1518, N1548,
         N1549, N1550, N1555, N1558, N1559, N1589, N1597, N1599, N1600, N1630,
         N1631, N1632, N1633, N1637, N1638, N1641, N1671, N1672, N1673, N1678,
         N1679, N1682, N1719, N1720, N1761, N1801, N1802, net10203, net10221,
         net10226, n315, n317, n318, n319, n320, n321, n322, n325, n346, n349,
         n350, n366, n369, n383, n386, n405, n408, n438, n440, n441, n442,
         n445, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n671, sub_398_S2_I10_aco_carry_5_, sub_398_S2_I9_aco_carry_5_, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n120, n121, n123, n124,
         n126, n128, n129, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n316, n323, n324, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n347, n348, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n367, n368, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n384, n385, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n406, n407,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n439, n443, n444, n446,
         n459, n460, n531, n532, n543, n544, n555, n556, n579, n580, n591,
         n604, n605, n616, n617, n618, n619, n620, n621, n622, n633, n634,
         n635, n636, n647, n648, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816;
  wire   [16:4] neg_dacis;
  wire   [5:3] sub_398_S2_I14_aco_carry;
  wire   [5:2] sub_398_S2_I11_aco_carry;
  wire   [5:2] sub_398_S2_I7_aco_carry;
  wire   [5:3] sub_398_S2_I6_aco_carry;
  wire   [5:2] sub_398_S2_I5_aco_carry;
  wire   [5:2] sub_398_S2_I4_aco_carry;
  wire   [5:2] sub_398_S2_I3_aco_carry;
  wire   [5:2] sub_398_S2_aco_carry;

  SNPS_CLOCK_GATE_LOW_shmux_00000005_00000012_00000012 clk_gate_neg_dacis_reg ( 
        .CLK(clk), .EN(N949), .ENCLK(net10203), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 clk_gate_r_dacis_reg ( 
        .CLK(clk), .EN(N971), .ENCLK(net10221), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 clk_gate_cs_mux_reg ( 
        .CLK(clk), .EN(N994), .ENCLK(net10226), .TE(1'b0) );
  FAD1X1 sub_398_S2_I7_aco_U2_4 ( .A(N1385), .B(n80), .CI(
        sub_398_S2_I7_aco_carry[4]), .CO(sub_398_S2_I7_aco_carry[5]), .SO(
        N1394) );
  FAD1X1 sub_398_S2_I5_aco_U2_4 ( .A(N1303), .B(n81), .CI(
        sub_398_S2_I5_aco_carry[4]), .CO(sub_398_S2_I5_aco_carry[5]), .SO(
        N1312) );
  FAD1X1 sub_398_S2_I4_aco_U2_4 ( .A(N1262), .B(n1), .CI(
        sub_398_S2_I4_aco_carry[4]), .CO(sub_398_S2_I4_aco_carry[5]), .SO(
        N1271) );
  FAD1X1 sub_398_S2_I3_aco_U2_4 ( .A(N1221), .B(n82), .CI(
        sub_398_S2_I3_aco_carry[4]), .CO(sub_398_S2_I3_aco_carry[5]), .SO(
        N1230) );
  FAD1X1 sub_398_S2_aco_U2_4 ( .A(N1139), .B(n79), .CI(sub_398_S2_aco_carry[4]), .CO(sub_398_S2_aco_carry[5]), .SO(N1148) );
  DFFQX1 cs_mux_reg_3_ ( .D(N998), .C(net10226), .Q(N1179) );
  DFFQX1 cs_mux_reg_4_ ( .D(N999), .C(net10226), .Q(N1181) );
  DFFQX1 cs_mux_reg_0_ ( .D(N995), .C(net10226), .Q(N1185) );
  DFFQX1 cs_mux_reg_2_ ( .D(N997), .C(net10226), .Q(N1178) );
  DFFQX1 cs_mux_reg_1_ ( .D(N996), .C(net10226), .Q(N1177) );
  DFFQX1 r_dacis_reg_17_ ( .D(N989), .C(net10221), .Q(pos_dacis[17]) );
  DFFQX1 r_dacis_reg_16_ ( .D(N988), .C(net10221), .Q(pos_dacis[16]) );
  DFFQX1 r_dacis_reg_15_ ( .D(N987), .C(net10221), .Q(pos_dacis[15]) );
  DFFQX1 r_dacis_reg_14_ ( .D(N986), .C(net10221), .Q(pos_dacis[14]) );
  DFFQX1 r_dacis_reg_12_ ( .D(N984), .C(net10221), .Q(pos_dacis[12]) );
  DFFQX1 cs_mux_reg_5_ ( .D(n671), .C(clk), .Q(cs_mux_5_) );
  DFFQX1 r_dacis_reg_13_ ( .D(N985), .C(net10221), .Q(pos_dacis[13]) );
  DFFQX1 r_dacis_reg_11_ ( .D(N983), .C(net10221), .Q(pos_dacis[11]) );
  DFFQX1 r_dacis_reg_10_ ( .D(N982), .C(net10221), .Q(pos_dacis[10]) );
  DFFQX1 r_dacis_reg_8_ ( .D(N980), .C(net10221), .Q(pos_dacis[8]) );
  DFFQX1 r_dacis_reg_9_ ( .D(N981), .C(net10221), .Q(pos_dacis[9]) );
  DFFQX1 r_dacis_reg_7_ ( .D(N979), .C(net10221), .Q(pos_dacis[7]) );
  DFFQX1 r_dacis_reg_6_ ( .D(N978), .C(net10221), .Q(pos_dacis[6]) );
  DFFQX1 r_dacis_reg_5_ ( .D(N977), .C(net10221), .Q(pos_dacis[5]) );
  DFFQX1 r_dacis_reg_4_ ( .D(N976), .C(net10221), .Q(pos_dacis[4]) );
  DFFQX1 r_dacis_reg_3_ ( .D(N975), .C(net10221), .Q(pos_dacis[3]) );
  DFFQX1 r_dacis_reg_1_ ( .D(N973), .C(net10221), .Q(pos_dacis[1]) );
  DFFQX1 r_dacis_reg_2_ ( .D(N974), .C(net10221), .Q(pos_dacis[2]) );
  DFFNQX4 neg_dacis_reg_9_ ( .D(N959), .XC(net10203), .Q(neg_dacis[9]) );
  DFFNQX4 neg_dacis_reg_16_ ( .D(N966), .XC(net10203), .Q(neg_dacis[16]) );
  DFFNQX4 neg_dacis_reg_4_ ( .D(N954), .XC(net10203), .Q(neg_dacis[4]) );
  DFFNQX4 neg_dacis_reg_12_ ( .D(N962), .XC(net10203), .Q(neg_dacis[12]) );
  DFFNQX4 neg_dacis_reg_13_ ( .D(N963), .XC(net10203), .Q(neg_dacis[13]) );
  DFFNQXX4 neg_dacis_reg_15_ ( .D(N965), .XC(net10203), .Q(n55), .XQ(n56) );
  DFFNQXX4 neg_dacis_reg_5_ ( .D(N955), .XC(net10203), .Q(n53), .XQ(n54) );
  DFFNQXX4 neg_dacis_reg_11_ ( .D(N961), .XC(net10203), .Q(), .XQ(n52) );
  DFFNQXX4 neg_dacis_reg_14_ ( .D(N964), .XC(net10203), .Q(n50), .XQ(n51) );
  DFFNQXX4 neg_dacis_reg_8_ ( .D(N958), .XC(net10203), .Q(n46), .XQ(n47) );
  DFFNQXX4 neg_dacis_reg_0_ ( .D(N950), .XC(net10203), .Q(), .XQ(n45) );
  DFFNQXX4 neg_dacis_reg_2_ ( .D(N952), .XC(net10203), .Q(), .XQ(n44) );
  DFFNQXX4 neg_dacis_reg_6_ ( .D(N956), .XC(net10203), .Q(n42), .XQ(n43) );
  DFFNQXX4 neg_dacis_reg_3_ ( .D(N953), .XC(net10203), .Q(), .XQ(n41) );
  DFFNQXX4 neg_dacis_reg_1_ ( .D(N951), .XC(net10203), .Q(), .XQ(n40) );
  DFFNQXX4 neg_dacis_reg_7_ ( .D(N957), .XC(net10203), .Q(n38), .XQ(n39) );
  DFFNQXX4 neg_dacis_reg_17_ ( .D(N967), .XC(net10203), .Q(n36), .XQ(n37) );
  DFFNQXX4 neg_dacis_reg_10_ ( .D(N960), .XC(net10203), .Q(), .XQ(n35) );
  DFFQX4 r_dacis_reg_0_ ( .D(N972), .C(net10221), .Q(pos_dacis[0]) );
  MUX2X1 U3 ( .D0(n582), .D1(n581), .S(n196), .Y(n195) );
  NAND21X1 U4 ( .B(n218), .A(n445), .Y(n357) );
  NAND6XL U5 ( .A(n288), .B(n287), .C(n286), .D(n285), .E(n8), .F(n136), .Y(
        n324) );
  AND2X1 U6 ( .A(n57), .B(n118), .Y(N963) );
  AND2X1 U7 ( .A(n58), .B(n118), .Y(N962) );
  AND2X1 U8 ( .A(n48), .B(n118), .Y(N954) );
  AND3X1 U9 ( .A(n66), .B(n118), .C(pos_dacis[16]), .Y(N966) );
  AND3X1 U10 ( .A(n556), .B(n118), .C(pos_dacis[9]), .Y(N959) );
  OA21X1 U11 ( .B(n410), .C(n409), .A(n720), .Y(n1) );
  OA22X1 U12 ( .A(N1425), .B(n282), .C(n169), .D(n168), .Y(n2) );
  INVX1 U13 ( .A(n244), .Y(n3) );
  INVX1 U14 ( .A(n245), .Y(n4) );
  INVX1 U15 ( .A(r_dac_en[0]), .Y(n5) );
  INVX1 U16 ( .A(n5), .Y(n6) );
  INVX1 U17 ( .A(n5), .Y(n7) );
  INVX1 U18 ( .A(r_dac_en[1]), .Y(n8) );
  INVX1 U19 ( .A(n8), .Y(n9) );
  INVX1 U20 ( .A(n8), .Y(n10) );
  INVX1 U21 ( .A(r_dac_en[9]), .Y(n11) );
  INVX1 U22 ( .A(n11), .Y(n12) );
  INVX1 U23 ( .A(n11), .Y(n13) );
  INVX1 U24 ( .A(r_dac_en[10]), .Y(n14) );
  INVX1 U25 ( .A(n14), .Y(n15) );
  INVX1 U26 ( .A(n14), .Y(n16) );
  INVX1 U27 ( .A(r_dac_en[11]), .Y(n17) );
  INVX1 U28 ( .A(n17), .Y(n18) );
  INVX1 U29 ( .A(n17), .Y(n19) );
  INVX1 U30 ( .A(r_dac_en[12]), .Y(n20) );
  INVX1 U31 ( .A(n20), .Y(n21) );
  INVX1 U32 ( .A(n20), .Y(n22) );
  INVX1 U33 ( .A(r_dac_en[13]), .Y(n23) );
  INVX1 U34 ( .A(n23), .Y(n24) );
  INVX1 U35 ( .A(n23), .Y(n25) );
  INVX1 U36 ( .A(r_dac_en[15]), .Y(n26) );
  INVX1 U37 ( .A(n26), .Y(n27) );
  INVX1 U38 ( .A(n26), .Y(n28) );
  INVX1 U39 ( .A(r_dac_en[8]), .Y(n29) );
  INVX1 U40 ( .A(n29), .Y(n30) );
  INVX1 U41 ( .A(n29), .Y(n31) );
  INVX1 U42 ( .A(r_dac_en[14]), .Y(n32) );
  INVX1 U43 ( .A(n32), .Y(n33) );
  INVX1 U44 ( .A(n32), .Y(n34) );
  OR3XL U45 ( .A(wr_dacv[0]), .B(n78), .C(n7), .Y(n258) );
  AND2X1 U46 ( .A(pos_dacis[4]), .B(n66), .Y(n48) );
  INVXL U47 ( .A(sampl_done), .Y(n49) );
  AND3X1 U48 ( .A(n66), .B(pos_dacis[11]), .C(n118), .Y(N961) );
  AND3X1 U49 ( .A(n66), .B(pos_dacis[14]), .C(n118), .Y(N964) );
  AND3X1 U50 ( .A(n66), .B(pos_dacis[5]), .C(n118), .Y(N955) );
  AND3X1 U51 ( .A(n66), .B(pos_dacis[15]), .C(n118), .Y(N965) );
  AND3XL U52 ( .A(n117), .B(pos_dacis[0]), .C(n556), .Y(N950) );
  AND3XL U53 ( .A(n117), .B(pos_dacis[3]), .C(n556), .Y(N953) );
  AND3XL U54 ( .A(n117), .B(pos_dacis[1]), .C(n556), .Y(N951) );
  AND3XL U55 ( .A(n117), .B(pos_dacis[2]), .C(n556), .Y(N952) );
  AND3XL U56 ( .A(n117), .B(pos_dacis[6]), .C(n556), .Y(N956) );
  AND2X1 U57 ( .A(pos_dacis[13]), .B(n66), .Y(n57) );
  AND2X1 U58 ( .A(pos_dacis[12]), .B(n66), .Y(n58) );
  AND3XL U59 ( .A(n117), .B(pos_dacis[17]), .C(n556), .Y(N967) );
  AND3XL U60 ( .A(n117), .B(pos_dacis[8]), .C(n556), .Y(N958) );
  AND3XL U61 ( .A(n117), .B(pos_dacis[7]), .C(n556), .Y(N957) );
  AND3XL U62 ( .A(n117), .B(pos_dacis[10]), .C(n556), .Y(N960) );
  INVX1 U63 ( .A(r_dac_en[7]), .Y(n59) );
  INVX1 U64 ( .A(n152), .Y(n60) );
  BUFX6 U65 ( .A(sampl_done), .Y(n117) );
  BUFX6 U66 ( .A(sampl_done), .Y(n118) );
  INVX1 U67 ( .A(n64), .Y(n61) );
  INVX1 U68 ( .A(r_dac_en[4]), .Y(n62) );
  INVX1 U69 ( .A(r_dac_en[5]), .Y(n63) );
  BUFX3 U70 ( .A(n713), .Y(n64) );
  INVX1 U71 ( .A(r_dac_en[6]), .Y(n65) );
  INVX1 U72 ( .A(n579), .Y(n66) );
  BUFX3 U73 ( .A(r_dac_en[3]), .Y(n67) );
  NOR2X1 U74 ( .A(r_semi), .B(auto_start), .Y(n78) );
  INVX1 U75 ( .A(n678), .Y(n371) );
  INVX1 U76 ( .A(n378), .Y(n345) );
  GEN2XL U77 ( .D(n329), .E(N1178), .C(n348), .B(n351), .A(n328), .Y(n296) );
  INVX1 U78 ( .A(n177), .Y(n229) );
  OR2XL U79 ( .A(stop), .B(n137), .Y(n416) );
  INVXL U80 ( .A(ps_ptr[4]), .Y(n684) );
  AND2XL U81 ( .A(n685), .B(ps_ptr[2]), .Y(N997) );
  AND2XL U82 ( .A(n685), .B(ps_ptr[4]), .Y(N999) );
  AND2XL U83 ( .A(n685), .B(ps_ptr[0]), .Y(N995) );
  OAI21AXL U84 ( .B(stop), .C(srstz), .A(n685), .Y(N994) );
  OAI211XL U85 ( .C(n70), .D(n378), .A(n377), .B(n376), .Y(ps_ptr[3]) );
  AOI32XL U86 ( .A(n95), .B(n373), .C(n372), .D(n371), .E(n370), .Y(n377) );
  AND2XL U87 ( .A(n374), .B(n378), .Y(n263) );
  NAND21XL U88 ( .B(n128), .A(ps_ptr[3]), .Y(n660) );
  AND2XL U89 ( .A(n685), .B(ps_ptr[1]), .Y(N996) );
  AND4XL U90 ( .A(n287), .B(n286), .C(n190), .D(n8), .Y(n235) );
  AOI211XL U91 ( .C(n291), .D(n186), .A(n293), .B(n327), .Y(n187) );
  AND3XL U92 ( .A(n290), .B(n289), .C(n32), .Y(n185) );
  NAND2XL U93 ( .A(n178), .B(n78), .Y(n374) );
  NAND2XL U94 ( .A(n230), .B(n229), .Y(n375) );
  NOR32XL U95 ( .B(n244), .C(n121), .A(wr_dacv[17]), .Y(n246) );
  NAND43XL U96 ( .B(n297), .C(n326), .D(n296), .A(n113), .Y(n309) );
  INVXL U97 ( .A(n353), .Y(n329) );
  INVXL U98 ( .A(n295), .Y(n351) );
  INVXL U99 ( .A(n243), .Y(n253) );
  AOI211XL U100 ( .C(n329), .D(n133), .A(n348), .B(n328), .Y(n330) );
  INVXL U101 ( .A(n293), .Y(n251) );
  OAI211XL U102 ( .C(n129), .D(n353), .A(n352), .B(n351), .Y(n372) );
  INVXL U103 ( .A(n348), .Y(n352) );
  AO21XL U104 ( .B(ps_ptr[1]), .C(n123), .A(ps_ptr[0]), .Y(n668) );
  OA21XL U105 ( .B(ps_ptr[1]), .C(n663), .A(n662), .Y(n667) );
  AO21XL U106 ( .B(ps_ptr[2]), .C(n126), .A(n664), .Y(n665) );
  AOI21XL U107 ( .B(n680), .C(n679), .A(n678), .Y(n681) );
  NAND21XL U108 ( .B(n33), .A(n290), .Y(n249) );
  AND3XL U109 ( .A(n289), .B(n26), .C(n247), .Y(n250) );
  NOR2XL U110 ( .A(n31), .B(wr_dacv[8]), .Y(n112) );
  OR4XL U111 ( .A(n30), .B(n187), .C(wr_dacv[8]), .D(n292), .Y(n188) );
  OAI32XL U112 ( .A(n664), .B(ps_ptr[2]), .C(n126), .D(ps_ptr[3]), .E(n129), 
        .Y(n661) );
  INVX1 U113 ( .A(srstz), .Y(n137) );
  INVX1 U114 ( .A(n501), .Y(n768) );
  INVX1 U115 ( .A(n525), .Y(n746) );
  INVX1 U116 ( .A(n181), .Y(n280) );
  INVX1 U117 ( .A(n627), .Y(n802) );
  INVX1 U118 ( .A(wr_dacv[1]), .Y(n286) );
  INVX1 U119 ( .A(n416), .Y(n687) );
  NAND2X1 U120 ( .A(N1392), .B(n770), .Y(n501) );
  NOR2X1 U121 ( .A(n770), .B(N1392), .Y(n499) );
  INVX1 U122 ( .A(n502), .Y(n769) );
  NAND2X1 U123 ( .A(N1228), .B(n748), .Y(n525) );
  NOR2X1 U124 ( .A(n748), .B(N1228), .Y(n523) );
  INVX1 U125 ( .A(n526), .Y(n747) );
  INVX1 U126 ( .A(n477), .Y(n757) );
  INVX1 U127 ( .A(N1270), .Y(n751) );
  INVX1 U128 ( .A(N1599), .Y(n788) );
  NOR2X1 U129 ( .A(n804), .B(N1720), .Y(n625) );
  INVX1 U130 ( .A(n68), .Y(n771) );
  INVX1 U131 ( .A(n610), .Y(n793) );
  INVX1 U132 ( .A(n573), .Y(n785) );
  NAND21X1 U133 ( .B(n702), .A(n160), .Y(n181) );
  NAND2X1 U134 ( .A(N1720), .B(n804), .Y(n627) );
  INVX1 U135 ( .A(n628), .Y(n803) );
  INVX1 U136 ( .A(n549), .Y(n776) );
  INVX1 U137 ( .A(n654), .Y(n811) );
  INVX1 U138 ( .A(n653), .Y(n810) );
  INVX1 U139 ( .A(N1391), .Y(n770) );
  INVX1 U140 ( .A(N1148), .Y(n735) );
  INVX1 U141 ( .A(N1219), .Y(n702) );
  NAND2X1 U142 ( .A(N1392), .B(N1391), .Y(n502) );
  INVX1 U143 ( .A(n268), .Y(n710) );
  NOR2XL U144 ( .A(N1391), .B(N1392), .Y(n500) );
  NOR2X1 U145 ( .A(n759), .B(N1310), .Y(n475) );
  INVX1 U146 ( .A(N1227), .Y(n748) );
  INVX1 U147 ( .A(N1147), .Y(n736) );
  INVX1 U148 ( .A(N1393), .Y(n767) );
  INVX1 U149 ( .A(N1271), .Y(n750) );
  NAND2X1 U150 ( .A(N1228), .B(N1227), .Y(n526) );
  NAND2X1 U151 ( .A(N1310), .B(n759), .Y(n477) );
  NOR2XL U152 ( .A(N1227), .B(N1228), .Y(n524) );
  INVX1 U153 ( .A(n478), .Y(n758) );
  INVX1 U154 ( .A(n454), .Y(n738) );
  INVX1 U155 ( .A(n513), .Y(n752) );
  INVX1 U156 ( .A(n453), .Y(n737) );
  XOR3X1 U157 ( .A(n698), .B(n403), .C(n402), .Y(N1599) );
  INVX1 U158 ( .A(n694), .Y(n760) );
  INVX1 U159 ( .A(n194), .Y(n270) );
  INVX1 U160 ( .A(n199), .Y(n276) );
  INVX1 U161 ( .A(n490), .Y(n763) );
  INVX1 U162 ( .A(n489), .Y(n762) );
  NAND21X1 U163 ( .B(N1425), .A(n272), .Y(n389) );
  XNOR3X1 U164 ( .A(n149), .B(n390), .C(n389), .Y(n68) );
  XNOR2XL U165 ( .A(N1219), .B(sub_398_S2_I11_aco_carry[2]), .Y(n69) );
  INVX1 U166 ( .A(n205), .Y(n267) );
  INVX1 U167 ( .A(N1719), .Y(n804) );
  INVX1 U168 ( .A(n693), .Y(n796) );
  INVX1 U169 ( .A(n711), .Y(n775) );
  NAND2X1 U170 ( .A(N1638), .B(n795), .Y(n610) );
  NAND2X1 U171 ( .A(n69), .B(n787), .Y(n573) );
  NAND2X1 U172 ( .A(N1474), .B(n778), .Y(n549) );
  INVX1 U173 ( .A(n281), .Y(n160) );
  NOR2X1 U174 ( .A(n795), .B(N1638), .Y(n608) );
  NOR2X1 U175 ( .A(n787), .B(n69), .Y(n571) );
  NOR2X1 U176 ( .A(n778), .B(N1474), .Y(n547) );
  INVX1 U177 ( .A(n611), .Y(n794) );
  INVX1 U178 ( .A(n586), .Y(n790) );
  INVX1 U179 ( .A(n585), .Y(n789) );
  NAND21X1 U180 ( .B(n180), .A(n280), .Y(n179) );
  AO21X1 U181 ( .B(n281), .C(n702), .A(n280), .Y(N1720) );
  INVX1 U182 ( .A(n812), .Y(N1801) );
  NAND2X1 U183 ( .A(N1720), .B(N1719), .Y(n628) );
  INVX1 U184 ( .A(n359), .Y(n196) );
  INVX1 U185 ( .A(n784), .Y(n692) );
  NOR2X1 U186 ( .A(n812), .B(N1802), .Y(n651) );
  NOR2X1 U187 ( .A(N1719), .B(N1720), .Y(n626) );
  NOR2X1 U188 ( .A(N1801), .B(N1802), .Y(n652) );
  INVX1 U189 ( .A(n174), .Y(n284) );
  INVX1 U190 ( .A(n538), .Y(n773) );
  INVX1 U191 ( .A(n599), .Y(n799) );
  INVX1 U192 ( .A(n550), .Y(n777) );
  INVX1 U193 ( .A(n466), .Y(n742) );
  INVX1 U194 ( .A(n574), .Y(n786) );
  INVX1 U195 ( .A(n537), .Y(n772) );
  INVX1 U196 ( .A(n598), .Y(n798) );
  NAND2X1 U197 ( .A(N1802), .B(n812), .Y(n653) );
  NAND2X1 U198 ( .A(N1802), .B(N1801), .Y(n654) );
  AOI21AX1 U199 ( .B(n181), .C(n180), .A(n179), .Y(n70) );
  INVX1 U200 ( .A(n641), .Y(n806) );
  INVX1 U201 ( .A(N1638), .Y(n305) );
  NAND21X1 U202 ( .B(n406), .A(n404), .Y(sub_398_S2_I10_aco_carry_5_) );
  AND2X1 U203 ( .A(n685), .B(ps_ptr[3]), .Y(N998) );
  AND2X1 U204 ( .A(n432), .B(n531), .Y(N986) );
  AND2X1 U205 ( .A(n432), .B(n532), .Y(N985) );
  AND2X1 U206 ( .A(n432), .B(n555), .Y(N984) );
  AND2X1 U207 ( .A(n531), .B(n544), .Y(N974) );
  AND2X1 U208 ( .A(n532), .B(n544), .Y(N973) );
  INVX1 U209 ( .A(N1309), .Y(n759) );
  INVX1 U210 ( .A(N1145), .Y(n739) );
  NAND21X1 U211 ( .B(n412), .A(n154), .Y(N1219) );
  NAND21X1 U212 ( .B(n278), .A(n279), .Y(n268) );
  INVX1 U213 ( .A(N1262), .Y(n410) );
  NAND2X1 U214 ( .A(N1140), .B(n411), .Y(N1139) );
  INVX1 U215 ( .A(N1394), .Y(n766) );
  INVX1 U216 ( .A(n203), .Y(n425) );
  INVX1 U217 ( .A(N1466), .Y(n712) );
  NOR2X1 U218 ( .A(N1309), .B(N1310), .Y(n476) );
  NOR2X1 U219 ( .A(N1145), .B(N1146), .Y(n452) );
  INVX1 U220 ( .A(n154), .Y(n414) );
  NOR2X1 U221 ( .A(n754), .B(N1269), .Y(n511) );
  NOR2X1 U222 ( .A(n739), .B(N1146), .Y(n451) );
  INVX1 U223 ( .A(n393), .Y(n412) );
  INVX1 U224 ( .A(n162), .Y(n397) );
  INVX1 U225 ( .A(n396), .Y(n413) );
  INVX1 U226 ( .A(N1312), .Y(n755) );
  INVX1 U227 ( .A(N1230), .Y(n744) );
  NAND2XL U228 ( .A(N1310), .B(N1309), .Y(n478) );
  NAND2XL U229 ( .A(N1146), .B(N1145), .Y(n454) );
  NAND2X1 U230 ( .A(N1269), .B(n754), .Y(n513) );
  NAND2X1 U231 ( .A(N1146), .B(n739), .Y(n453) );
  INVX1 U232 ( .A(N1548), .Y(N1220) );
  INVX1 U233 ( .A(N1589), .Y(n697) );
  INVX1 U234 ( .A(N1630), .Y(n696) );
  INVX1 U235 ( .A(n407), .Y(n391) );
  INVX1 U236 ( .A(n514), .Y(n753) );
  XOR3X1 U237 ( .A(sub_398_S2_I6_aco_carry[4]), .B(n335), .C(n334), .Y(n694)
         );
  NAND21X1 U238 ( .B(N1589), .A(n270), .Y(n402) );
  NAND21X1 U239 ( .B(N1630), .A(n276), .Y(n399) );
  NAND21X1 U240 ( .B(n403), .A(n409), .Y(n194) );
  NAND21X1 U241 ( .B(n714), .A(n198), .Y(n199) );
  NAND21X1 U242 ( .B(n394), .A(n278), .Y(sub_398_S2_I6_aco_carry[3]) );
  INVX1 U243 ( .A(n415), .Y(n433) );
  INVX1 U244 ( .A(N1350), .Y(n764) );
  INVX1 U245 ( .A(n695), .Y(n792) );
  INVX1 U246 ( .A(n277), .Y(n198) );
  NAND2X1 U247 ( .A(N1351), .B(N1350), .Y(n490) );
  NAND2X1 U248 ( .A(N1351), .B(n764), .Y(n489) );
  INVX1 U249 ( .A(n146), .Y(n698) );
  NOR2X1 U250 ( .A(n764), .B(N1351), .Y(n487) );
  NOR2X1 U251 ( .A(N1350), .B(N1351), .Y(n488) );
  INVX1 U252 ( .A(N1344), .Y(n335) );
  INVX1 U253 ( .A(n363), .Y(n339) );
  INVX1 U254 ( .A(n269), .Y(n403) );
  INVX1 U255 ( .A(n334), .Y(n394) );
  XOR3X1 U256 ( .A(sub_398_S2_I14_aco_carry[4]), .B(n316), .C(n314), .Y(n693)
         );
  XNOR3X1 U257 ( .A(N1469), .B(N1467), .C(n380), .Y(n711) );
  AO21X1 U258 ( .B(n277), .C(n714), .A(n276), .Y(N1638) );
  NAND21X1 U259 ( .B(n204), .A(N1469), .Y(n205) );
  AO21X1 U260 ( .B(n161), .C(n64), .A(n160), .Y(N1719) );
  INVX1 U261 ( .A(n159), .Y(n161) );
  NAND21X1 U262 ( .B(n142), .A(n191), .Y(n266) );
  NAND21X1 U263 ( .B(n387), .A(n166), .Y(N1425) );
  XOR2X1 U264 ( .A(sub_398_S2_I6_aco_carry[3]), .B(N1671), .Y(N1352) );
  NAND21X1 U265 ( .B(N1466), .A(n267), .Y(n380) );
  OR2X1 U266 ( .A(n267), .B(n71), .Y(N1474) );
  AOI21X1 U267 ( .B(N1469), .C(n64), .A(n714), .Y(n71) );
  NAND21X1 U268 ( .B(n64), .A(n159), .Y(n281) );
  NAND21X1 U269 ( .B(n384), .A(n278), .Y(sub_398_S2_I14_aco_carry[3]) );
  INVX1 U270 ( .A(N1633), .Y(n400) );
  INVX1 U271 ( .A(n791), .Y(n701) );
  INVX1 U272 ( .A(N1637), .Y(n795) );
  INVX1 U273 ( .A(N1558), .Y(n783) );
  INVX1 U274 ( .A(N1555), .Y(n787) );
  INVX1 U275 ( .A(N1678), .Y(n800) );
  INVX1 U276 ( .A(N1473), .Y(n778) );
  NAND2X1 U277 ( .A(N1597), .B(n791), .Y(n585) );
  NAND2X1 U278 ( .A(N1638), .B(N1637), .Y(n611) );
  NAND2X1 U279 ( .A(n69), .B(N1555), .Y(n574) );
  NAND2X1 U280 ( .A(N1474), .B(N1473), .Y(n550) );
  NAND2X1 U281 ( .A(N1597), .B(n701), .Y(n586) );
  INVX1 U282 ( .A(N1384), .Y(n180) );
  INVX1 U283 ( .A(N1426), .Y(n149) );
  INVX1 U284 ( .A(n365), .Y(n675) );
  NOR2X1 U285 ( .A(n791), .B(N1597), .Y(n583) );
  NOR2X1 U286 ( .A(n774), .B(N1433), .Y(n535) );
  NOR2X1 U287 ( .A(n800), .B(N1679), .Y(n596) );
  NOR2X1 U288 ( .A(N1637), .B(N1638), .Y(n609) );
  NOR2X1 U289 ( .A(N1555), .B(n69), .Y(n572) );
  NOR2X1 U290 ( .A(N1473), .B(N1474), .Y(n548) );
  NOR2X1 U291 ( .A(N1678), .B(N1679), .Y(n597) );
  NOR2X1 U292 ( .A(n700), .B(N1433), .Y(n536) );
  NOR2X1 U293 ( .A(N1186), .B(N1187), .Y(n464) );
  NOR2X1 U294 ( .A(n701), .B(N1597), .Y(n584) );
  INVX1 U295 ( .A(n150), .Y(n272) );
  INVX1 U296 ( .A(n147), .Y(n387) );
  INVX1 U297 ( .A(n139), .Y(n142) );
  INVX1 U298 ( .A(n271), .Y(n390) );
  INVX1 U299 ( .A(n314), .Y(n384) );
  OR2X1 U300 ( .A(n284), .B(n72), .Y(N1802) );
  AOI21X1 U301 ( .B(n283), .C(n64), .A(n714), .Y(n72) );
  XOR2X1 U302 ( .A(n283), .B(n64), .Y(n812) );
  XOR2X1 U303 ( .A(sub_398_S2_I14_aco_carry[3]), .B(N1671), .Y(n797) );
  XOR2X1 U304 ( .A(N1548), .B(sub_398_S2_I11_aco_carry[3]), .Y(n784) );
  NAND21X1 U305 ( .B(n406), .A(n191), .Y(n273) );
  OAI21BBX1 U306 ( .A(N1589), .B(n194), .C(n402), .Y(n359) );
  NAND2X1 U307 ( .A(n283), .B(n173), .Y(n174) );
  INVX1 U308 ( .A(n774), .Y(n700) );
  INVX1 U309 ( .A(N1514), .Y(n782) );
  INVX1 U310 ( .A(n715), .Y(n779) );
  NAND2X1 U311 ( .A(N1433), .B(n774), .Y(n537) );
  NAND2X1 U312 ( .A(N1679), .B(N1678), .Y(n599) );
  NAND2X1 U313 ( .A(N1679), .B(n800), .Y(n598) );
  NAND2X1 U314 ( .A(N1187), .B(N1186), .Y(n466) );
  NAND2X1 U315 ( .A(N1433), .B(n700), .Y(n538) );
  INVX1 U316 ( .A(n153), .Y(n404) );
  NAND21X1 U317 ( .B(n433), .A(n203), .Y(n153) );
  AOI21AX1 U318 ( .B(N1630), .C(n199), .A(n399), .Y(n73) );
  AOI21AX1 U319 ( .B(n150), .C(N1425), .A(n389), .Y(n74) );
  INVX1 U320 ( .A(n204), .Y(n173) );
  INVX1 U321 ( .A(n275), .Y(n406) );
  OAI21BBX1 U322 ( .A(n205), .B(N1466), .C(n380), .Y(n358) );
  INVX1 U323 ( .A(n562), .Y(n781) );
  INVX1 U324 ( .A(n561), .Y(n780) );
  INVX1 U325 ( .A(n465), .Y(n741) );
  NOR2X1 U326 ( .A(n808), .B(N1761), .Y(n639) );
  OA22X1 U327 ( .A(N1466), .B(n284), .C(n712), .D(n174), .Y(n75) );
  NAND2X1 U328 ( .A(N1761), .B(n808), .Y(n641) );
  INVX1 U329 ( .A(n801), .Y(n344) );
  INVX1 U330 ( .A(n642), .Y(n807) );
  INVX1 U331 ( .A(N1679), .Y(n304) );
  INVX1 U332 ( .A(N1433), .Y(n303) );
  XOR2X1 U333 ( .A(N1263), .B(sub_398_S2_I4_aco_carry[5]), .Y(n76) );
  AO21X1 U334 ( .B(sub_398_S2_I6_aco_carry[4]), .C(N1344), .A(n395), .Y(
        sub_398_S2_I6_aco_carry[5]) );
  OA21X1 U335 ( .B(sub_398_S2_I6_aco_carry[4]), .C(N1344), .A(n394), .Y(n395)
         );
  XOR2X1 U336 ( .A(N1427), .B(n77), .Y(N1436) );
  OAI21X1 U337 ( .B(N1426), .C(n390), .A(n389), .Y(n77) );
  OA21X1 U338 ( .B(N1467), .C(n381), .A(n380), .Y(sub_398_S2_I9_aco_carry_5_)
         );
  INVX1 U339 ( .A(N1469), .Y(n381) );
  INVX1 U340 ( .A(n436), .Y(n555) );
  OAI221X1 U341 ( .A(n805), .B(n375), .C(n809), .D(n374), .E(n347), .Y(
        ps_ptr[4]) );
  AOI211X1 U342 ( .C(n345), .D(n344), .A(n343), .B(n342), .Y(n347) );
  OA21X1 U343 ( .B(n341), .C(n340), .A(n371), .Y(n342) );
  AND4X1 U344 ( .A(n95), .B(n332), .C(n331), .D(n330), .Y(n343) );
  OAI221X1 U345 ( .A(n313), .B(n375), .C(n312), .D(n374), .E(n311), .Y(
        ps_ptr[2]) );
  INVX1 U346 ( .A(N1761), .Y(n313) );
  INVX1 U347 ( .A(N1802), .Y(n312) );
  AOI222XL U348 ( .A(n310), .B(n309), .C(n371), .D(n308), .E(n345), .F(N1720), 
        .Y(n311) );
  INVX1 U349 ( .A(n324), .Y(n310) );
  OA22X1 U350 ( .A(n2), .B(n375), .C(n75), .D(n374), .Y(n376) );
  NAND21X1 U351 ( .B(n368), .A(n367), .Y(n370) );
  NAND21X1 U352 ( .B(n265), .A(n264), .Y(ps_ptr[0]) );
  MUX2X1 U353 ( .D0(n263), .D1(n375), .S(cs_ptr[0]), .Y(n264) );
  GEN2XL U354 ( .D(n361), .E(n262), .C(n261), .B(n371), .A(n260), .Y(n265) );
  INVX1 U355 ( .A(n660), .Y(n664) );
  INVX1 U356 ( .A(n237), .Y(n685) );
  OAI31XL U357 ( .A(semi_start), .B(mxcyc_done), .C(auto_start), .D(n687), .Y(
        n237) );
  AND2X1 U358 ( .A(n432), .B(n460), .Y(N987) );
  AND2X1 U359 ( .A(n460), .B(n544), .Y(N975) );
  INVX1 U360 ( .A(n459), .Y(n544) );
  INVX1 U361 ( .A(n427), .Y(n432) );
  NAND21X1 U362 ( .B(n426), .A(n433), .Y(n427) );
  INVX1 U363 ( .A(n434), .Y(n443) );
  NAND21X1 U364 ( .B(n128), .A(cs_ptr[4]), .Y(n203) );
  NAND21X1 U365 ( .B(n663), .A(cs_ptr[2]), .Y(n154) );
  XOR2X1 U366 ( .A(n162), .B(n128), .Y(N1466) );
  XOR2X1 U367 ( .A(n407), .B(cs_ptr[4]), .Y(N1262) );
  XOR2X1 U368 ( .A(n154), .B(n128), .Y(N1384) );
  AO21X1 U369 ( .B(n397), .C(N1179), .A(n131), .Y(N1140) );
  NAND21X1 U370 ( .B(n274), .A(N1185), .Y(n162) );
  NAND21X1 U371 ( .B(N1178), .A(n662), .Y(n396) );
  NAND21X1 U372 ( .B(cs_ptr[2]), .A(n663), .Y(n393) );
  NAND21X1 U373 ( .B(n1), .A(cs_ptr[1]), .Y(sub_398_S2_I4_aco_carry[2]) );
  NAND21X1 U374 ( .B(cs_ptr[3]), .A(n191), .Y(n407) );
  INVX1 U375 ( .A(N1136), .Y(n713) );
  AO21X1 U376 ( .B(n414), .C(n131), .A(n690), .Y(N1386) );
  AND2X1 U377 ( .A(n717), .B(n716), .Y(n79) );
  AND2X1 U378 ( .A(n725), .B(n724), .Y(n80) );
  AND2X1 U379 ( .A(n722), .B(n721), .Y(n81) );
  NAND21X1 U380 ( .B(n307), .A(n306), .Y(n308) );
  OA2222XL U381 ( .A(n305), .B(n365), .C(n304), .D(n364), .E(n303), .F(n363), 
        .G(n302), .H(n362), .Y(n306) );
  AO2222XL U382 ( .A(n69), .B(n672), .C(n361), .D(n301), .E(n674), .F(N1597), 
        .G(n102), .H(N1474), .Y(n307) );
  INVX1 U383 ( .A(N1515), .Y(n302) );
  INVX1 U384 ( .A(n350), .Y(n749) );
  INVX1 U385 ( .A(n144), .Y(n191) );
  INVX1 U386 ( .A(n138), .Y(n278) );
  NAND21X1 U387 ( .B(N1177), .A(cs_ptr[2]), .Y(n138) );
  AND3X1 U388 ( .A(n425), .B(n532), .C(n426), .Y(N989) );
  AND3X1 U389 ( .A(n425), .B(n555), .C(n426), .Y(N988) );
  INVX1 U390 ( .A(n689), .Y(n325) );
  AND2X1 U391 ( .A(n443), .B(n460), .Y(N983) );
  AND2X1 U392 ( .A(n446), .B(n460), .Y(N979) );
  AND2X1 U393 ( .A(n446), .B(n531), .Y(N978) );
  NOR2X1 U394 ( .A(N1268), .B(N1269), .Y(n512) );
  INVX1 U395 ( .A(n424), .Y(n663) );
  OAI22X1 U396 ( .A(n765), .B(n770), .C(n754), .D(n350), .Y(n408) );
  AOI22XL U397 ( .A(n325), .B(N1227), .C(n98), .D(N1145), .Y(n405) );
  INVX1 U398 ( .A(n145), .Y(n409) );
  NAND21X1 U399 ( .B(n710), .A(cs_ptr[1]), .Y(n145) );
  AOI22X1 U400 ( .A(n325), .B(N1228), .C(n98), .D(N1146), .Y(n383) );
  INVX1 U401 ( .A(n143), .Y(n417) );
  NAND21X1 U402 ( .B(cs_ptr[1]), .A(N1185), .Y(n143) );
  AOI22X1 U403 ( .A(n325), .B(N1230), .C(n98), .D(N1148), .Y(n346) );
  NAND21X1 U404 ( .B(n131), .A(cs_ptr[3]), .Y(n415) );
  NAND21X1 U405 ( .B(n162), .A(n690), .Y(n411) );
  XOR2X1 U406 ( .A(n393), .B(n128), .Y(N1548) );
  XOR2X1 U407 ( .A(n144), .B(n128), .Y(N1589) );
  XOR2X1 U408 ( .A(n396), .B(n128), .Y(N1630) );
  NAND21X1 U409 ( .B(N1178), .A(cs_ptr[1]), .Y(n279) );
  AO21X1 U410 ( .B(n131), .C(n393), .A(n690), .Y(N1222) );
  AO21X1 U411 ( .B(n131), .C(n396), .A(n690), .Y(N1304) );
  AND2X1 U412 ( .A(n719), .B(n718), .Y(n82) );
  INVX1 U413 ( .A(N1268), .Y(n754) );
  NAND2X1 U414 ( .A(N1269), .B(N1268), .Y(n514) );
  INVX1 U415 ( .A(N1137), .Y(n714) );
  OAI22X1 U416 ( .A(n765), .B(n766), .C(n750), .D(n350), .Y(n349) );
  INVX1 U417 ( .A(n354), .Y(n706) );
  AOI22X1 U418 ( .A(n325), .B(N1229), .C(n98), .D(N1147), .Y(n366) );
  INVX1 U419 ( .A(n392), .Y(N1263) );
  NAND21X1 U420 ( .B(n391), .A(cs_ptr[4]), .Y(n392) );
  XNOR3X1 U421 ( .A(N1633), .B(N1631), .C(n399), .Y(n695) );
  NAND21X1 U422 ( .B(N1136), .A(N1633), .Y(n277) );
  OAI211X1 U423 ( .C(N1178), .D(n334), .A(sub_398_S2_I6_aco_carry[3]), .B(n279), .Y(N1351) );
  XOR2X1 U424 ( .A(n334), .B(N1177), .Y(N1350) );
  NAND21X1 U425 ( .B(n709), .A(n670), .Y(n363) );
  OR2X1 U426 ( .A(n433), .B(n83), .Y(N1344) );
  MUX2IX1 U427 ( .D0(n203), .D1(N1181), .S(cs_ptr[2]), .Y(n83) );
  NAND21X1 U428 ( .B(n191), .A(cs_ptr[3]), .Y(n401) );
  XOR2X1 U429 ( .A(n401), .B(cs_ptr[4]), .Y(n146) );
  OAI21X1 U430 ( .B(n278), .C(n335), .A(n723), .Y(n334) );
  OAI21X1 U431 ( .B(n409), .C(n146), .A(n731), .Y(n269) );
  AO2222XL U432 ( .A(n102), .B(n711), .C(n672), .D(N1558), .E(n339), .F(n68), 
        .G(n674), .H(N1599), .Y(n340) );
  AO21X1 U433 ( .B(N1178), .C(n131), .A(n690), .Y(N1345) );
  INVX1 U434 ( .A(n333), .Y(n704) );
  OAI22X1 U435 ( .A(n765), .B(n767), .C(n751), .D(n350), .Y(n369) );
  XOR3X1 U436 ( .A(sub_398_S2_I11_aco_carry[4]), .B(n87), .C(N1549), .Y(N1558)
         );
  OAI21X1 U437 ( .B(n149), .C(n167), .A(n726), .Y(n271) );
  OR2X1 U438 ( .A(n272), .B(n84), .Y(N1433) );
  AOI21X1 U439 ( .B(N1177), .C(n271), .A(n710), .Y(n84) );
  XOR2X1 U440 ( .A(n61), .B(N1469), .Y(N1473) );
  XOR2X1 U441 ( .A(n61), .B(n87), .Y(N1555) );
  XOR2X1 U442 ( .A(n314), .B(cs_ptr[1]), .Y(N1678) );
  AO21X1 U443 ( .B(n61), .C(n400), .A(n198), .Y(N1637) );
  NAND21X1 U444 ( .B(n212), .A(n364), .Y(n365) );
  AO21X1 U445 ( .B(n155), .C(n156), .A(n60), .Y(n159) );
  NAND32X1 U446 ( .B(n64), .C(n180), .A(N1219), .Y(n155) );
  OAI211X1 U447 ( .C(N1178), .D(n314), .A(sub_398_S2_I14_aco_carry[3]), .B(
        n279), .Y(N1679) );
  XOR2X1 U448 ( .A(n269), .B(N1177), .Y(n791) );
  NAND21X1 U449 ( .B(n274), .A(n128), .Y(n166) );
  OR2X1 U450 ( .A(n433), .B(n85), .Y(N1467) );
  MUX2IX1 U451 ( .D0(n203), .D1(N1181), .S(n397), .Y(n85) );
  XOR2X1 U452 ( .A(n147), .B(cs_ptr[4]), .Y(N1426) );
  OR2X1 U453 ( .A(n270), .B(n86), .Y(N1597) );
  AOI21X1 U454 ( .B(N1177), .C(n269), .A(n268), .Y(n86) );
  NAND2X1 U455 ( .A(n274), .B(n266), .Y(N1187) );
  NAND21X1 U456 ( .B(n128), .A(n274), .Y(n147) );
  NAND21X1 U457 ( .B(N1137), .A(n713), .Y(n204) );
  OAI21X1 U458 ( .B(n278), .C(n316), .A(n734), .Y(n314) );
  NAND21X1 U459 ( .B(n390), .A(n167), .Y(n150) );
  NAND21X1 U460 ( .B(cs_ptr[4]), .A(n391), .Y(n139) );
  AO21X1 U461 ( .B(n397), .C(n131), .A(n690), .Y(N1468) );
  AND2X1 U462 ( .A(n730), .B(n729), .Y(n87) );
  INVX1 U463 ( .A(n240), .Y(n674) );
  NOR2X1 U464 ( .A(n743), .B(N1187), .Y(n463) );
  INVX1 U465 ( .A(n362), .Y(n676) );
  INVX1 U466 ( .A(N1672), .Y(n316) );
  INVX1 U467 ( .A(n398), .Y(N1632) );
  NAND21X1 U468 ( .B(n413), .A(n690), .Y(n398) );
  INVX1 U469 ( .A(n388), .Y(N1427) );
  NAND21X1 U470 ( .B(n387), .A(cs_ptr[4]), .Y(n388) );
  INVX1 U471 ( .A(n379), .Y(N1550) );
  NAND21X1 U472 ( .B(n412), .A(n690), .Y(n379) );
  NOR2X1 U473 ( .A(n128), .B(n266), .Y(n88) );
  AND2X1 U474 ( .A(n192), .B(n89), .Y(n715) );
  XNOR2XL U475 ( .A(n275), .B(n404), .Y(n89) );
  XOR2X1 U476 ( .A(n275), .B(cs_ptr[1]), .Y(N1514) );
  OA2222XL U477 ( .A(n73), .B(n365), .C(n364), .D(n797), .E(n74), .F(n363), 
        .G(n109), .H(n362), .Y(n367) );
  XOR2X1 U478 ( .A(n271), .B(cs_ptr[1]), .Y(n774) );
  OR2X1 U479 ( .A(n690), .B(n90), .Y(n275) );
  AOI21X1 U480 ( .B(n191), .C(N1179), .A(n404), .Y(n90) );
  NAND21X1 U481 ( .B(n165), .A(n164), .Y(n283) );
  INVX1 U482 ( .A(n411), .Y(n165) );
  AO21X1 U483 ( .B(n173), .C(N1466), .A(n163), .Y(n164) );
  INVX1 U484 ( .A(n172), .Y(n163) );
  NAND21X1 U485 ( .B(n158), .A(n179), .Y(n801) );
  XOR2X1 U486 ( .A(n159), .B(n157), .Y(n158) );
  INVX1 U487 ( .A(n156), .Y(n157) );
  NAND2X1 U488 ( .A(N1187), .B(n743), .Y(n465) );
  NAND2X1 U489 ( .A(N1515), .B(N1514), .Y(n562) );
  NAND2X1 U490 ( .A(N1515), .B(n782), .Y(n561) );
  INVX1 U491 ( .A(N1343), .Y(N1671) );
  INVX1 U492 ( .A(n743), .Y(N1186) );
  AOI21X1 U493 ( .B(N1179), .C(n266), .A(n88), .Y(n91) );
  NOR2X1 U494 ( .A(n782), .B(N1515), .Y(n559) );
  NOR2X1 U495 ( .A(N1514), .B(N1515), .Y(n560) );
  OR2X1 U496 ( .A(n282), .B(n92), .Y(N1761) );
  AOI21X1 U497 ( .B(N1177), .C(N1181), .A(n710), .Y(n92) );
  NAND21X1 U498 ( .B(n283), .A(n172), .Y(n809) );
  MUX2BXL U499 ( .D0(n242), .D1(n241), .S(n120), .Y(n261) );
  NAND32X1 U500 ( .B(n672), .C(n102), .A(n365), .Y(n242) );
  AND4X1 U501 ( .A(n240), .B(n364), .C(n362), .D(n363), .Y(n241) );
  INVX1 U502 ( .A(n168), .Y(n282) );
  NAND2X1 U503 ( .A(N1761), .B(n699), .Y(n642) );
  NOR2X1 U504 ( .A(n699), .B(N1761), .Y(n640) );
  OR2X1 U505 ( .A(n131), .B(n166), .Y(n805) );
  INVX1 U506 ( .A(n699), .Y(n808) );
  INVX1 U507 ( .A(N1425), .Y(n169) );
  NAND3X1 U508 ( .A(n319), .B(n320), .C(n321), .Y(n317) );
  AOI21BBXL U509 ( .B(n76), .C(n350), .A(n116), .Y(n321) );
  AOI22X1 U510 ( .A(N1354), .B(n704), .C(N1231), .D(n325), .Y(n320) );
  AOI22X1 U511 ( .A(N1149), .B(n98), .C(N1313), .D(n707), .Y(n319) );
  XOR2X1 U512 ( .A(N1632), .B(n93), .Y(N1641) );
  OAI21X1 U513 ( .B(N1631), .C(n400), .A(n399), .Y(n93) );
  XOR2X1 U514 ( .A(n106), .B(n94), .Y(N1600) );
  OAI21X1 U515 ( .B(n698), .C(n403), .A(n402), .Y(n94) );
  AO21X1 U516 ( .B(sub_398_S2_I14_aco_carry[4]), .C(N1672), .A(n385), .Y(
        sub_398_S2_I14_aco_carry[5]) );
  OA21X1 U517 ( .B(sub_398_S2_I14_aco_carry[4]), .C(N1672), .A(n384), .Y(n385)
         );
  NAND21X1 U518 ( .B(n424), .A(n428), .Y(n436) );
  INVX1 U519 ( .A(n419), .Y(n532) );
  NAND21X1 U520 ( .B(n418), .A(n417), .Y(n419) );
  INVX1 U521 ( .A(n418), .Y(n428) );
  INVX1 U522 ( .A(n435), .Y(n531) );
  NAND21X1 U523 ( .B(n579), .A(n49), .Y(N949) );
  OAI221X1 U524 ( .A(n808), .B(n375), .C(n812), .D(n374), .E(n236), .Y(
        ps_ptr[1]) );
  AOI211X1 U525 ( .C(n345), .D(N1719), .A(n235), .B(n234), .Y(n236) );
  OA21X1 U526 ( .B(n233), .C(n232), .A(n371), .Y(n234) );
  NAND32X1 U527 ( .B(n231), .C(n230), .A(n229), .Y(n678) );
  INVX1 U528 ( .A(wr_dacv[2]), .Y(n285) );
  NAND21X1 U529 ( .B(n178), .A(n78), .Y(n177) );
  OAI211X1 U530 ( .C(n123), .D(n353), .A(n26), .B(n185), .Y(n186) );
  INVX1 U531 ( .A(n258), .Y(n287) );
  NOR3XL U532 ( .A(n326), .B(n324), .C(n323), .Y(n95) );
  NAND32X1 U533 ( .B(n183), .C(n230), .A(n229), .Y(n378) );
  INVX1 U534 ( .A(n231), .Y(n183) );
  NAND5XL U535 ( .A(n291), .B(n290), .C(n289), .D(n32), .E(n26), .Y(n348) );
  INVX1 U536 ( .A(n294), .Y(n332) );
  NAND32X1 U537 ( .B(n293), .C(n292), .A(n112), .Y(n294) );
  INVX1 U538 ( .A(n184), .Y(n291) );
  NAND32XL U539 ( .B(wr_dacv[13]), .C(n243), .A(n23), .Y(n184) );
  NAND21X1 U540 ( .B(n327), .A(n332), .Y(n295) );
  NAND32XL U541 ( .B(wr_dacv[16]), .C(n246), .A(n245), .Y(n247) );
  AOI31X1 U542 ( .A(n286), .B(n8), .C(n259), .D(n258), .Y(n260) );
  NAND32X1 U543 ( .B(n135), .C(wr_dacv[2]), .A(n257), .Y(n259) );
  GEN3XL U544 ( .F(n112), .G(n256), .E(n328), .D(n255), .C(n297), .B(n113), 
        .A(n254), .Y(n257) );
  GEN2XL U545 ( .D(n253), .E(n252), .C(n327), .B(n251), .A(n292), .Y(n256) );
  INVX1 U546 ( .A(n327), .Y(n331) );
  NAND21X1 U547 ( .B(n297), .A(n113), .Y(n323) );
  INVX1 U548 ( .A(n254), .Y(n288) );
  INVX1 U549 ( .A(n328), .Y(n373) );
  INVX1 U550 ( .A(n326), .Y(n255) );
  AOI31X1 U551 ( .A(n669), .B(n668), .C(n667), .D(n666), .Y(n683) );
  AO22XL U552 ( .A(ps_ptr[4]), .B(n133), .C(n669), .D(n665), .Y(n666) );
  AOI222XL U553 ( .A(N1682), .B(n677), .C(N1518), .D(n676), .E(N1641), .F(n675), .Y(n679) );
  AOI221XL U554 ( .A(N1477), .B(n102), .C(N1600), .D(n674), .E(n673), .Y(n680)
         );
  NAND21X1 U555 ( .B(n437), .A(n433), .Y(n434) );
  NAND32X1 U556 ( .B(n131), .C(n437), .A(n129), .Y(n459) );
  INVX1 U557 ( .A(n579), .Y(n556) );
  INVX1 U558 ( .A(n126), .Y(cs_ptr[2]) );
  INVX1 U559 ( .A(n124), .Y(cs_ptr[1]) );
  AND3X1 U560 ( .A(n555), .B(n544), .C(n543), .Y(N972) );
  INVX1 U561 ( .A(n121), .Y(cs_ptr[0]) );
  AND2X1 U562 ( .A(n532), .B(n444), .Y(N981) );
  AND2X1 U563 ( .A(n555), .B(n444), .Y(N980) );
  INVX1 U564 ( .A(n439), .Y(n446) );
  NAND32X1 U565 ( .B(n131), .C(N1179), .A(n437), .Y(n439) );
  OAI32X1 U566 ( .A(n459), .B(n436), .C(n543), .D(n435), .E(n434), .Y(N982) );
  INVX1 U567 ( .A(n437), .Y(n426) );
  NAND31X1 U568 ( .C(n703), .A(n440), .B(n438), .Y(n442) );
  AO21X1 U569 ( .B(N1177), .C(n121), .A(n417), .Y(N1136) );
  NAND21X1 U570 ( .B(n124), .A(cs_ptr[2]), .Y(n274) );
  NAND21X1 U571 ( .B(n442), .A(n708), .Y(n689) );
  NAND3X1 U572 ( .A(n438), .B(n440), .C(n703), .Y(n350) );
  NAND21X1 U573 ( .B(cs_ptr[2]), .A(n123), .Y(n144) );
  NAND21X1 U574 ( .B(N1177), .A(n121), .Y(n424) );
  INVX1 U575 ( .A(n221), .Y(n707) );
  NAND21X1 U576 ( .B(n438), .A(n440), .Y(n221) );
  AO22X1 U577 ( .A(n322), .B(N1392), .C(N1269), .D(n749), .Y(n386) );
  NAND2X1 U578 ( .A(n96), .B(n415), .Y(N1385) );
  MUX2IX1 U579 ( .D0(n425), .D1(n132), .S(n414), .Y(n96) );
  MUX2IX1 U580 ( .D0(n447), .D1(n448), .S(cs_ptr[0]), .Y(n218) );
  NAND21X1 U581 ( .B(n123), .A(N1185), .Y(n662) );
  NAND2X1 U582 ( .A(n97), .B(n415), .Y(N1303) );
  MUX2IX1 U583 ( .D0(n132), .D1(n425), .S(n413), .Y(n97) );
  NOR2X1 U584 ( .A(n322), .B(n705), .Y(n440) );
  INVX1 U585 ( .A(n322), .Y(n765) );
  AO2222XL U586 ( .A(n676), .B(n715), .C(n361), .D(n338), .E(n693), .F(n677), 
        .G(n675), .H(n695), .Y(n341) );
  OAI211X1 U587 ( .C(n133), .D(n357), .A(n337), .B(n336), .Y(n338) );
  AOI221XL U588 ( .A(n704), .B(n694), .C(N1312), .D(n707), .E(n349), .Y(n336)
         );
  OA21X1 U589 ( .B(n740), .C(n354), .A(n346), .Y(n337) );
  OAI211X1 U590 ( .C(n300), .D(n333), .A(n299), .B(n298), .Y(n301) );
  INVX1 U591 ( .A(N1351), .Y(n300) );
  AOI221XL U592 ( .A(n706), .B(N1187), .C(N1310), .D(n707), .E(n386), .Y(n298)
         );
  OA21X1 U593 ( .B(n126), .C(n357), .A(n383), .Y(n299) );
  NOR3XL U594 ( .A(n442), .B(n708), .C(n441), .Y(n445) );
  INVX1 U595 ( .A(n133), .Y(cs_ptr[4]) );
  AND3X1 U596 ( .A(n446), .B(n532), .C(n543), .Y(N977) );
  AND3X1 U597 ( .A(n446), .B(n555), .C(n543), .Y(N976) );
  INVX1 U598 ( .A(n129), .Y(n128) );
  AND2X1 U599 ( .A(n99), .B(n445), .Y(n98) );
  MUX2IX1 U600 ( .D0(n447), .D1(n448), .S(cs_ptr[0]), .Y(n99) );
  AO2222XL U601 ( .A(n672), .B(N1555), .C(n361), .D(n228), .E(n674), .F(n701), 
        .G(n102), .H(N1473), .Y(n232) );
  OAI211X1 U602 ( .C(n764), .D(n333), .A(n223), .B(n222), .Y(n228) );
  AOI221XL U603 ( .A(n706), .B(N1186), .C(N1309), .D(n707), .E(n408), .Y(n222)
         );
  OA21X1 U604 ( .B(n123), .C(n357), .A(n405), .Y(n223) );
  OAI21BBX1 U605 ( .A(n1), .B(n123), .C(sub_398_S2_I4_aco_carry[2]), .Y(N1268)
         );
  NAND32X1 U606 ( .B(n220), .C(n708), .A(n219), .Y(n354) );
  INVX1 U607 ( .A(n441), .Y(n220) );
  INVX1 U608 ( .A(n442), .Y(n219) );
  OR2X1 U609 ( .A(n278), .B(n100), .Y(N1137) );
  MUX2IX1 U610 ( .D0(n126), .D1(n279), .S(cs_ptr[0]), .Y(n100) );
  INVX1 U611 ( .A(n152), .Y(n690) );
  NAND21X1 U612 ( .B(n133), .A(cs_ptr[3]), .Y(n152) );
  NAND2X1 U613 ( .A(n101), .B(n415), .Y(N1221) );
  MUX2IX1 U614 ( .D0(n132), .D1(n425), .S(n412), .Y(n101) );
  AO2222XL U615 ( .A(n672), .B(n692), .C(n361), .D(n360), .E(n674), .F(n359), 
        .G(n102), .H(n358), .Y(n368) );
  OAI211X1 U616 ( .C(n129), .D(n357), .A(n356), .B(n355), .Y(n360) );
  AOI221XL U617 ( .A(n704), .B(N1352), .C(n707), .D(N1311), .E(n369), .Y(n355)
         );
  OA21X1 U618 ( .B(n91), .C(n354), .A(n366), .Y(n356) );
  INVX1 U619 ( .A(n129), .Y(cs_ptr[3]) );
  INVX1 U620 ( .A(n133), .Y(n131) );
  NAND21X1 U621 ( .B(n322), .A(n705), .Y(n333) );
  XOR2X1 U622 ( .A(n129), .B(cs_ptr[2]), .Y(N1343) );
  INVX1 U623 ( .A(n202), .Y(n208) );
  NAND32X1 U624 ( .B(n213), .C(n677), .A(n214), .Y(n202) );
  INVX1 U625 ( .A(n210), .Y(n227) );
  NAND21X1 U626 ( .B(n209), .A(n208), .Y(n210) );
  AND2X1 U627 ( .A(n226), .B(n227), .Y(n102) );
  OR2X1 U628 ( .A(n425), .B(n103), .Y(N1631) );
  MUX2IX1 U629 ( .D0(n415), .D1(n132), .S(n413), .Y(n103) );
  AO2222XL U630 ( .A(n676), .B(N1514), .C(n339), .D(n700), .E(n677), .F(N1678), 
        .G(n675), .H(N1637), .Y(n233) );
  INVX1 U631 ( .A(n225), .Y(n212) );
  INVX1 U632 ( .A(n211), .Y(n670) );
  NAND21X1 U633 ( .B(n226), .A(n227), .Y(n211) );
  INVX1 U634 ( .A(n201), .Y(n214) );
  NAND21X1 U635 ( .B(n224), .A(n212), .Y(n201) );
  INVX1 U636 ( .A(n217), .Y(n361) );
  NAND21X1 U637 ( .B(n318), .A(n670), .Y(n217) );
  AO21X1 U638 ( .B(n132), .C(n139), .A(n88), .Y(n740) );
  NAND2X1 U639 ( .A(n209), .B(n208), .Y(n362) );
  OR2X1 U640 ( .A(n425), .B(n104), .Y(N1672) );
  MUX2IX1 U641 ( .D0(n132), .D1(n415), .S(cs_ptr[2]), .Y(n104) );
  NAND32X1 U642 ( .B(n677), .C(n225), .A(n224), .Y(n240) );
  INVX1 U643 ( .A(n148), .Y(n167) );
  NAND21X1 U644 ( .B(n124), .A(n710), .Y(n148) );
  OR2X1 U645 ( .A(n425), .B(n105), .Y(N1549) );
  MUX2IX1 U646 ( .D0(n415), .D1(n132), .S(n412), .Y(n105) );
  MUX2BXL U647 ( .D0(n239), .D1(n238), .S(n120), .Y(n262) );
  NAND43X1 U648 ( .B(n707), .C(n98), .D(n322), .A(n689), .Y(n239) );
  AND4X1 U649 ( .A(n333), .B(n354), .C(n350), .D(n357), .Y(n238) );
  INVX1 U650 ( .A(n216), .Y(n672) );
  NAND32X1 U651 ( .B(n215), .C(n677), .A(n214), .Y(n216) );
  INVX1 U652 ( .A(n213), .Y(n215) );
  INVX1 U653 ( .A(n318), .Y(n709) );
  NOR2X1 U654 ( .A(n133), .B(n401), .Y(n106) );
  OAI211X1 U655 ( .C(n126), .D(n275), .A(n274), .B(n273), .Y(N1515) );
  NAND21X1 U656 ( .B(n142), .A(n123), .Y(n743) );
  OR2X1 U657 ( .A(n425), .B(n107), .Y(n172) );
  MUX2IX1 U658 ( .D0(n133), .D1(n415), .S(n397), .Y(n107) );
  OR2X1 U659 ( .A(n129), .B(n273), .Y(n192) );
  OR2X1 U660 ( .A(n425), .B(n108), .Y(n156) );
  MUX2IX1 U661 ( .D0(n132), .D1(n415), .S(n414), .Y(n108) );
  INVX1 U662 ( .A(n677), .Y(n364) );
  INVX1 U663 ( .A(n382), .Y(N1673) );
  NAND21X1 U664 ( .B(n126), .A(n690), .Y(n382) );
  NAND21X1 U665 ( .B(n133), .A(n167), .Y(n168) );
  AOI21AX1 U666 ( .B(n273), .C(n129), .A(n192), .Y(n109) );
  INVX1 U667 ( .A(n136), .Y(n134) );
  INVX1 U668 ( .A(n136), .Y(n135) );
  XOR2X1 U669 ( .A(n132), .B(cs_ptr[1]), .Y(n699) );
  INVX1 U670 ( .A(n121), .Y(n120) );
  MUX2IX1 U671 ( .D0(n245), .D1(n244), .S(cs_ptr[0]), .Y(n110) );
  MUX2IX1 U672 ( .D0(n244), .D1(n245), .S(cs_ptr[0]), .Y(n111) );
  AO22AXL U673 ( .A(N1559), .B(n672), .C(n670), .D(n315), .Y(n673) );
  AOI22X1 U674 ( .A(n709), .B(n317), .C(N1436), .D(n318), .Y(n315) );
  AND2X1 U675 ( .A(N1395), .B(n322), .Y(n116) );
  NAND21X1 U676 ( .B(n137), .A(sampl_begn), .Y(n418) );
  NAND2X1 U677 ( .A(n121), .B(n431), .Y(n435) );
  INVX1 U678 ( .A(n430), .Y(n460) );
  NAND21X1 U679 ( .B(n121), .A(n431), .Y(n430) );
  INVX1 U680 ( .A(n429), .Y(n431) );
  NAND21X1 U681 ( .B(n123), .A(n428), .Y(n429) );
  NAND43X1 U682 ( .B(wr_dacv[16]), .C(wr_dacv[17]), .D(n4), .A(n244), .Y(n353)
         );
  NAND43X1 U683 ( .B(n135), .C(n189), .D(wr_dacv[2]), .A(n288), .Y(n190) );
  AOI31X1 U684 ( .A(n373), .B(n255), .C(n188), .D(n323), .Y(n189) );
  OR2XL U685 ( .A(wr_dacv[10]), .B(n16), .Y(n293) );
  OR2XL U686 ( .A(wr_dacv[11]), .B(n19), .Y(n327) );
  OR2XL U687 ( .A(wr_dacv[12]), .B(n21), .Y(n243) );
  OR2XL U688 ( .A(wr_dacv[9]), .B(n13), .Y(n292) );
  OAI211X1 U689 ( .C(n250), .D(n249), .A(n248), .B(n23), .Y(n252) );
  INVXL U690 ( .A(wr_dacv[13]), .Y(n248) );
  INVX1 U691 ( .A(cs_mux_5_), .Y(busy) );
  OR2X1 U692 ( .A(wr_dacv[7]), .B(r_dac_en[7]), .Y(n328) );
  OR2X1 U693 ( .A(wr_dacv[6]), .B(r_dac_en[6]), .Y(n326) );
  OR2X1 U694 ( .A(wr_dacv[3]), .B(n67), .Y(n254) );
  OR2X1 U695 ( .A(wr_dacv[5]), .B(r_dac_en[5]), .Y(n297) );
  NOR2X1 U696 ( .A(wr_dacv[4]), .B(r_dac_en[4]), .Y(n113) );
  NAND21X1 U697 ( .B(pos_dacis[11]), .A(n52), .Y(app_dacis[11]) );
  NAND21XL U698 ( .B(pos_dacis[5]), .A(n54), .Y(app_dacis[5]) );
  NAND21XL U699 ( .B(pos_dacis[2]), .A(n44), .Y(app_dacis[2]) );
  NAND21X1 U700 ( .B(pos_dacis[12]), .A(n604), .Y(app_dacis[12]) );
  NAND21X1 U701 ( .B(pos_dacis[14]), .A(n51), .Y(app_dacis[14]) );
  NAND21XL U702 ( .B(pos_dacis[4]), .A(n580), .Y(app_dacis[4]) );
  INVX1 U703 ( .A(neg_dacis[4]), .Y(n580) );
  NAND21X1 U704 ( .B(pos_dacis[6]), .A(n43), .Y(app_dacis[6]) );
  NAND21X1 U705 ( .B(pos_dacis[7]), .A(n39), .Y(app_dacis[7]) );
  NAND21X1 U706 ( .B(pos_dacis[16]), .A(n616), .Y(app_dacis[16]) );
  INVX1 U707 ( .A(neg_dacis[16]), .Y(n616) );
  NAND21XL U708 ( .B(pos_dacis[1]), .A(n40), .Y(app_dacis[1]) );
  NAND21XL U709 ( .B(pos_dacis[3]), .A(n41), .Y(app_dacis[3]) );
  NAND21X1 U710 ( .B(pos_dacis[13]), .A(n605), .Y(app_dacis[13]) );
  NAND21X1 U711 ( .B(pos_dacis[15]), .A(n56), .Y(app_dacis[15]) );
  NAND21X1 U712 ( .B(pos_dacis[9]), .A(n591), .Y(app_dacis[9]) );
  NAND21X1 U713 ( .B(pos_dacis[8]), .A(n47), .Y(app_dacis[8]) );
  NAND21XL U714 ( .B(pos_dacis[0]), .A(n45), .Y(app_dacis[0]) );
  NAND21X1 U715 ( .B(pos_dacis[17]), .A(n37), .Y(app_dacis[17]) );
  NAND21X1 U716 ( .B(n688), .A(n687), .Y(n671) );
  MUX2X1 U717 ( .D0(cs_mux_5_), .D1(n686), .S(n685), .Y(n688) );
  GEN3XL U718 ( .F(N1181), .G(n684), .E(n683), .D(n682), .C(r_semi), .B(busy), 
        .A(n681), .Y(n686) );
  INVX1 U719 ( .A(r_loop), .Y(n682) );
  NAND21X1 U720 ( .B(pos_dacis[10]), .A(n35), .Y(app_dacis[10]) );
  INVX1 U721 ( .A(neg_dacis[13]), .Y(n605) );
  INVX1 U722 ( .A(neg_dacis[9]), .Y(n591) );
  INVX1 U723 ( .A(neg_dacis[12]), .Y(n604) );
  INVX1 U724 ( .A(n661), .Y(n669) );
  NAND21X1 U725 ( .B(n420), .A(n126), .Y(n437) );
  AND3X1 U726 ( .A(ps_md4ch), .B(n132), .C(n129), .Y(n420) );
  NAND6XL U727 ( .A(n41), .B(n44), .C(n40), .D(n45), .E(n423), .F(n422), .Y(
        n579) );
  NOR5X1 U728 ( .A(neg_dacis[4]), .B(n53), .C(n42), .D(n38), .E(n46), .Y(n423)
         );
  NOR6XL U729 ( .A(n421), .B(n50), .C(n55), .D(neg_dacis[16]), .E(n36), .F(
        n137), .Y(n422) );
  NAND5XL U730 ( .A(n605), .B(n604), .C(n52), .D(n35), .E(n591), .Y(n421) );
  AO21X1 U731 ( .B(r_comp_swtch), .C(n446), .A(n443), .Y(n444) );
  INVX1 U732 ( .A(N1177), .Y(n124) );
  INVX1 U733 ( .A(N1178), .Y(n126) );
  INVX1 U734 ( .A(N1185), .Y(n121) );
  MUX2IX1 U735 ( .D0(n495), .D1(n496), .S(N1185), .Y(n322) );
  AOI222XL U736 ( .A(N1394), .B(r_dac_en[16]), .C(n497), .D(n767), .E(N1393), 
        .F(n498), .Y(n496) );
  AOI222XL U737 ( .A(N1394), .B(r_dac_en[17]), .C(n504), .D(n767), .E(N1393), 
        .F(n505), .Y(n495) );
  AO2222XL U738 ( .A(n769), .B(n33), .C(n768), .D(n21), .E(n499), .F(n15), .G(
        n500), .H(n30), .Y(n498) );
  MUX2IX1 U739 ( .D0(n508), .D1(n507), .S(N1185), .Y(n703) );
  AOI222XL U740 ( .A(N1271), .B(r_dac_en[17]), .C(n516), .D(n751), .E(N1270), 
        .F(n517), .Y(n507) );
  AOI222XL U741 ( .A(N1271), .B(r_dac_en[16]), .C(n509), .D(n751), .E(N1270), 
        .F(n510), .Y(n508) );
  AO2222XL U742 ( .A(n753), .B(n27), .C(n752), .D(n25), .E(n511), .F(n19), .G(
        n512), .H(n13), .Y(n517) );
  MUX2AXL U743 ( .D0(n471), .D1(n472), .S(cs_ptr[0]), .Y(n438) );
  AOI222XL U744 ( .A(N1312), .B(r_dac_en[16]), .C(n473), .D(n756), .E(N1311), 
        .F(n474), .Y(n472) );
  AO222X1 U745 ( .A(N1312), .B(r_dac_en[17]), .C(n480), .D(n756), .E(N1311), 
        .F(n481), .Y(n471) );
  INVX1 U746 ( .A(N1311), .Y(n756) );
  AO2222XL U747 ( .A(n769), .B(n28), .C(n768), .D(n24), .E(n499), .F(n18), .G(
        n500), .H(n12), .Y(n505) );
  OAI221X1 U748 ( .A(n816), .B(n513), .C(n814), .D(n514), .E(n515), .Y(n509)
         );
  AOI32X1 U749 ( .A(n6), .B(n750), .C(n512), .D(n511), .E(n134), .Y(n515) );
  AOI222XL U750 ( .A(N1148), .B(n4), .C(n449), .D(n736), .E(N1147), .F(n450), 
        .Y(n448) );
  AO2222XL U751 ( .A(n738), .B(n33), .C(n737), .D(n21), .E(n451), .F(n15), .G(
        n452), .H(n30), .Y(n450) );
  OAI221X1 U752 ( .A(n816), .B(n453), .C(n814), .D(n454), .E(n455), .Y(n449)
         );
  AOI32X1 U753 ( .A(n7), .B(n735), .C(n452), .D(n451), .E(n134), .Y(n455) );
  OAI221X1 U754 ( .A(n816), .B(n501), .C(n814), .D(n502), .E(n503), .Y(n497)
         );
  AOI32X1 U755 ( .A(n7), .B(n766), .C(n500), .D(n499), .E(n134), .Y(n503) );
  OAI221X1 U756 ( .A(n815), .B(n477), .C(n813), .D(n478), .E(n482), .Y(n480)
         );
  AOI32X1 U757 ( .A(n9), .B(n755), .C(n476), .D(n475), .E(r_dac_en[3]), .Y(
        n482) );
  OAI221X1 U758 ( .A(n815), .B(n513), .C(n813), .D(n514), .E(n518), .Y(n516)
         );
  AOI32X1 U759 ( .A(n9), .B(n750), .C(n512), .D(n511), .E(r_dac_en[3]), .Y(
        n518) );
  AOI222XL U760 ( .A(N1148), .B(n3), .C(n456), .D(n736), .E(N1147), .F(n457), 
        .Y(n447) );
  AO2222XL U761 ( .A(n738), .B(n27), .C(n737), .D(n24), .E(n451), .F(n18), .G(
        n452), .H(n12), .Y(n457) );
  OAI221X1 U762 ( .A(n815), .B(n453), .C(n813), .D(n454), .E(n458), .Y(n456)
         );
  AOI32X1 U763 ( .A(n9), .B(n735), .C(n452), .D(n451), .E(r_dac_en[3]), .Y(
        n458) );
  OAI221X1 U764 ( .A(n815), .B(n501), .C(n813), .D(n502), .E(n506), .Y(n504)
         );
  AOI32X1 U765 ( .A(n10), .B(n766), .C(n500), .D(n499), .E(r_dac_en[3]), .Y(
        n506) );
  INVX1 U766 ( .A(N1181), .Y(n133) );
  AO2222XL U767 ( .A(n753), .B(n34), .C(n752), .D(n22), .E(n511), .F(n16), .G(
        n512), .H(n31), .Y(n510) );
  AO2222XL U768 ( .A(n758), .B(n33), .C(n757), .D(n21), .E(n475), .F(n15), .G(
        n476), .H(n30), .Y(n474) );
  AO2222XL U769 ( .A(n747), .B(n34), .C(n746), .D(n22), .E(n523), .F(n16), .G(
        n524), .H(n31), .Y(n522) );
  AO2222XL U770 ( .A(n747), .B(n28), .C(n746), .D(n25), .E(n523), .F(n19), .G(
        n524), .H(n13), .Y(n529) );
  AO2222XL U771 ( .A(n758), .B(n27), .C(n757), .D(n24), .E(n475), .F(n18), .G(
        n476), .H(n12), .Y(n481) );
  MUX2IX1 U772 ( .D0(n519), .D1(n520), .S(N1185), .Y(n708) );
  AOI222XL U773 ( .A(N1230), .B(r_dac_en[16]), .C(n521), .D(n745), .E(N1229), 
        .F(n522), .Y(n520) );
  AOI222XL U774 ( .A(N1230), .B(r_dac_en[17]), .C(n528), .D(n745), .E(N1229), 
        .F(n529), .Y(n519) );
  INVX1 U775 ( .A(N1229), .Y(n745) );
  OAI221X1 U776 ( .A(n816), .B(n477), .C(n814), .D(n478), .E(n479), .Y(n473)
         );
  AOI32X1 U777 ( .A(n7), .B(n755), .C(n476), .D(n475), .E(n134), .Y(n479) );
  OAI221X1 U778 ( .A(n816), .B(n525), .C(n814), .D(n526), .E(n527), .Y(n521)
         );
  AOI32X1 U779 ( .A(n6), .B(n744), .C(n524), .D(n523), .E(n134), .Y(n527) );
  OAI221X1 U780 ( .A(n815), .B(n525), .C(n813), .D(n526), .E(n530), .Y(n528)
         );
  AOI32X1 U781 ( .A(n9), .B(n744), .C(n524), .D(n523), .E(r_dac_en[3]), .Y(
        n530) );
  INVX1 U782 ( .A(N1177), .Y(n123) );
  INVX1 U783 ( .A(N1179), .Y(n129) );
  MUX2IX1 U784 ( .D0(n484), .D1(n483), .S(N1185), .Y(n705) );
  AOI222XL U785 ( .A(n694), .B(r_dac_en[16]), .C(n485), .D(n761), .E(N1352), 
        .F(n486), .Y(n484) );
  AOI222XL U786 ( .A(n694), .B(r_dac_en[17]), .C(n492), .D(n761), .E(N1352), 
        .F(n493), .Y(n483) );
  INVX1 U787 ( .A(N1352), .Y(n761) );
  AO21X1 U788 ( .B(n695), .C(n111), .A(n200), .Y(n225) );
  MUX4X1 U789 ( .D0(n614), .D1(n613), .D2(n607), .D3(n606), .S0(n73), .S1(n120), .Y(n200) );
  AO2222XL U790 ( .A(n794), .B(n34), .C(n793), .D(n22), .E(n608), .F(n16), .G(
        n609), .H(n31), .Y(n607) );
  AO2222XL U791 ( .A(n794), .B(n28), .C(n793), .D(n25), .E(n608), .F(n19), .G(
        n609), .H(n13), .Y(n614) );
  AO2222XL U792 ( .A(n763), .B(n34), .C(n762), .D(n22), .E(n487), .F(n16), .G(
        n488), .H(n31), .Y(n486) );
  AO2222XL U793 ( .A(n763), .B(n28), .C(n762), .D(n25), .E(n487), .F(n19), .G(
        n488), .H(n13), .Y(n493) );
  MUX2IX1 U794 ( .D0(n114), .D1(n115), .S(cs_ptr[0]), .Y(n224) );
  AOI21X1 U795 ( .B(n4), .C(N1599), .A(n195), .Y(n114) );
  AOI21X1 U796 ( .B(n3), .C(N1599), .A(n197), .Y(n115) );
  OAI221X1 U797 ( .A(n815), .B(n489), .C(n813), .D(n490), .E(n494), .Y(n492)
         );
  AOI32X1 U798 ( .A(n10), .B(n760), .C(n488), .D(n487), .E(r_dac_en[3]), .Y(
        n494) );
  OAI221X1 U799 ( .A(n816), .B(n489), .C(n814), .D(n490), .E(n491), .Y(n485)
         );
  AOI32X1 U800 ( .A(n6), .B(n760), .C(n488), .D(n487), .E(n134), .Y(n491) );
  OAI221X1 U801 ( .A(n815), .B(n610), .C(n813), .D(n611), .E(n615), .Y(n613)
         );
  AOI32X1 U802 ( .A(n9), .B(n792), .C(n609), .D(n608), .E(r_dac_en[3]), .Y(
        n615) );
  OAI221X1 U803 ( .A(n816), .B(n585), .C(n814), .D(n586), .E(n587), .Y(n581)
         );
  AOI32X1 U804 ( .A(n7), .B(n788), .C(n584), .D(n583), .E(n135), .Y(n587) );
  OAI221X1 U805 ( .A(n816), .B(n610), .C(n814), .D(n611), .E(n612), .Y(n606)
         );
  AOI32X1 U806 ( .A(n6), .B(n792), .C(n609), .D(n608), .E(n135), .Y(n612) );
  MUX2X1 U807 ( .D0(n589), .D1(n588), .S(n196), .Y(n197) );
  AO2222XL U808 ( .A(n790), .B(n28), .C(n789), .D(n25), .E(n583), .F(n19), .G(
        n584), .H(n13), .Y(n589) );
  OAI221X1 U809 ( .A(n815), .B(n585), .C(n813), .D(n586), .E(n590), .Y(n588)
         );
  AOI32X1 U810 ( .A(n10), .B(n788), .C(n584), .D(n583), .E(r_dac_en[3]), .Y(
        n590) );
  INVX1 U811 ( .A(N1181), .Y(n132) );
  MUX2IX1 U812 ( .D0(n593), .D1(n592), .S(N1185), .Y(n677) );
  AOI222XL U813 ( .A(n693), .B(n3), .C(n601), .D(n797), .E(n691), .F(n602), 
        .Y(n592) );
  AOI222XL U814 ( .A(n693), .B(n4), .C(n594), .D(n797), .E(n691), .F(n595), 
        .Y(n593) );
  INVX1 U815 ( .A(n797), .Y(n691) );
  AO21X1 U816 ( .B(n68), .C(n110), .A(n151), .Y(n318) );
  MUX4X1 U817 ( .D0(n534), .D1(n533), .D2(n541), .D3(n540), .S0(n74), .S1(n120), .Y(n151) );
  AO2222XL U818 ( .A(n773), .B(n28), .C(n772), .D(n25), .E(n535), .F(n19), .G(
        n536), .H(n13), .Y(n541) );
  AO2222XL U819 ( .A(n773), .B(n34), .C(n772), .D(n22), .E(n535), .F(n16), .G(
        n536), .H(n31), .Y(n534) );
  AO21X1 U820 ( .B(n711), .C(n111), .A(n207), .Y(n226) );
  MUX4X1 U821 ( .D0(n553), .D1(n552), .D2(n546), .D3(n545), .S0(n206), .S1(
        n120), .Y(n207) );
  INVX1 U822 ( .A(n358), .Y(n206) );
  AO2222XL U823 ( .A(n777), .B(n34), .C(n776), .D(n22), .E(n547), .F(n16), .G(
        n548), .H(n31), .Y(n546) );
  AO21X1 U824 ( .B(n141), .C(n110), .A(n140), .Y(n441) );
  INVX1 U825 ( .A(n740), .Y(n141) );
  MUX4X1 U826 ( .D0(n462), .D1(n461), .D2(n469), .D3(n468), .S0(n91), .S1(n120), .Y(n140) );
  AO2222XL U827 ( .A(n742), .B(n27), .C(n741), .D(n24), .E(n463), .F(n18), .G(
        n464), .H(n12), .Y(n469) );
  AO21X1 U828 ( .B(n111), .C(n344), .A(n182), .Y(n231) );
  MUX4X1 U829 ( .D0(n631), .D1(n630), .D2(n624), .D3(n623), .S0(n70), .S1(n120), .Y(n182) );
  AO2222XL U830 ( .A(n803), .B(n34), .C(n802), .D(n22), .E(n625), .F(n15), .G(
        n626), .H(n30), .Y(n624) );
  AO2222XL U831 ( .A(n803), .B(n27), .C(n802), .D(n24), .E(n625), .F(n18), .G(
        n626), .H(n12), .Y(n631) );
  AO2222XL U832 ( .A(n799), .B(n33), .C(n798), .D(n21), .E(n596), .F(n15), .G(
        n597), .H(n30), .Y(n595) );
  AO2222XL U833 ( .A(n790), .B(n34), .C(n789), .D(n22), .E(n583), .F(n16), .G(
        n584), .H(n31), .Y(n582) );
  AO2222XL U834 ( .A(n786), .B(n27), .C(n785), .D(n24), .E(n571), .F(n18), .G(
        n572), .H(n12), .Y(n577) );
  AO2222XL U835 ( .A(n799), .B(n27), .C(n798), .D(n24), .E(n596), .F(n18), .G(
        n597), .H(n12), .Y(n602) );
  MUX2IX1 U836 ( .D0(n567), .D1(n568), .S(N1185), .Y(n213) );
  AOI222XL U837 ( .A(N1558), .B(n4), .C(n569), .D(n784), .E(n692), .F(n570), 
        .Y(n568) );
  AOI222XL U838 ( .A(N1558), .B(n3), .C(n576), .D(n784), .E(n692), .F(n577), 
        .Y(n567) );
  AO2222XL U839 ( .A(n786), .B(n33), .C(n785), .D(n21), .E(n571), .F(n15), .G(
        n572), .H(n30), .Y(n570) );
  OAI221X1 U840 ( .A(n63), .B(n573), .C(n59), .D(n574), .E(n578), .Y(n576) );
  AOI32X1 U841 ( .A(n10), .B(n783), .C(n572), .D(n571), .E(n67), .Y(n578) );
  OAI221X1 U842 ( .A(n62), .B(n573), .C(n65), .D(n574), .E(n575), .Y(n569) );
  AOI32X1 U843 ( .A(n7), .B(n783), .C(n572), .D(n571), .E(n135), .Y(n575) );
  OAI221X1 U844 ( .A(n816), .B(n598), .C(n814), .D(n599), .E(n600), .Y(n594)
         );
  AOI32X1 U845 ( .A(n7), .B(n796), .C(n597), .D(n596), .E(n135), .Y(n600) );
  OAI221X1 U846 ( .A(n815), .B(n598), .C(n813), .D(n599), .E(n603), .Y(n601)
         );
  AOI32X1 U847 ( .A(n10), .B(n796), .C(n597), .D(n596), .E(n67), .Y(n603) );
  OAI221X1 U848 ( .A(n63), .B(n549), .C(n59), .D(n550), .E(n554), .Y(n552) );
  AOI32X1 U849 ( .A(n9), .B(n775), .C(n548), .D(n547), .E(n67), .Y(n554) );
  OAI221X1 U850 ( .A(n816), .B(n465), .C(n814), .D(n466), .E(n467), .Y(n461)
         );
  AOI32X1 U851 ( .A(n6), .B(n740), .C(n464), .D(n463), .E(n134), .Y(n467) );
  OAI221X1 U852 ( .A(n63), .B(n627), .C(n59), .D(n628), .E(n632), .Y(n630) );
  AOI32X1 U853 ( .A(n9), .B(n801), .C(n626), .D(n625), .E(n67), .Y(n632) );
  OAI221X1 U854 ( .A(n62), .B(n537), .C(n65), .D(n538), .E(n539), .Y(n533) );
  AOI32X1 U855 ( .A(n6), .B(n771), .C(n536), .D(n535), .E(n134), .Y(n539) );
  OAI221X1 U856 ( .A(n62), .B(n549), .C(n65), .D(n550), .E(n551), .Y(n545) );
  AOI32X1 U857 ( .A(n6), .B(n775), .C(n548), .D(n547), .E(n134), .Y(n551) );
  OAI221X1 U858 ( .A(n815), .B(n465), .C(n813), .D(n466), .E(n470), .Y(n468)
         );
  AOI32X1 U859 ( .A(n10), .B(n740), .C(n464), .D(n463), .E(r_dac_en[3]), .Y(
        n470) );
  OAI221X1 U860 ( .A(n63), .B(n537), .C(n59), .D(n538), .E(n542), .Y(n540) );
  AOI32X1 U861 ( .A(n9), .B(n771), .C(n536), .D(n535), .E(n67), .Y(n542) );
  OAI221X1 U862 ( .A(n62), .B(n627), .C(n65), .D(n628), .E(n629), .Y(n623) );
  AOI32X1 U863 ( .A(n6), .B(n801), .C(n626), .D(n625), .E(n135), .Y(n629) );
  AO21X1 U864 ( .B(n715), .C(n110), .A(n193), .Y(n209) );
  MUX4X1 U865 ( .D0(n558), .D1(n557), .D2(n565), .D3(n564), .S0(n109), .S1(
        n120), .Y(n193) );
  AO2222XL U866 ( .A(n781), .B(n28), .C(n780), .D(n25), .E(n559), .F(n18), .G(
        n560), .H(n13), .Y(n565) );
  AO2222XL U867 ( .A(n781), .B(n33), .C(n780), .D(n21), .E(n559), .F(n15), .G(
        n560), .H(n30), .Y(n558) );
  AO21X1 U868 ( .B(n111), .C(n176), .A(n175), .Y(n178) );
  INVX1 U869 ( .A(n809), .Y(n176) );
  MUX4X1 U870 ( .D0(n657), .D1(n656), .D2(n650), .D3(n649), .S0(n75), .S1(n120), .Y(n175) );
  AO2222XL U871 ( .A(n811), .B(n33), .C(n810), .D(n21), .E(n651), .F(n15), .G(
        n652), .H(n31), .Y(n650) );
  AO2222XL U872 ( .A(n742), .B(n33), .C(n741), .D(n21), .E(n463), .F(n15), .G(
        n464), .H(n30), .Y(n462) );
  AO2222XL U873 ( .A(n777), .B(n27), .C(n776), .D(n24), .E(n547), .F(n19), .G(
        n548), .H(n12), .Y(n553) );
  OAI221X1 U874 ( .A(n63), .B(n653), .C(n59), .D(n654), .E(n658), .Y(n656) );
  AOI32X1 U875 ( .A(n10), .B(n809), .C(n652), .D(n651), .E(n67), .Y(n658) );
  OAI221X1 U876 ( .A(n63), .B(n561), .C(n59), .D(n562), .E(n566), .Y(n564) );
  AOI32X1 U877 ( .A(n10), .B(n779), .C(n560), .D(n559), .E(n67), .Y(n566) );
  OAI221X1 U878 ( .A(n62), .B(n561), .C(n65), .D(n562), .E(n563), .Y(n557) );
  AOI32X1 U879 ( .A(n7), .B(n779), .C(n560), .D(n559), .E(n135), .Y(n563) );
  OAI221X1 U880 ( .A(n62), .B(n653), .C(n65), .D(n654), .E(n655), .Y(n649) );
  AOI32X1 U881 ( .A(n6), .B(n809), .C(n652), .D(n651), .E(n135), .Y(n655) );
  AO21X1 U882 ( .B(n110), .C(n171), .A(n170), .Y(n230) );
  INVX1 U883 ( .A(n805), .Y(n171) );
  MUX4X1 U884 ( .D0(n638), .D1(n637), .D2(n645), .D3(n644), .S0(n2), .S1(n120), 
        .Y(n170) );
  AO2222XL U885 ( .A(n28), .B(n807), .C(n25), .D(n806), .E(n19), .F(n639), .G(
        n12), .H(n640), .Y(n645) );
  AO2222XL U886 ( .A(n811), .B(n27), .C(n810), .D(n24), .E(n651), .F(n18), .G(
        n652), .H(n13), .Y(n657) );
  OAI221X1 U887 ( .A(n641), .B(n62), .C(n642), .D(n65), .E(n643), .Y(n637) );
  AOI32X1 U888 ( .A(n640), .B(n805), .C(n7), .D(n134), .E(n639), .Y(n643) );
  OAI221X1 U889 ( .A(n641), .B(n63), .C(n642), .D(n59), .E(n646), .Y(n644) );
  AOI32X1 U890 ( .A(n640), .B(n805), .C(n9), .D(n67), .E(n639), .Y(n646) );
  INVX1 U891 ( .A(r_dac_en[2]), .Y(n136) );
  AO2222XL U892 ( .A(n34), .B(n807), .C(n22), .D(n806), .E(n16), .F(n639), .G(
        n30), .H(n640), .Y(n638) );
  INVX1 U893 ( .A(r_dac_en[5]), .Y(n815) );
  INVX1 U894 ( .A(r_dac_en[7]), .Y(n813) );
  INVX1 U895 ( .A(r_dac_en[4]), .Y(n816) );
  INVX1 U896 ( .A(r_dac_en[6]), .Y(n814) );
  INVX1 U897 ( .A(r_dac_en[17]), .Y(n244) );
  INVX1 U898 ( .A(r_dac_en[16]), .Y(n245) );
  NOR32XL U899 ( .B(n633), .C(n622), .A(n621), .Y(n634) );
  NAND31X1 U900 ( .C(pos_dacis[14]), .A(n620), .B(n619), .Y(n621) );
  INVX1 U901 ( .A(pos_dacis[16]), .Y(n633) );
  INVX1 U902 ( .A(pos_dacis[17]), .Y(n622) );
  NOR32XL U903 ( .B(n659), .C(n648), .A(n647), .Y(sh_hold) );
  INVX1 U904 ( .A(pos_dacis[9]), .Y(n659) );
  NOR21XL U905 ( .B(n618), .A(n617), .Y(n648) );
  NAND31X1 U906 ( .C(n636), .A(n635), .B(n634), .Y(n647) );
  OR3XL U907 ( .A(pos_dacis[7]), .B(pos_dacis[6]), .C(pos_dacis[8]), .Y(n636)
         );
  OR2X1 U908 ( .A(pos_dacis[10]), .B(pos_dacis[11]), .Y(n617) );
  NOR6XL U909 ( .A(pos_dacis[5]), .B(pos_dacis[4]), .C(pos_dacis[3]), .D(
        pos_dacis[2]), .E(pos_dacis[1]), .F(pos_dacis[0]), .Y(n635) );
  INVX1 U910 ( .A(pos_dacis[15]), .Y(n619) );
  INVX1 U911 ( .A(pos_dacis[13]), .Y(n620) );
  INVX1 U912 ( .A(pos_dacis[12]), .Y(n618) );
  INVX1 U913 ( .A(r_comp_swtch), .Y(n543) );
  INVXL U914 ( .A(wr_dacv[14]), .Y(n290) );
  INVXL U915 ( .A(wr_dacv[15]), .Y(n289) );
  NAND32XL U916 ( .B(n428), .C(n416), .A(n49), .Y(N971) );
  MAJ3X1 U917 ( .A(sub_398_S2_I11_aco_carry[4]), .B(n87), .C(N1549), .Y(
        sub_398_S2_I11_aco_carry[5]) );
  XNOR2XL U918 ( .A(N1550), .B(sub_398_S2_I11_aco_carry[5]), .Y(N1559) );
  XNOR2XL U919 ( .A(N1468), .B(sub_398_S2_I9_aco_carry_5_), .Y(N1477) );
  XNOR2XL U920 ( .A(N1673), .B(sub_398_S2_I14_aco_carry[5]), .Y(N1682) );
  XNOR2XL U921 ( .A(N1386), .B(sub_398_S2_I7_aco_carry[5]), .Y(N1395) );
  XNOR2XL U922 ( .A(N1222), .B(sub_398_S2_I3_aco_carry[5]), .Y(N1231) );
  XNOR2XL U923 ( .A(N1345), .B(sub_398_S2_I6_aco_carry[5]), .Y(N1354) );
  XNOR2XL U924 ( .A(N1304), .B(sub_398_S2_I5_aco_carry[5]), .Y(N1313) );
  XNOR2XL U925 ( .A(N1140), .B(sub_398_S2_aco_carry[5]), .Y(N1149) );
  XNOR2XL U926 ( .A(n60), .B(sub_398_S2_I10_aco_carry_5_), .Y(N1518) );
  OR2X1 U927 ( .A(sub_398_S2_aco_carry[3]), .B(n712), .Y(
        sub_398_S2_aco_carry[4]) );
  XNOR2XL U928 ( .A(sub_398_S2_aco_carry[3]), .B(n712), .Y(N1147) );
  OR2X1 U929 ( .A(sub_398_S2_aco_carry[2]), .B(N1137), .Y(
        sub_398_S2_aco_carry[3]) );
  XNOR2XL U930 ( .A(sub_398_S2_aco_carry[2]), .B(N1137), .Y(N1146) );
  OR2X1 U931 ( .A(N1136), .B(n79), .Y(sub_398_S2_aco_carry[2]) );
  XNOR2XL U932 ( .A(N1136), .B(n79), .Y(N1145) );
  OR2X1 U933 ( .A(sub_398_S2_I5_aco_carry[3]), .B(n696), .Y(
        sub_398_S2_I5_aco_carry[4]) );
  XNOR2XL U934 ( .A(sub_398_S2_I5_aco_carry[3]), .B(n696), .Y(N1311) );
  OR2X1 U935 ( .A(sub_398_S2_I5_aco_carry[2]), .B(n714), .Y(
        sub_398_S2_I5_aco_carry[3]) );
  XNOR2XL U936 ( .A(sub_398_S2_I5_aco_carry[2]), .B(n714), .Y(N1310) );
  OR2X1 U937 ( .A(N1136), .B(n81), .Y(sub_398_S2_I5_aco_carry[2]) );
  XNOR2XL U938 ( .A(N1136), .B(n81), .Y(N1309) );
  OR2X1 U939 ( .A(sub_398_S2_I6_aco_carry[3]), .B(N1343), .Y(
        sub_398_S2_I6_aco_carry[4]) );
  OR2X1 U940 ( .A(sub_398_S2_I7_aco_carry[3]), .B(N1384), .Y(
        sub_398_S2_I7_aco_carry[4]) );
  XNOR2XL U941 ( .A(sub_398_S2_I7_aco_carry[3]), .B(N1384), .Y(N1393) );
  OR2X1 U942 ( .A(sub_398_S2_I7_aco_carry[2]), .B(n702), .Y(
        sub_398_S2_I7_aco_carry[3]) );
  XNOR2XL U943 ( .A(sub_398_S2_I7_aco_carry[2]), .B(n702), .Y(N1392) );
  OR2X1 U944 ( .A(n713), .B(n80), .Y(sub_398_S2_I7_aco_carry[2]) );
  XNOR2XL U945 ( .A(n713), .B(n80), .Y(N1391) );
  OR2X1 U946 ( .A(sub_398_S2_I4_aco_carry[3]), .B(n697), .Y(
        sub_398_S2_I4_aco_carry[4]) );
  XNOR2XL U947 ( .A(sub_398_S2_I4_aco_carry[3]), .B(n697), .Y(N1270) );
  OR2X1 U948 ( .A(sub_398_S2_I4_aco_carry[2]), .B(n710), .Y(
        sub_398_S2_I4_aco_carry[3]) );
  XNOR2XL U949 ( .A(sub_398_S2_I4_aco_carry[2]), .B(n710), .Y(N1269) );
  OR2X1 U950 ( .A(sub_398_S2_I3_aco_carry[3]), .B(N1220), .Y(
        sub_398_S2_I3_aco_carry[4]) );
  XNOR2XL U951 ( .A(sub_398_S2_I3_aco_carry[3]), .B(N1220), .Y(N1229) );
  OR2X1 U952 ( .A(sub_398_S2_I3_aco_carry[2]), .B(N1219), .Y(
        sub_398_S2_I3_aco_carry[3]) );
  XNOR2XL U953 ( .A(sub_398_S2_I3_aco_carry[2]), .B(N1219), .Y(N1228) );
  OR2X1 U954 ( .A(n713), .B(n82), .Y(sub_398_S2_I3_aco_carry[2]) );
  XNOR2XL U955 ( .A(n713), .B(n82), .Y(N1227) );
  OR2X1 U956 ( .A(sub_398_S2_I11_aco_carry[3]), .B(N1548), .Y(
        sub_398_S2_I11_aco_carry[4]) );
  OR2X1 U957 ( .A(sub_398_S2_I11_aco_carry[2]), .B(N1219), .Y(
        sub_398_S2_I11_aco_carry[3]) );
  OR2X1 U958 ( .A(n713), .B(n87), .Y(sub_398_S2_I11_aco_carry[2]) );
  OR2X1 U959 ( .A(sub_398_S2_I14_aco_carry[3]), .B(N1671), .Y(
        sub_398_S2_I14_aco_carry[4]) );
  AOI21X1 U960 ( .B(N1139), .C(n712), .A(N1140), .Y(n717) );
  OAI21X1 U961 ( .B(N1137), .C(N1136), .A(N1139), .Y(n716) );
  AOI21X1 U962 ( .B(N1221), .C(N1220), .A(N1222), .Y(n719) );
  OAI21X1 U963 ( .B(N1219), .C(n713), .A(N1221), .Y(n718) );
  AOI21X1 U964 ( .B(N1262), .C(n697), .A(N1263), .Y(n720) );
  AOI21X1 U965 ( .B(N1303), .C(n696), .A(N1304), .Y(n722) );
  OAI21X1 U966 ( .B(n714), .C(N1136), .A(N1303), .Y(n721) );
  AOI21X1 U967 ( .B(N1344), .C(N1343), .A(N1345), .Y(n723) );
  AOI21X1 U968 ( .B(N1385), .C(N1384), .A(N1386), .Y(n725) );
  OAI21X1 U969 ( .B(n702), .C(n713), .A(N1385), .Y(n724) );
  AOI21X1 U970 ( .B(N1426), .C(N1425), .A(N1427), .Y(n726) );
  AOI21X1 U971 ( .B(N1467), .C(N1466), .A(N1468), .Y(n728) );
  OAI21X1 U972 ( .B(N1137), .C(N1136), .A(N1467), .Y(n727) );
  NAND2X1 U973 ( .A(n728), .B(n727), .Y(N1469) );
  AOI21X1 U974 ( .B(N1549), .C(N1548), .A(N1550), .Y(n730) );
  OAI21X1 U975 ( .B(N1219), .C(n713), .A(N1549), .Y(n729) );
  AOI21X1 U976 ( .B(n698), .C(N1589), .A(n106), .Y(n731) );
  AOI21X1 U977 ( .B(N1631), .C(N1630), .A(N1632), .Y(n733) );
  OAI21X1 U978 ( .B(n714), .C(N1136), .A(N1631), .Y(n732) );
  NAND2X1 U979 ( .A(n733), .B(n732), .Y(N1633) );
  AOI21X1 U980 ( .B(N1672), .C(N1671), .A(N1673), .Y(n734) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_LOW_shmux_00000005_00000012_00000012 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLNXL latch ( .CKN(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dac2sar_a0 ( r_dac_t, r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, 
        auto_sar, busy, stop, sync_i, ps_sample, sampl_begn, sampl_done, 
        sh_rst, dacyc_done, sacyc_done, dac_v, rpt_v, clk, srstz );
  input [1:0] r_dac_t;
  output [9:0] dac_v;
  output [9:0] rpt_v;
  input r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, auto_sar, busy, stop,
         sync_i, ps_sample, clk, srstz;
  output sampl_begn, sampl_done, sh_rst, dacyc_done, sacyc_done;
  wire   n117, N31, N32, N33, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N71, N72, N73, N74, N75, N79, updlo, updup,
         upd1v, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, net10243, net10249, n87,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n126, n127, n128, n129, net96943, net96947, net96949, net121241,
         net146888, net146896, net146899, net146965, net146968, net146970,
         net146971, net146973, net146976, net146978, net146980, net146984,
         net146989, net146992, net146995, net146996, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n111, n112, n113, n114, n115, n116,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3;
  wire   [3:0] sarcyc;
  wire   [6:0] dacnt;
  wire   [9:0] r_lt_lo;
  wire   [9:0] r_lt_up;
  wire   [9:0] r_avg00;
  wire   [9:0] r_avgup;
  wire   [9:0] r_dacvo;

  glreg_WIDTH10_2 u0_dac1v ( .clk(clk), .arstz(n47), .we(upd1v), .wdat(r_dacvo), .rdat({dac_v[9:1], n117}) );
  glreg_WIDTH10_1 u0_lt_lo ( .clk(clk), .arstz(n46), .we(updlo), .wdat({n41, 
        n40, n39, n38, n37, n36, n35, n34, n32, n33}), .rdat(r_lt_lo) );
  glreg_WIDTH10_0 u0_lt_up ( .clk(clk), .arstz(n45), .we(updup), .wdat(r_avgup), .rdat(r_lt_up) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 clk_gate_dacnt_reg ( .CLK(clk), .EN(N54), 
        .ENCLK(net10243), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 clk_gate_sarcyc_reg ( .CLK(clk), .EN(N71), 
        .ENCLK(net10249), .TE(1'b0) );
  dac2sar_a0_DW01_add_0 add_312 ( .A({1'b0, n85, n86, n89, n91, n93, n95, n97, 
        n111, n113, n115}), .B({1'b0, n84, n88, n90, n92, n94, n96, n98, n112, 
        n114, n116}), .CI(1'b0), .SUM({N102, N101, N100, N99, N98, N97, N96, 
        N95, N94, N93, SYNOPSYS_UNCONNECTED_1}), .CO() );
  dac2sar_a0_DW01_add_1 add_310 ( .A({1'b0, n41, n40, n39, n38, n37, n36, n35, 
        n34, n32, n33}), .B({1'b0, r_avgup}), .CI(1'b0), .SUM({N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, SYNOPSYS_UNCONNECTED_2}), .CO() );
  dac2sar_a0_DW01_add_2 add_305 ( .A({1'b0, r_lt_lo}), .B({1'b0, r_lt_up}), 
        .CI(1'b0), .SUM({r_avg00, SYNOPSYS_UNCONNECTED_3}), .CO() );
  dac2sar_a0_DW01_inc_0 add_285 ( .A(dacnt), .SUM({N53, N52, N51, N50, N49, 
        N48, N47}) );
  DFFQX1 dacnt_reg_0_ ( .D(N55), .C(net10243), .Q(dacnt[0]) );
  DFFQX1 dacnt_reg_1_ ( .D(N56), .C(net10243), .Q(dacnt[1]) );
  DFFQX1 dacnt_reg_3_ ( .D(N58), .C(net10243), .Q(dacnt[3]) );
  DFFQX1 sarcyc_reg_3_ ( .D(N75), .C(net10249), .Q(sarcyc[3]) );
  DFFQX1 sarcyc_reg_0_ ( .D(N72), .C(net10249), .Q(sarcyc[0]) );
  DFFQX1 dacnt_reg_2_ ( .D(N57), .C(net10243), .Q(dacnt[2]) );
  DFFQX1 dacnt_reg_4_ ( .D(N59), .C(net10243), .Q(dacnt[4]) );
  DFFQX1 dacnt_reg_5_ ( .D(N60), .C(net10243), .Q(dacnt[5]) );
  DFFQX1 dacnt_reg_6_ ( .D(N61), .C(net10243), .Q(dacnt[6]) );
  DFFQX1 sarcyc_reg_1_ ( .D(N73), .C(net10249), .Q(sarcyc[1]) );
  DFFQX1 sarcyc_reg_2_ ( .D(N74), .C(net10249), .Q(sarcyc[2]) );
  DFFNQX1 sh_rst_n_reg ( .D(N79), .XC(clk), .Q(sh_rst) );
  MUX2IX2 U3 ( .D0(n5), .D1(n6), .S(ps_sample), .Y(n4) );
  NOR32X4 U4 ( .B(net121241), .C(dacnt[1]), .A(n4), .Y(sampl_done) );
  NOR43XL U5 ( .B(n7), .C(n8), .D(n9), .A(n10), .Y(n6) );
  NAND31X1 U6 ( .C(n11), .A(n12), .B(n13), .Y(n10) );
  XOR2X1 U7 ( .A(n26), .B(r_dacyc), .Y(n13) );
  INVX1 U8 ( .A(dacnt[2]), .Y(n26) );
  NAND4X1 U9 ( .A(net96943), .B(n26), .C(n109), .D(n110), .Y(n87) );
  XOR2X1 U10 ( .A(r_dacyc), .B(dacnt[3]), .Y(n12) );
  NAND31X1 U14 ( .C(n14), .A(n25), .B(sarcyc[0]), .Y(n11) );
  INVX1 U15 ( .A(net146888), .Y(n8) );
  XOR2X1 U16 ( .A(n15), .B(r_dacyc), .Y(n7) );
  INVX1 U17 ( .A(dacnt[4]), .Y(n15) );
  XOR2X1 U18 ( .A(n15), .B(n126), .Y(net146992) );
  NOR43XL U19 ( .B(n16), .C(n17), .D(n18), .A(n19), .Y(n5) );
  NAND21X1 U20 ( .B(n20), .A(n21), .Y(n19) );
  XOR2X1 U21 ( .A(net146896), .B(dacnt[6]), .Y(n21) );
  XOR2X1 U22 ( .A(N32), .B(dacnt[3]), .Y(n20) );
  XNOR2XL U23 ( .A(N31), .B(dacnt[2]), .Y(n18) );
  XNOR2XL U24 ( .A(N33), .B(dacnt[4]), .Y(n17) );
  XNOR2XL U25 ( .A(net146896), .B(dacnt[5]), .Y(n16) );
  XOR2X1 U26 ( .A(n23), .B(r_sar10), .Y(n9) );
  NAND5XL U27 ( .A(dacyc_done), .B(sarcyc[0]), .C(n25), .D(n9), .E(n24), .Y(
        net146980) );
  INVX1 U28 ( .A(sarcyc[3]), .Y(n23) );
  MUX2X1 U29 ( .D0(n23), .D1(net146973), .S(sarcyc[2]), .Y(n22) );
  OAI22X1 U30 ( .A(n22), .B(net146970), .C(net146971), .D(n23), .Y(N75) );
  XOR2X1 U31 ( .A(dacnt[2]), .B(n129), .Y(net146989) );
  XNOR2XL U32 ( .A(sarcyc[2]), .B(r_sar10), .Y(n14) );
  INVX1 U33 ( .A(n14), .Y(n24) );
  XNOR2XL U34 ( .A(net146984), .B(r_sar10), .Y(n25) );
  INVX1 U35 ( .A(sarcyc[1]), .Y(net146984) );
  BUFX3 U36 ( .A(semi_nxt), .Y(n27) );
  BUFX3 U37 ( .A(sar_ini), .Y(n28) );
  INVX1 U38 ( .A(n117), .Y(n29) );
  INVX1 U39 ( .A(n29), .Y(dac_v[0]) );
  INVX1 U40 ( .A(n29), .Y(n31) );
  INVX1 U41 ( .A(sar_ini), .Y(n61) );
  OR2XL U42 ( .A(stop), .B(n48), .Y(n60) );
  NOR2XL U43 ( .A(sar_ini), .B(n107), .Y(n32) );
  NOR2XL U44 ( .A(sar_ini), .B(n106), .Y(n34) );
  NOR2XL U45 ( .A(sar_ini), .B(n108), .Y(n33) );
  NAND2XL U46 ( .A(n76), .B(n61), .Y(r_avgup[2]) );
  NOR2XL U47 ( .A(sar_ini), .B(n105), .Y(n35) );
  NOR2XL U48 ( .A(sar_ini), .B(n104), .Y(n36) );
  NOR2XL U49 ( .A(sar_ini), .B(n103), .Y(n37) );
  NOR2XL U50 ( .A(sar_ini), .B(n102), .Y(n38) );
  NOR2XL U51 ( .A(sar_ini), .B(n101), .Y(n39) );
  NOR2XL U52 ( .A(n28), .B(n100), .Y(n40) );
  NOR2XL U53 ( .A(n28), .B(n99), .Y(n41) );
  AO21XL U54 ( .B(sar_nxt), .C(sync_i), .A(n28), .Y(updlo) );
  INVX1 U55 ( .A(n48), .Y(n46) );
  INVX1 U56 ( .A(n48), .Y(n47) );
  INVX1 U57 ( .A(srstz), .Y(n48) );
  INVX1 U58 ( .A(n48), .Y(n45) );
  NAND32X1 U59 ( .B(dacyc_done), .C(n60), .A(n59), .Y(N54) );
  OR2X1 U60 ( .A(net146965), .B(n58), .Y(N71) );
  INVX1 U61 ( .A(n59), .Y(n53) );
  INVX1 U62 ( .A(net146970), .Y(net146965) );
  INVX1 U63 ( .A(net146971), .Y(net146976) );
  INVX1 U64 ( .A(net146896), .Y(net146899) );
  NAND2X1 U65 ( .A(n75), .B(n61), .Y(r_avgup[1]) );
  MUX2X1 U66 ( .D0(N91), .D1(r_avg00[9]), .S(n27), .Y(r_dacvo[9]) );
  MUX2X1 U67 ( .D0(N90), .D1(r_avg00[8]), .S(n27), .Y(r_dacvo[8]) );
  MUX2X1 U68 ( .D0(N89), .D1(r_avg00[7]), .S(semi_nxt), .Y(r_dacvo[7]) );
  NAND2X1 U69 ( .A(n74), .B(n61), .Y(r_avgup[0]) );
  NAND2XL U70 ( .A(n77), .B(n61), .Y(r_avgup[3]) );
  MUX2X1 U71 ( .D0(N87), .D1(r_avg00[5]), .S(semi_nxt), .Y(r_dacvo[5]) );
  MUX2X1 U72 ( .D0(N88), .D1(r_avg00[6]), .S(semi_nxt), .Y(r_dacvo[6]) );
  NAND2XL U73 ( .A(n78), .B(n61), .Y(r_avgup[4]) );
  NAND2XL U74 ( .A(n79), .B(n61), .Y(r_avgup[5]) );
  MUX2X1 U75 ( .D0(N86), .D1(r_avg00[4]), .S(semi_nxt), .Y(r_dacvo[4]) );
  NAND2XL U76 ( .A(n80), .B(n61), .Y(r_avgup[6]) );
  MUX2X1 U77 ( .D0(N84), .D1(r_avg00[2]), .S(semi_nxt), .Y(r_dacvo[2]) );
  MUX2X1 U78 ( .D0(N85), .D1(r_avg00[3]), .S(semi_nxt), .Y(r_dacvo[3]) );
  NAND2XL U79 ( .A(n81), .B(n61), .Y(r_avgup[7]) );
  NAND2XL U80 ( .A(n82), .B(n61), .Y(r_avgup[8]) );
  MUX2X1 U81 ( .D0(N83), .D1(r_avg00[1]), .S(semi_nxt), .Y(r_dacvo[1]) );
  NAND2XL U82 ( .A(n83), .B(n61), .Y(r_avgup[9]) );
  MUX2X1 U83 ( .D0(N82), .D1(r_avg00[0]), .S(semi_nxt), .Y(r_dacvo[0]) );
  OR3XL U84 ( .A(sar_nxt), .B(n28), .C(semi_nxt), .Y(upd1v) );
  NAND31X1 U85 ( .C(n60), .A(busy), .B(net146978), .Y(n59) );
  NAND21X1 U86 ( .B(n57), .A(net146965), .Y(net146971) );
  NAND32X1 U87 ( .B(net146978), .C(n58), .A(auto_sar), .Y(net146970) );
  OR2X1 U88 ( .A(sacyc_done), .B(n60), .Y(n58) );
  AND2X1 U89 ( .A(net146976), .B(n55), .Y(N73) );
  AND2X1 U90 ( .A(N52), .B(n53), .Y(N60) );
  AND2X1 U91 ( .A(N51), .B(n53), .Y(N59) );
  AND2X1 U92 ( .A(N50), .B(n53), .Y(N58) );
  AND2X1 U93 ( .A(N49), .B(n53), .Y(N57) );
  AND2X1 U94 ( .A(N48), .B(n53), .Y(N56) );
  AND2X1 U95 ( .A(net146965), .B(net146968), .Y(N72) );
  NAND21X1 U96 ( .B(N32), .A(n73), .Y(net146896) );
  INVX1 U97 ( .A(n127), .Y(n73) );
  NOR32XL U98 ( .B(busy), .C(net121241), .A(n87), .Y(N79) );
  INVX1 U99 ( .A(net96947), .Y(n109) );
  INVX1 U100 ( .A(net146978), .Y(dacyc_done) );
  INVX1 U101 ( .A(n82), .Y(n88) );
  INVX1 U102 ( .A(n100), .Y(n86) );
  INVX1 U103 ( .A(n99), .Y(n85) );
  INVX1 U104 ( .A(n83), .Y(n84) );
  INVX1 U105 ( .A(r_avg00[8]), .Y(n63) );
  INVX1 U106 ( .A(n106), .Y(n111) );
  INVX1 U107 ( .A(n76), .Y(n112) );
  INVX1 U108 ( .A(n105), .Y(n97) );
  INVX1 U109 ( .A(n77), .Y(n98) );
  INVX1 U110 ( .A(n104), .Y(n95) );
  INVX1 U111 ( .A(n78), .Y(n96) );
  INVX1 U112 ( .A(n103), .Y(n93) );
  INVX1 U113 ( .A(n79), .Y(n94) );
  INVX1 U114 ( .A(n102), .Y(n91) );
  INVX1 U115 ( .A(n80), .Y(n92) );
  INVX1 U116 ( .A(n81), .Y(n90) );
  INVX1 U117 ( .A(n101), .Y(n89) );
  INVX1 U118 ( .A(n107), .Y(n113) );
  INVX1 U119 ( .A(n75), .Y(n114) );
  INVX1 U120 ( .A(r_avg00[9]), .Y(n62) );
  INVX1 U121 ( .A(r_avg00[0]), .Y(n71) );
  INVX1 U122 ( .A(r_avg00[1]), .Y(n70) );
  INVX1 U123 ( .A(r_avg00[2]), .Y(n69) );
  INVX1 U124 ( .A(r_avg00[3]), .Y(n68) );
  INVX1 U125 ( .A(r_avg00[4]), .Y(n67) );
  INVX1 U126 ( .A(r_avg00[5]), .Y(n66) );
  INVX1 U127 ( .A(r_avg00[6]), .Y(n65) );
  INVX1 U128 ( .A(r_avg00[7]), .Y(n64) );
  INVX1 U129 ( .A(n74), .Y(n116) );
  INVX1 U130 ( .A(n108), .Y(n115) );
  INVX1 U131 ( .A(n44), .Y(n42) );
  INVX1 U132 ( .A(n44), .Y(n43) );
  NOR2X1 U133 ( .A(net121241), .B(n87), .Y(sampl_begn) );
  AO21XL U134 ( .B(sar_nxt), .C(n44), .A(n28), .Y(updup) );
  ENOX1 U135 ( .A(n31), .B(n80), .C(N99), .D(n31), .Y(rpt_v[6]) );
  MUX2X1 U136 ( .D0(n56), .D1(net146976), .S(sarcyc[2]), .Y(N74) );
  AND2X1 U137 ( .A(n57), .B(net146965), .Y(n56) );
  AND2X1 U138 ( .A(N53), .B(n53), .Y(N61) );
  AND2X1 U139 ( .A(N47), .B(n53), .Y(N55) );
  NAND21X1 U140 ( .B(sarcyc[3]), .A(n57), .Y(net146973) );
  ENOX1 U141 ( .A(n31), .B(n82), .C(N101), .D(n31), .Y(rpt_v[8]) );
  ENOX1 U142 ( .A(n117), .B(n83), .C(n117), .D(N102), .Y(rpt_v[9]) );
  ENOX1 U143 ( .A(n117), .B(n81), .C(N100), .D(n117), .Y(rpt_v[7]) );
  ENOX1 U144 ( .A(n31), .B(n76), .C(N95), .D(n31), .Y(rpt_v[2]) );
  ENOX1 U145 ( .A(n117), .B(n78), .C(N97), .D(dac_v[0]), .Y(rpt_v[4]) );
  ENOX1 U146 ( .A(n31), .B(n79), .C(N98), .D(n31), .Y(rpt_v[5]) );
  ENOX1 U147 ( .A(n31), .B(n74), .C(N93), .D(n31), .Y(rpt_v[0]) );
  AO21X1 U148 ( .B(n73), .C(n72), .A(net146899), .Y(N33) );
  INVX1 U149 ( .A(r_dac_t[0]), .Y(n72) );
  ENOX1 U150 ( .A(n117), .B(n75), .C(N94), .D(n117), .Y(rpt_v[1]) );
  ENOX1 U151 ( .A(n117), .B(n77), .C(N96), .D(n117), .Y(rpt_v[3]) );
  NOR2X1 U152 ( .A(r_dac_t[1]), .B(r_dac_t[0]), .Y(n127) );
  AOI21X1 U153 ( .B(r_dac_t[0]), .C(r_dac_t[1]), .A(n127), .Y(N32) );
  NOR2X1 U154 ( .A(n127), .B(r_dac_t[1]), .Y(N31) );
  OR3XL U155 ( .A(sarcyc[2]), .B(sarcyc[3]), .C(n55), .Y(net96947) );
  NAND21X1 U156 ( .B(sarcyc[0]), .A(net146984), .Y(n55) );
  NAND21X1 U157 ( .B(dacnt[6]), .A(net146995), .Y(net146888) );
  INVX1 U158 ( .A(dacnt[1]), .Y(net96943) );
  NOR4XL U159 ( .A(dacnt[6]), .B(dacnt[5]), .C(dacnt[4]), .D(dacnt[3]), .Y(
        n110) );
  INVX1 U160 ( .A(dacnt[5]), .Y(net146995) );
  INVX1 U161 ( .A(dacnt[0]), .Y(net121241) );
  NAND5XL U162 ( .A(dacnt[1]), .B(dacnt[0]), .C(n52), .D(net146989), .E(n51), 
        .Y(net146978) );
  XOR2X1 U163 ( .A(dacnt[3]), .B(n128), .Y(n52) );
  AOI211X1 U164 ( .C(dacnt[6]), .D(dacnt[5]), .A(n50), .B(net146992), .Y(n51)
         );
  AOI22X1 U165 ( .A(n109), .B(N33), .C(net96947), .D(r_dacyc), .Y(n126) );
  INVX1 U166 ( .A(net146980), .Y(sacyc_done) );
  MUX2X1 U167 ( .D0(net146888), .D1(n49), .S(n109), .Y(n50) );
  MUX2X1 U168 ( .D0(net146995), .D1(net146996), .S(net146899), .Y(n49) );
  INVX1 U169 ( .A(dacnt[6]), .Y(net146996) );
  AOI22X1 U170 ( .A(N31), .B(n109), .C(net96947), .D(r_dacyc), .Y(n129) );
  AOI22X1 U171 ( .A(N32), .B(n109), .C(net96947), .D(net96949), .Y(n128) );
  INVX1 U172 ( .A(r_dacyc), .Y(net96949) );
  MUX2AXL U173 ( .D0(r_lt_lo[8]), .D1(n63), .S(n42), .Y(n100) );
  MUX2BXL U174 ( .D0(n69), .D1(r_lt_up[2]), .S(n43), .Y(n76) );
  MUX2BXL U175 ( .D0(n68), .D1(r_lt_up[3]), .S(n43), .Y(n77) );
  MUX2BXL U176 ( .D0(n67), .D1(r_lt_up[4]), .S(n43), .Y(n78) );
  MUX2BXL U177 ( .D0(n66), .D1(r_lt_up[5]), .S(n43), .Y(n79) );
  MUX2BXL U178 ( .D0(n65), .D1(r_lt_up[6]), .S(n43), .Y(n80) );
  MUX2BXL U179 ( .D0(n64), .D1(r_lt_up[7]), .S(n43), .Y(n81) );
  MUX2BXL U180 ( .D0(n63), .D1(r_lt_up[8]), .S(n43), .Y(n82) );
  MUX2BXL U181 ( .D0(n62), .D1(r_lt_up[9]), .S(n42), .Y(n83) );
  MUX2BXL U182 ( .D0(n71), .D1(r_lt_up[0]), .S(n43), .Y(n74) );
  MUX2BXL U183 ( .D0(n70), .D1(r_lt_up[1]), .S(n43), .Y(n75) );
  MUX2AXL U184 ( .D0(r_lt_lo[0]), .D1(n71), .S(n43), .Y(n108) );
  MUX2AXL U185 ( .D0(r_lt_lo[1]), .D1(n70), .S(n42), .Y(n107) );
  MUX2AXL U186 ( .D0(r_lt_lo[2]), .D1(n69), .S(n42), .Y(n106) );
  MUX2AXL U187 ( .D0(r_lt_lo[3]), .D1(n68), .S(n42), .Y(n105) );
  MUX2AXL U188 ( .D0(r_lt_lo[4]), .D1(n67), .S(n42), .Y(n104) );
  MUX2AXL U189 ( .D0(r_lt_lo[5]), .D1(n66), .S(n42), .Y(n103) );
  MUX2AXL U190 ( .D0(r_lt_lo[6]), .D1(n65), .S(n42), .Y(n102) );
  MUX2AXL U191 ( .D0(r_lt_lo[7]), .D1(n64), .S(n42), .Y(n101) );
  MUX2AXL U192 ( .D0(r_lt_lo[9]), .D1(n62), .S(n42), .Y(n99) );
  INVX1 U193 ( .A(sync_i), .Y(n44) );
  INVX1 U194 ( .A(n54), .Y(n57) );
  NAND21X1 U195 ( .B(net146968), .A(sarcyc[1]), .Y(n54) );
  INVX1 U196 ( .A(sarcyc[0]), .Y(net146968) );
endmodule


module dac2sar_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module dac2sar_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module dac2sar_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module dac2sar_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_0 ( clk, arstz, we, wdat, rdat );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we;
  wire   net10266;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10266), .TE(1'b0) );
  DFFRQX1 mem_reg_9_ ( .D(wdat[9]), .C(net10266), .XR(arstz), .Q(rdat[9]) );
  DFFRQX1 mem_reg_8_ ( .D(wdat[8]), .C(net10266), .XR(arstz), .Q(rdat[8]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10266), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10266), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10266), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10266), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10266), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10266), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10266), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10266), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_1 ( clk, arstz, we, wdat, rdat );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we;
  wire   net10284;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10284), .TE(1'b0) );
  DFFRQX1 mem_reg_9_ ( .D(wdat[9]), .C(net10284), .XR(arstz), .Q(rdat[9]) );
  DFFRQX1 mem_reg_8_ ( .D(wdat[8]), .C(net10284), .XR(arstz), .Q(rdat[8]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10284), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10284), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10284), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10284), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10284), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10284), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10284), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10284), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_2 ( clk, arstz, we, wdat, rdat );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we;
  wire   net10302;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10302), .TE(1'b0) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10302), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10302), .XR(arstz), .Q(rdat[0]) );
  DFFRQXL mem_reg_9_ ( .D(wdat[9]), .C(net10302), .XR(arstz), .Q(rdat[9]) );
  DFFRQXL mem_reg_8_ ( .D(wdat[8]), .C(net10302), .XR(arstz), .Q(rdat[8]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10302), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10302), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10302), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10302), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10302), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10302), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_00000012 ( clk, arstz, we, wdat, rdat );
  input [17:0] wdat;
  output [17:0] rdat;
  input clk, arstz, we;
  wire   net10320, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_glreg_00000012 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10320), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10320), .XR(n2), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10320), .XR(n2), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10320), .XR(n2), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10320), .XR(n2), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10320), .XR(n2), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10320), .XR(n2), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10320), .XR(n2), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10320), .XR(n2), .Q(rdat[0]) );
  DFFRQX1 mem_reg_13_ ( .D(wdat[13]), .C(net10320), .XR(n1), .Q(rdat[13]) );
  DFFRQX1 mem_reg_11_ ( .D(wdat[11]), .C(net10320), .XR(n1), .Q(rdat[11]) );
  DFFRQX1 mem_reg_9_ ( .D(wdat[9]), .C(net10320), .XR(n1), .Q(rdat[9]) );
  DFFRQX1 mem_reg_17_ ( .D(wdat[17]), .C(net10320), .XR(n1), .Q(rdat[17]) );
  DFFRQX1 mem_reg_14_ ( .D(wdat[14]), .C(net10320), .XR(n1), .Q(rdat[14]) );
  DFFRQX1 mem_reg_12_ ( .D(wdat[12]), .C(net10320), .XR(n1), .Q(rdat[12]) );
  DFFRQX1 mem_reg_10_ ( .D(wdat[10]), .C(net10320), .XR(n1), .Q(rdat[10]) );
  DFFRQX1 mem_reg_8_ ( .D(wdat[8]), .C(net10320), .XR(n1), .Q(rdat[8]) );
  DFFRQX1 mem_reg_16_ ( .D(wdat[16]), .C(net10320), .XR(n1), .Q(rdat[16]) );
  DFFRQX1 mem_reg_15_ ( .D(wdat[15]), .C(net10320), .XR(n1), .Q(rdat[15]) );
  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(arstz), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_00000012 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( i_cc, i_cc_49, i_sqlch, r_sqlch, 
        r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, 
        r_fiforst, r_unlock, r_first, r_last, r_set_cpmsgid, r_rdy, r_wdat, 
        r_rdat, r_txnumk, r_txendk, r_txshrt, r_auto_discard, r_txauto, 
        r_rxords_ena, r_spec, r_dat_spec, r_auto_gdcrc, r_rxdb_opt, r_pshords, 
        r_dat_portrole, r_dat_datarole, r_discard, pid_goidle, pid_gobusy, 
        pff_ack, pff_rdat, pff_rxpart, prx_rcvinf, pff_obsd, pff_ptr, 
        pff_empty, pff_full, ptx_ack, ptx_cc, ptx_oe, prx_setsta, prx_rst, 
        prl_c0set, prl_cany0, prl_cany0r, prl_cany0w, prl_discard, 
        prl_GCTxDone, prl_cany0adr, prl_cpmsgid, prx_fifowdat, ptx_fsm, 
        prl_fsm, prx_fsm, prx_adpn, dbgpo, clk, srstz );
  input [1:0] r_sqlch;
  input [7:0] r_wdat;
  input [7:0] r_rdat;
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [6:0] r_rxords_ena;
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [1:0] r_auto_gdcrc;
  input [1:0] r_rxdb_opt;
  output [1:0] pff_ack;
  output [7:0] pff_rdat;
  output [15:0] pff_rxpart;
  output [4:0] prx_rcvinf;
  output [5:0] pff_ptr;
  output [6:0] prx_setsta;
  output [1:0] prx_rst;
  output [7:0] prl_cany0adr;
  output [2:0] prl_cpmsgid;
  output [7:0] prx_fifowdat;
  output [2:0] ptx_fsm;
  output [3:0] prl_fsm;
  output [3:0] prx_fsm;
  output [5:0] prx_adpn;
  output [31:0] dbgpo;
  input i_cc, i_cc_49, i_sqlch, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4,
         r_fifopsh, r_fifopop, r_fiforst, r_unlock, r_first, r_last,
         r_set_cpmsgid, r_rdy, r_txendk, r_txshrt, r_auto_discard, r_pshords,
         r_dat_portrole, r_dat_datarole, r_discard, clk, srstz;
  output pid_goidle, pid_gobusy, pff_obsd, pff_empty, pff_full, ptx_ack,
         ptx_cc, ptx_oe, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_discard, prl_GCTxDone;
  wire   n66, dbgpo_29, rx_pshords, auto_rx_gdcrc, prx_trans, prx_fiforst,
         pcc_rxgood, prx_crcstart, prx_crcshfi4, prx_eoprcvd, x_trans,
         ptx_goidle, c0_txendk, mux_one, ptx_crcstart, ptx_crcshfi4,
         ptx_crcshfo4, crcstart, crcshfi4, crcshfo4, prl_idle, lockena,
         fifosrstz, fifopop_pff, fifopsh_pff, pff_txreq, pff_one, obsd,
         prl_last, prl_txreq, fifopop_prl, fifopsh_prl, prx_gdmsgrcvd, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, d_sqlch, net10338, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n3, n4, n5, n6, n7, n9, n10, n11,
         n13, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4;
  wire   [1:0] prx_cccnt;
  wire   [3:0] prx_crcsidat;
  wire   [4:0] c0_txnumk;
  wire   [6:0] c0_txauto;
  wire   [7:0] mux_rdat;
  wire   [3:0] ptx_crcsidat;
  wire   [3:0] crc32_3_0;
  wire   [3:0] crcsidat;
  wire   [55:0] pff_dat_7_1;
  wire   [47:16] pff_c0dat;
  wire   [7:0] prl_rdat;
  wire   [4:0] prl_txauto;
  wire   [1:0] d_cc;
  wire   [8:0] cclow_cnt;

  phyrx_a0 u0_phyrx ( .i_cc(i_cc), .ptx_txact(ptx_oe), .r_adprx_en(r_adprx_en), 
        .r_adp2nd(r_adp2nd), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), 
        .r_rxdb_opt(r_rxdb_opt), .r_ords_ena(r_rxords_ena), .r_pshords(
        rx_pshords), .r_rgdcrc(auto_rx_gdcrc), .prx_cccnt(prx_cccnt), 
        .prx_rst(prx_rst), .prx_setsta({prx_setsta[6:1], 
        SYNOPSYS_UNCONNECTED_1}), .prx_idle(), .prx_d_cc(dbgpo[17]), .prx_bmc(
        dbgpo[18]), .prx_trans(prx_trans), .prx_fiforst(prx_fiforst), 
        .prx_fifopsh(dbgpo_29), .prx_fifowdat(prx_fifowdat), .pff_txreq(n13), 
        .pid_gobusy(pid_gobusy), .pid_goidle(pid_goidle), .pid_ccidle(
        prx_rcvinf[4]), .pcc_rxgood(pcc_rxgood), .prx_crcstart(prx_crcstart), 
        .prx_crcshfi4(prx_crcshfi4), .prx_crcsidat(prx_crcsidat), .prx_rxcode(
        dbgpo[28:24]), .prx_adpn(prx_adpn), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_eoprcvd(prx_eoprcvd), .prx_fsm(prx_fsm), .clk(clk), .srstz(n47)
         );
  phyidd_a0 u0_phyidd ( .i_trans(x_trans), .i_goidle(ptx_goidle), .o_ccidle(
        prx_rcvinf[4]), .o_goidle(pid_goidle), .o_gobusy(pid_gobusy), .clk(clk), .srstz(n47) );
  phytx_a0 u0_phytx ( .r_txnumk(c0_txnumk), .r_txendk(c0_txendk), .r_txshrt(
        r_txshrt), .r_txauto(c0_txauto), .prx_cccnt(prx_cccnt), .ptx_txact(n66), .ptx_cc(ptx_cc), .ptx_goidle(ptx_goidle), .ptx_fifopop(dbgpo[30]), 
        .ptx_pspyld(), .i_rdat(mux_rdat), .i_txreq(n13), .i_one(mux_one), 
        .ptx_crcstart(ptx_crcstart), .ptx_crcshfi4(ptx_crcshfi4), 
        .ptx_crcshfo4(ptx_crcshfo4), .ptx_crcsidat(ptx_crcsidat), .ptx_fsm(
        ptx_fsm), .pcc_crc30(crc32_3_0), .clk(clk), .srstz(n47) );
  phycrc_a0 u0_phycrc ( .crc32_3_0(crc32_3_0), .rx_good(pcc_rxgood), 
        .i_shfidat(crcsidat), .i_start(crcstart), .i_shfi4(crcshfi4), 
        .i_shfo4(crcshfo4), .clk(clk) );
  phyff_DEPTH_NUM34_DEPTH_NBT6 u0_phyff ( .r_psh(r_fifopsh), .r_pop(r_fifopop), 
        .prx_psh(fifopsh_pff), .ptx_pop(fifopop_pff), .r_last(r_last), 
        .r_unlock(r_unlock), .i_lockena(lockena), .r_fiforst(r_fiforst), 
        .i_ccidle(prx_rcvinf[4]), .r_wdat(r_wdat), .prx_wdat(prx_fifowdat), 
        .txreq(pff_txreq), .ffack(pff_ack), .rdat0(pff_rdat), .full(pff_full), 
        .empty(pff_empty), .one(pff_one), .half(), .obsd(obsd), .dat_7_1(
        pff_dat_7_1), .ptr(pff_ptr), .fifowdat(dbgpo[7:0]), .fifopsh(dbgpo[16]), .clk(clk), .srstz(fifosrstz) );
  updprl_a0 u0_updprl ( .r_spec(r_spec), .r_dat_spec(r_dat_spec), 
        .r_auto_txgdcrc(r_auto_gdcrc[0]), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_auto_discard(r_auto_discard), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_dat_cpmsgid(r_wdat[2:0]), .r_rdat(
        r_rdat), .r_rdy(r_rdy), .pid_ccidle(prx_rcvinf[4]), .r_discard(
        r_discard), .ptx_ack(ptx_goidle), .ptx_txact(ptx_oe), .ptx_fifopop(
        fifopop_prl), .prx_fifopsh(fifopsh_prl), .prx_gdmsgrcvd(prx_gdmsgrcvd), 
        .prx_eoprcvd(prx_eoprcvd), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_fifowdat(prx_fifowdat), .pff_c0dat({pff_c0dat, pff_rxpart}), 
        .prl_rdat(prl_rdat), .prl_txauto({SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, prl_txauto[4], SYNOPSYS_UNCONNECTED_4, 
        prl_txauto[2:0]}), .prl_last(prl_last), .prl_txreq(prl_txreq), 
        .prl_c0set(prl_c0set), .prl_cany0(prl_cany0), .prl_cany0r(prl_cany0r), 
        .prl_cany0w(prl_cany0w), .prl_idle(prl_idle), .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_fsm(prl_fsm), .prl_cpmsgid(prl_cpmsgid), 
        .prl_cany0adr(prl_cany0adr), .clk(clk), .srstz(n46) );
  dbnc_WIDTH3 u0_sqlch_db ( .o_dbc(d_sqlch), .o_chg(), .i_org(i_sqlch), .clk(
        clk), .rstz(n46) );
  SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 clk_gate_cclow_cnt_reg ( 
        .CLK(clk), .EN(N34), .ENCLK(net10338), .TE(1'b0) );
  DFFSQX1 d_cc_reg_1_ ( .D(d_cc[0]), .C(clk), .XS(n47), .Q(d_cc[1]) );
  DFFSQX1 d_cc_reg_0_ ( .D(i_cc_49), .C(clk), .XS(n47), .Q(d_cc[0]) );
  DFFQX1 cclow_cnt_reg_2_ ( .D(N37), .C(net10338), .Q(cclow_cnt[2]) );
  DFFQX1 cclow_cnt_reg_3_ ( .D(N38), .C(net10338), .Q(cclow_cnt[3]) );
  DFFQX1 cclow_cnt_reg_4_ ( .D(N39), .C(net10338), .Q(cclow_cnt[4]) );
  DFFQX1 cclow_cnt_reg_5_ ( .D(N40), .C(net10338), .Q(cclow_cnt[5]) );
  DFFQX1 cclow_cnt_reg_6_ ( .D(N41), .C(net10338), .Q(cclow_cnt[6]) );
  DFFQX1 cclow_cnt_reg_8_ ( .D(N43), .C(net10338), .Q(cclow_cnt[8]) );
  DFFQX1 cclow_cnt_reg_7_ ( .D(N42), .C(net10338), .Q(cclow_cnt[7]) );
  DFFQX1 cclow_cnt_reg_1_ ( .D(N36), .C(net10338), .Q(cclow_cnt[1]) );
  DFFQX1 cclow_cnt_reg_0_ ( .D(N35), .C(net10338), .Q(cclow_cnt[0]) );
  INVX1 U3 ( .A(1'b1), .Y(dbgpo[31]) );
  MUX2X2 U5 ( .D0(prl_rdat[7]), .D1(pff_rdat[7]), .S(n41), .Y(mux_rdat[7]) );
  AND2X2 U6 ( .A(r_txnumk[1]), .B(n42), .Y(c0_txnumk[1]) );
  BUFX3 U7 ( .A(n43), .Y(n3) );
  INVXL U8 ( .A(n45), .Y(n43) );
  MUX2X2 U9 ( .D0(prl_last), .D1(pff_one), .S(n3), .Y(mux_one) );
  NAND2X1 U10 ( .A(n10), .B(n11), .Y(mux_rdat[0]) );
  AND2X1 U11 ( .A(r_txnumk[2]), .B(n42), .Y(c0_txnumk[2]) );
  INVX1 U12 ( .A(n54), .Y(n53) );
  NAND2X1 U13 ( .A(prl_rdat[3]), .B(n4), .Y(n5) );
  NAND2X1 U14 ( .A(pff_rdat[3]), .B(n42), .Y(n6) );
  NAND2X1 U15 ( .A(n5), .B(n6), .Y(mux_rdat[3]) );
  INVX1 U16 ( .A(n42), .Y(n4) );
  MUX2X1 U17 ( .D0(prl_rdat[6]), .D1(pff_rdat[6]), .S(n41), .Y(mux_rdat[6]) );
  MUX2X1 U18 ( .D0(prl_rdat[2]), .D1(pff_rdat[2]), .S(n41), .Y(mux_rdat[2]) );
  INVX1 U19 ( .A(r_pshords), .Y(n54) );
  INVX1 U20 ( .A(n66), .Y(n7) );
  INVX1 U21 ( .A(n7), .Y(ptx_oe) );
  INVX3 U22 ( .A(n45), .Y(n42) );
  INVX4 U23 ( .A(n44), .Y(n41) );
  NAND2X1 U24 ( .A(prl_rdat[0]), .B(n9), .Y(n10) );
  NAND2XL U25 ( .A(pff_rdat[0]), .B(n42), .Y(n11) );
  INVXL U26 ( .A(n42), .Y(n9) );
  MUX2X2 U27 ( .D0(prl_rdat[4]), .D1(pff_rdat[4]), .S(n42), .Y(mux_rdat[4]) );
  MUX2X2 U28 ( .D0(prl_rdat[1]), .D1(pff_rdat[1]), .S(n3), .Y(mux_rdat[1]) );
  BUFXL U29 ( .A(dbgpo_29), .Y(dbgpo[29]) );
  AND2X2 U30 ( .A(dbgpo[30]), .B(n44), .Y(fifopop_prl) );
  AO22XL U31 ( .A(ptx_crcstart), .B(n66), .C(prx_crcstart), .D(n7), .Y(
        crcstart) );
  BUFX3 U32 ( .A(prx_rcvinf[4]), .Y(dbgpo[19]) );
  BUFXL U33 ( .A(pff_rdat[0]), .Y(dbgpo[8]) );
  BUFXL U34 ( .A(pff_rdat[2]), .Y(dbgpo[10]) );
  BUFXL U35 ( .A(pff_rdat[3]), .Y(dbgpo[11]) );
  BUFXL U36 ( .A(pff_rdat[5]), .Y(dbgpo[13]) );
  BUFXL U37 ( .A(pff_rdat[6]), .Y(dbgpo[14]) );
  BUFXL U38 ( .A(pff_rdat[7]), .Y(dbgpo[15]) );
  BUFXL U39 ( .A(pff_rdat[1]), .Y(dbgpo[9]) );
  BUFXL U40 ( .A(pff_rdat[4]), .Y(dbgpo[12]) );
  BUFX3 U41 ( .A(prx_fsm[3]), .Y(dbgpo[23]) );
  BUFXL U42 ( .A(prx_fsm[0]), .Y(dbgpo[20]) );
  BUFXL U43 ( .A(prx_fsm[1]), .Y(dbgpo[21]) );
  BUFXL U44 ( .A(prx_fsm[2]), .Y(dbgpo[22]) );
  INVX2 U45 ( .A(prl_idle), .Y(n44) );
  AND2X2 U46 ( .A(dbgpo_29), .B(n44), .Y(fifopsh_prl) );
  AND2XL U47 ( .A(dbgpo[30]), .B(n3), .Y(fifopop_pff) );
  INVX2 U48 ( .A(prl_idle), .Y(n45) );
  AND2XL U49 ( .A(n53), .B(n3), .Y(rx_pshords) );
  MUX2XL U50 ( .D0(prl_txreq), .D1(pff_txreq), .S(n41), .Y(n13) );
  INVXL U51 ( .A(n54), .Y(n51) );
  INVXL U52 ( .A(n54), .Y(n52) );
  AND2X1 U53 ( .A(r_txnumk[3]), .B(n42), .Y(c0_txnumk[3]) );
  AND2X1 U54 ( .A(prx_setsta[3]), .B(n28), .Y(prx_gdmsgrcvd) );
  NOR21XL U55 ( .B(ptx_crcshfo4), .A(n7), .Y(crcshfo4) );
  NOR2X1 U56 ( .A(prx_fiforst), .B(n48), .Y(fifosrstz) );
  AO22X1 U57 ( .A(ptx_crcshfi4), .B(n66), .C(prx_crcshfi4), .D(n7), .Y(
        crcshfi4) );
  NOR21XL U58 ( .B(obsd), .A(prx_setsta[6]), .Y(pff_obsd) );
  NAND42X1 U59 ( .C(pff_rxpart[1]), .D(pff_rxpart[15]), .A(n29), .B(n30), .Y(
        n28) );
  NOR3XL U60 ( .A(pff_rxpart[2]), .B(pff_rxpart[4]), .C(pff_rxpart[3]), .Y(n29) );
  NOR41XL U61 ( .D(pff_rxpart[0]), .A(pff_rxpart[14]), .B(pff_rxpart[13]), .C(
        pff_rxpart[12]), .Y(n30) );
  INVX1 U62 ( .A(n54), .Y(n49) );
  INVX1 U63 ( .A(n54), .Y(n50) );
  INVX1 U64 ( .A(n48), .Y(n47) );
  INVX1 U65 ( .A(n48), .Y(n46) );
  NAND21X1 U66 ( .B(n36), .A(n35), .Y(n33) );
  INVX1 U67 ( .A(n34), .Y(n63) );
  NAND3X1 U68 ( .A(n34), .B(n33), .C(n35), .Y(N34) );
  MUX2X2 U69 ( .D0(prl_rdat[5]), .D1(pff_rdat[5]), .S(n3), .Y(mux_rdat[5]) );
  AND2X2 U70 ( .A(r_txnumk[0]), .B(n42), .Y(c0_txnumk[0]) );
  AND2XL U71 ( .A(r_txendk), .B(n3), .Y(c0_txendk) );
  AND2XL U72 ( .A(r_txnumk[4]), .B(n3), .Y(c0_txnumk[4]) );
  AND2XL U73 ( .A(r_txauto[6]), .B(n3), .Y(c0_txauto[6]) );
  AOI21AXL U74 ( .B(n66), .C(n3), .A(r_first), .Y(lockena) );
  NAND21XL U75 ( .B(r_txauto[5]), .A(n41), .Y(c0_txauto[5]) );
  MUX2X1 U76 ( .D0(pff_dat_7_1[8]), .D1(pff_dat_7_1[24]), .S(n49), .Y(
        pff_c0dat[16]) );
  MUX2X1 U77 ( .D0(pff_dat_7_1[10]), .D1(pff_dat_7_1[26]), .S(n49), .Y(
        pff_c0dat[18]) );
  MUX2X1 U78 ( .D0(pff_dat_7_1[16]), .D1(pff_dat_7_1[32]), .S(n50), .Y(
        pff_c0dat[24]) );
  MUX2X1 U79 ( .D0(pff_dat_7_1[13]), .D1(pff_dat_7_1[29]), .S(n50), .Y(
        pff_c0dat[21]) );
  AO22XL U80 ( .A(ptx_crcsidat[1]), .B(n66), .C(prx_crcsidat[1]), .D(n7), .Y(
        crcsidat[1]) );
  AO22XL U81 ( .A(ptx_crcsidat[0]), .B(n66), .C(prx_crcsidat[0]), .D(n7), .Y(
        crcsidat[0]) );
  MUX2XL U82 ( .D0(pff_dat_7_1[0]), .D1(pff_dat_7_1[16]), .S(n53), .Y(
        pff_rxpart[8]) );
  MUX2XL U83 ( .D0(pff_rdat[5]), .D1(pff_dat_7_1[13]), .S(n53), .Y(
        pff_rxpart[5]) );
  MUX2XL U84 ( .D0(pff_rdat[6]), .D1(pff_dat_7_1[14]), .S(n53), .Y(
        pff_rxpart[6]) );
  MUX2XL U85 ( .D0(pff_rdat[7]), .D1(pff_dat_7_1[15]), .S(n53), .Y(
        pff_rxpart[7]) );
  AO22XL U86 ( .A(ptx_crcsidat[3]), .B(n66), .C(prx_crcsidat[3]), .D(n7), .Y(
        crcsidat[3]) );
  AO22XL U87 ( .A(ptx_crcsidat[2]), .B(ptx_oe), .C(prx_crcsidat[2]), .D(n7), 
        .Y(crcsidat[2]) );
  MUX2X1 U88 ( .D0(pff_dat_7_1[4]), .D1(pff_dat_7_1[20]), .S(n49), .Y(
        pff_rxpart[12]) );
  MUX2X1 U89 ( .D0(pff_dat_7_1[5]), .D1(pff_dat_7_1[21]), .S(n49), .Y(
        pff_rxpart[13]) );
  MUX2XL U90 ( .D0(pff_rdat[3]), .D1(pff_dat_7_1[11]), .S(n52), .Y(
        pff_rxpart[3]) );
  MUX2XL U91 ( .D0(pff_rdat[2]), .D1(pff_dat_7_1[10]), .S(n51), .Y(
        pff_rxpart[2]) );
  MUX2XL U92 ( .D0(pff_rdat[0]), .D1(pff_dat_7_1[8]), .S(n49), .Y(
        pff_rxpart[0]) );
  MUX2XL U93 ( .D0(pff_rdat[4]), .D1(pff_dat_7_1[12]), .S(n53), .Y(
        pff_rxpart[4]) );
  NOR21XL U94 ( .B(r_auto_gdcrc[1]), .A(n28), .Y(auto_rx_gdcrc) );
  MUX2X1 U95 ( .D0(pff_dat_7_1[6]), .D1(pff_dat_7_1[22]), .S(n49), .Y(
        pff_rxpart[14]) );
  MUX2XL U96 ( .D0(pff_rdat[1]), .D1(pff_dat_7_1[9]), .S(n50), .Y(
        pff_rxpart[1]) );
  MUX2X1 U97 ( .D0(pff_dat_7_1[7]), .D1(pff_dat_7_1[23]), .S(n49), .Y(
        pff_rxpart[15]) );
  MUX2X1 U98 ( .D0(pff_dat_7_1[27]), .D1(pff_dat_7_1[43]), .S(n51), .Y(
        pff_c0dat[35]) );
  MUX2X1 U99 ( .D0(pff_dat_7_1[29]), .D1(pff_dat_7_1[45]), .S(n52), .Y(
        pff_c0dat[37]) );
  MUX2X1 U100 ( .D0(pff_dat_7_1[32]), .D1(pff_dat_7_1[48]), .S(n52), .Y(
        pff_c0dat[40]) );
  MUX2X1 U101 ( .D0(pff_dat_7_1[9]), .D1(pff_dat_7_1[25]), .S(n49), .Y(
        pff_c0dat[17]) );
  MUX2X1 U102 ( .D0(pff_dat_7_1[11]), .D1(pff_dat_7_1[27]), .S(n50), .Y(
        pff_c0dat[19]) );
  MUX2X1 U103 ( .D0(pff_dat_7_1[23]), .D1(pff_dat_7_1[39]), .S(n51), .Y(
        pff_c0dat[31]) );
  MUX2X1 U104 ( .D0(pff_dat_7_1[21]), .D1(pff_dat_7_1[37]), .S(n51), .Y(
        pff_c0dat[29]) );
  MUX2X1 U105 ( .D0(pff_dat_7_1[24]), .D1(pff_dat_7_1[40]), .S(n51), .Y(
        pff_c0dat[32]) );
  MUX2X1 U106 ( .D0(pff_dat_7_1[20]), .D1(pff_dat_7_1[36]), .S(n51), .Y(
        pff_c0dat[28]) );
  MUX2X1 U107 ( .D0(pff_dat_7_1[19]), .D1(pff_dat_7_1[35]), .S(n50), .Y(
        pff_c0dat[27]) );
  MUX2X1 U108 ( .D0(pff_dat_7_1[25]), .D1(pff_dat_7_1[41]), .S(n51), .Y(
        pff_c0dat[33]) );
  MUX2X1 U109 ( .D0(pff_dat_7_1[22]), .D1(pff_dat_7_1[38]), .S(n51), .Y(
        pff_c0dat[30]) );
  MUX2X1 U110 ( .D0(pff_dat_7_1[18]), .D1(pff_dat_7_1[34]), .S(n50), .Y(
        pff_c0dat[26]) );
  MUX2X1 U111 ( .D0(pff_dat_7_1[17]), .D1(pff_dat_7_1[33]), .S(n50), .Y(
        pff_c0dat[25]) );
  MUX2X1 U112 ( .D0(pff_dat_7_1[15]), .D1(pff_dat_7_1[31]), .S(n50), .Y(
        pff_c0dat[23]) );
  MUX2X1 U113 ( .D0(pff_dat_7_1[33]), .D1(pff_dat_7_1[49]), .S(n52), .Y(
        pff_c0dat[41]) );
  MUX2X1 U114 ( .D0(pff_dat_7_1[31]), .D1(pff_dat_7_1[47]), .S(n52), .Y(
        pff_c0dat[39]) );
  MUX2X1 U115 ( .D0(pff_dat_7_1[30]), .D1(pff_dat_7_1[46]), .S(n52), .Y(
        pff_c0dat[38]) );
  MUX2XL U116 ( .D0(pff_dat_7_1[38]), .D1(pff_dat_7_1[54]), .S(n53), .Y(
        pff_c0dat[46]) );
  MUX2X1 U117 ( .D0(pff_dat_7_1[14]), .D1(pff_dat_7_1[30]), .S(n50), .Y(
        pff_c0dat[22]) );
  MUX2X1 U118 ( .D0(pff_dat_7_1[12]), .D1(pff_dat_7_1[28]), .S(n50), .Y(
        pff_c0dat[20]) );
  MUX2X1 U119 ( .D0(pff_dat_7_1[35]), .D1(pff_dat_7_1[51]), .S(n52), .Y(
        pff_c0dat[43]) );
  MUX2X1 U120 ( .D0(pff_dat_7_1[28]), .D1(pff_dat_7_1[44]), .S(n51), .Y(
        pff_c0dat[36]) );
  MUX2X1 U121 ( .D0(pff_dat_7_1[34]), .D1(pff_dat_7_1[50]), .S(n52), .Y(
        pff_c0dat[42]) );
  MUX2X1 U122 ( .D0(pff_dat_7_1[26]), .D1(pff_dat_7_1[42]), .S(n51), .Y(
        pff_c0dat[34]) );
  MUX2X1 U123 ( .D0(pff_dat_7_1[36]), .D1(pff_dat_7_1[52]), .S(n52), .Y(
        pff_c0dat[44]) );
  MUX2XL U124 ( .D0(pff_dat_7_1[39]), .D1(pff_dat_7_1[55]), .S(n53), .Y(
        pff_c0dat[47]) );
  MUX2X1 U125 ( .D0(pff_dat_7_1[37]), .D1(pff_dat_7_1[53]), .S(n52), .Y(
        pff_c0dat[45]) );
  INVX1 U126 ( .A(srstz), .Y(n48) );
  MUX2XL U127 ( .D0(prl_txauto[0]), .D1(r_txauto[0]), .S(n41), .Y(c0_txauto[0]) );
  MUX2XL U128 ( .D0(prl_txauto[2]), .D1(r_txauto[2]), .S(n41), .Y(c0_txauto[2]) );
  MUX2XL U129 ( .D0(prl_txauto[1]), .D1(r_txauto[1]), .S(n41), .Y(c0_txauto[1]) );
  AOI31X1 U130 ( .A(d_sqlch), .B(n27), .C(r_sqlch[0]), .D(n62), .Y(x_trans) );
  OAI21X1 U131 ( .B(prx_fsm[3]), .C(n66), .A(r_sqlch[1]), .Y(n27) );
  INVX1 U132 ( .A(prx_trans), .Y(n62) );
  NAND21XL U133 ( .B(r_txauto[3]), .A(n41), .Y(c0_txauto[3]) );
  MUX2XL U134 ( .D0(prl_txauto[4]), .D1(r_txauto[4]), .S(n41), .Y(c0_txauto[4]) );
  NOR21XL U135 ( .B(ptx_goidle), .A(prl_cany0), .Y(ptx_ack) );
  OAI21BBX1 U136 ( .A(N33), .B(n63), .C(n33), .Y(N43) );
  NOR4XL U137 ( .A(n31), .B(n32), .C(cclow_cnt[5]), .D(cclow_cnt[4]), .Y(
        prx_setsta[0]) );
  OR3XL U138 ( .A(cclow_cnt[7]), .B(cclow_cnt[8]), .C(cclow_cnt[6]), .Y(n32)
         );
  NAND43X1 U139 ( .B(cclow_cnt[1]), .C(cclow_cnt[3]), .D(cclow_cnt[2]), .A(
        cclow_cnt[0]), .Y(n31) );
  AND2X1 U140 ( .A(N32), .B(n63), .Y(N42) );
  OAI21BBX1 U141 ( .A(N31), .B(n63), .C(n33), .Y(N41) );
  AOI21BBXL U142 ( .B(d_cc[1]), .C(n64), .A(n48), .Y(n35) );
  OAI211X1 U143 ( .C(n37), .D(n38), .A(n36), .B(n35), .Y(n34) );
  OR4X1 U144 ( .A(cclow_cnt[0]), .B(cclow_cnt[1]), .C(cclow_cnt[2]), .D(
        cclow_cnt[3]), .Y(n38) );
  NAND43X1 U145 ( .B(cclow_cnt[4]), .C(cclow_cnt[5]), .D(cclow_cnt[6]), .A(n39), .Y(n37) );
  NOR2X1 U146 ( .A(cclow_cnt[8]), .B(cclow_cnt[7]), .Y(n39) );
  MUX2XL U147 ( .D0(pff_dat_7_1[1]), .D1(pff_dat_7_1[17]), .S(n53), .Y(
        pff_rxpart[9]) );
  MUX2X1 U148 ( .D0(pff_dat_7_1[2]), .D1(pff_dat_7_1[18]), .S(n49), .Y(
        pff_rxpart[10]) );
  MUX2X1 U149 ( .D0(pff_dat_7_1[3]), .D1(pff_dat_7_1[19]), .S(n49), .Y(
        pff_rxpart[11]) );
  AND2X1 U150 ( .A(N25), .B(n63), .Y(N35) );
  AND2X1 U151 ( .A(N28), .B(n63), .Y(N38) );
  AND2X1 U152 ( .A(N27), .B(n63), .Y(N37) );
  OAI21BBX1 U153 ( .A(N30), .B(n63), .C(n33), .Y(N40) );
  OAI21BBX1 U154 ( .A(N29), .B(n63), .C(n33), .Y(N39) );
  OAI21BBX1 U155 ( .A(N26), .B(n63), .C(n33), .Y(N36) );
  NAND2X1 U156 ( .A(d_cc[1]), .B(n64), .Y(n36) );
  INVX1 U157 ( .A(d_cc[0]), .Y(n64) );
  BUFXL U158 ( .A(dbgpo[17]), .Y(prx_rcvinf[3]) );
  AND2XL U159 ( .A(dbgpo[29]), .B(n3), .Y(fifopsh_pff) );
  INVX1 U160 ( .A(cclow_cnt[0]), .Y(N25) );
  OR2X1 U161 ( .A(cclow_cnt[1]), .B(cclow_cnt[0]), .Y(n55) );
  OAI21BBX1 U162 ( .A(cclow_cnt[0]), .B(cclow_cnt[1]), .C(n55), .Y(N26) );
  OR2X1 U163 ( .A(n55), .B(cclow_cnt[2]), .Y(n56) );
  OAI21BBX1 U164 ( .A(n55), .B(cclow_cnt[2]), .C(n56), .Y(N27) );
  OR2X1 U165 ( .A(n56), .B(cclow_cnt[3]), .Y(n57) );
  OAI21BBX1 U166 ( .A(n56), .B(cclow_cnt[3]), .C(n57), .Y(N28) );
  OR2X1 U167 ( .A(n57), .B(cclow_cnt[4]), .Y(n58) );
  OAI21BBX1 U168 ( .A(n57), .B(cclow_cnt[4]), .C(n58), .Y(N29) );
  OR2X1 U169 ( .A(n58), .B(cclow_cnt[5]), .Y(n59) );
  OAI21BBX1 U170 ( .A(n58), .B(cclow_cnt[5]), .C(n59), .Y(N30) );
  OR2X1 U171 ( .A(n59), .B(cclow_cnt[6]), .Y(n60) );
  OAI21BBX1 U172 ( .A(n59), .B(cclow_cnt[6]), .C(n60), .Y(N31) );
  XNOR2XL U173 ( .A(n60), .B(cclow_cnt[7]), .Y(N32) );
  OR2X1 U174 ( .A(cclow_cnt[7]), .B(n60), .Y(n61) );
  XNOR2XL U175 ( .A(cclow_cnt[8]), .B(n61), .Y(N33) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N14, N15, N16, N17, net10356, n4, n5, n6, n7, n8, n1, n2,
         n3;
  wire   [2:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N14), 
        .ENCLK(net10356), .TE(1'b0) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N17), .C(net10356), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N16), .C(net10356), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N15), .C(net10356), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n8), .C(net10356), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n5), .A(n4), .Y(n6) );
  OAI32X1 U4 ( .A(n6), .B(n1), .C(n2), .D(n6), .E(n3), .Y(N17) );
  NOR2X1 U5 ( .A(n7), .B(n6), .Y(N16) );
  XNOR2XL U6 ( .A(n2), .B(n1), .Y(n7) );
  NAND4X1 U7 ( .A(n5), .B(n1), .C(n2), .D(n3), .Y(N14) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  AO22AXL U9 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n8) );
  NOR2X1 U10 ( .A(n4), .B(n5), .Y(o_chg) );
  NAND3X1 U11 ( .A(db_cnt[1]), .B(db_cnt[0]), .C(db_cnt[2]), .Y(n4) );
  NOR2X1 U12 ( .A(db_cnt[0]), .B(n6), .Y(N15) );
  INVX1 U13 ( .A(db_cnt[0]), .Y(n1) );
  INVX1 U14 ( .A(db_cnt[1]), .Y(n2) );
  INVX1 U15 ( .A(db_cnt[2]), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updprl_a0 ( r_spec, r_dat_spec, r_auto_txgdcrc, r_dat_portrole, 
        r_dat_datarole, r_auto_discard, r_set_cpmsgid, r_dat_cpmsgid, r_rdat, 
        r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact, ptx_fifopop, 
        prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, prx_rcvdords, prx_fifowdat, 
        pff_c0dat, prl_rdat, prl_txauto, prl_last, prl_txreq, prl_c0set, 
        prl_cany0, prl_cany0r, prl_cany0w, prl_idle, prl_discard, prl_GCTxDone, 
        prl_fsm, prl_cpmsgid, prl_cany0adr, clk, srstz );
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [2:0] r_dat_cpmsgid;
  input [7:0] r_rdat;
  input [2:0] prx_rcvdords;
  input [7:0] prx_fifowdat;
  input [47:0] pff_c0dat;
  output [7:0] prl_rdat;
  output [6:0] prl_txauto;
  output [3:0] prl_fsm;
  output [2:0] prl_cpmsgid;
  output [7:0] prl_cany0adr;
  input r_auto_txgdcrc, r_dat_portrole, r_dat_datarole, r_auto_discard,
         r_set_cpmsgid, r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact,
         ptx_fifopop, prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, clk, srstz;
  output prl_last, prl_txreq, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_idle, prl_discard, prl_GCTxDone;
  wire   sendgdcrc, stoptimer, N40, N41, c0_iop, N113, N114, N115, N116, N117,
         N118, N119, N120, N151, N152, N153, N154, N155, N156, N157, N158,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N189, N190,
         N191, N192, N193, N194, N196, N203, N204, N205, N206, net10379,
         net10385, net10390, net10395, net10400, n6, n8, n23, n26, n30, n37,
         n62, n77, n78, n79, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n99, n100, net147299, net147301, net147313, net147314, net147315,
         net147316, net147317, net147318, net147322, net147324, net147339,
         net147374, net147387, net160754, net166386, net166630, net166864,
         net167948, net168085, net168105, net169142, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n27, n28, n31,
         n32, n33, n34, n35, n36, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61,
         n63, n64, n65, n66, n67, n71, n72, n73, n74, n75, n76, n80, n81, n93,
         n94, n95, n96, n97, n98, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151;
  wire   [1:0] PrlTo;
  wire   [8:0] c0_cnt;
  wire   [7:0] txbuf;

  PrlTimer_1112a0 u0_PrlTimer ( .to(PrlTo), .restart(sendgdcrc), .stop(
        stoptimer), .clk(clk), .srstz(srstz) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_0 clk_gate_txbuf_reg ( .CLK(clk), .EN(N41), 
        .ENCLK(net10379), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_4 clk_gate_c0_adr_reg ( .CLK(clk), .EN(N194), 
        .ENCLK(net10385), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_3 clk_gate_cs_prcl_reg ( .CLK(clk), .EN(N189), 
        .ENCLK(net10390), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_2 clk_gate_c0_cnt_reg ( .CLK(clk), .EN(N196), 
        .ENCLK(net10395), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_1 clk_gate_CpMsgId_reg ( .CLK(clk), .EN(N203), 
        .ENCLK(net10400), .TE(1'b0) );
  updprl_a0_DW01_inc_0 r328 ( .A(prl_cany0adr), .SUM({N120, N119, N118, N117, 
        N116, N115, N114, N113}) );
  DFFQX1 c0_cnt_reg_3_ ( .D(N168), .C(net10395), .Q(c0_cnt[3]) );
  DFFQX1 c0_iop_reg ( .D(n99), .C(net10390), .Q(c0_iop) );
  DFFQX1 canyon_m0_reg ( .D(n100), .C(clk), .Q(prl_cany0) );
  DFFQX1 c0_adr_reg_1_ ( .D(N152), .C(net10385), .Q(prl_cany0adr[1]) );
  DFFQX1 c0_adr_reg_2_ ( .D(N153), .C(net10385), .Q(prl_cany0adr[2]) );
  DFFQX1 c0_adr_reg_3_ ( .D(N154), .C(net10385), .Q(prl_cany0adr[3]) );
  DFFQX1 c0_adr_reg_5_ ( .D(N156), .C(net10385), .Q(prl_cany0adr[5]) );
  DFFQX1 c0_adr_reg_6_ ( .D(N157), .C(net10385), .Q(prl_cany0adr[6]) );
  DFFQX1 c0_adr_reg_0_ ( .D(N151), .C(net10385), .Q(prl_cany0adr[0]) );
  DFFQX1 c0_adr_reg_7_ ( .D(N158), .C(net10385), .Q(prl_cany0adr[7]) );
  DFFQX1 txbuf_reg_7_ ( .D(r_rdat[7]), .C(net10379), .Q(txbuf[7]) );
  DFFQX1 txbuf_reg_4_ ( .D(r_rdat[4]), .C(net10379), .Q(txbuf[4]) );
  DFFQX1 txbuf_reg_3_ ( .D(r_rdat[3]), .C(net10379), .Q(txbuf[3]) );
  DFFQX1 c0_cnt_reg_8_ ( .D(N173), .C(net10395), .Q(c0_cnt[8]) );
  DFFQX1 c0_cnt_reg_4_ ( .D(N169), .C(net10395), .Q(c0_cnt[4]) );
  DFFQX1 c0_cnt_reg_5_ ( .D(N170), .C(net10395), .Q(c0_cnt[5]) );
  DFFQX1 c0_cnt_reg_6_ ( .D(N171), .C(net10395), .Q(c0_cnt[6]) );
  DFFQX1 c0_cnt_reg_7_ ( .D(N172), .C(net10395), .Q(c0_cnt[7]) );
  DFFQX1 CpMsgId_reg_1_ ( .D(N205), .C(net10400), .Q(prl_cpmsgid[1]) );
  DFFQX1 CpMsgId_reg_0_ ( .D(N204), .C(net10400), .Q(prl_cpmsgid[0]) );
  DFFQX1 CpMsgId_reg_2_ ( .D(N206), .C(net10400), .Q(prl_cpmsgid[2]) );
  DFFQXX2 cs_prcl_reg_3_ ( .D(N193), .C(net10390), .Q(prl_fsm[3]), .XQ(n54) );
  DFFQXX2 cs_prcl_reg_0_ ( .D(N190), .C(net10390), .Q(prl_fsm[0]), .XQ(
        net168085) );
  DFFQX2 c0_cnt_reg_0_ ( .D(N165), .C(net10395), .Q(c0_cnt[0]) );
  DFFQX2 cs_prcl_reg_1_ ( .D(N191), .C(net10390), .Q(prl_fsm[1]) );
  DFFQX2 c0_cnt_reg_1_ ( .D(N166), .C(net10395), .Q(n52) );
  DFFQX1 txbuf_reg_5_ ( .D(r_rdat[5]), .C(net10379), .Q(txbuf[5]) );
  DFFQX1 c0_cnt_reg_2_ ( .D(N167), .C(net10395), .Q(c0_cnt[2]) );
  DFFQX1 c0_adr_reg_4_ ( .D(N155), .C(net10385), .Q(prl_cany0adr[4]) );
  DFFQX1 txbuf_reg_2_ ( .D(r_rdat[2]), .C(net10379), .Q(txbuf[2]) );
  DFFQX1 txbuf_reg_1_ ( .D(r_rdat[1]), .C(net10379), .Q(txbuf[1]) );
  DFFQX1 txbuf_reg_0_ ( .D(r_rdat[0]), .C(net10379), .Q(txbuf[0]) );
  DFFQX1 txbuf_reg_6_ ( .D(r_rdat[6]), .C(net10379), .Q(txbuf[6]) );
  DFFQX2 cs_prcl_reg_2_ ( .D(N192), .C(net10390), .Q(prl_fsm[2]) );
  INVX1 U3 ( .A(1'b0), .Y(prl_txauto[3]) );
  INVX1 U5 ( .A(1'b0), .Y(prl_txauto[5]) );
  INVX1 U7 ( .A(1'b1), .Y(prl_txauto[6]) );
  NAND2X2 U9 ( .A(prl_fsm[1]), .B(net168085), .Y(net147314) );
  INVX3 U10 ( .A(prl_fsm[1]), .Y(net166630) );
  INVX2 U11 ( .A(n110), .Y(n108) );
  NAND21X2 U12 ( .B(c0_cnt[3]), .A(n105), .Y(n110) );
  NAND21X2 U13 ( .B(c0_cnt[4]), .A(n108), .Y(n113) );
  INVXL U14 ( .A(n141), .Y(n19) );
  NAND2XL U15 ( .A(prl_cpmsgid[2]), .B(n141), .Y(n10) );
  NAND32X2 U16 ( .B(net166630), .C(net147374), .A(net147316), .Y(n48) );
  INVX12 U17 ( .A(prl_fsm[2]), .Y(net147316) );
  NAND21X2 U18 ( .B(c0_cnt[6]), .A(n58), .Y(n118) );
  NOR21X2 U19 ( .B(n59), .A(n113), .Y(n58) );
  NOR2X2 U20 ( .A(c0_cnt[0]), .B(n52), .Y(n34) );
  AND2X2 U21 ( .A(n28), .B(net168105), .Y(n27) );
  NOR21X2 U22 ( .B(n51), .A(n118), .Y(net168105) );
  INVX1 U23 ( .A(r_dat_portrole), .Y(n55) );
  NAND2X2 U24 ( .A(n36), .B(n46), .Y(prl_cany0r) );
  INVX1 U25 ( .A(prx_rcvdords[0]), .Y(n142) );
  AND2X1 U26 ( .A(r_spec[1]), .B(r_spec[0]), .Y(n66) );
  INVX1 U27 ( .A(net147313), .Y(n44) );
  NAND21X1 U28 ( .B(prl_fsm[3]), .A(prl_fsm[0]), .Y(net147374) );
  INVX1 U29 ( .A(c0_cnt[5]), .Y(n59) );
  INVX1 U30 ( .A(c0_cnt[7]), .Y(n51) );
  INVX1 U31 ( .A(n107), .Y(n105) );
  NAND21X1 U32 ( .B(c0_cnt[2]), .A(n34), .Y(n107) );
  INVX1 U33 ( .A(ptx_txact), .Y(n40) );
  NAND21X1 U34 ( .B(net147315), .A(n42), .Y(n41) );
  NAND31X1 U35 ( .C(n39), .A(n45), .B(n25), .Y(n42) );
  INVX1 U36 ( .A(net147322), .Y(n39) );
  NAND21X1 U37 ( .B(n20), .A(n35), .Y(prl_txreq) );
  INVX1 U38 ( .A(n41), .Y(net147318) );
  NAND2XL U39 ( .A(txbuf[3]), .B(n145), .Y(n9) );
  NAND2X1 U40 ( .A(n9), .B(n10), .Y(prl_rdat[3]) );
  INVX1 U41 ( .A(n48), .Y(n141) );
  NAND2X1 U42 ( .A(txbuf[7]), .B(n145), .Y(n11) );
  NAND2X1 U43 ( .A(n146), .B(n56), .Y(n12) );
  NAND2X1 U44 ( .A(n11), .B(n12), .Y(prl_rdat[7]) );
  NAND2XL U45 ( .A(r_spec[1]), .B(n13), .Y(n14) );
  NAND2XL U46 ( .A(r_dat_spec[1]), .B(n66), .Y(n15) );
  NAND2X1 U47 ( .A(n14), .B(n15), .Y(n56) );
  INVXL U48 ( .A(n66), .Y(n13) );
  NAND2XL U49 ( .A(txbuf[5]), .B(n145), .Y(n16) );
  INVXL U50 ( .A(n144), .Y(n17) );
  NAND2X1 U51 ( .A(n16), .B(n17), .Y(prl_rdat[5]) );
  NOR5X1 U52 ( .A(n21), .B(prx_rcvdords[2]), .C(prx_rcvdords[1]), .D(
        r_dat_datarole), .E(n142), .Y(n144) );
  NAND2X1 U53 ( .A(n27), .B(net147299), .Y(n18) );
  NAND2X1 U54 ( .A(n18), .B(n19), .Y(prl_last) );
  INVXL U55 ( .A(n27), .Y(n43) );
  NAND32X2 U56 ( .B(prl_fsm[2]), .C(prl_fsm[0]), .A(n80), .Y(n137) );
  NOR2X1 U57 ( .A(n8), .B(n124), .Y(n20) );
  INVX1 U58 ( .A(c0_cnt[8]), .Y(n28) );
  INVX1 U59 ( .A(n22), .Y(n104) );
  NAND32X1 U60 ( .B(net147314), .C(prl_fsm[2]), .A(n54), .Y(n21) );
  NAND32X1 U61 ( .B(net147314), .C(prl_fsm[2]), .A(n54), .Y(n143) );
  BUFXL U62 ( .A(n34), .Y(n22) );
  NAND31X4 U63 ( .C(prl_txauto[4]), .A(ptx_fifopop), .B(n43), .Y(n46) );
  INVX1 U64 ( .A(prl_txauto[4]), .Y(net147299) );
  INVX1 U65 ( .A(n50), .Y(n24) );
  INVXL U66 ( .A(prl_cany0w), .Y(n25) );
  NAND21X1 U67 ( .B(n140), .A(txbuf[0]), .Y(n138) );
  INVX1 U68 ( .A(n33), .Y(n38) );
  BUFXL U69 ( .A(net147374), .Y(n31) );
  BUFXL U70 ( .A(n108), .Y(n32) );
  NAND31XL U71 ( .C(n31), .A(prl_fsm[1]), .B(prl_fsm[2]), .Y(net147313) );
  INVX3 U72 ( .A(n140), .Y(n145) );
  AOI21BBXL U73 ( .B(net169142), .C(n28), .A(n27), .Y(net160754) );
  BUFXL U74 ( .A(prx_fifopsh), .Y(n33) );
  OAI2B11X1 U75 ( .D(n55), .C(n48), .A(n138), .B(n21), .Y(prl_rdat[0]) );
  INVX3 U76 ( .A(net147301), .Y(prl_cany0w) );
  NAND21X2 U77 ( .B(net147324), .A(prx_fifopsh), .Y(net147301) );
  NAND2X2 U78 ( .A(prx_fifopsh), .B(n44), .Y(n36) );
  NAND21XL U79 ( .B(prl_txauto[4]), .A(ptx_fifopop), .Y(n45) );
  NAND21XL U80 ( .B(prl_txauto[4]), .A(n40), .Y(n35) );
  BUFXL U81 ( .A(net168105), .Y(net169142) );
  AO22X1 U82 ( .A(txbuf[1]), .B(n145), .C(prl_cpmsgid[0]), .D(n141), .Y(
        prl_rdat[1]) );
  INVXL U83 ( .A(n118), .Y(n116) );
  BUFXL U84 ( .A(n58), .Y(n47) );
  NAND32X1 U85 ( .B(prl_fsm[2]), .C(n54), .A(net166630), .Y(n98) );
  NAND32X1 U86 ( .B(net166630), .C(net147374), .A(net147316), .Y(n139) );
  NAND32XL U87 ( .B(n31), .C(net147316), .A(net166630), .Y(n132) );
  NAND2X2 U88 ( .A(n143), .B(n139), .Y(n140) );
  NAND21XL U89 ( .B(c0_cnt[4]), .A(n32), .Y(n49) );
  INVXL U90 ( .A(n49), .Y(n111) );
  AO22AX1 U91 ( .A(txbuf[6]), .B(n145), .C(n146), .D(n57), .Y(prl_rdat[6]) );
  INVX1 U92 ( .A(n21), .Y(n146) );
  BUFXL U93 ( .A(n105), .Y(n50) );
  INVXL U94 ( .A(n47), .Y(n115) );
  BUFXL U95 ( .A(net147314), .Y(net167948) );
  MUX2IXL U96 ( .D0(r_spec[0]), .D1(r_dat_spec[0]), .S(n66), .Y(n57) );
  AO22X1 U97 ( .A(txbuf[2]), .B(n145), .C(prl_cpmsgid[1]), .D(n141), .Y(
        prl_rdat[2]) );
  NAND32XL U98 ( .B(net167948), .C(net147316), .A(n54), .Y(n125) );
  INVXL U99 ( .A(n98), .Y(n60) );
  NAND21XL U100 ( .B(prl_fsm[0]), .A(n131), .Y(net147324) );
  INVXL U101 ( .A(n98), .Y(n131) );
  BUFX1 U102 ( .A(net147313), .Y(net166864) );
  BUFXL U103 ( .A(prl_cany0r), .Y(net166386) );
  OAI211XL U104 ( .C(n48), .D(n71), .A(n93), .B(n128), .Y(N192) );
  NAND21XL U105 ( .B(n131), .A(net147313), .Y(n134) );
  OR4X1 U106 ( .A(net147315), .B(n127), .C(n126), .D(n61), .Y(N189) );
  AOI21XL U107 ( .B(n125), .C(n132), .A(n38), .Y(n61) );
  OAI211XL U108 ( .C(net147315), .D(net166864), .A(n93), .B(n81), .Y(N190) );
  INVXL U109 ( .A(net147324), .Y(net147387) );
  AOI21AXL U110 ( .B(net166864), .C(n67), .A(net147339), .Y(N193) );
  NAND21XL U111 ( .B(net147313), .A(pid_ccidle), .Y(net147322) );
  INVX1 U112 ( .A(r_discard), .Y(n120) );
  NOR21XL U113 ( .B(prx_gdmsgrcvd), .A(r_set_cpmsgid), .Y(n37) );
  INVX1 U114 ( .A(n23), .Y(prl_c0set) );
  NAND32X1 U115 ( .B(r_set_cpmsgid), .C(prx_gdmsgrcvd), .A(srstz), .Y(N203) );
  NAND21X1 U116 ( .B(n132), .A(net147339), .Y(n128) );
  INVX1 U117 ( .A(srstz), .Y(n71) );
  INVX1 U118 ( .A(n125), .Y(n97) );
  INVX1 U119 ( .A(n132), .Y(n133) );
  INVX3 U120 ( .A(n137), .Y(prl_idle) );
  NAND6XL U121 ( .A(n79), .B(n83), .C(n78), .D(n77), .E(n135), .F(n72), .Y(n23) );
  NOR3XL U122 ( .A(pff_c0dat[42]), .B(pff_c0dat[44]), .C(pff_c0dat[43]), .Y(
        n83) );
  NOR5X1 U123 ( .A(pff_c0dat[47]), .B(pff_c0dat[45]), .C(pff_c0dat[36]), .D(
        pff_c0dat[34]), .E(n82), .Y(n72) );
  NOR4XL U124 ( .A(n84), .B(n85), .C(pff_c0dat[22]), .D(pff_c0dat[20]), .Y(n79) );
  NAND31X1 U125 ( .C(prl_discard), .A(n8), .B(n120), .Y(n6) );
  AO21XL U126 ( .B(ptx_fifopop), .C(n140), .A(n136), .Y(n127) );
  OAI221XL U127 ( .A(n148), .B(n124), .C(n123), .D(n137), .E(net147322), .Y(
        n126) );
  OAI211X1 U128 ( .C(n96), .D(n71), .A(n95), .B(n128), .Y(N191) );
  AOI31XL U129 ( .A(n119), .B(n120), .C(n20), .D(n146), .Y(n96) );
  OAI21BBX1 U130 ( .A(r_dat_cpmsgid[0]), .B(r_set_cpmsgid), .C(n63), .Y(N204)
         );
  AOI21X1 U131 ( .B(pff_c0dat[9]), .C(n37), .A(n71), .Y(n63) );
  OAI21BBX1 U132 ( .A(r_dat_cpmsgid[1]), .B(r_set_cpmsgid), .C(n64), .Y(N205)
         );
  AOI21X1 U133 ( .B(pff_c0dat[10]), .C(n37), .A(n71), .Y(n64) );
  OAI21BBX1 U134 ( .A(r_dat_cpmsgid[2]), .B(r_set_cpmsgid), .C(n65), .Y(N206)
         );
  AOI21X1 U135 ( .B(pff_c0dat[11]), .C(n37), .A(n71), .Y(n65) );
  INVX1 U136 ( .A(sendgdcrc), .Y(n123) );
  AO21XL U137 ( .B(n137), .C(n21), .A(n71), .Y(n81) );
  INVX1 U138 ( .A(n76), .Y(n93) );
  OAI31XL U139 ( .A(n121), .B(n71), .C(n135), .D(n95), .Y(n76) );
  INVX1 U140 ( .A(net147315), .Y(net147339) );
  AO22X1 U141 ( .A(N118), .B(n134), .C(prx_fifowdat[5]), .D(n133), .Y(N156) );
  AO22X1 U142 ( .A(N119), .B(n134), .C(prx_fifowdat[6]), .D(n133), .Y(N157) );
  AO22X1 U143 ( .A(N117), .B(n134), .C(n133), .D(prx_fifowdat[4]), .Y(N155) );
  INVX1 U144 ( .A(n122), .Y(n136) );
  NAND21X1 U145 ( .B(n121), .A(ptx_ack), .Y(n122) );
  AND2X1 U146 ( .A(n136), .B(n135), .Y(prl_GCTxDone) );
  INVX1 U147 ( .A(n119), .Y(prl_discard) );
  AO22X1 U148 ( .A(N116), .B(n134), .C(n133), .D(prx_fifowdat[3]), .Y(N154) );
  NAND2XL U149 ( .A(prl_fsm[0]), .B(n60), .Y(prl_txauto[4]) );
  AND2XL U150 ( .A(txbuf[4]), .B(n145), .Y(prl_rdat[4]) );
  NAND42X1 U151 ( .C(pff_c0dat[14]), .D(pff_c0dat[13]), .A(prx_gdmsgrcvd), .B(
        n89), .Y(n87) );
  NOR3XL U152 ( .A(pff_c0dat[15]), .B(pff_c0dat[18]), .C(pff_c0dat[16]), .Y(
        n89) );
  NOR42XL U153 ( .C(pff_c0dat[24]), .D(pff_c0dat[21]), .A(n87), .B(n88), .Y(
        n78) );
  NAND3X1 U154 ( .A(pff_c0dat[17]), .B(pff_c0dat[12]), .C(pff_c0dat[19]), .Y(
        n88) );
  OAI21BX1 U155 ( .C(PrlTo[0]), .B(r_auto_discard), .A(n148), .Y(stoptimer) );
  INVX1 U156 ( .A(n6), .Y(n148) );
  NAND21X1 U157 ( .B(r_rdy), .A(net147317), .Y(N41) );
  AO21X1 U158 ( .B(prx_gdmsgrcvd), .C(r_auto_txgdcrc), .A(prl_c0set), .Y(
        sendgdcrc) );
  NAND42X1 U159 ( .C(prx_fifowdat[0]), .D(net147315), .A(n30), .B(n97), .Y(n95) );
  NAND32X1 U160 ( .B(n74), .C(n71), .A(n73), .Y(net147315) );
  OA21X1 U161 ( .B(prx_eoprcvd), .C(pid_ccidle), .A(net147387), .Y(n74) );
  OA21X1 U162 ( .B(prl_cany0), .C(prl_c0set), .A(net147339), .Y(n100) );
  ENOX1 U163 ( .A(n26), .B(n151), .C(n26), .D(c0_iop), .Y(n99) );
  INVX1 U164 ( .A(prx_fifowdat[1]), .Y(n151) );
  NAND43X1 U165 ( .B(net167948), .C(net147315), .D(net147316), .A(n30), .Y(n26) );
  NAND3X1 U166 ( .A(n30), .B(prx_fifowdat[0]), .C(n97), .Y(n67) );
  INVX1 U167 ( .A(c0_iop), .Y(n130) );
  INVX1 U168 ( .A(n128), .Y(n129) );
  NAND32X1 U169 ( .B(pff_c0dat[28]), .C(pff_c0dat[27]), .A(n86), .Y(n84) );
  NOR3XL U170 ( .A(pff_c0dat[29]), .B(pff_c0dat[32]), .C(pff_c0dat[31]), .Y(
        n86) );
  AND2X1 U171 ( .A(pff_c0dat[33]), .B(pff_c0dat[30]), .Y(n92) );
  OR3XL U172 ( .A(pff_c0dat[26]), .B(pff_c0dat[25]), .C(pff_c0dat[23]), .Y(n85) );
  OR3XL U173 ( .A(pff_c0dat[41]), .B(pff_c0dat[39]), .C(pff_c0dat[38]), .Y(n82) );
  NOR42XL U174 ( .C(pff_c0dat[3]), .D(pff_c0dat[2]), .A(n90), .B(n91), .Y(n77)
         );
  NAND3X1 U175 ( .A(pff_c0dat[0]), .B(pff_c0dat[46]), .C(pff_c0dat[1]), .Y(n91) );
  NAND4X1 U176 ( .A(pff_c0dat[40]), .B(pff_c0dat[37]), .C(n92), .D(
        pff_c0dat[35]), .Y(n90) );
  NOR43XL U177 ( .B(n150), .C(n149), .D(n62), .A(prx_fifowdat[2]), .Y(n30) );
  INVX1 U178 ( .A(prx_fifowdat[3]), .Y(n150) );
  INVX1 U179 ( .A(prx_fifowdat[4]), .Y(n149) );
  NOR3XL U180 ( .A(prx_fifowdat[5]), .B(prx_fifowdat[7]), .C(prx_fifowdat[6]), 
        .Y(n62) );
  INVX1 U181 ( .A(prl_cany0), .Y(n135) );
  GEN2XL U182 ( .D(c0_cnt[7]), .E(n118), .C(net169142), .B(n131), .A(n117), 
        .Y(N172) );
  NOR21XL U183 ( .B(prx_fifowdat[7]), .A(net166864), .Y(n117) );
  GEN2XL U184 ( .D(c0_cnt[5]), .E(n49), .C(n47), .B(n131), .A(n112), .Y(N170)
         );
  NOR21XL U185 ( .B(prx_fifowdat[5]), .A(net166864), .Y(n112) );
  AO22X1 U186 ( .A(N120), .B(n134), .C(prx_fifowdat[7]), .D(n133), .Y(N158) );
  GEN2XL U187 ( .D(c0_cnt[6]), .E(n115), .C(n116), .B(n131), .A(n114), .Y(N171) );
  NOR21XL U188 ( .B(prx_fifowdat[6]), .A(net166864), .Y(n114) );
  GEN2XL U189 ( .D(c0_cnt[4]), .E(n110), .C(n111), .B(n131), .A(n109), .Y(N169) );
  NOR21XL U190 ( .B(prx_fifowdat[4]), .A(net166864), .Y(n109) );
  NAND2X1 U191 ( .A(pid_ccidle), .B(PrlTo[0]), .Y(n8) );
  NAND32XL U192 ( .B(prl_fsm[2]), .C(n31), .A(net166630), .Y(n124) );
  NAND32X1 U193 ( .B(n94), .C(n124), .A(PrlTo[1]), .Y(n119) );
  INVX1 U194 ( .A(r_auto_discard), .Y(n94) );
  NOR21XL U195 ( .B(n131), .A(net160754), .Y(N173) );
  GEN2XL U196 ( .D(n52), .E(c0_cnt[0]), .C(n22), .B(n131), .A(n102), .Y(N166)
         );
  NOR21XL U197 ( .B(prx_fifowdat[1]), .A(net147313), .Y(n102) );
  GEN2XL U198 ( .D(c0_cnt[2]), .E(n104), .C(n50), .B(n131), .A(n103), .Y(N167)
         );
  NOR21XL U199 ( .B(prx_fifowdat[2]), .A(net166864), .Y(n103) );
  GEN2XL U200 ( .D(c0_cnt[3]), .E(n24), .C(n32), .B(n131), .A(n106), .Y(N168)
         );
  NOR21XL U201 ( .B(prx_fifowdat[3]), .A(net166864), .Y(n106) );
  AO22X1 U202 ( .A(N115), .B(n134), .C(prx_fifowdat[2]), .D(n133), .Y(N153) );
  AO22X1 U203 ( .A(N113), .B(n134), .C(prx_fifowdat[0]), .D(n133), .Y(N151) );
  AO22X1 U204 ( .A(N114), .B(n134), .C(n133), .D(prx_fifowdat[1]), .Y(N152) );
  OAI22XL U205 ( .A(n101), .B(net166864), .C(c0_cnt[0]), .D(n98), .Y(N165) );
  INVX1 U206 ( .A(prx_fifowdat[0]), .Y(n101) );
  BUFXL U207 ( .A(prx_rcvdords[2]), .Y(prl_txauto[2]) );
  BUFXL U208 ( .A(prx_rcvdords[1]), .Y(prl_txauto[1]) );
  BUFXL U209 ( .A(prx_rcvdords[0]), .Y(prl_txauto[0]) );
  AND2XL U210 ( .A(net147339), .B(net166386), .Y(N196) );
  INVXL U211 ( .A(net166386), .Y(net147317) );
  NAND21X2 U212 ( .B(prl_fsm[3]), .A(net166630), .Y(n75) );
  INVX3 U213 ( .A(n75), .Y(n80) );
  NAND32XL U214 ( .B(prl_fsm[0]), .C(net147316), .A(n80), .Y(n121) );
  AO22XL U215 ( .A(net147318), .B(n130), .C(n129), .D(n33), .Y(N194) );
  AOI32XL U216 ( .A(N40), .B(n33), .C(n97), .D(ptx_ack), .E(net147299), .Y(n73) );
  NOR3XL U217 ( .A(prx_fifowdat[5]), .B(prx_fifowdat[7]), .C(prx_fifowdat[6]), 
        .Y(n147) );
  NAND43X1 U218 ( .B(prx_fifowdat[4]), .C(prx_fifowdat[3]), .D(prx_fifowdat[2]), .A(n147), .Y(N40) );
endmodule


module updprl_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module PrlTimer_1112a0 ( to, restart, stop, clk, srstz );
  output [1:0] to;
  input restart, stop, clk, srstz;
  wire   ena, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, net10417, n12,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [11:0] timer;

  SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 clk_gate_timer_reg ( .CLK(clk), .EN(N18), .ENCLK(net10417), .TE(1'b0) );
  PrlTimer_1112a0_DW01_inc_0 add_25 ( .A(timer), .SUM({N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}) );
  DFFQX1 ena_reg ( .D(n12), .C(clk), .Q(ena) );
  DFFQX1 timer_reg_1_ ( .D(N20), .C(net10417), .Q(timer[1]) );
  DFFQX1 timer_reg_2_ ( .D(N21), .C(net10417), .Q(timer[2]) );
  DFFQX1 timer_reg_0_ ( .D(N19), .C(net10417), .Q(timer[0]) );
  DFFQX1 timer_reg_11_ ( .D(N30), .C(net10417), .Q(timer[11]) );
  DFFQX1 timer_reg_9_ ( .D(N28), .C(net10417), .Q(timer[9]) );
  DFFQX1 timer_reg_10_ ( .D(N29), .C(net10417), .Q(timer[10]) );
  DFFQX1 timer_reg_5_ ( .D(N24), .C(net10417), .Q(timer[5]) );
  DFFQX1 timer_reg_6_ ( .D(N25), .C(net10417), .Q(timer[6]) );
  DFFQX1 timer_reg_7_ ( .D(N26), .C(net10417), .Q(timer[7]) );
  DFFQX1 timer_reg_8_ ( .D(N27), .C(net10417), .Q(timer[8]) );
  DFFQX1 timer_reg_4_ ( .D(N23), .C(net10417), .Q(timer[4]) );
  DFFQX1 timer_reg_3_ ( .D(N22), .C(net10417), .Q(timer[3]) );
  BUFX3 U3 ( .A(n8), .Y(n1) );
  NAND3X1 U4 ( .A(srstz), .B(ena), .C(n9), .Y(n8) );
  INVX1 U5 ( .A(n2), .Y(to[0]) );
  AOI211X1 U6 ( .C(n3), .D(timer[9]), .A(timer[10]), .B(timer[11]), .Y(n2) );
  INVX1 U7 ( .A(n4), .Y(n3) );
  AOI211X1 U8 ( .C(timer[6]), .D(n5), .A(timer[8]), .B(timer[7]), .Y(n4) );
  AO21X1 U9 ( .B(timer[4]), .C(timer[3]), .A(timer[5]), .Y(n5) );
  INVX1 U10 ( .A(n6), .Y(n12) );
  AOI31X1 U11 ( .A(srstz), .B(n7), .C(ena), .D(restart), .Y(n6) );
  INVX1 U12 ( .A(stop), .Y(n7) );
  NOR21XL U13 ( .B(N15), .A(n1), .Y(N30) );
  NOR21XL U14 ( .B(N14), .A(n1), .Y(N29) );
  NOR21XL U15 ( .B(N13), .A(n1), .Y(N28) );
  NOR21XL U16 ( .B(N12), .A(n1), .Y(N27) );
  NOR21XL U17 ( .B(N11), .A(n8), .Y(N26) );
  NOR21XL U18 ( .B(N10), .A(n8), .Y(N25) );
  NOR21XL U19 ( .B(N9), .A(n8), .Y(N24) );
  NOR21XL U20 ( .B(N8), .A(n8), .Y(N23) );
  NOR21XL U21 ( .B(N7), .A(n8), .Y(N22) );
  NOR21XL U22 ( .B(N6), .A(n8), .Y(N21) );
  NOR21XL U23 ( .B(N5), .A(n8), .Y(N20) );
  NOR21XL U24 ( .B(N4), .A(n8), .Y(N19) );
  NAND31X1 U25 ( .C(restart), .A(n8), .B(srstz), .Y(N18) );
  NOR3XL U26 ( .A(to[1]), .B(stop), .C(restart), .Y(n9) );
  INVX1 U27 ( .A(n10), .Y(to[1]) );
  OAI31XL U28 ( .A(timer[10]), .B(timer[9]), .C(timer[8]), .D(timer[11]), .Y(
        n10) );
endmodule


module PrlTimer_1112a0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyff_DEPTH_NUM34_DEPTH_NBT6 ( r_psh, r_pop, prx_psh, ptx_pop, r_last, 
        r_unlock, i_lockena, r_fiforst, i_ccidle, r_wdat, prx_wdat, txreq, 
        ffack, rdat0, full, empty, one, half, obsd, dat_7_1, ptr, fifowdat, 
        fifopsh, clk, srstz );
  input [7:0] r_wdat;
  input [7:0] prx_wdat;
  output [1:0] ffack;
  output [7:0] rdat0;
  output [55:0] dat_7_1;
  output [5:0] ptr;
  output [7:0] fifowdat;
  input r_psh, r_pop, prx_psh, ptx_pop, r_last, r_unlock, i_lockena, r_fiforst,
         i_ccidle, clk, srstz;
  output txreq, full, empty, one, half, obsd, fifopsh;
  wire   ps_locked, locked, mem_8__7_, mem_8__6_, mem_8__5_, mem_8__4_,
         mem_8__3_, mem_8__2_, mem_8__1_, mem_8__0_, mem_9__7_, mem_9__6_,
         mem_9__5_, mem_9__4_, mem_9__3_, mem_9__2_, mem_9__1_, mem_9__0_,
         mem_10__7_, mem_10__6_, mem_10__5_, mem_10__4_, mem_10__3_,
         mem_10__2_, mem_10__1_, mem_10__0_, mem_11__7_, mem_11__6_,
         mem_11__5_, mem_11__4_, mem_11__3_, mem_11__2_, mem_11__1_,
         mem_11__0_, mem_12__7_, mem_12__6_, mem_12__5_, mem_12__4_,
         mem_12__3_, mem_12__2_, mem_12__1_, mem_12__0_, mem_13__7_,
         mem_13__6_, mem_13__5_, mem_13__4_, mem_13__3_, mem_13__2_,
         mem_13__1_, mem_13__0_, mem_14__7_, mem_14__6_, mem_14__5_,
         mem_14__4_, mem_14__3_, mem_14__2_, mem_14__1_, mem_14__0_,
         mem_15__7_, mem_15__6_, mem_15__5_, mem_15__4_, mem_15__3_,
         mem_15__2_, mem_15__1_, mem_15__0_, mem_16__7_, mem_16__6_,
         mem_16__5_, mem_16__4_, mem_16__3_, mem_16__2_, mem_16__1_,
         mem_16__0_, mem_17__7_, mem_17__6_, mem_17__5_, mem_17__4_,
         mem_17__3_, mem_17__2_, mem_17__1_, mem_17__0_, mem_18__7_,
         mem_18__6_, mem_18__5_, mem_18__4_, mem_18__3_, mem_18__2_,
         mem_18__1_, mem_18__0_, mem_19__7_, mem_19__6_, mem_19__5_,
         mem_19__4_, mem_19__3_, mem_19__2_, mem_19__1_, mem_19__0_,
         mem_20__7_, mem_20__6_, mem_20__5_, mem_20__4_, mem_20__3_,
         mem_20__2_, mem_20__1_, mem_20__0_, mem_21__7_, mem_21__6_,
         mem_21__5_, mem_21__4_, mem_21__3_, mem_21__2_, mem_21__1_,
         mem_21__0_, mem_22__7_, mem_22__6_, mem_22__5_, mem_22__4_,
         mem_22__3_, mem_22__2_, mem_22__1_, mem_22__0_, mem_23__7_,
         mem_23__6_, mem_23__5_, mem_23__4_, mem_23__3_, mem_23__2_,
         mem_23__1_, mem_23__0_, mem_24__7_, mem_24__6_, mem_24__5_,
         mem_24__4_, mem_24__3_, mem_24__2_, mem_24__1_, mem_24__0_,
         mem_25__7_, mem_25__6_, mem_25__5_, mem_25__4_, mem_25__3_,
         mem_25__2_, mem_25__1_, mem_25__0_, mem_26__7_, mem_26__6_,
         mem_26__5_, mem_26__4_, mem_26__3_, mem_26__2_, mem_26__1_,
         mem_26__0_, mem_27__7_, mem_27__6_, mem_27__5_, mem_27__4_,
         mem_27__3_, mem_27__2_, mem_27__1_, mem_27__0_, mem_28__7_,
         mem_28__6_, mem_28__5_, mem_28__4_, mem_28__3_, mem_28__2_,
         mem_28__1_, mem_28__0_, mem_29__7_, mem_29__6_, mem_29__5_,
         mem_29__4_, mem_29__3_, mem_29__2_, mem_29__1_, mem_29__0_,
         mem_30__7_, mem_30__6_, mem_30__5_, mem_30__4_, mem_30__3_,
         mem_30__2_, mem_30__1_, mem_30__0_, mem_31__7_, mem_31__6_,
         mem_31__5_, mem_31__4_, mem_31__3_, mem_31__2_, mem_31__1_,
         mem_31__0_, mem_32__7_, mem_32__6_, mem_32__5_, mem_32__4_,
         mem_32__3_, mem_32__2_, mem_32__1_, mem_32__0_, mem_33__7_,
         mem_33__6_, mem_33__5_, mem_33__4_, mem_33__3_, mem_33__2_,
         mem_33__1_, mem_33__0_, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1053, N1054, N1055,
         N1056, N1057, N1058, N1059, net10435, net10441, net10446, net10451,
         net10456, net10461, net10466, net10471, net10476, net10481, net10486,
         net10491, net10496, net10501, net10506, net10511, net10516, net10521,
         net10526, net10531, net10536, net10541, net10546, net10551, net10556,
         net10561, net10566, net10571, net10576, net10581, net10586, net10591,
         net10596, net10601, net10606, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n43, n44, n45, n47, n48, n49, n51, n52, n53, n55, n56, n57,
         n59, n60, n61, n63, n64, n65, n67, n68, n69, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639;

  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 clk_gate_mem_reg_0_ ( 
        .CLK(clk), .EN(N1022), .ENCLK(net10435), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 clk_gate_mem_reg_1_ ( 
        .CLK(clk), .EN(N1013), .ENCLK(net10441), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 clk_gate_mem_reg_2_ ( 
        .CLK(clk), .EN(N1004), .ENCLK(net10446), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 clk_gate_mem_reg_3_ ( 
        .CLK(clk), .EN(N995), .ENCLK(net10451), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 clk_gate_mem_reg_4_ ( 
        .CLK(clk), .EN(N986), .ENCLK(net10456), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 clk_gate_mem_reg_5_ ( 
        .CLK(clk), .EN(N977), .ENCLK(net10461), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 clk_gate_mem_reg_6_ ( 
        .CLK(clk), .EN(N968), .ENCLK(net10466), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 clk_gate_mem_reg_7_ ( 
        .CLK(clk), .EN(N959), .ENCLK(net10471), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 clk_gate_mem_reg_8_ ( 
        .CLK(clk), .EN(N950), .ENCLK(net10476), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 clk_gate_mem_reg_9_ ( 
        .CLK(clk), .EN(N941), .ENCLK(net10481), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 clk_gate_mem_reg_10_ ( 
        .CLK(clk), .EN(N932), .ENCLK(net10486), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 clk_gate_mem_reg_11_ ( 
        .CLK(clk), .EN(N923), .ENCLK(net10491), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 clk_gate_mem_reg_12_ ( 
        .CLK(clk), .EN(N914), .ENCLK(net10496), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 clk_gate_mem_reg_13_ ( 
        .CLK(clk), .EN(N905), .ENCLK(net10501), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 clk_gate_mem_reg_14_ ( 
        .CLK(clk), .EN(N896), .ENCLK(net10506), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 clk_gate_mem_reg_15_ ( 
        .CLK(clk), .EN(N887), .ENCLK(net10511), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 clk_gate_mem_reg_16_ ( 
        .CLK(clk), .EN(N878), .ENCLK(net10516), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 clk_gate_mem_reg_17_ ( 
        .CLK(clk), .EN(N869), .ENCLK(net10521), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 clk_gate_mem_reg_18_ ( 
        .CLK(clk), .EN(N860), .ENCLK(net10526), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 clk_gate_mem_reg_19_ ( 
        .CLK(clk), .EN(N851), .ENCLK(net10531), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 clk_gate_mem_reg_20_ ( 
        .CLK(clk), .EN(N842), .ENCLK(net10536), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 clk_gate_mem_reg_21_ ( 
        .CLK(clk), .EN(N833), .ENCLK(net10541), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 clk_gate_mem_reg_22_ ( 
        .CLK(clk), .EN(N824), .ENCLK(net10546), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 clk_gate_mem_reg_23_ ( 
        .CLK(clk), .EN(N815), .ENCLK(net10551), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 clk_gate_mem_reg_24_ ( 
        .CLK(clk), .EN(N806), .ENCLK(net10556), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 clk_gate_mem_reg_25_ ( 
        .CLK(clk), .EN(N797), .ENCLK(net10561), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 clk_gate_mem_reg_26_ ( 
        .CLK(clk), .EN(N788), .ENCLK(net10566), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 clk_gate_mem_reg_27_ ( 
        .CLK(clk), .EN(N779), .ENCLK(net10571), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 clk_gate_mem_reg_28_ ( 
        .CLK(clk), .EN(N770), .ENCLK(net10576), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 clk_gate_mem_reg_29_ ( 
        .CLK(clk), .EN(N761), .ENCLK(net10581), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 clk_gate_mem_reg_30_ ( 
        .CLK(clk), .EN(N752), .ENCLK(net10586), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 clk_gate_mem_reg_31_ ( 
        .CLK(clk), .EN(N743), .ENCLK(net10591), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 clk_gate_mem_reg_32_ ( 
        .CLK(clk), .EN(N734), .ENCLK(net10596), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 clk_gate_mem_reg_33_ ( 
        .CLK(clk), .EN(N733), .ENCLK(net10601), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 clk_gate_pshptr_reg ( 
        .CLK(clk), .EN(N1053), .ENCLK(net10606), .TE(1'b0) );
  DFFQX1 mem_reg_33__7_ ( .D(fifowdat[7]), .C(net10601), .Q(mem_33__7_) );
  DFFQX1 mem_reg_32__7_ ( .D(N742), .C(net10596), .Q(mem_32__7_) );
  DFFQX1 mem_reg_31__7_ ( .D(N751), .C(net10591), .Q(mem_31__7_) );
  DFFQX1 mem_reg_30__7_ ( .D(N760), .C(net10586), .Q(mem_30__7_) );
  DFFQX1 mem_reg_29__7_ ( .D(N769), .C(net10581), .Q(mem_29__7_) );
  DFFQX1 mem_reg_28__7_ ( .D(N778), .C(net10576), .Q(mem_28__7_) );
  DFFQX1 mem_reg_33__6_ ( .D(fifowdat[6]), .C(net10601), .Q(mem_33__6_) );
  DFFQX1 mem_reg_32__6_ ( .D(N741), .C(net10596), .Q(mem_32__6_) );
  DFFQX1 mem_reg_31__6_ ( .D(N750), .C(net10591), .Q(mem_31__6_) );
  DFFQX1 mem_reg_30__6_ ( .D(N759), .C(net10586), .Q(mem_30__6_) );
  DFFQX1 mem_reg_29__6_ ( .D(N768), .C(net10581), .Q(mem_29__6_) );
  DFFQX1 mem_reg_28__6_ ( .D(N777), .C(net10576), .Q(mem_28__6_) );
  DFFQX1 mem_reg_33__5_ ( .D(fifowdat[5]), .C(net10601), .Q(mem_33__5_) );
  DFFQX1 mem_reg_32__5_ ( .D(N740), .C(net10596), .Q(mem_32__5_) );
  DFFQX1 mem_reg_31__5_ ( .D(N749), .C(net10591), .Q(mem_31__5_) );
  DFFQX1 mem_reg_30__5_ ( .D(N758), .C(net10586), .Q(mem_30__5_) );
  DFFQX1 mem_reg_29__5_ ( .D(N767), .C(net10581), .Q(mem_29__5_) );
  DFFQX1 mem_reg_28__5_ ( .D(N776), .C(net10576), .Q(mem_28__5_) );
  DFFQX1 mem_reg_33__4_ ( .D(fifowdat[4]), .C(net10601), .Q(mem_33__4_) );
  DFFQX1 mem_reg_32__4_ ( .D(N739), .C(net10596), .Q(mem_32__4_) );
  DFFQX1 mem_reg_31__4_ ( .D(N748), .C(net10591), .Q(mem_31__4_) );
  DFFQX1 mem_reg_30__4_ ( .D(N757), .C(net10586), .Q(mem_30__4_) );
  DFFQX1 mem_reg_29__4_ ( .D(N766), .C(net10581), .Q(mem_29__4_) );
  DFFQX1 mem_reg_28__4_ ( .D(N775), .C(net10576), .Q(mem_28__4_) );
  DFFQX1 mem_reg_33__3_ ( .D(fifowdat[3]), .C(net10601), .Q(mem_33__3_) );
  DFFQX1 mem_reg_32__3_ ( .D(N738), .C(net10596), .Q(mem_32__3_) );
  DFFQX1 mem_reg_31__3_ ( .D(N747), .C(net10591), .Q(mem_31__3_) );
  DFFQX1 mem_reg_30__3_ ( .D(N756), .C(net10586), .Q(mem_30__3_) );
  DFFQX1 mem_reg_29__3_ ( .D(N765), .C(net10581), .Q(mem_29__3_) );
  DFFQX1 mem_reg_28__3_ ( .D(N774), .C(net10576), .Q(mem_28__3_) );
  DFFQX1 mem_reg_33__2_ ( .D(fifowdat[2]), .C(net10601), .Q(mem_33__2_) );
  DFFQX1 mem_reg_32__2_ ( .D(N737), .C(net10596), .Q(mem_32__2_) );
  DFFQX1 mem_reg_31__2_ ( .D(N746), .C(net10591), .Q(mem_31__2_) );
  DFFQX1 mem_reg_30__2_ ( .D(N755), .C(net10586), .Q(mem_30__2_) );
  DFFQX1 mem_reg_29__2_ ( .D(N764), .C(net10581), .Q(mem_29__2_) );
  DFFQX1 mem_reg_28__2_ ( .D(N773), .C(net10576), .Q(mem_28__2_) );
  DFFQX1 mem_reg_33__1_ ( .D(fifowdat[1]), .C(net10601), .Q(mem_33__1_) );
  DFFQX1 mem_reg_32__1_ ( .D(N736), .C(net10596), .Q(mem_32__1_) );
  DFFQX1 mem_reg_31__1_ ( .D(N745), .C(net10591), .Q(mem_31__1_) );
  DFFQX1 mem_reg_30__1_ ( .D(N754), .C(net10586), .Q(mem_30__1_) );
  DFFQX1 mem_reg_29__1_ ( .D(N763), .C(net10581), .Q(mem_29__1_) );
  DFFQX1 mem_reg_28__1_ ( .D(N772), .C(net10576), .Q(mem_28__1_) );
  DFFQX1 mem_reg_33__0_ ( .D(fifowdat[0]), .C(net10601), .Q(mem_33__0_) );
  DFFQX1 mem_reg_32__0_ ( .D(N735), .C(net10596), .Q(mem_32__0_) );
  DFFQX1 mem_reg_31__0_ ( .D(N744), .C(net10591), .Q(mem_31__0_) );
  DFFQX1 mem_reg_30__0_ ( .D(N753), .C(net10586), .Q(mem_30__0_) );
  DFFQX1 mem_reg_29__0_ ( .D(N762), .C(net10581), .Q(mem_29__0_) );
  DFFQX1 mem_reg_28__0_ ( .D(N771), .C(net10576), .Q(mem_28__0_) );
  DFFQX1 mem_reg_27__7_ ( .D(N787), .C(net10571), .Q(mem_27__7_) );
  DFFQX1 mem_reg_26__7_ ( .D(N796), .C(net10566), .Q(mem_26__7_) );
  DFFQX1 mem_reg_25__7_ ( .D(N805), .C(net10561), .Q(mem_25__7_) );
  DFFQX1 mem_reg_24__7_ ( .D(N814), .C(net10556), .Q(mem_24__7_) );
  DFFQX1 mem_reg_23__7_ ( .D(N823), .C(net10551), .Q(mem_23__7_) );
  DFFQX1 mem_reg_22__7_ ( .D(N832), .C(net10546), .Q(mem_22__7_) );
  DFFQX1 mem_reg_21__7_ ( .D(N841), .C(net10541), .Q(mem_21__7_) );
  DFFQX1 mem_reg_20__7_ ( .D(N850), .C(net10536), .Q(mem_20__7_) );
  DFFQX1 mem_reg_19__7_ ( .D(N859), .C(net10531), .Q(mem_19__7_) );
  DFFQX1 mem_reg_18__7_ ( .D(N868), .C(net10526), .Q(mem_18__7_) );
  DFFQX1 mem_reg_17__7_ ( .D(N877), .C(net10521), .Q(mem_17__7_) );
  DFFQX1 mem_reg_16__7_ ( .D(N886), .C(net10516), .Q(mem_16__7_) );
  DFFQX1 mem_reg_15__7_ ( .D(N895), .C(net10511), .Q(mem_15__7_) );
  DFFQX1 mem_reg_14__7_ ( .D(N904), .C(net10506), .Q(mem_14__7_) );
  DFFQX1 mem_reg_13__7_ ( .D(N913), .C(net10501), .Q(mem_13__7_) );
  DFFQX1 mem_reg_12__7_ ( .D(N922), .C(net10496), .Q(mem_12__7_) );
  DFFQX1 mem_reg_11__7_ ( .D(N931), .C(net10491), .Q(mem_11__7_) );
  DFFQX1 mem_reg_10__7_ ( .D(N940), .C(net10486), .Q(mem_10__7_) );
  DFFQX1 mem_reg_9__7_ ( .D(N949), .C(net10481), .Q(mem_9__7_) );
  DFFQX1 mem_reg_8__7_ ( .D(N958), .C(net10476), .Q(mem_8__7_) );
  DFFQX1 mem_reg_27__6_ ( .D(N786), .C(net10571), .Q(mem_27__6_) );
  DFFQX1 mem_reg_26__6_ ( .D(N795), .C(net10566), .Q(mem_26__6_) );
  DFFQX1 mem_reg_25__6_ ( .D(N804), .C(net10561), .Q(mem_25__6_) );
  DFFQX1 mem_reg_24__6_ ( .D(N813), .C(net10556), .Q(mem_24__6_) );
  DFFQX1 mem_reg_23__6_ ( .D(N822), .C(net10551), .Q(mem_23__6_) );
  DFFQX1 mem_reg_22__6_ ( .D(N831), .C(net10546), .Q(mem_22__6_) );
  DFFQX1 mem_reg_21__6_ ( .D(N840), .C(net10541), .Q(mem_21__6_) );
  DFFQX1 mem_reg_20__6_ ( .D(N849), .C(net10536), .Q(mem_20__6_) );
  DFFQX1 mem_reg_19__6_ ( .D(N858), .C(net10531), .Q(mem_19__6_) );
  DFFQX1 mem_reg_18__6_ ( .D(N867), .C(net10526), .Q(mem_18__6_) );
  DFFQX1 mem_reg_17__6_ ( .D(N876), .C(net10521), .Q(mem_17__6_) );
  DFFQX1 mem_reg_16__6_ ( .D(N885), .C(net10516), .Q(mem_16__6_) );
  DFFQX1 mem_reg_15__6_ ( .D(N894), .C(net10511), .Q(mem_15__6_) );
  DFFQX1 mem_reg_14__6_ ( .D(N903), .C(net10506), .Q(mem_14__6_) );
  DFFQX1 mem_reg_13__6_ ( .D(N912), .C(net10501), .Q(mem_13__6_) );
  DFFQX1 mem_reg_12__6_ ( .D(N921), .C(net10496), .Q(mem_12__6_) );
  DFFQX1 mem_reg_11__6_ ( .D(N930), .C(net10491), .Q(mem_11__6_) );
  DFFQX1 mem_reg_10__6_ ( .D(N939), .C(net10486), .Q(mem_10__6_) );
  DFFQX1 mem_reg_9__6_ ( .D(N948), .C(net10481), .Q(mem_9__6_) );
  DFFQX1 mem_reg_8__6_ ( .D(N957), .C(net10476), .Q(mem_8__6_) );
  DFFQX1 mem_reg_27__5_ ( .D(N785), .C(net10571), .Q(mem_27__5_) );
  DFFQX1 mem_reg_26__5_ ( .D(N794), .C(net10566), .Q(mem_26__5_) );
  DFFQX1 mem_reg_25__5_ ( .D(N803), .C(net10561), .Q(mem_25__5_) );
  DFFQX1 mem_reg_24__5_ ( .D(N812), .C(net10556), .Q(mem_24__5_) );
  DFFQX1 mem_reg_23__5_ ( .D(N821), .C(net10551), .Q(mem_23__5_) );
  DFFQX1 mem_reg_22__5_ ( .D(N830), .C(net10546), .Q(mem_22__5_) );
  DFFQX1 mem_reg_21__5_ ( .D(N839), .C(net10541), .Q(mem_21__5_) );
  DFFQX1 mem_reg_20__5_ ( .D(N848), .C(net10536), .Q(mem_20__5_) );
  DFFQX1 mem_reg_19__5_ ( .D(N857), .C(net10531), .Q(mem_19__5_) );
  DFFQX1 mem_reg_18__5_ ( .D(N866), .C(net10526), .Q(mem_18__5_) );
  DFFQX1 mem_reg_17__5_ ( .D(N875), .C(net10521), .Q(mem_17__5_) );
  DFFQX1 mem_reg_16__5_ ( .D(N884), .C(net10516), .Q(mem_16__5_) );
  DFFQX1 mem_reg_15__5_ ( .D(N893), .C(net10511), .Q(mem_15__5_) );
  DFFQX1 mem_reg_14__5_ ( .D(N902), .C(net10506), .Q(mem_14__5_) );
  DFFQX1 mem_reg_13__5_ ( .D(N911), .C(net10501), .Q(mem_13__5_) );
  DFFQX1 mem_reg_12__5_ ( .D(N920), .C(net10496), .Q(mem_12__5_) );
  DFFQX1 mem_reg_11__5_ ( .D(N929), .C(net10491), .Q(mem_11__5_) );
  DFFQX1 mem_reg_10__5_ ( .D(N938), .C(net10486), .Q(mem_10__5_) );
  DFFQX1 mem_reg_9__5_ ( .D(N947), .C(net10481), .Q(mem_9__5_) );
  DFFQX1 mem_reg_8__5_ ( .D(N956), .C(net10476), .Q(mem_8__5_) );
  DFFQX1 mem_reg_27__4_ ( .D(N784), .C(net10571), .Q(mem_27__4_) );
  DFFQX1 mem_reg_26__4_ ( .D(N793), .C(net10566), .Q(mem_26__4_) );
  DFFQX1 mem_reg_25__4_ ( .D(N802), .C(net10561), .Q(mem_25__4_) );
  DFFQX1 mem_reg_24__4_ ( .D(N811), .C(net10556), .Q(mem_24__4_) );
  DFFQX1 mem_reg_23__4_ ( .D(N820), .C(net10551), .Q(mem_23__4_) );
  DFFQX1 mem_reg_22__4_ ( .D(N829), .C(net10546), .Q(mem_22__4_) );
  DFFQX1 mem_reg_21__4_ ( .D(N838), .C(net10541), .Q(mem_21__4_) );
  DFFQX1 mem_reg_20__4_ ( .D(N847), .C(net10536), .Q(mem_20__4_) );
  DFFQX1 mem_reg_19__4_ ( .D(N856), .C(net10531), .Q(mem_19__4_) );
  DFFQX1 mem_reg_18__4_ ( .D(N865), .C(net10526), .Q(mem_18__4_) );
  DFFQX1 mem_reg_17__4_ ( .D(N874), .C(net10521), .Q(mem_17__4_) );
  DFFQX1 mem_reg_16__4_ ( .D(N883), .C(net10516), .Q(mem_16__4_) );
  DFFQX1 mem_reg_15__4_ ( .D(N892), .C(net10511), .Q(mem_15__4_) );
  DFFQX1 mem_reg_14__4_ ( .D(N901), .C(net10506), .Q(mem_14__4_) );
  DFFQX1 mem_reg_13__4_ ( .D(N910), .C(net10501), .Q(mem_13__4_) );
  DFFQX1 mem_reg_12__4_ ( .D(N919), .C(net10496), .Q(mem_12__4_) );
  DFFQX1 mem_reg_11__4_ ( .D(N928), .C(net10491), .Q(mem_11__4_) );
  DFFQX1 mem_reg_10__4_ ( .D(N937), .C(net10486), .Q(mem_10__4_) );
  DFFQX1 mem_reg_9__4_ ( .D(N946), .C(net10481), .Q(mem_9__4_) );
  DFFQX1 mem_reg_8__4_ ( .D(N955), .C(net10476), .Q(mem_8__4_) );
  DFFQX1 mem_reg_27__3_ ( .D(N783), .C(net10571), .Q(mem_27__3_) );
  DFFQX1 mem_reg_26__3_ ( .D(N792), .C(net10566), .Q(mem_26__3_) );
  DFFQX1 mem_reg_25__3_ ( .D(N801), .C(net10561), .Q(mem_25__3_) );
  DFFQX1 mem_reg_24__3_ ( .D(N810), .C(net10556), .Q(mem_24__3_) );
  DFFQX1 mem_reg_23__3_ ( .D(N819), .C(net10551), .Q(mem_23__3_) );
  DFFQX1 mem_reg_22__3_ ( .D(N828), .C(net10546), .Q(mem_22__3_) );
  DFFQX1 mem_reg_21__3_ ( .D(N837), .C(net10541), .Q(mem_21__3_) );
  DFFQX1 mem_reg_20__3_ ( .D(N846), .C(net10536), .Q(mem_20__3_) );
  DFFQX1 mem_reg_19__3_ ( .D(N855), .C(net10531), .Q(mem_19__3_) );
  DFFQX1 mem_reg_18__3_ ( .D(N864), .C(net10526), .Q(mem_18__3_) );
  DFFQX1 mem_reg_17__3_ ( .D(N873), .C(net10521), .Q(mem_17__3_) );
  DFFQX1 mem_reg_16__3_ ( .D(N882), .C(net10516), .Q(mem_16__3_) );
  DFFQX1 mem_reg_15__3_ ( .D(N891), .C(net10511), .Q(mem_15__3_) );
  DFFQX1 mem_reg_14__3_ ( .D(N900), .C(net10506), .Q(mem_14__3_) );
  DFFQX1 mem_reg_13__3_ ( .D(N909), .C(net10501), .Q(mem_13__3_) );
  DFFQX1 mem_reg_12__3_ ( .D(N918), .C(net10496), .Q(mem_12__3_) );
  DFFQX1 mem_reg_11__3_ ( .D(N927), .C(net10491), .Q(mem_11__3_) );
  DFFQX1 mem_reg_10__3_ ( .D(N936), .C(net10486), .Q(mem_10__3_) );
  DFFQX1 mem_reg_9__3_ ( .D(N945), .C(net10481), .Q(mem_9__3_) );
  DFFQX1 mem_reg_8__3_ ( .D(N954), .C(net10476), .Q(mem_8__3_) );
  DFFQX1 mem_reg_27__2_ ( .D(N782), .C(net10571), .Q(mem_27__2_) );
  DFFQX1 mem_reg_26__2_ ( .D(N791), .C(net10566), .Q(mem_26__2_) );
  DFFQX1 mem_reg_25__2_ ( .D(N800), .C(net10561), .Q(mem_25__2_) );
  DFFQX1 mem_reg_24__2_ ( .D(N809), .C(net10556), .Q(mem_24__2_) );
  DFFQX1 mem_reg_23__2_ ( .D(N818), .C(net10551), .Q(mem_23__2_) );
  DFFQX1 mem_reg_22__2_ ( .D(N827), .C(net10546), .Q(mem_22__2_) );
  DFFQX1 mem_reg_21__2_ ( .D(N836), .C(net10541), .Q(mem_21__2_) );
  DFFQX1 mem_reg_20__2_ ( .D(N845), .C(net10536), .Q(mem_20__2_) );
  DFFQX1 mem_reg_19__2_ ( .D(N854), .C(net10531), .Q(mem_19__2_) );
  DFFQX1 mem_reg_18__2_ ( .D(N863), .C(net10526), .Q(mem_18__2_) );
  DFFQX1 mem_reg_17__2_ ( .D(N872), .C(net10521), .Q(mem_17__2_) );
  DFFQX1 mem_reg_16__2_ ( .D(N881), .C(net10516), .Q(mem_16__2_) );
  DFFQX1 mem_reg_15__2_ ( .D(N890), .C(net10511), .Q(mem_15__2_) );
  DFFQX1 mem_reg_14__2_ ( .D(N899), .C(net10506), .Q(mem_14__2_) );
  DFFQX1 mem_reg_13__2_ ( .D(N908), .C(net10501), .Q(mem_13__2_) );
  DFFQX1 mem_reg_12__2_ ( .D(N917), .C(net10496), .Q(mem_12__2_) );
  DFFQX1 mem_reg_11__2_ ( .D(N926), .C(net10491), .Q(mem_11__2_) );
  DFFQX1 mem_reg_10__2_ ( .D(N935), .C(net10486), .Q(mem_10__2_) );
  DFFQX1 mem_reg_9__2_ ( .D(N944), .C(net10481), .Q(mem_9__2_) );
  DFFQX1 mem_reg_8__2_ ( .D(N953), .C(net10476), .Q(mem_8__2_) );
  DFFQX1 mem_reg_27__1_ ( .D(N781), .C(net10571), .Q(mem_27__1_) );
  DFFQX1 mem_reg_26__1_ ( .D(N790), .C(net10566), .Q(mem_26__1_) );
  DFFQX1 mem_reg_25__1_ ( .D(N799), .C(net10561), .Q(mem_25__1_) );
  DFFQX1 mem_reg_24__1_ ( .D(N808), .C(net10556), .Q(mem_24__1_) );
  DFFQX1 mem_reg_23__1_ ( .D(N817), .C(net10551), .Q(mem_23__1_) );
  DFFQX1 mem_reg_22__1_ ( .D(N826), .C(net10546), .Q(mem_22__1_) );
  DFFQX1 mem_reg_21__1_ ( .D(N835), .C(net10541), .Q(mem_21__1_) );
  DFFQX1 mem_reg_20__1_ ( .D(N844), .C(net10536), .Q(mem_20__1_) );
  DFFQX1 mem_reg_19__1_ ( .D(N853), .C(net10531), .Q(mem_19__1_) );
  DFFQX1 mem_reg_18__1_ ( .D(N862), .C(net10526), .Q(mem_18__1_) );
  DFFQX1 mem_reg_17__1_ ( .D(N871), .C(net10521), .Q(mem_17__1_) );
  DFFQX1 mem_reg_16__1_ ( .D(N880), .C(net10516), .Q(mem_16__1_) );
  DFFQX1 mem_reg_15__1_ ( .D(N889), .C(net10511), .Q(mem_15__1_) );
  DFFQX1 mem_reg_14__1_ ( .D(N898), .C(net10506), .Q(mem_14__1_) );
  DFFQX1 mem_reg_13__1_ ( .D(N907), .C(net10501), .Q(mem_13__1_) );
  DFFQX1 mem_reg_12__1_ ( .D(N916), .C(net10496), .Q(mem_12__1_) );
  DFFQX1 mem_reg_11__1_ ( .D(N925), .C(net10491), .Q(mem_11__1_) );
  DFFQX1 mem_reg_10__1_ ( .D(N934), .C(net10486), .Q(mem_10__1_) );
  DFFQX1 mem_reg_9__1_ ( .D(N943), .C(net10481), .Q(mem_9__1_) );
  DFFQX1 mem_reg_8__1_ ( .D(N952), .C(net10476), .Q(mem_8__1_) );
  DFFQX1 mem_reg_27__0_ ( .D(N780), .C(net10571), .Q(mem_27__0_) );
  DFFQX1 mem_reg_26__0_ ( .D(N789), .C(net10566), .Q(mem_26__0_) );
  DFFQX1 mem_reg_25__0_ ( .D(N798), .C(net10561), .Q(mem_25__0_) );
  DFFQX1 mem_reg_24__0_ ( .D(N807), .C(net10556), .Q(mem_24__0_) );
  DFFQX1 mem_reg_23__0_ ( .D(N816), .C(net10551), .Q(mem_23__0_) );
  DFFQX1 mem_reg_22__0_ ( .D(N825), .C(net10546), .Q(mem_22__0_) );
  DFFQX1 mem_reg_21__0_ ( .D(N834), .C(net10541), .Q(mem_21__0_) );
  DFFQX1 mem_reg_20__0_ ( .D(N843), .C(net10536), .Q(mem_20__0_) );
  DFFQX1 mem_reg_19__0_ ( .D(N852), .C(net10531), .Q(mem_19__0_) );
  DFFQX1 mem_reg_18__0_ ( .D(N861), .C(net10526), .Q(mem_18__0_) );
  DFFQX1 mem_reg_17__0_ ( .D(N870), .C(net10521), .Q(mem_17__0_) );
  DFFQX1 mem_reg_16__0_ ( .D(N879), .C(net10516), .Q(mem_16__0_) );
  DFFQX1 mem_reg_15__0_ ( .D(N888), .C(net10511), .Q(mem_15__0_) );
  DFFQX1 mem_reg_14__0_ ( .D(N897), .C(net10506), .Q(mem_14__0_) );
  DFFQX1 mem_reg_13__0_ ( .D(N906), .C(net10501), .Q(mem_13__0_) );
  DFFQX1 mem_reg_12__0_ ( .D(N915), .C(net10496), .Q(mem_12__0_) );
  DFFQX1 mem_reg_11__0_ ( .D(N924), .C(net10491), .Q(mem_11__0_) );
  DFFQX1 mem_reg_10__0_ ( .D(N933), .C(net10486), .Q(mem_10__0_) );
  DFFQX1 mem_reg_9__0_ ( .D(N942), .C(net10481), .Q(mem_9__0_) );
  DFFQX1 mem_reg_8__0_ ( .D(N951), .C(net10476), .Q(mem_8__0_) );
  DFFQX1 mem_reg_1__0_ ( .D(N1014), .C(net10441), .Q(dat_7_1[0]) );
  DFFQX1 mem_reg_1__3_ ( .D(N1017), .C(net10441), .Q(dat_7_1[3]) );
  DFFQX1 mem_reg_1__2_ ( .D(N1016), .C(net10441), .Q(dat_7_1[2]) );
  DFFQX1 mem_reg_1__1_ ( .D(N1015), .C(net10441), .Q(dat_7_1[1]) );
  DFFQX1 locked_reg ( .D(ps_locked), .C(clk), .Q(locked) );
  DFFQX1 mem_reg_7__7_ ( .D(N967), .C(net10471), .Q(dat_7_1[55]) );
  DFFQX1 mem_reg_7__5_ ( .D(N965), .C(net10471), .Q(dat_7_1[53]) );
  DFFQX1 mem_reg_7__4_ ( .D(N964), .C(net10471), .Q(dat_7_1[52]) );
  DFFQX1 mem_reg_6__4_ ( .D(N973), .C(net10466), .Q(dat_7_1[44]) );
  DFFQX1 mem_reg_7__3_ ( .D(N963), .C(net10471), .Q(dat_7_1[51]) );
  DFFQX1 mem_reg_7__2_ ( .D(N962), .C(net10471), .Q(dat_7_1[50]) );
  DFFQX1 mem_reg_6__2_ ( .D(N971), .C(net10466), .Q(dat_7_1[42]) );
  DFFQX1 mem_reg_2__6_ ( .D(N1011), .C(net10446), .Q(dat_7_1[14]) );
  DFFQX1 mem_reg_6__7_ ( .D(N976), .C(net10466), .Q(dat_7_1[47]) );
  DFFQX1 mem_reg_7__6_ ( .D(N966), .C(net10471), .Q(dat_7_1[54]) );
  DFFQX1 mem_reg_6__6_ ( .D(N975), .C(net10466), .Q(dat_7_1[46]) );
  DFFQX1 mem_reg_6__5_ ( .D(N974), .C(net10466), .Q(dat_7_1[45]) );
  DFFQX1 mem_reg_6__3_ ( .D(N972), .C(net10466), .Q(dat_7_1[43]) );
  DFFQX1 mem_reg_7__1_ ( .D(N961), .C(net10471), .Q(dat_7_1[49]) );
  DFFQX1 mem_reg_6__1_ ( .D(N970), .C(net10466), .Q(dat_7_1[41]) );
  DFFQX1 mem_reg_7__0_ ( .D(N960), .C(net10471), .Q(dat_7_1[48]) );
  DFFQX1 mem_reg_6__0_ ( .D(N969), .C(net10466), .Q(dat_7_1[40]) );
  DFFQX1 mem_reg_5__7_ ( .D(N985), .C(net10461), .Q(dat_7_1[39]) );
  DFFQX1 mem_reg_4__7_ ( .D(N994), .C(net10456), .Q(dat_7_1[31]) );
  DFFQX1 mem_reg_5__6_ ( .D(N984), .C(net10461), .Q(dat_7_1[38]) );
  DFFQX1 mem_reg_4__6_ ( .D(N993), .C(net10456), .Q(dat_7_1[30]) );
  DFFQX1 mem_reg_5__5_ ( .D(N983), .C(net10461), .Q(dat_7_1[37]) );
  DFFQX1 mem_reg_4__5_ ( .D(N992), .C(net10456), .Q(dat_7_1[29]) );
  DFFQX1 mem_reg_5__4_ ( .D(N982), .C(net10461), .Q(dat_7_1[36]) );
  DFFQX1 mem_reg_4__4_ ( .D(N991), .C(net10456), .Q(dat_7_1[28]) );
  DFFQX1 mem_reg_5__3_ ( .D(N981), .C(net10461), .Q(dat_7_1[35]) );
  DFFQX1 mem_reg_4__3_ ( .D(N990), .C(net10456), .Q(dat_7_1[27]) );
  DFFQX1 mem_reg_5__2_ ( .D(N980), .C(net10461), .Q(dat_7_1[34]) );
  DFFQX1 mem_reg_4__2_ ( .D(N989), .C(net10456), .Q(dat_7_1[26]) );
  DFFQX1 mem_reg_5__1_ ( .D(N979), .C(net10461), .Q(dat_7_1[33]) );
  DFFQX1 mem_reg_4__1_ ( .D(N988), .C(net10456), .Q(dat_7_1[25]) );
  DFFQX1 mem_reg_5__0_ ( .D(N978), .C(net10461), .Q(dat_7_1[32]) );
  DFFQX1 mem_reg_4__0_ ( .D(N987), .C(net10456), .Q(dat_7_1[24]) );
  DFFQX1 mem_reg_3__3_ ( .D(N999), .C(net10451), .Q(dat_7_1[19]) );
  DFFQX1 mem_reg_3__2_ ( .D(N998), .C(net10451), .Q(dat_7_1[18]) );
  DFFQX1 mem_reg_3__1_ ( .D(N997), .C(net10451), .Q(dat_7_1[17]) );
  DFFQX1 mem_reg_3__0_ ( .D(N996), .C(net10451), .Q(dat_7_1[16]) );
  DFFQX1 mem_reg_2__7_ ( .D(N1012), .C(net10446), .Q(dat_7_1[15]) );
  DFFQX1 mem_reg_2__5_ ( .D(N1010), .C(net10446), .Q(dat_7_1[13]) );
  DFFQX1 mem_reg_1__7_ ( .D(N1021), .C(net10441), .Q(dat_7_1[7]) );
  DFFQX1 mem_reg_1__6_ ( .D(N1020), .C(net10441), .Q(dat_7_1[6]) );
  DFFQX1 mem_reg_1__5_ ( .D(N1019), .C(net10441), .Q(dat_7_1[5]) );
  DFFQX1 mem_reg_3__7_ ( .D(N1003), .C(net10451), .Q(dat_7_1[23]) );
  DFFQX1 mem_reg_3__6_ ( .D(N1002), .C(net10451), .Q(dat_7_1[22]) );
  DFFQX1 mem_reg_2__3_ ( .D(N1008), .C(net10446), .Q(dat_7_1[11]) );
  DFFQX1 mem_reg_2__1_ ( .D(N1006), .C(net10446), .Q(dat_7_1[9]) );
  DFFQX1 mem_reg_1__4_ ( .D(N1018), .C(net10441), .Q(dat_7_1[4]) );
  DFFQX1 mem_reg_3__5_ ( .D(N1001), .C(net10451), .Q(dat_7_1[21]) );
  DFFQX1 mem_reg_3__4_ ( .D(N1000), .C(net10451), .Q(dat_7_1[20]) );
  DFFQX1 mem_reg_2__4_ ( .D(N1009), .C(net10446), .Q(dat_7_1[12]) );
  DFFQX1 mem_reg_2__2_ ( .D(N1007), .C(net10446), .Q(dat_7_1[10]) );
  DFFQX1 mem_reg_2__0_ ( .D(N1005), .C(net10446), .Q(dat_7_1[8]) );
  DFFQX1 mem_reg_0__4_ ( .D(N1027), .C(net10435), .Q(rdat0[4]) );
  DFFQX1 mem_reg_0__1_ ( .D(N1024), .C(net10435), .Q(rdat0[1]) );
  DFFQX1 mem_reg_0__0_ ( .D(N1023), .C(net10435), .Q(rdat0[0]) );
  DFFQX1 mem_reg_0__7_ ( .D(N1030), .C(net10435), .Q(rdat0[7]) );
  DFFQX1 mem_reg_0__6_ ( .D(N1029), .C(net10435), .Q(rdat0[6]) );
  DFFQX1 mem_reg_0__5_ ( .D(N1028), .C(net10435), .Q(rdat0[5]) );
  DFFQX1 mem_reg_0__3_ ( .D(N1026), .C(net10435), .Q(rdat0[3]) );
  DFFQX1 mem_reg_0__2_ ( .D(N1025), .C(net10435), .Q(rdat0[2]) );
  DFFQX1 pshptr_reg_5_ ( .D(N1059), .C(net10606), .Q(ptr[5]) );
  DFFQX1 pshptr_reg_1_ ( .D(N1055), .C(net10606), .Q(ptr[1]) );
  DFFQX1 pshptr_reg_0_ ( .D(N1054), .C(net10606), .Q(ptr[0]) );
  DFFQX1 pshptr_reg_4_ ( .D(N1058), .C(net10606), .Q(ptr[4]) );
  DFFQX1 pshptr_reg_2_ ( .D(N1056), .C(net10606), .Q(ptr[2]) );
  DFFQX1 pshptr_reg_3_ ( .D(N1057), .C(net10606), .Q(ptr[3]) );
  NOR3X1 U3 ( .A(n300), .B(n299), .C(ptr[4]), .Y(one) );
  INVX1 U4 ( .A(ptr[3]), .Y(n103) );
  INVX1 U5 ( .A(ptr[0]), .Y(n299) );
  OR3XL U6 ( .A(ptr[5]), .B(ptr[1]), .C(n107), .Y(n300) );
  INVX1 U7 ( .A(n162), .Y(n1) );
  INVX1 U8 ( .A(n193), .Y(n2) );
  AND3XL U9 ( .A(ptr[4]), .B(ptr[0]), .C(n298), .Y(half) );
  NAND21X1 U10 ( .B(ptr[2]), .A(n103), .Y(n107) );
  OAI31XL U11 ( .A(n107), .B(ptr[4]), .C(ptr[1]), .D(ptr[5]), .Y(n230) );
  INVX1 U12 ( .A(n74), .Y(n72) );
  INVX1 U13 ( .A(n102), .Y(n101) );
  INVX1 U14 ( .A(n102), .Y(n100) );
  INVX1 U15 ( .A(n98), .Y(n97) );
  INVX1 U16 ( .A(n98), .Y(n96) );
  INVX1 U17 ( .A(n94), .Y(n93) );
  INVX1 U18 ( .A(n94), .Y(n92) );
  INVX1 U19 ( .A(n74), .Y(n73) );
  INVX1 U20 ( .A(n74), .Y(n71) );
  INVX1 U21 ( .A(n367), .Y(n74) );
  INVX1 U22 ( .A(n86), .Y(n84) );
  INVX1 U23 ( .A(n82), .Y(n80) );
  INVX1 U24 ( .A(n78), .Y(n76) );
  INVX1 U25 ( .A(n86), .Y(n85) );
  INVX1 U26 ( .A(n82), .Y(n81) );
  INVX1 U27 ( .A(n78), .Y(n77) );
  INVX1 U28 ( .A(n102), .Y(n99) );
  INVX1 U29 ( .A(n382), .Y(n102) );
  INVX1 U30 ( .A(n98), .Y(n95) );
  INVX1 U31 ( .A(n380), .Y(n98) );
  INVX1 U32 ( .A(n94), .Y(n91) );
  INVX1 U33 ( .A(n378), .Y(n94) );
  INVX1 U34 ( .A(n90), .Y(n88) );
  INVX1 U35 ( .A(n90), .Y(n87) );
  INVX1 U36 ( .A(n90), .Y(n89) );
  NAND21X1 U37 ( .B(n359), .A(n31), .Y(n367) );
  NAND21X1 U38 ( .B(n350), .A(n31), .Y(n382) );
  NAND21X1 U39 ( .B(n351), .A(n31), .Y(n380) );
  NAND21X1 U40 ( .B(n49), .A(n31), .Y(n378) );
  INVX1 U41 ( .A(n82), .Y(n79) );
  INVX1 U42 ( .A(n371), .Y(n82) );
  INVX1 U43 ( .A(n78), .Y(n75) );
  INVX1 U44 ( .A(n369), .Y(n78) );
  INVX1 U45 ( .A(n373), .Y(n86) );
  INVX1 U46 ( .A(n86), .Y(n83) );
  INVX1 U47 ( .A(n131), .Y(n275) );
  AND2X1 U48 ( .A(n287), .B(n284), .Y(n3) );
  INVX1 U49 ( .A(n133), .Y(n360) );
  NAND21X1 U50 ( .B(n225), .A(n282), .Y(n133) );
  AND2X1 U51 ( .A(n283), .B(n280), .Y(n4) );
  INVX1 U52 ( .A(n138), .Y(n349) );
  NAND21X1 U53 ( .B(n137), .A(n278), .Y(n138) );
  INVX1 U54 ( .A(n143), .Y(n345) );
  NAND21X1 U55 ( .B(n275), .A(n273), .Y(n143) );
  INVX1 U56 ( .A(n179), .Y(n322) );
  NAND21X1 U57 ( .B(n247), .A(n244), .Y(n179) );
  AND2X1 U58 ( .A(n267), .B(n265), .Y(n5) );
  AND2X1 U59 ( .A(n241), .B(n239), .Y(n6) );
  INVX1 U60 ( .A(n140), .Y(n347) );
  NAND21X1 U61 ( .B(n294), .A(n279), .Y(n140) );
  INVX1 U62 ( .A(n224), .Y(n305) );
  NAND21X1 U63 ( .B(n31), .A(n306), .Y(n224) );
  INVX1 U64 ( .A(n228), .Y(n304) );
  NAND21X1 U65 ( .B(n31), .A(n3), .Y(n228) );
  INVX1 U66 ( .A(n134), .Y(n358) );
  NAND21X1 U67 ( .B(n31), .A(n360), .Y(n134) );
  INVX1 U68 ( .A(n136), .Y(n353) );
  NAND21X1 U69 ( .B(n34), .A(n4), .Y(n136) );
  INVX1 U70 ( .A(n139), .Y(n348) );
  NAND21X1 U71 ( .B(n34), .A(n349), .Y(n139) );
  INVX1 U72 ( .A(n141), .Y(n346) );
  NAND21X1 U73 ( .B(n33), .A(n347), .Y(n141) );
  INVX1 U74 ( .A(n144), .Y(n344) );
  NAND21X1 U75 ( .B(n34), .A(n345), .Y(n144) );
  INVX1 U76 ( .A(n145), .Y(n343) );
  NAND21X1 U77 ( .B(n34), .A(n16), .Y(n145) );
  INVX1 U78 ( .A(n148), .Y(n342) );
  NAND21X1 U79 ( .B(n34), .A(n7), .Y(n148) );
  INVX1 U80 ( .A(n149), .Y(n341) );
  NAND21X1 U81 ( .B(n34), .A(n8), .Y(n149) );
  INVX1 U82 ( .A(n153), .Y(n338) );
  NAND21X1 U83 ( .B(n34), .A(n5), .Y(n153) );
  INVX1 U84 ( .A(n156), .Y(n336) );
  NAND21X1 U85 ( .B(n34), .A(n337), .Y(n156) );
  INVX1 U86 ( .A(n161), .Y(n334) );
  NAND21X1 U87 ( .B(n33), .A(n335), .Y(n161) );
  INVX1 U88 ( .A(n164), .Y(n332) );
  NAND21X1 U89 ( .B(n33), .A(n333), .Y(n164) );
  INVX1 U90 ( .A(n168), .Y(n330) );
  NAND21X1 U91 ( .B(n33), .A(n331), .Y(n168) );
  INVX1 U92 ( .A(n169), .Y(n329) );
  NAND21X1 U93 ( .B(n33), .A(n9), .Y(n169) );
  INVX1 U94 ( .A(n170), .Y(n328) );
  NAND21X1 U95 ( .B(n33), .A(n10), .Y(n170) );
  INVX1 U96 ( .A(n171), .Y(n327) );
  NAND21X1 U97 ( .B(n33), .A(n11), .Y(n171) );
  INVX1 U98 ( .A(n173), .Y(n326) );
  NAND21X1 U99 ( .B(n33), .A(n12), .Y(n173) );
  INVX1 U100 ( .A(n174), .Y(n325) );
  NAND21X1 U101 ( .B(n33), .A(n13), .Y(n174) );
  INVX1 U102 ( .A(n177), .Y(n323) );
  NAND21X1 U103 ( .B(n33), .A(n324), .Y(n177) );
  INVX1 U104 ( .A(n180), .Y(n321) );
  NAND21X1 U105 ( .B(n32), .A(n322), .Y(n180) );
  INVX1 U106 ( .A(n186), .Y(n319) );
  NAND21X1 U107 ( .B(n32), .A(n320), .Y(n186) );
  INVX1 U108 ( .A(n188), .Y(n318) );
  NAND21X1 U109 ( .B(n32), .A(n14), .Y(n188) );
  INVX1 U110 ( .A(n190), .Y(n317) );
  NAND21X1 U111 ( .B(n32), .A(n6), .Y(n190) );
  INVX1 U112 ( .A(n199), .Y(n314) );
  NAND21X1 U113 ( .B(n32), .A(n15), .Y(n199) );
  INVX1 U114 ( .A(n208), .Y(n310) );
  NAND21X1 U115 ( .B(n32), .A(n311), .Y(n208) );
  INVX1 U116 ( .A(n220), .Y(n307) );
  NAND21X1 U117 ( .B(n32), .A(n17), .Y(n220) );
  INVX1 U118 ( .A(n376), .Y(n90) );
  INVX1 U119 ( .A(n154), .Y(n263) );
  NAND21X1 U120 ( .B(n200), .A(n159), .Y(n154) );
  INVX1 U121 ( .A(n201), .Y(n234) );
  NAND21X1 U122 ( .B(n200), .A(n206), .Y(n201) );
  NAND21X1 U123 ( .B(n226), .A(n225), .Y(n287) );
  INVX1 U124 ( .A(n130), .Y(n127) );
  NAND21X1 U125 ( .B(n204), .A(n275), .Y(n279) );
  INVX1 U126 ( .A(n281), .Y(n137) );
  INVX1 U127 ( .A(fifowdat[3]), .Y(n67) );
  INVX1 U128 ( .A(fifowdat[3]), .Y(n68) );
  INVX1 U129 ( .A(fifowdat[3]), .Y(n69) );
  INVX1 U130 ( .A(n126), .Y(n124) );
  INVX1 U131 ( .A(n302), .Y(n303) );
  NAND21X1 U132 ( .B(n301), .A(n18), .Y(n302) );
  NAND21X1 U133 ( .B(n355), .A(n31), .Y(n373) );
  NAND21X1 U134 ( .B(n356), .A(n31), .Y(n371) );
  NAND21X1 U135 ( .B(n65), .A(n31), .Y(n369) );
  INVX1 U136 ( .A(n129), .Y(n120) );
  INVX1 U137 ( .A(n36), .Y(n31) );
  INVX1 U138 ( .A(n614), .Y(n106) );
  OR2X1 U139 ( .A(n277), .B(n227), .Y(n284) );
  OR2X1 U140 ( .A(n277), .B(n191), .Y(n282) );
  OR2X1 U141 ( .A(n277), .B(n198), .Y(n280) );
  OR2X1 U142 ( .A(n277), .B(n200), .Y(n278) );
  NAND21X1 U143 ( .B(n210), .A(n159), .Y(n273) );
  NAND21X1 U144 ( .B(n210), .A(n175), .Y(n260) );
  NAND21X1 U145 ( .B(n210), .A(n206), .Y(n244) );
  NAND21X1 U146 ( .B(n227), .A(n159), .Y(n268) );
  NAND21X1 U147 ( .B(n198), .A(n159), .Y(n265) );
  NAND21X1 U148 ( .B(n227), .A(n175), .Y(n254) );
  NAND21X1 U149 ( .B(n191), .A(n175), .Y(n252) );
  NAND21X1 U150 ( .B(n198), .A(n175), .Y(n250) );
  NAND21X1 U151 ( .B(n200), .A(n175), .Y(n248) );
  NAND21X1 U152 ( .B(n227), .A(n206), .Y(n239) );
  NAND21X1 U153 ( .B(n198), .A(n206), .Y(n236) );
  AO21X1 U154 ( .B(n158), .C(n147), .A(n272), .Y(n274) );
  NAND21X1 U155 ( .B(n158), .A(n261), .Y(n131) );
  INVX1 U156 ( .A(n176), .Y(n324) );
  NAND21X1 U157 ( .B(n175), .A(n249), .Y(n176) );
  INVX1 U158 ( .A(n223), .Y(n306) );
  NAND21X1 U159 ( .B(n293), .A(n286), .Y(n223) );
  INVX1 U160 ( .A(n155), .Y(n337) );
  NAND21X1 U161 ( .B(n263), .A(n23), .Y(n155) );
  INVX1 U162 ( .A(n167), .Y(n331) );
  NAND21X1 U163 ( .B(n258), .A(n24), .Y(n167) );
  INVX1 U164 ( .A(n185), .Y(n320) );
  NAND21X1 U165 ( .B(n242), .A(n245), .Y(n185) );
  INVX1 U166 ( .A(n163), .Y(n333) );
  NAND21X1 U167 ( .B(n261), .A(n260), .Y(n163) );
  INVX1 U168 ( .A(n262), .Y(n159) );
  INVX1 U169 ( .A(n233), .Y(n206) );
  NAND21X1 U170 ( .B(n36), .A(fifowdat[7]), .Y(n376) );
  AO21X1 U171 ( .B(n295), .C(n294), .A(n18), .Y(N1022) );
  AND2X1 U172 ( .A(n272), .B(n269), .Y(n7) );
  AND2X1 U173 ( .A(n270), .B(n268), .Y(n8) );
  AND2X1 U174 ( .A(n259), .B(n256), .Y(n9) );
  AND2X1 U175 ( .A(n257), .B(n254), .Y(n10) );
  AND2X1 U176 ( .A(n255), .B(n252), .Y(n11) );
  AND2X1 U177 ( .A(n253), .B(n250), .Y(n12) );
  AND2X1 U178 ( .A(n251), .B(n248), .Y(n13) );
  AND2X1 U179 ( .A(n243), .B(n240), .Y(n14) );
  AND2X1 U180 ( .A(n238), .B(n236), .Y(n15) );
  AND2X1 U181 ( .A(n274), .B(n271), .Y(n16) );
  INVX1 U182 ( .A(n160), .Y(n335) );
  NAND21X1 U183 ( .B(n159), .A(n264), .Y(n160) );
  INVX1 U184 ( .A(n207), .Y(n311) );
  NAND21X1 U185 ( .B(n206), .A(n235), .Y(n207) );
  AND2X1 U186 ( .A(n229), .B(n25), .Y(n17) );
  INVX1 U187 ( .A(n277), .Y(n294) );
  INVX1 U188 ( .A(n152), .Y(n339) );
  NAND21X1 U189 ( .B(n34), .A(n340), .Y(n152) );
  INVX1 U190 ( .A(n195), .Y(n315) );
  NAND21X1 U191 ( .B(n32), .A(n316), .Y(n195) );
  INVX1 U192 ( .A(n203), .Y(n312) );
  NAND21X1 U193 ( .B(n32), .A(n313), .Y(n203) );
  INVX1 U194 ( .A(n216), .Y(n308) );
  NAND21X1 U195 ( .B(n32), .A(n309), .Y(n216) );
  INVX1 U196 ( .A(n35), .Y(n33) );
  INVX1 U197 ( .A(n36), .Y(n32) );
  INVX1 U198 ( .A(n35), .Y(n34) );
  OAI22X1 U199 ( .A(n277), .B(n276), .C(n275), .D(n291), .Y(N959) );
  OAI22X1 U200 ( .A(n276), .B(n262), .C(n261), .D(n291), .Y(N887) );
  INVX1 U201 ( .A(n150), .Y(n266) );
  NAND21X1 U202 ( .B(n191), .A(n159), .Y(n150) );
  INVX1 U203 ( .A(n192), .Y(n237) );
  NAND21X1 U204 ( .B(n191), .A(n206), .Y(n192) );
  INVX1 U205 ( .A(n214), .Y(n231) );
  NAND21X1 U206 ( .B(n218), .A(n217), .Y(n214) );
  NAND21X1 U207 ( .B(n158), .A(n115), .Y(n130) );
  AO21X1 U208 ( .B(n158), .C(n197), .A(n23), .Y(n267) );
  AO21X1 U209 ( .B(n38), .C(n290), .A(n301), .Y(N1013) );
  OAI21BBX1 U210 ( .A(n37), .B(n287), .C(n286), .Y(N1004) );
  OAI21BBX1 U211 ( .A(n37), .B(n285), .C(n284), .Y(N995) );
  OAI21BBX1 U212 ( .A(n37), .B(n283), .C(n282), .Y(N986) );
  OAI21BBX1 U213 ( .A(n37), .B(n281), .C(n280), .Y(N977) );
  OAI21BBX1 U214 ( .A(n38), .B(n279), .C(n278), .Y(N968) );
  AO21X1 U215 ( .B(n38), .C(n264), .A(n263), .Y(N896) );
  OAI21BBX1 U216 ( .A(n35), .B(n249), .C(n248), .Y(N824) );
  AO21X1 U217 ( .B(n35), .C(n235), .A(n234), .Y(N752) );
  OAI21BBX1 U218 ( .A(n37), .B(n274), .C(n273), .Y(N950) );
  OAI21BBX1 U219 ( .A(n38), .B(n272), .C(n271), .Y(N941) );
  OAI21BBX1 U220 ( .A(n35), .B(n270), .C(n269), .Y(N932) );
  OAI21BBX1 U221 ( .A(n23), .B(n37), .C(n265), .Y(N905) );
  OAI21BBX1 U222 ( .A(n24), .B(n37), .C(n260), .Y(N878) );
  OAI21BBX1 U223 ( .A(n37), .B(n257), .C(n256), .Y(N860) );
  OAI21BBX1 U224 ( .A(n38), .B(n255), .C(n254), .Y(N851) );
  OAI21BBX1 U225 ( .A(n38), .B(n253), .C(n252), .Y(N842) );
  OAI21BBX1 U226 ( .A(n38), .B(n251), .C(n250), .Y(N833) );
  OAI21BBX1 U227 ( .A(n245), .B(n37), .C(n244), .Y(N806) );
  OAI21BBX1 U228 ( .A(n36), .B(n241), .C(n240), .Y(N788) );
  AO21X1 U229 ( .B(n38), .C(n267), .A(n266), .Y(N914) );
  AO21X1 U230 ( .B(n35), .C(n259), .A(n258), .Y(N869) );
  AO21X1 U231 ( .B(n35), .C(n243), .A(n242), .Y(N797) );
  AO21X1 U232 ( .B(n35), .C(n238), .A(n237), .Y(N770) );
  AO21X1 U233 ( .B(n25), .C(n38), .A(n231), .Y(N734) );
  INVX1 U234 ( .A(n132), .Y(n142) );
  INVX1 U235 ( .A(n112), .Y(n226) );
  INVX1 U236 ( .A(n178), .Y(n205) );
  INVX1 U237 ( .A(n285), .Y(n225) );
  INVX1 U238 ( .A(n182), .Y(n247) );
  INVX1 U239 ( .A(n210), .Y(n295) );
  INVX1 U240 ( .A(n118), .Y(n115) );
  INVX1 U241 ( .A(n290), .Y(n293) );
  NAND21X1 U242 ( .B(n147), .A(n172), .Y(n200) );
  AO21X1 U243 ( .B(n205), .C(n226), .A(n189), .Y(n241) );
  NAND21X1 U244 ( .B(n197), .A(n137), .Y(n283) );
  NAND21X1 U245 ( .B(n172), .A(n275), .Y(n281) );
  INVX1 U246 ( .A(n184), .Y(n245) );
  NAND21X1 U247 ( .B(n183), .A(n182), .Y(n184) );
  INVX1 U248 ( .A(n276), .Y(n204) );
  INVX1 U249 ( .A(n359), .Y(fifowdat[3]) );
  INVX1 U250 ( .A(fifowdat[6]), .Y(n49) );
  INVX1 U251 ( .A(fifowdat[4]), .Y(n39) );
  INVX1 U252 ( .A(fifowdat[4]), .Y(n40) );
  INVX1 U253 ( .A(fifowdat[5]), .Y(n43) );
  INVX1 U254 ( .A(fifowdat[5]), .Y(n44) );
  INVX1 U255 ( .A(fifowdat[6]), .Y(n47) );
  INVX1 U256 ( .A(fifowdat[6]), .Y(n48) );
  INVX1 U257 ( .A(fifowdat[7]), .Y(n52) );
  INVX1 U258 ( .A(fifowdat[4]), .Y(n41) );
  INVX1 U259 ( .A(fifowdat[5]), .Y(n45) );
  INVX1 U260 ( .A(fifowdat[7]), .Y(n51) );
  NAND21X1 U261 ( .B(n613), .A(n612), .Y(n129) );
  OR2X1 U262 ( .A(n612), .B(n613), .Y(n126) );
  INVX1 U263 ( .A(n612), .Y(n361) );
  OAI22X1 U264 ( .A(n109), .B(n126), .C(n108), .D(n129), .Y(N1058) );
  XOR2X1 U265 ( .A(n130), .B(n1), .Y(n108) );
  XOR2X1 U266 ( .A(n122), .B(n1), .Y(n109) );
  AOI21X1 U267 ( .B(n293), .C(n292), .A(n291), .Y(n18) );
  OAI22BX1 U268 ( .B(n120), .A(n19), .D(n124), .C(n20), .Y(N1057) );
  AOI21X1 U269 ( .B(n158), .C(n118), .A(n127), .Y(n19) );
  XNOR2XL U270 ( .A(n158), .B(n119), .Y(n20) );
  OAI22BX1 U271 ( .B(n120), .A(n21), .D(n124), .C(n22), .Y(N1056) );
  AOI21X1 U272 ( .B(n2), .C(n116), .A(n115), .Y(n21) );
  XNOR2XL U273 ( .A(n2), .B(n117), .Y(n22) );
  OAI32X1 U274 ( .A(n129), .B(empty), .C(n147), .D(n121), .E(n126), .Y(N1054)
         );
  XOR2X1 U275 ( .A(full), .B(n147), .Y(n121) );
  INVX1 U276 ( .A(n291), .Y(n35) );
  INVX1 U277 ( .A(n291), .Y(n36) );
  OR2X1 U278 ( .A(n131), .B(n212), .Y(n277) );
  OR2X1 U279 ( .A(n277), .B(n222), .Y(n286) );
  NAND21X1 U280 ( .B(n222), .A(n159), .Y(n269) );
  NAND21X1 U281 ( .B(n222), .A(n175), .Y(n256) );
  NAND21X1 U282 ( .B(n222), .A(n206), .Y(n240) );
  NAND21X1 U283 ( .B(n288), .A(n159), .Y(n271) );
  AO21X1 U284 ( .B(n158), .C(n221), .A(n27), .Y(n272) );
  NAND21X1 U285 ( .B(n288), .A(n217), .Y(n229) );
  NAND21X1 U286 ( .B(n212), .A(n205), .Y(n233) );
  NAND32X1 U287 ( .B(n157), .C(n212), .A(n158), .Y(n262) );
  INVX1 U288 ( .A(n151), .Y(n340) );
  NAND21X1 U289 ( .B(n266), .A(n27), .Y(n151) );
  INVX1 U290 ( .A(n194), .Y(n316) );
  NAND21X1 U291 ( .B(n237), .A(n29), .Y(n194) );
  INVX1 U292 ( .A(n202), .Y(n313) );
  NAND21X1 U293 ( .B(n234), .A(n28), .Y(n202) );
  INVX1 U294 ( .A(n215), .Y(n309) );
  NAND21X1 U295 ( .B(n231), .A(n219), .Y(n215) );
  INVX1 U296 ( .A(n246), .Y(n175) );
  INVX1 U297 ( .A(n157), .Y(n261) );
  INVX1 U298 ( .A(n213), .Y(n217) );
  NAND21X1 U299 ( .B(n212), .A(n219), .Y(n213) );
  OAI22X1 U300 ( .A(n247), .B(n291), .C(n276), .D(n246), .Y(N815) );
  INVX1 U301 ( .A(n165), .Y(n258) );
  NAND21X1 U302 ( .B(n288), .A(n175), .Y(n165) );
  INVX1 U303 ( .A(n181), .Y(n242) );
  NAND21X1 U304 ( .B(n288), .A(n206), .Y(n181) );
  INVX1 U305 ( .A(n289), .Y(n301) );
  NAND21X1 U306 ( .B(n288), .A(n294), .Y(n289) );
  NAND32X1 U307 ( .B(n211), .C(n210), .A(n209), .Y(n218) );
  NAND21X1 U308 ( .B(n221), .A(n292), .Y(n132) );
  NAND21X1 U309 ( .B(n219), .A(n178), .Y(n182) );
  NAND21X1 U310 ( .B(n187), .A(n142), .Y(n210) );
  NAND21X1 U311 ( .B(n209), .A(n211), .Y(n178) );
  AO21X1 U312 ( .B(n211), .C(n187), .A(n182), .Y(n255) );
  NAND21X1 U313 ( .B(n132), .A(n187), .Y(n191) );
  AO21X1 U314 ( .B(n211), .C(n172), .A(n182), .Y(n251) );
  NAND21X1 U315 ( .B(n209), .A(n119), .Y(n122) );
  NAND21X1 U316 ( .B(empty), .A(n142), .Y(n116) );
  AO21X1 U317 ( .B(n158), .C(n226), .A(n27), .Y(n270) );
  AO21X1 U318 ( .B(n211), .C(n197), .A(n251), .Y(n253) );
  AO21X1 U319 ( .B(n205), .C(n197), .A(n28), .Y(n238) );
  AO21X1 U320 ( .B(n211), .C(n221), .A(n255), .Y(n259) );
  AO21X1 U321 ( .B(n211), .C(n226), .A(n255), .Y(n257) );
  INVX1 U322 ( .A(n209), .Y(n158) );
  NAND21X1 U323 ( .B(n292), .A(n221), .Y(n112) );
  NAND21X1 U324 ( .B(n187), .A(n275), .Y(n285) );
  NAND21X1 U325 ( .B(n221), .A(n225), .Y(n290) );
  OAI21BBX1 U326 ( .A(n27), .B(n37), .C(n268), .Y(N923) );
  OAI21BBX1 U327 ( .A(n29), .B(n38), .C(n239), .Y(N779) );
  OAI21BBX1 U328 ( .A(n28), .B(n35), .C(n236), .Y(N761) );
  AOI21X1 U329 ( .B(n261), .C(n196), .A(n275), .Y(n23) );
  AOI21X1 U330 ( .B(n183), .C(n209), .A(n261), .Y(n24) );
  AND2X1 U331 ( .A(n218), .B(n219), .Y(n25) );
  INVX1 U332 ( .A(n104), .Y(n117) );
  NAND21X1 U333 ( .B(full), .A(n226), .Y(n104) );
  OR2X1 U334 ( .A(n187), .B(n116), .Y(n118) );
  INVX1 U335 ( .A(n291), .Y(n37) );
  INVX1 U336 ( .A(n291), .Y(n38) );
  INVX1 U337 ( .A(n166), .Y(n183) );
  NAND21X1 U338 ( .B(n219), .A(n295), .Y(n166) );
  NAND21X1 U339 ( .B(n292), .A(n172), .Y(n276) );
  NAND21X1 U340 ( .B(n187), .A(n226), .Y(n227) );
  NAND21X1 U341 ( .B(n221), .A(n197), .Y(n198) );
  AO21X1 U342 ( .B(n205), .C(n221), .A(n189), .Y(n243) );
  INVX1 U343 ( .A(n135), .Y(n197) );
  NAND21X1 U344 ( .B(n292), .A(n187), .Y(n135) );
  INVX1 U345 ( .A(n292), .Y(n147) );
  AO21X1 U346 ( .B(n158), .C(n204), .A(n157), .Y(n264) );
  AO21X1 U347 ( .B(n211), .C(n204), .A(n182), .Y(n249) );
  AO21X1 U348 ( .B(n205), .C(n204), .A(n219), .Y(n235) );
  AO21X1 U349 ( .B(n205), .C(n187), .A(n219), .Y(n189) );
  INVX1 U350 ( .A(n196), .Y(n172) );
  MUX2IX1 U351 ( .D0(r_wdat[3]), .D1(prx_wdat[3]), .S(prx_psh), .Y(n359) );
  INVX1 U352 ( .A(n350), .Y(fifowdat[4]) );
  INVX1 U353 ( .A(n351), .Y(fifowdat[5]) );
  INVX1 U354 ( .A(n352), .Y(fifowdat[6]) );
  INVX1 U355 ( .A(fifowdat[2]), .Y(n65) );
  INVX1 U356 ( .A(fifowdat[0]), .Y(n55) );
  INVX1 U357 ( .A(fifowdat[0]), .Y(n56) );
  INVX1 U358 ( .A(fifowdat[1]), .Y(n59) );
  INVX1 U359 ( .A(fifowdat[1]), .Y(n60) );
  INVX1 U360 ( .A(fifowdat[2]), .Y(n63) );
  INVX1 U361 ( .A(fifowdat[2]), .Y(n64) );
  INVX1 U362 ( .A(fifowdat[7]), .Y(n53) );
  INVX1 U363 ( .A(fifowdat[0]), .Y(n57) );
  INVX1 U364 ( .A(fifowdat[1]), .Y(n61) );
  INVX1 U365 ( .A(n354), .Y(fifowdat[7]) );
  NAND21X1 U366 ( .B(n114), .A(n113), .Y(N1055) );
  AO21X1 U367 ( .B(n116), .C(n112), .A(n129), .Y(n113) );
  MUX2BXL U368 ( .D0(n111), .D1(n110), .S(n221), .Y(n114) );
  AO21X1 U369 ( .B(n147), .C(n230), .A(n126), .Y(n110) );
  AND3X1 U370 ( .A(n124), .B(n147), .C(n230), .Y(n111) );
  OAI31XL U371 ( .A(n130), .B(n157), .C(n129), .D(n128), .Y(N1059) );
  GEN2XL U372 ( .D(n127), .E(n162), .C(n129), .B(n126), .A(n125), .Y(n128) );
  AOI31X1 U373 ( .A(n124), .B(n123), .C(n211), .D(n219), .Y(n125) );
  INVX1 U374 ( .A(n122), .Y(n123) );
  NAND21X1 U375 ( .B(n361), .A(n297), .Y(n291) );
  NAND21X1 U376 ( .B(n211), .A(n232), .Y(n157) );
  NAND32X1 U377 ( .B(n212), .C(n162), .A(n209), .Y(n246) );
  NAND21X1 U378 ( .B(n611), .A(n230), .Y(n212) );
  AO2222XL U379 ( .A(r_psh), .B(full), .C(r_pop), .D(empty), .E(n365), .F(n363), .G(n362), .H(n366), .Y(ffack[1]) );
  NOR2X1 U380 ( .A(n26), .B(n363), .Y(ffack[0]) );
  AOI21X1 U381 ( .B(one), .C(r_pop), .A(n366), .Y(n26) );
  INVX1 U382 ( .A(n162), .Y(n211) );
  AOI21X1 U383 ( .B(n261), .C(n193), .A(n275), .Y(n27) );
  OAI22X1 U384 ( .A(n276), .B(n233), .C(n34), .D(n232), .Y(N743) );
  OAI31XL U385 ( .A(n611), .B(n230), .C(n291), .D(n229), .Y(N733) );
  NAND21X1 U386 ( .B(n103), .A(n614), .Y(n209) );
  NAND21X1 U387 ( .B(n299), .A(n614), .Y(n292) );
  INVX1 U388 ( .A(n232), .Y(n219) );
  NAND21X1 U389 ( .B(n146), .A(n187), .Y(n196) );
  INVX1 U390 ( .A(n193), .Y(n187) );
  INVX1 U391 ( .A(n146), .Y(n221) );
  AOI21X1 U392 ( .B(n196), .C(n232), .A(n247), .Y(n28) );
  INVX1 U393 ( .A(n105), .Y(n119) );
  NAND21X1 U394 ( .B(n193), .A(n117), .Y(n105) );
  NAND32X1 U395 ( .B(n147), .C(n146), .A(n193), .Y(n222) );
  NAND32X1 U396 ( .B(n187), .C(n292), .A(n146), .Y(n288) );
  AOI21X1 U397 ( .B(n193), .C(n232), .A(n247), .Y(n29) );
  MUX2IX1 U398 ( .D0(r_wdat[7]), .D1(prx_wdat[7]), .S(prx_psh), .Y(n354) );
  MUX2IX1 U399 ( .D0(r_wdat[4]), .D1(prx_wdat[4]), .S(prx_psh), .Y(n350) );
  MUX2IX1 U400 ( .D0(r_wdat[5]), .D1(prx_wdat[5]), .S(prx_psh), .Y(n351) );
  MUX2IX1 U401 ( .D0(r_wdat[6]), .D1(prx_wdat[6]), .S(prx_psh), .Y(n352) );
  INVX1 U402 ( .A(n355), .Y(fifowdat[0]) );
  INVX1 U403 ( .A(n356), .Y(fifowdat[1]) );
  INVX1 U404 ( .A(n357), .Y(fifowdat[2]) );
  AND2X1 U405 ( .A(n297), .B(n296), .Y(obsd) );
  INVX1 U406 ( .A(srstz), .Y(n296) );
  INVX1 U407 ( .A(n297), .Y(empty) );
  INVX1 U408 ( .A(n230), .Y(full) );
  INVX1 U409 ( .A(n300), .Y(n298) );
  MUX2X1 U410 ( .D0(fifowdat[0]), .D1(dat_7_1[0]), .S(n303), .Y(N1023) );
  MUX2X1 U411 ( .D0(fifowdat[1]), .D1(dat_7_1[1]), .S(n303), .Y(N1024) );
  MUX2X1 U412 ( .D0(fifowdat[2]), .D1(dat_7_1[2]), .S(n303), .Y(N1025) );
  MUX2X1 U413 ( .D0(fifowdat[3]), .D1(dat_7_1[3]), .S(n303), .Y(N1026) );
  MUX2X1 U414 ( .D0(fifowdat[4]), .D1(dat_7_1[4]), .S(n303), .Y(N1027) );
  MUX2X1 U415 ( .D0(fifowdat[5]), .D1(dat_7_1[5]), .S(n303), .Y(N1028) );
  MUX2X1 U416 ( .D0(fifowdat[6]), .D1(dat_7_1[6]), .S(n303), .Y(N1029) );
  MUX2X1 U417 ( .D0(fifowdat[7]), .D1(dat_7_1[7]), .S(n303), .Y(N1030) );
  NAND21XL U418 ( .B(n106), .A(ptr[4]), .Y(n162) );
  NAND2XL U419 ( .A(ptr[5]), .B(n614), .Y(n232) );
  NAND21XL U420 ( .B(n106), .A(ptr[2]), .Y(n193) );
  NAND21XL U421 ( .B(n106), .A(ptr[1]), .Y(n146) );
  MUX2IX1 U422 ( .D0(r_wdat[0]), .D1(prx_wdat[0]), .S(prx_psh), .Y(n355) );
  MUX2IX1 U423 ( .D0(r_wdat[1]), .D1(prx_wdat[1]), .S(prx_psh), .Y(n356) );
  MUX2IX1 U424 ( .D0(r_wdat[2]), .D1(prx_wdat[2]), .S(prx_psh), .Y(n357) );
  NAND32XL U425 ( .B(ptr[4]), .C(n300), .A(n299), .Y(n297) );
  NOR3XL U426 ( .A(n362), .B(n363), .C(n364), .Y(txreq) );
  INVX1 U427 ( .A(i_ccidle), .Y(n362) );
  INVX1 U428 ( .A(n364), .Y(n366) );
  NAND2X1 U429 ( .A(r_psh), .B(r_last), .Y(n364) );
  OAI211X1 U430 ( .C(n360), .D(n67), .A(n71), .B(n368), .Y(N999) );
  NAND2X1 U431 ( .A(dat_7_1[27]), .B(n358), .Y(n368) );
  OAI211X1 U432 ( .C(n360), .D(n63), .A(n75), .B(n370), .Y(N998) );
  NAND2X1 U433 ( .A(dat_7_1[26]), .B(n358), .Y(n370) );
  OAI211X1 U434 ( .C(n360), .D(n59), .A(n79), .B(n372), .Y(N997) );
  NAND2X1 U435 ( .A(dat_7_1[25]), .B(n358), .Y(n372) );
  OAI211X1 U436 ( .C(n360), .D(n55), .A(n83), .B(n374), .Y(N996) );
  NAND2X1 U437 ( .A(dat_7_1[24]), .B(n358), .Y(n374) );
  OAI211X1 U438 ( .C(n4), .D(n354), .A(n375), .B(n89), .Y(N994) );
  NAND2X1 U439 ( .A(dat_7_1[39]), .B(n353), .Y(n375) );
  OAI211X1 U440 ( .C(n4), .D(n47), .A(n377), .B(n378), .Y(N993) );
  NAND2X1 U441 ( .A(dat_7_1[38]), .B(n353), .Y(n377) );
  OAI211X1 U442 ( .C(n4), .D(n43), .A(n379), .B(n380), .Y(N992) );
  NAND2X1 U443 ( .A(dat_7_1[37]), .B(n353), .Y(n379) );
  OAI211X1 U444 ( .C(n4), .D(n39), .A(n381), .B(n382), .Y(N991) );
  NAND2X1 U445 ( .A(dat_7_1[36]), .B(n353), .Y(n381) );
  OAI211X1 U446 ( .C(n4), .D(n67), .A(n383), .B(n71), .Y(N990) );
  NAND2X1 U447 ( .A(dat_7_1[35]), .B(n353), .Y(n383) );
  OAI211X1 U448 ( .C(n4), .D(n63), .A(n384), .B(n75), .Y(N989) );
  NAND2X1 U449 ( .A(dat_7_1[34]), .B(n353), .Y(n384) );
  OAI211X1 U450 ( .C(n4), .D(n59), .A(n385), .B(n79), .Y(N988) );
  NAND2X1 U451 ( .A(dat_7_1[33]), .B(n353), .Y(n385) );
  OAI211X1 U452 ( .C(n4), .D(n55), .A(n386), .B(n83), .Y(N987) );
  NAND2X1 U453 ( .A(dat_7_1[32]), .B(n353), .Y(n386) );
  OAI211X1 U454 ( .C(n349), .D(n354), .A(n387), .B(n89), .Y(N985) );
  NAND2X1 U455 ( .A(dat_7_1[47]), .B(n348), .Y(n387) );
  OAI211X1 U456 ( .C(n349), .D(n47), .A(n388), .B(n378), .Y(N984) );
  NAND2X1 U457 ( .A(dat_7_1[46]), .B(n348), .Y(n388) );
  OAI211X1 U458 ( .C(n349), .D(n43), .A(n389), .B(n380), .Y(N983) );
  NAND2X1 U459 ( .A(dat_7_1[45]), .B(n348), .Y(n389) );
  OAI211X1 U460 ( .C(n349), .D(n39), .A(n390), .B(n382), .Y(N982) );
  NAND2X1 U461 ( .A(dat_7_1[44]), .B(n348), .Y(n390) );
  OAI211X1 U462 ( .C(n349), .D(n67), .A(n391), .B(n71), .Y(N981) );
  NAND2X1 U463 ( .A(dat_7_1[43]), .B(n348), .Y(n391) );
  OAI211X1 U464 ( .C(n349), .D(n63), .A(n392), .B(n75), .Y(N980) );
  NAND2X1 U465 ( .A(dat_7_1[42]), .B(n348), .Y(n392) );
  OAI211X1 U466 ( .C(n349), .D(n59), .A(n393), .B(n79), .Y(N979) );
  NAND2X1 U467 ( .A(dat_7_1[41]), .B(n348), .Y(n393) );
  OAI211X1 U468 ( .C(n349), .D(n55), .A(n394), .B(n83), .Y(N978) );
  NAND2X1 U469 ( .A(dat_7_1[40]), .B(n348), .Y(n394) );
  OAI211X1 U470 ( .C(n347), .D(n53), .A(n395), .B(n88), .Y(N976) );
  NAND2X1 U471 ( .A(dat_7_1[55]), .B(n346), .Y(n395) );
  OAI211X1 U472 ( .C(n347), .D(n47), .A(n396), .B(n93), .Y(N975) );
  NAND2X1 U473 ( .A(dat_7_1[54]), .B(n346), .Y(n396) );
  OAI211X1 U474 ( .C(n347), .D(n43), .A(n397), .B(n97), .Y(N974) );
  NAND2X1 U475 ( .A(dat_7_1[53]), .B(n346), .Y(n397) );
  OAI211X1 U476 ( .C(n347), .D(n39), .A(n398), .B(n101), .Y(N973) );
  NAND2X1 U477 ( .A(dat_7_1[52]), .B(n346), .Y(n398) );
  OAI211X1 U478 ( .C(n347), .D(n67), .A(n399), .B(n71), .Y(N972) );
  NAND2X1 U479 ( .A(dat_7_1[51]), .B(n346), .Y(n399) );
  OAI211X1 U480 ( .C(n347), .D(n63), .A(n400), .B(n75), .Y(N971) );
  NAND2X1 U481 ( .A(dat_7_1[50]), .B(n346), .Y(n400) );
  OAI211X1 U482 ( .C(n347), .D(n59), .A(n401), .B(n79), .Y(N970) );
  NAND2X1 U483 ( .A(dat_7_1[49]), .B(n346), .Y(n401) );
  OAI211X1 U484 ( .C(n347), .D(n55), .A(n402), .B(n83), .Y(N969) );
  NAND2X1 U485 ( .A(dat_7_1[48]), .B(n346), .Y(n402) );
  OAI211X1 U486 ( .C(n345), .D(n53), .A(n403), .B(n88), .Y(N967) );
  NAND2X1 U487 ( .A(mem_8__7_), .B(n344), .Y(n403) );
  OAI211X1 U488 ( .C(n345), .D(n47), .A(n404), .B(n93), .Y(N966) );
  NAND2X1 U489 ( .A(mem_8__6_), .B(n344), .Y(n404) );
  OAI211X1 U490 ( .C(n345), .D(n43), .A(n405), .B(n97), .Y(N965) );
  NAND2X1 U491 ( .A(mem_8__5_), .B(n344), .Y(n405) );
  OAI211X1 U492 ( .C(n345), .D(n39), .A(n406), .B(n101), .Y(N964) );
  NAND2X1 U493 ( .A(mem_8__4_), .B(n344), .Y(n406) );
  OAI211X1 U494 ( .C(n345), .D(n67), .A(n407), .B(n71), .Y(N963) );
  NAND2X1 U495 ( .A(mem_8__3_), .B(n344), .Y(n407) );
  OAI211X1 U496 ( .C(n345), .D(n63), .A(n408), .B(n75), .Y(N962) );
  NAND2X1 U497 ( .A(mem_8__2_), .B(n344), .Y(n408) );
  OAI211X1 U498 ( .C(n345), .D(n59), .A(n409), .B(n79), .Y(N961) );
  NAND2X1 U499 ( .A(mem_8__1_), .B(n344), .Y(n409) );
  OAI211X1 U500 ( .C(n345), .D(n55), .A(n410), .B(n83), .Y(N960) );
  NAND2X1 U501 ( .A(mem_8__0_), .B(n344), .Y(n410) );
  OAI211X1 U502 ( .C(n16), .D(n53), .A(n411), .B(n88), .Y(N958) );
  NAND2X1 U503 ( .A(mem_9__7_), .B(n343), .Y(n411) );
  OAI211X1 U504 ( .C(n16), .D(n47), .A(n412), .B(n93), .Y(N957) );
  NAND2X1 U505 ( .A(mem_9__6_), .B(n343), .Y(n412) );
  OAI211X1 U506 ( .C(n16), .D(n43), .A(n413), .B(n97), .Y(N956) );
  NAND2X1 U507 ( .A(mem_9__5_), .B(n343), .Y(n413) );
  OAI211X1 U508 ( .C(n16), .D(n39), .A(n414), .B(n101), .Y(N955) );
  NAND2X1 U509 ( .A(mem_9__4_), .B(n343), .Y(n414) );
  OAI211X1 U510 ( .C(n16), .D(n67), .A(n415), .B(n71), .Y(N954) );
  NAND2X1 U511 ( .A(mem_9__3_), .B(n343), .Y(n415) );
  OAI211X1 U512 ( .C(n16), .D(n63), .A(n416), .B(n75), .Y(N953) );
  NAND2X1 U513 ( .A(mem_9__2_), .B(n343), .Y(n416) );
  OAI211X1 U514 ( .C(n16), .D(n59), .A(n417), .B(n79), .Y(N952) );
  NAND2X1 U515 ( .A(mem_9__1_), .B(n343), .Y(n417) );
  OAI211X1 U516 ( .C(n16), .D(n55), .A(n418), .B(n83), .Y(N951) );
  NAND2X1 U517 ( .A(mem_9__0_), .B(n343), .Y(n418) );
  OAI211X1 U518 ( .C(n7), .D(n53), .A(n419), .B(n88), .Y(N949) );
  NAND2X1 U519 ( .A(mem_10__7_), .B(n342), .Y(n419) );
  OAI211X1 U520 ( .C(n7), .D(n47), .A(n420), .B(n93), .Y(N948) );
  NAND2X1 U521 ( .A(mem_10__6_), .B(n342), .Y(n420) );
  OAI211X1 U522 ( .C(n7), .D(n43), .A(n421), .B(n97), .Y(N947) );
  NAND2X1 U523 ( .A(mem_10__5_), .B(n342), .Y(n421) );
  OAI211X1 U524 ( .C(n7), .D(n39), .A(n422), .B(n101), .Y(N946) );
  NAND2X1 U525 ( .A(mem_10__4_), .B(n342), .Y(n422) );
  OAI211X1 U526 ( .C(n7), .D(n67), .A(n423), .B(n71), .Y(N945) );
  NAND2X1 U527 ( .A(mem_10__3_), .B(n342), .Y(n423) );
  OAI211X1 U528 ( .C(n7), .D(n63), .A(n424), .B(n75), .Y(N944) );
  NAND2X1 U529 ( .A(mem_10__2_), .B(n342), .Y(n424) );
  OAI211X1 U530 ( .C(n7), .D(n59), .A(n425), .B(n79), .Y(N943) );
  NAND2X1 U531 ( .A(mem_10__1_), .B(n342), .Y(n425) );
  OAI211X1 U532 ( .C(n7), .D(n55), .A(n426), .B(n83), .Y(N942) );
  NAND2X1 U533 ( .A(mem_10__0_), .B(n342), .Y(n426) );
  OAI211X1 U534 ( .C(n8), .D(n53), .A(n427), .B(n88), .Y(N940) );
  NAND2X1 U535 ( .A(mem_11__7_), .B(n341), .Y(n427) );
  OAI211X1 U536 ( .C(n8), .D(n47), .A(n428), .B(n93), .Y(N939) );
  NAND2X1 U537 ( .A(mem_11__6_), .B(n341), .Y(n428) );
  OAI211X1 U538 ( .C(n8), .D(n43), .A(n429), .B(n97), .Y(N938) );
  NAND2X1 U539 ( .A(mem_11__5_), .B(n341), .Y(n429) );
  OAI211X1 U540 ( .C(n8), .D(n39), .A(n430), .B(n101), .Y(N937) );
  NAND2X1 U541 ( .A(mem_11__4_), .B(n341), .Y(n430) );
  OAI211X1 U542 ( .C(n8), .D(n67), .A(n431), .B(n71), .Y(N936) );
  NAND2X1 U543 ( .A(mem_11__3_), .B(n341), .Y(n431) );
  OAI211X1 U544 ( .C(n8), .D(n63), .A(n432), .B(n75), .Y(N935) );
  NAND2X1 U545 ( .A(mem_11__2_), .B(n341), .Y(n432) );
  OAI211X1 U546 ( .C(n8), .D(n59), .A(n433), .B(n79), .Y(N934) );
  NAND2X1 U547 ( .A(mem_11__1_), .B(n341), .Y(n433) );
  OAI211X1 U548 ( .C(n8), .D(n55), .A(n434), .B(n83), .Y(N933) );
  NAND2X1 U549 ( .A(mem_11__0_), .B(n341), .Y(n434) );
  OAI211X1 U550 ( .C(n340), .D(n53), .A(n435), .B(n88), .Y(N931) );
  NAND2X1 U551 ( .A(mem_12__7_), .B(n339), .Y(n435) );
  OAI211X1 U552 ( .C(n340), .D(n47), .A(n436), .B(n93), .Y(N930) );
  NAND2X1 U553 ( .A(mem_12__6_), .B(n339), .Y(n436) );
  OAI211X1 U554 ( .C(n340), .D(n43), .A(n437), .B(n97), .Y(N929) );
  NAND2X1 U555 ( .A(mem_12__5_), .B(n339), .Y(n437) );
  OAI211X1 U556 ( .C(n340), .D(n39), .A(n438), .B(n101), .Y(N928) );
  NAND2X1 U557 ( .A(mem_12__4_), .B(n339), .Y(n438) );
  OAI211X1 U558 ( .C(n340), .D(n67), .A(n439), .B(n72), .Y(N927) );
  NAND2X1 U559 ( .A(mem_12__3_), .B(n339), .Y(n439) );
  OAI211X1 U560 ( .C(n340), .D(n63), .A(n440), .B(n76), .Y(N926) );
  NAND2X1 U561 ( .A(mem_12__2_), .B(n339), .Y(n440) );
  OAI211X1 U562 ( .C(n340), .D(n59), .A(n441), .B(n80), .Y(N925) );
  NAND2X1 U563 ( .A(mem_12__1_), .B(n339), .Y(n441) );
  OAI211X1 U564 ( .C(n340), .D(n55), .A(n442), .B(n83), .Y(N924) );
  NAND2X1 U565 ( .A(mem_12__0_), .B(n339), .Y(n442) );
  OAI211X1 U566 ( .C(n5), .D(n53), .A(n443), .B(n88), .Y(N922) );
  NAND2X1 U567 ( .A(mem_13__7_), .B(n338), .Y(n443) );
  OAI211X1 U568 ( .C(n5), .D(n47), .A(n444), .B(n93), .Y(N921) );
  NAND2X1 U569 ( .A(mem_13__6_), .B(n338), .Y(n444) );
  OAI211X1 U570 ( .C(n5), .D(n43), .A(n445), .B(n97), .Y(N920) );
  NAND2X1 U571 ( .A(mem_13__5_), .B(n338), .Y(n445) );
  OAI211X1 U572 ( .C(n5), .D(n39), .A(n446), .B(n101), .Y(N919) );
  NAND2X1 U573 ( .A(mem_13__4_), .B(n338), .Y(n446) );
  OAI211X1 U574 ( .C(n5), .D(n67), .A(n447), .B(n72), .Y(N918) );
  NAND2X1 U575 ( .A(mem_13__3_), .B(n338), .Y(n447) );
  OAI211X1 U576 ( .C(n5), .D(n63), .A(n448), .B(n76), .Y(N917) );
  NAND2X1 U577 ( .A(mem_13__2_), .B(n338), .Y(n448) );
  OAI211X1 U578 ( .C(n5), .D(n59), .A(n449), .B(n80), .Y(N916) );
  NAND2X1 U579 ( .A(mem_13__1_), .B(n338), .Y(n449) );
  OAI211X1 U580 ( .C(n5), .D(n55), .A(n450), .B(n83), .Y(N915) );
  NAND2X1 U581 ( .A(mem_13__0_), .B(n338), .Y(n450) );
  OAI211X1 U582 ( .C(n337), .D(n53), .A(n451), .B(n88), .Y(N913) );
  NAND2X1 U583 ( .A(mem_14__7_), .B(n336), .Y(n451) );
  OAI211X1 U584 ( .C(n337), .D(n47), .A(n452), .B(n93), .Y(N912) );
  NAND2X1 U585 ( .A(mem_14__6_), .B(n336), .Y(n452) );
  OAI211X1 U586 ( .C(n337), .D(n43), .A(n453), .B(n97), .Y(N911) );
  NAND2X1 U587 ( .A(mem_14__5_), .B(n336), .Y(n453) );
  OAI211X1 U588 ( .C(n337), .D(n39), .A(n454), .B(n101), .Y(N910) );
  NAND2X1 U589 ( .A(mem_14__4_), .B(n336), .Y(n454) );
  OAI211X1 U590 ( .C(n337), .D(n68), .A(n455), .B(n72), .Y(N909) );
  NAND2X1 U591 ( .A(mem_14__3_), .B(n336), .Y(n455) );
  OAI211X1 U592 ( .C(n337), .D(n64), .A(n456), .B(n76), .Y(N908) );
  NAND2X1 U593 ( .A(mem_14__2_), .B(n336), .Y(n456) );
  OAI211X1 U594 ( .C(n337), .D(n60), .A(n457), .B(n80), .Y(N907) );
  NAND2X1 U595 ( .A(mem_14__1_), .B(n336), .Y(n457) );
  OAI211X1 U596 ( .C(n337), .D(n56), .A(n458), .B(n84), .Y(N906) );
  NAND2X1 U597 ( .A(mem_14__0_), .B(n336), .Y(n458) );
  OAI211X1 U598 ( .C(n335), .D(n53), .A(n459), .B(n88), .Y(N904) );
  NAND2X1 U599 ( .A(mem_15__7_), .B(n334), .Y(n459) );
  OAI211X1 U600 ( .C(n335), .D(n48), .A(n460), .B(n93), .Y(N903) );
  NAND2X1 U601 ( .A(mem_15__6_), .B(n334), .Y(n460) );
  OAI211X1 U602 ( .C(n335), .D(n44), .A(n461), .B(n97), .Y(N902) );
  NAND2X1 U603 ( .A(mem_15__5_), .B(n334), .Y(n461) );
  OAI211X1 U604 ( .C(n335), .D(n40), .A(n462), .B(n101), .Y(N901) );
  NAND2X1 U605 ( .A(mem_15__4_), .B(n334), .Y(n462) );
  OAI211X1 U606 ( .C(n335), .D(n68), .A(n463), .B(n72), .Y(N900) );
  NAND2X1 U607 ( .A(mem_15__3_), .B(n334), .Y(n463) );
  OAI211X1 U608 ( .C(n335), .D(n64), .A(n464), .B(n76), .Y(N899) );
  NAND2X1 U609 ( .A(mem_15__2_), .B(n334), .Y(n464) );
  OAI211X1 U610 ( .C(n335), .D(n60), .A(n465), .B(n80), .Y(N898) );
  NAND2X1 U611 ( .A(mem_15__1_), .B(n334), .Y(n465) );
  OAI211X1 U612 ( .C(n335), .D(n56), .A(n466), .B(n84), .Y(N897) );
  NAND2X1 U613 ( .A(mem_15__0_), .B(n334), .Y(n466) );
  OAI211X1 U614 ( .C(n333), .D(n53), .A(n467), .B(n88), .Y(N895) );
  NAND2X1 U615 ( .A(mem_16__7_), .B(n332), .Y(n467) );
  OAI211X1 U616 ( .C(n333), .D(n48), .A(n468), .B(n93), .Y(N894) );
  NAND2X1 U617 ( .A(mem_16__6_), .B(n332), .Y(n468) );
  OAI211X1 U618 ( .C(n333), .D(n44), .A(n469), .B(n97), .Y(N893) );
  NAND2X1 U619 ( .A(mem_16__5_), .B(n332), .Y(n469) );
  OAI211X1 U620 ( .C(n333), .D(n40), .A(n470), .B(n101), .Y(N892) );
  NAND2X1 U621 ( .A(mem_16__4_), .B(n332), .Y(n470) );
  OAI211X1 U622 ( .C(n333), .D(n68), .A(n471), .B(n72), .Y(N891) );
  NAND2X1 U623 ( .A(mem_16__3_), .B(n332), .Y(n471) );
  OAI211X1 U624 ( .C(n333), .D(n64), .A(n472), .B(n76), .Y(N890) );
  NAND2X1 U625 ( .A(mem_16__2_), .B(n332), .Y(n472) );
  OAI211X1 U626 ( .C(n333), .D(n60), .A(n473), .B(n80), .Y(N889) );
  NAND2X1 U627 ( .A(mem_16__1_), .B(n332), .Y(n473) );
  OAI211X1 U628 ( .C(n333), .D(n56), .A(n474), .B(n84), .Y(N888) );
  NAND2X1 U629 ( .A(mem_16__0_), .B(n332), .Y(n474) );
  OAI211X1 U630 ( .C(n331), .D(n52), .A(n475), .B(n87), .Y(N886) );
  NAND2X1 U631 ( .A(mem_17__7_), .B(n330), .Y(n475) );
  OAI211X1 U632 ( .C(n331), .D(n48), .A(n476), .B(n92), .Y(N885) );
  NAND2X1 U633 ( .A(mem_17__6_), .B(n330), .Y(n476) );
  OAI211X1 U634 ( .C(n331), .D(n44), .A(n477), .B(n96), .Y(N884) );
  NAND2X1 U635 ( .A(mem_17__5_), .B(n330), .Y(n477) );
  OAI211X1 U636 ( .C(n331), .D(n40), .A(n478), .B(n100), .Y(N883) );
  NAND2X1 U637 ( .A(mem_17__4_), .B(n330), .Y(n478) );
  OAI211X1 U638 ( .C(n331), .D(n68), .A(n479), .B(n72), .Y(N882) );
  NAND2X1 U639 ( .A(mem_17__3_), .B(n330), .Y(n479) );
  OAI211X1 U640 ( .C(n331), .D(n64), .A(n480), .B(n76), .Y(N881) );
  NAND2X1 U641 ( .A(mem_17__2_), .B(n330), .Y(n480) );
  OAI211X1 U642 ( .C(n331), .D(n60), .A(n481), .B(n80), .Y(N880) );
  NAND2X1 U643 ( .A(mem_17__1_), .B(n330), .Y(n481) );
  OAI211X1 U644 ( .C(n331), .D(n56), .A(n482), .B(n84), .Y(N879) );
  NAND2X1 U645 ( .A(mem_17__0_), .B(n330), .Y(n482) );
  OAI211X1 U646 ( .C(n9), .D(n52), .A(n483), .B(n87), .Y(N877) );
  NAND2X1 U647 ( .A(mem_18__7_), .B(n329), .Y(n483) );
  OAI211X1 U648 ( .C(n9), .D(n48), .A(n484), .B(n92), .Y(N876) );
  NAND2X1 U649 ( .A(mem_18__6_), .B(n329), .Y(n484) );
  OAI211X1 U650 ( .C(n9), .D(n44), .A(n485), .B(n96), .Y(N875) );
  NAND2X1 U651 ( .A(mem_18__5_), .B(n329), .Y(n485) );
  OAI211X1 U652 ( .C(n9), .D(n40), .A(n486), .B(n100), .Y(N874) );
  NAND2X1 U653 ( .A(mem_18__4_), .B(n329), .Y(n486) );
  OAI211X1 U654 ( .C(n9), .D(n68), .A(n487), .B(n72), .Y(N873) );
  NAND2X1 U655 ( .A(mem_18__3_), .B(n329), .Y(n487) );
  OAI211X1 U656 ( .C(n9), .D(n64), .A(n488), .B(n76), .Y(N872) );
  NAND2X1 U657 ( .A(mem_18__2_), .B(n329), .Y(n488) );
  OAI211X1 U658 ( .C(n9), .D(n60), .A(n489), .B(n80), .Y(N871) );
  NAND2X1 U659 ( .A(mem_18__1_), .B(n329), .Y(n489) );
  OAI211X1 U660 ( .C(n9), .D(n56), .A(n490), .B(n84), .Y(N870) );
  NAND2X1 U661 ( .A(mem_18__0_), .B(n329), .Y(n490) );
  OAI211X1 U662 ( .C(n10), .D(n52), .A(n491), .B(n87), .Y(N868) );
  NAND2X1 U663 ( .A(mem_19__7_), .B(n328), .Y(n491) );
  OAI211X1 U664 ( .C(n10), .D(n48), .A(n492), .B(n92), .Y(N867) );
  NAND2X1 U665 ( .A(mem_19__6_), .B(n328), .Y(n492) );
  OAI211X1 U666 ( .C(n10), .D(n44), .A(n493), .B(n96), .Y(N866) );
  NAND2X1 U667 ( .A(mem_19__5_), .B(n328), .Y(n493) );
  OAI211X1 U668 ( .C(n10), .D(n40), .A(n494), .B(n100), .Y(N865) );
  NAND2X1 U669 ( .A(mem_19__4_), .B(n328), .Y(n494) );
  OAI211X1 U670 ( .C(n10), .D(n68), .A(n495), .B(n72), .Y(N864) );
  NAND2X1 U671 ( .A(mem_19__3_), .B(n328), .Y(n495) );
  OAI211X1 U672 ( .C(n10), .D(n64), .A(n496), .B(n76), .Y(N863) );
  NAND2X1 U673 ( .A(mem_19__2_), .B(n328), .Y(n496) );
  OAI211X1 U674 ( .C(n10), .D(n60), .A(n497), .B(n80), .Y(N862) );
  NAND2X1 U675 ( .A(mem_19__1_), .B(n328), .Y(n497) );
  OAI211X1 U676 ( .C(n10), .D(n56), .A(n498), .B(n84), .Y(N861) );
  NAND2X1 U677 ( .A(mem_19__0_), .B(n328), .Y(n498) );
  OAI211X1 U678 ( .C(n11), .D(n52), .A(n499), .B(n87), .Y(N859) );
  NAND2X1 U679 ( .A(mem_20__7_), .B(n327), .Y(n499) );
  OAI211X1 U680 ( .C(n11), .D(n48), .A(n500), .B(n92), .Y(N858) );
  NAND2X1 U681 ( .A(mem_20__6_), .B(n327), .Y(n500) );
  OAI211X1 U682 ( .C(n11), .D(n44), .A(n501), .B(n96), .Y(N857) );
  NAND2X1 U683 ( .A(mem_20__5_), .B(n327), .Y(n501) );
  OAI211X1 U684 ( .C(n11), .D(n40), .A(n502), .B(n100), .Y(N856) );
  NAND2X1 U685 ( .A(mem_20__4_), .B(n327), .Y(n502) );
  OAI211X1 U686 ( .C(n11), .D(n68), .A(n503), .B(n72), .Y(N855) );
  NAND2X1 U687 ( .A(mem_20__3_), .B(n327), .Y(n503) );
  OAI211X1 U688 ( .C(n11), .D(n64), .A(n504), .B(n76), .Y(N854) );
  NAND2X1 U689 ( .A(mem_20__2_), .B(n327), .Y(n504) );
  OAI211X1 U690 ( .C(n11), .D(n60), .A(n505), .B(n80), .Y(N853) );
  NAND2X1 U691 ( .A(mem_20__1_), .B(n327), .Y(n505) );
  OAI211X1 U692 ( .C(n11), .D(n56), .A(n506), .B(n84), .Y(N852) );
  NAND2X1 U693 ( .A(mem_20__0_), .B(n327), .Y(n506) );
  OAI211X1 U694 ( .C(n12), .D(n52), .A(n507), .B(n87), .Y(N850) );
  NAND2X1 U695 ( .A(mem_21__7_), .B(n326), .Y(n507) );
  OAI211X1 U696 ( .C(n12), .D(n48), .A(n508), .B(n92), .Y(N849) );
  NAND2X1 U697 ( .A(mem_21__6_), .B(n326), .Y(n508) );
  OAI211X1 U698 ( .C(n12), .D(n44), .A(n509), .B(n96), .Y(N848) );
  NAND2X1 U699 ( .A(mem_21__5_), .B(n326), .Y(n509) );
  OAI211X1 U700 ( .C(n12), .D(n40), .A(n510), .B(n100), .Y(N847) );
  NAND2X1 U701 ( .A(mem_21__4_), .B(n326), .Y(n510) );
  OAI211X1 U702 ( .C(n12), .D(n68), .A(n511), .B(n72), .Y(N846) );
  NAND2X1 U703 ( .A(mem_21__3_), .B(n326), .Y(n511) );
  OAI211X1 U704 ( .C(n12), .D(n64), .A(n512), .B(n76), .Y(N845) );
  NAND2X1 U705 ( .A(mem_21__2_), .B(n326), .Y(n512) );
  OAI211X1 U706 ( .C(n12), .D(n60), .A(n513), .B(n80), .Y(N844) );
  NAND2X1 U707 ( .A(mem_21__1_), .B(n326), .Y(n513) );
  OAI211X1 U708 ( .C(n12), .D(n56), .A(n514), .B(n84), .Y(N843) );
  NAND2X1 U709 ( .A(mem_21__0_), .B(n326), .Y(n514) );
  OAI211X1 U710 ( .C(n13), .D(n52), .A(n515), .B(n87), .Y(N841) );
  NAND2X1 U711 ( .A(mem_22__7_), .B(n325), .Y(n515) );
  OAI211X1 U712 ( .C(n13), .D(n48), .A(n516), .B(n92), .Y(N840) );
  NAND2X1 U713 ( .A(mem_22__6_), .B(n325), .Y(n516) );
  OAI211X1 U714 ( .C(n13), .D(n44), .A(n517), .B(n96), .Y(N839) );
  NAND2X1 U715 ( .A(mem_22__5_), .B(n325), .Y(n517) );
  OAI211X1 U716 ( .C(n13), .D(n40), .A(n518), .B(n100), .Y(N838) );
  NAND2X1 U717 ( .A(mem_22__4_), .B(n325), .Y(n518) );
  OAI211X1 U718 ( .C(n13), .D(n68), .A(n519), .B(n73), .Y(N837) );
  NAND2X1 U719 ( .A(mem_22__3_), .B(n325), .Y(n519) );
  OAI211X1 U720 ( .C(n13), .D(n64), .A(n520), .B(n77), .Y(N836) );
  NAND2X1 U721 ( .A(mem_22__2_), .B(n325), .Y(n520) );
  OAI211X1 U722 ( .C(n13), .D(n60), .A(n521), .B(n81), .Y(N835) );
  NAND2X1 U723 ( .A(mem_22__1_), .B(n325), .Y(n521) );
  OAI211X1 U724 ( .C(n13), .D(n56), .A(n522), .B(n84), .Y(N834) );
  NAND2X1 U725 ( .A(mem_22__0_), .B(n325), .Y(n522) );
  OAI211X1 U726 ( .C(n324), .D(n52), .A(n523), .B(n87), .Y(N832) );
  NAND2X1 U727 ( .A(mem_23__7_), .B(n323), .Y(n523) );
  OAI211X1 U728 ( .C(n324), .D(n48), .A(n524), .B(n92), .Y(N831) );
  NAND2X1 U729 ( .A(mem_23__6_), .B(n323), .Y(n524) );
  OAI211X1 U730 ( .C(n324), .D(n44), .A(n525), .B(n96), .Y(N830) );
  NAND2X1 U731 ( .A(mem_23__5_), .B(n323), .Y(n525) );
  OAI211X1 U732 ( .C(n324), .D(n40), .A(n526), .B(n100), .Y(N829) );
  NAND2X1 U733 ( .A(mem_23__4_), .B(n323), .Y(n526) );
  OAI211X1 U734 ( .C(n324), .D(n68), .A(n527), .B(n73), .Y(N828) );
  NAND2X1 U735 ( .A(mem_23__3_), .B(n323), .Y(n527) );
  OAI211X1 U736 ( .C(n324), .D(n64), .A(n528), .B(n77), .Y(N827) );
  NAND2X1 U737 ( .A(mem_23__2_), .B(n323), .Y(n528) );
  OAI211X1 U738 ( .C(n324), .D(n60), .A(n529), .B(n81), .Y(N826) );
  NAND2X1 U739 ( .A(mem_23__1_), .B(n323), .Y(n529) );
  OAI211X1 U740 ( .C(n324), .D(n56), .A(n530), .B(n84), .Y(N825) );
  NAND2X1 U741 ( .A(mem_23__0_), .B(n323), .Y(n530) );
  OAI211X1 U742 ( .C(n322), .D(n52), .A(n531), .B(n87), .Y(N823) );
  NAND2X1 U743 ( .A(mem_24__7_), .B(n321), .Y(n531) );
  OAI211X1 U744 ( .C(n322), .D(n48), .A(n532), .B(n92), .Y(N822) );
  NAND2X1 U745 ( .A(mem_24__6_), .B(n321), .Y(n532) );
  OAI211X1 U746 ( .C(n322), .D(n44), .A(n533), .B(n96), .Y(N821) );
  NAND2X1 U747 ( .A(mem_24__5_), .B(n321), .Y(n533) );
  OAI211X1 U748 ( .C(n322), .D(n40), .A(n534), .B(n100), .Y(N820) );
  NAND2X1 U749 ( .A(mem_24__4_), .B(n321), .Y(n534) );
  OAI211X1 U750 ( .C(n322), .D(n69), .A(n535), .B(n73), .Y(N819) );
  NAND2X1 U751 ( .A(mem_24__3_), .B(n321), .Y(n535) );
  OAI211X1 U752 ( .C(n322), .D(n357), .A(n536), .B(n77), .Y(N818) );
  NAND2X1 U753 ( .A(mem_24__2_), .B(n321), .Y(n536) );
  OAI211X1 U754 ( .C(n322), .D(n61), .A(n537), .B(n81), .Y(N817) );
  NAND2X1 U755 ( .A(mem_24__1_), .B(n321), .Y(n537) );
  OAI211X1 U756 ( .C(n322), .D(n57), .A(n538), .B(n85), .Y(N816) );
  NAND2X1 U757 ( .A(mem_24__0_), .B(n321), .Y(n538) );
  OAI211X1 U758 ( .C(n320), .D(n52), .A(n539), .B(n87), .Y(N814) );
  NAND2X1 U759 ( .A(mem_25__7_), .B(n319), .Y(n539) );
  OAI211X1 U760 ( .C(n320), .D(n49), .A(n540), .B(n92), .Y(N813) );
  NAND2X1 U761 ( .A(mem_25__6_), .B(n319), .Y(n540) );
  OAI211X1 U762 ( .C(n320), .D(n45), .A(n541), .B(n96), .Y(N812) );
  NAND2X1 U763 ( .A(mem_25__5_), .B(n319), .Y(n541) );
  OAI211X1 U764 ( .C(n320), .D(n41), .A(n542), .B(n100), .Y(N811) );
  NAND2X1 U765 ( .A(mem_25__4_), .B(n319), .Y(n542) );
  OAI211X1 U766 ( .C(n320), .D(n69), .A(n543), .B(n73), .Y(N810) );
  NAND2X1 U767 ( .A(mem_25__3_), .B(n319), .Y(n543) );
  OAI211X1 U768 ( .C(n320), .D(n357), .A(n544), .B(n77), .Y(N809) );
  NAND2X1 U769 ( .A(mem_25__2_), .B(n319), .Y(n544) );
  OAI211X1 U770 ( .C(n320), .D(n61), .A(n545), .B(n81), .Y(N808) );
  NAND2X1 U771 ( .A(mem_25__1_), .B(n319), .Y(n545) );
  OAI211X1 U772 ( .C(n320), .D(n57), .A(n546), .B(n85), .Y(N807) );
  NAND2X1 U773 ( .A(mem_25__0_), .B(n319), .Y(n546) );
  OAI211X1 U774 ( .C(n14), .D(n52), .A(n547), .B(n87), .Y(N805) );
  NAND2X1 U775 ( .A(mem_26__7_), .B(n318), .Y(n547) );
  OAI211X1 U776 ( .C(n14), .D(n49), .A(n548), .B(n92), .Y(N804) );
  NAND2X1 U777 ( .A(mem_26__6_), .B(n318), .Y(n548) );
  OAI211X1 U778 ( .C(n14), .D(n45), .A(n549), .B(n96), .Y(N803) );
  NAND2X1 U779 ( .A(mem_26__5_), .B(n318), .Y(n549) );
  OAI211X1 U780 ( .C(n14), .D(n41), .A(n550), .B(n100), .Y(N802) );
  NAND2X1 U781 ( .A(mem_26__4_), .B(n318), .Y(n550) );
  OAI211X1 U782 ( .C(n14), .D(n69), .A(n551), .B(n73), .Y(N801) );
  NAND2X1 U783 ( .A(mem_26__3_), .B(n318), .Y(n551) );
  OAI211X1 U784 ( .C(n14), .D(n357), .A(n552), .B(n77), .Y(N800) );
  NAND2X1 U785 ( .A(mem_26__2_), .B(n318), .Y(n552) );
  OAI211X1 U786 ( .C(n14), .D(n61), .A(n553), .B(n81), .Y(N799) );
  NAND2X1 U787 ( .A(mem_26__1_), .B(n318), .Y(n553) );
  OAI211X1 U788 ( .C(n14), .D(n57), .A(n554), .B(n85), .Y(N798) );
  NAND2X1 U789 ( .A(mem_26__0_), .B(n318), .Y(n554) );
  OAI211X1 U790 ( .C(n6), .D(n51), .A(n555), .B(n89), .Y(N796) );
  NAND2X1 U791 ( .A(mem_27__7_), .B(n317), .Y(n555) );
  OAI211X1 U792 ( .C(n6), .D(n352), .A(n556), .B(n91), .Y(N795) );
  NAND2X1 U793 ( .A(mem_27__6_), .B(n317), .Y(n556) );
  OAI211X1 U794 ( .C(n6), .D(n45), .A(n557), .B(n95), .Y(N794) );
  NAND2X1 U795 ( .A(mem_27__5_), .B(n317), .Y(n557) );
  OAI211X1 U796 ( .C(n6), .D(n41), .A(n558), .B(n99), .Y(N793) );
  NAND2X1 U797 ( .A(mem_27__4_), .B(n317), .Y(n558) );
  OAI211X1 U798 ( .C(n6), .D(n69), .A(n559), .B(n73), .Y(N792) );
  NAND2X1 U799 ( .A(mem_27__3_), .B(n317), .Y(n559) );
  OAI211X1 U800 ( .C(n6), .D(n357), .A(n560), .B(n77), .Y(N791) );
  NAND2X1 U801 ( .A(mem_27__2_), .B(n317), .Y(n560) );
  OAI211X1 U802 ( .C(n6), .D(n61), .A(n561), .B(n81), .Y(N790) );
  NAND2X1 U803 ( .A(mem_27__1_), .B(n317), .Y(n561) );
  OAI211X1 U804 ( .C(n6), .D(n57), .A(n562), .B(n85), .Y(N789) );
  NAND2X1 U805 ( .A(mem_27__0_), .B(n317), .Y(n562) );
  OAI211X1 U806 ( .C(n316), .D(n51), .A(n563), .B(n89), .Y(N787) );
  NAND2X1 U807 ( .A(mem_28__7_), .B(n315), .Y(n563) );
  OAI211X1 U808 ( .C(n316), .D(n352), .A(n564), .B(n91), .Y(N786) );
  NAND2X1 U809 ( .A(mem_28__6_), .B(n315), .Y(n564) );
  OAI211X1 U810 ( .C(n316), .D(n45), .A(n565), .B(n95), .Y(N785) );
  NAND2X1 U811 ( .A(mem_28__5_), .B(n315), .Y(n565) );
  OAI211X1 U812 ( .C(n316), .D(n41), .A(n566), .B(n99), .Y(N784) );
  NAND2X1 U813 ( .A(mem_28__4_), .B(n315), .Y(n566) );
  OAI211X1 U814 ( .C(n316), .D(n69), .A(n567), .B(n73), .Y(N783) );
  NAND2X1 U815 ( .A(mem_28__3_), .B(n315), .Y(n567) );
  OAI211X1 U816 ( .C(n316), .D(n357), .A(n568), .B(n77), .Y(N782) );
  NAND2X1 U817 ( .A(mem_28__2_), .B(n315), .Y(n568) );
  OAI211X1 U818 ( .C(n316), .D(n61), .A(n569), .B(n81), .Y(N781) );
  NAND2X1 U819 ( .A(mem_28__1_), .B(n315), .Y(n569) );
  OAI211X1 U820 ( .C(n316), .D(n57), .A(n570), .B(n85), .Y(N780) );
  NAND2X1 U821 ( .A(mem_28__0_), .B(n315), .Y(n570) );
  OAI211X1 U822 ( .C(n15), .D(n51), .A(n571), .B(n89), .Y(N778) );
  NAND2X1 U823 ( .A(mem_29__7_), .B(n314), .Y(n571) );
  OAI211X1 U824 ( .C(n15), .D(n352), .A(n572), .B(n91), .Y(N777) );
  NAND2X1 U825 ( .A(mem_29__6_), .B(n314), .Y(n572) );
  OAI211X1 U826 ( .C(n15), .D(n45), .A(n573), .B(n95), .Y(N776) );
  NAND2X1 U827 ( .A(mem_29__5_), .B(n314), .Y(n573) );
  OAI211X1 U828 ( .C(n15), .D(n41), .A(n574), .B(n99), .Y(N775) );
  NAND2X1 U829 ( .A(mem_29__4_), .B(n314), .Y(n574) );
  OAI211X1 U830 ( .C(n15), .D(n69), .A(n575), .B(n73), .Y(N774) );
  NAND2X1 U831 ( .A(mem_29__3_), .B(n314), .Y(n575) );
  OAI211X1 U832 ( .C(n15), .D(n357), .A(n576), .B(n77), .Y(N773) );
  NAND2X1 U833 ( .A(mem_29__2_), .B(n314), .Y(n576) );
  OAI211X1 U834 ( .C(n15), .D(n61), .A(n577), .B(n81), .Y(N772) );
  NAND2X1 U835 ( .A(mem_29__1_), .B(n314), .Y(n577) );
  OAI211X1 U836 ( .C(n15), .D(n57), .A(n578), .B(n85), .Y(N771) );
  NAND2X1 U837 ( .A(mem_29__0_), .B(n314), .Y(n578) );
  OAI211X1 U838 ( .C(n313), .D(n51), .A(n579), .B(n89), .Y(N769) );
  NAND2X1 U839 ( .A(mem_30__7_), .B(n312), .Y(n579) );
  OAI211X1 U840 ( .C(n313), .D(n352), .A(n580), .B(n91), .Y(N768) );
  NAND2X1 U841 ( .A(mem_30__6_), .B(n312), .Y(n580) );
  OAI211X1 U842 ( .C(n313), .D(n45), .A(n581), .B(n95), .Y(N767) );
  NAND2X1 U843 ( .A(mem_30__5_), .B(n312), .Y(n581) );
  OAI211X1 U844 ( .C(n313), .D(n41), .A(n582), .B(n99), .Y(N766) );
  NAND2X1 U845 ( .A(mem_30__4_), .B(n312), .Y(n582) );
  OAI211X1 U846 ( .C(n313), .D(n69), .A(n583), .B(n73), .Y(N765) );
  NAND2X1 U847 ( .A(mem_30__3_), .B(n312), .Y(n583) );
  OAI211X1 U848 ( .C(n313), .D(n65), .A(n584), .B(n77), .Y(N764) );
  NAND2X1 U849 ( .A(mem_30__2_), .B(n312), .Y(n584) );
  OAI211X1 U850 ( .C(n313), .D(n61), .A(n585), .B(n81), .Y(N763) );
  NAND2X1 U851 ( .A(mem_30__1_), .B(n312), .Y(n585) );
  OAI211X1 U852 ( .C(n313), .D(n57), .A(n586), .B(n85), .Y(N762) );
  NAND2X1 U853 ( .A(mem_30__0_), .B(n312), .Y(n586) );
  OAI211X1 U854 ( .C(n311), .D(n51), .A(n587), .B(n89), .Y(N760) );
  NAND2X1 U855 ( .A(mem_31__7_), .B(n310), .Y(n587) );
  OAI211X1 U856 ( .C(n311), .D(n352), .A(n588), .B(n91), .Y(N759) );
  NAND2X1 U857 ( .A(mem_31__6_), .B(n310), .Y(n588) );
  OAI211X1 U858 ( .C(n311), .D(n45), .A(n589), .B(n95), .Y(N758) );
  NAND2X1 U859 ( .A(mem_31__5_), .B(n310), .Y(n589) );
  OAI211X1 U860 ( .C(n311), .D(n41), .A(n590), .B(n99), .Y(N757) );
  NAND2X1 U861 ( .A(mem_31__4_), .B(n310), .Y(n590) );
  OAI211X1 U862 ( .C(n311), .D(n69), .A(n591), .B(n73), .Y(N756) );
  NAND2X1 U863 ( .A(mem_31__3_), .B(n310), .Y(n591) );
  OAI211X1 U864 ( .C(n311), .D(n65), .A(n592), .B(n77), .Y(N755) );
  NAND2X1 U865 ( .A(mem_31__2_), .B(n310), .Y(n592) );
  OAI211X1 U866 ( .C(n311), .D(n61), .A(n593), .B(n81), .Y(N754) );
  NAND2X1 U867 ( .A(mem_31__1_), .B(n310), .Y(n593) );
  OAI211X1 U868 ( .C(n311), .D(n57), .A(n594), .B(n85), .Y(N753) );
  NAND2X1 U869 ( .A(mem_31__0_), .B(n310), .Y(n594) );
  OAI211X1 U870 ( .C(n309), .D(n51), .A(n595), .B(n89), .Y(N751) );
  NAND2X1 U871 ( .A(mem_32__7_), .B(n308), .Y(n595) );
  OAI211X1 U872 ( .C(n309), .D(n352), .A(n596), .B(n91), .Y(N750) );
  NAND2X1 U873 ( .A(mem_32__6_), .B(n308), .Y(n596) );
  OAI211X1 U874 ( .C(n309), .D(n45), .A(n597), .B(n95), .Y(N749) );
  NAND2X1 U875 ( .A(mem_32__5_), .B(n308), .Y(n597) );
  OAI211X1 U876 ( .C(n309), .D(n41), .A(n598), .B(n99), .Y(N748) );
  NAND2X1 U877 ( .A(mem_32__4_), .B(n308), .Y(n598) );
  OAI211X1 U878 ( .C(n309), .D(n69), .A(n599), .B(n367), .Y(N747) );
  NAND2X1 U879 ( .A(mem_32__3_), .B(n308), .Y(n599) );
  OAI211X1 U880 ( .C(n309), .D(n357), .A(n600), .B(n369), .Y(N746) );
  NAND2X1 U881 ( .A(mem_32__2_), .B(n308), .Y(n600) );
  OAI211X1 U882 ( .C(n309), .D(n61), .A(n601), .B(n371), .Y(N745) );
  NAND2X1 U883 ( .A(mem_32__1_), .B(n308), .Y(n601) );
  OAI211X1 U884 ( .C(n309), .D(n57), .A(n602), .B(n85), .Y(N744) );
  NAND2X1 U885 ( .A(mem_32__0_), .B(n308), .Y(n602) );
  OAI211X1 U886 ( .C(n17), .D(n51), .A(n603), .B(n89), .Y(N742) );
  NAND2X1 U887 ( .A(mem_33__7_), .B(n307), .Y(n603) );
  OAI211X1 U888 ( .C(n17), .D(n352), .A(n604), .B(n91), .Y(N741) );
  NAND2X1 U889 ( .A(mem_33__6_), .B(n307), .Y(n604) );
  OAI211X1 U890 ( .C(n17), .D(n45), .A(n605), .B(n95), .Y(N740) );
  NAND2X1 U891 ( .A(mem_33__5_), .B(n307), .Y(n605) );
  OAI211X1 U892 ( .C(n17), .D(n41), .A(n606), .B(n99), .Y(N739) );
  NAND2X1 U893 ( .A(mem_33__4_), .B(n307), .Y(n606) );
  OAI211X1 U894 ( .C(n17), .D(n69), .A(n607), .B(n367), .Y(N738) );
  NAND2X1 U895 ( .A(mem_33__3_), .B(n307), .Y(n607) );
  OAI211X1 U896 ( .C(n17), .D(n357), .A(n608), .B(n369), .Y(N737) );
  NAND2X1 U897 ( .A(mem_33__2_), .B(n307), .Y(n608) );
  OAI211X1 U898 ( .C(n17), .D(n61), .A(n609), .B(n371), .Y(N736) );
  NAND2X1 U899 ( .A(mem_33__1_), .B(n307), .Y(n609) );
  OAI211X1 U900 ( .C(n17), .D(n57), .A(n610), .B(n85), .Y(N735) );
  NAND2X1 U901 ( .A(mem_33__0_), .B(n307), .Y(n610) );
  NAND2X1 U902 ( .A(n613), .B(n614), .Y(N1053) );
  XNOR2XL U903 ( .A(n611), .B(n361), .Y(n613) );
  OAI211X1 U904 ( .C(n306), .D(n51), .A(n615), .B(n89), .Y(N1021) );
  NAND2X1 U905 ( .A(dat_7_1[15]), .B(n305), .Y(n615) );
  OAI211X1 U906 ( .C(n306), .D(n352), .A(n616), .B(n91), .Y(N1020) );
  NAND2X1 U907 ( .A(dat_7_1[14]), .B(n305), .Y(n616) );
  OAI211X1 U908 ( .C(n306), .D(n45), .A(n617), .B(n95), .Y(N1019) );
  NAND2X1 U909 ( .A(dat_7_1[13]), .B(n305), .Y(n617) );
  OAI211X1 U910 ( .C(n306), .D(n41), .A(n618), .B(n99), .Y(N1018) );
  NAND2X1 U911 ( .A(dat_7_1[12]), .B(n305), .Y(n618) );
  OAI211X1 U912 ( .C(n306), .D(n359), .A(n619), .B(n71), .Y(N1017) );
  NAND2X1 U913 ( .A(dat_7_1[11]), .B(n305), .Y(n619) );
  OAI211X1 U914 ( .C(n306), .D(n65), .A(n620), .B(n75), .Y(N1016) );
  NAND2X1 U915 ( .A(dat_7_1[10]), .B(n305), .Y(n620) );
  OAI211X1 U916 ( .C(n306), .D(n356), .A(n621), .B(n79), .Y(N1015) );
  NAND2X1 U917 ( .A(dat_7_1[9]), .B(n305), .Y(n621) );
  OAI211X1 U918 ( .C(n306), .D(n355), .A(n622), .B(n373), .Y(N1014) );
  NAND2X1 U919 ( .A(dat_7_1[8]), .B(n305), .Y(n622) );
  OAI211X1 U920 ( .C(n3), .D(n51), .A(n623), .B(n376), .Y(N1012) );
  NAND2X1 U921 ( .A(dat_7_1[23]), .B(n304), .Y(n623) );
  OAI211X1 U922 ( .C(n3), .D(n49), .A(n624), .B(n91), .Y(N1011) );
  NAND2X1 U923 ( .A(dat_7_1[22]), .B(n304), .Y(n624) );
  OAI211X1 U924 ( .C(n3), .D(n351), .A(n625), .B(n95), .Y(N1010) );
  NAND2X1 U925 ( .A(dat_7_1[21]), .B(n304), .Y(n625) );
  OAI211X1 U926 ( .C(n3), .D(n350), .A(n626), .B(n99), .Y(N1009) );
  NAND2X1 U927 ( .A(dat_7_1[20]), .B(n304), .Y(n626) );
  OAI211X1 U928 ( .C(n3), .D(n359), .A(n71), .B(n627), .Y(N1008) );
  NAND2X1 U929 ( .A(dat_7_1[19]), .B(n304), .Y(n627) );
  OAI211X1 U930 ( .C(n3), .D(n65), .A(n75), .B(n628), .Y(N1007) );
  NAND2X1 U931 ( .A(dat_7_1[18]), .B(n304), .Y(n628) );
  OAI211X1 U932 ( .C(n3), .D(n356), .A(n79), .B(n629), .Y(N1006) );
  NAND2X1 U933 ( .A(dat_7_1[17]), .B(n304), .Y(n629) );
  OAI211X1 U934 ( .C(n3), .D(n355), .A(n630), .B(n373), .Y(N1005) );
  NAND2X1 U935 ( .A(dat_7_1[16]), .B(n304), .Y(n630) );
  OAI211X1 U936 ( .C(n360), .D(n51), .A(n376), .B(n631), .Y(N1003) );
  NAND2X1 U937 ( .A(dat_7_1[31]), .B(n358), .Y(n631) );
  OAI211X1 U938 ( .C(n360), .D(n49), .A(n91), .B(n632), .Y(N1002) );
  NAND2X1 U939 ( .A(dat_7_1[30]), .B(n358), .Y(n632) );
  OAI211X1 U940 ( .C(n360), .D(n351), .A(n95), .B(n633), .Y(N1001) );
  NAND2X1 U941 ( .A(dat_7_1[29]), .B(n358), .Y(n633) );
  OAI211X1 U942 ( .C(n360), .D(n350), .A(n634), .B(n99), .Y(N1000) );
  NAND2X1 U943 ( .A(dat_7_1[28]), .B(n358), .Y(n634) );
  OAI21X1 U944 ( .B(n363), .C(n635), .A(n636), .Y(n612) );
  INVX1 U945 ( .A(fifopsh), .Y(n611) );
  OAI21X1 U946 ( .B(n363), .C(n637), .A(n638), .Y(fifopsh) );
  NOR2X1 U947 ( .A(r_unlock), .B(ps_locked), .Y(n363) );
  NOR43XL U948 ( .B(n636), .C(n614), .D(n638), .A(n639), .Y(ps_locked) );
  AOI21X1 U949 ( .B(i_lockena), .C(n365), .A(locked), .Y(n639) );
  NAND2X1 U950 ( .A(n637), .B(n635), .Y(n365) );
  INVX1 U951 ( .A(r_pop), .Y(n635) );
  INVX1 U952 ( .A(r_psh), .Y(n637) );
  INVX1 U953 ( .A(prx_psh), .Y(n638) );
  NOR21XL U954 ( .B(srstz), .A(r_fiforst), .Y(n614) );
  INVX1 U955 ( .A(ptx_pop), .Y(n636) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phycrc_a0 ( crc32_3_0, rx_good, i_shfidat, i_start, i_shfi4, i_shfo4, 
        clk );
  output [3:0] crc32_3_0;
  input [3:0] i_shfidat;
  input i_start, i_shfi4, i_shfo4, clk;
  output rx_good;
  wire   N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         net10623, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n56, n57, n58, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n55, n59, n118, n120, n121,
         n122, n123, n125, n126, n127, n128;
  wire   [31:0] crc32_r;

  SNPS_CLOCK_GATE_HIGH_phycrc_a0 clk_gate_crc32_r_reg ( .CLK(clk), .EN(N188), 
        .ENCLK(net10623), .TE(1'b0) );
  DFFQX1 crc32_r_reg_26_ ( .D(N215), .C(net10623), .Q(crc32_r[26]) );
  DFFQX1 crc32_r_reg_16_ ( .D(N205), .C(net10623), .Q(crc32_r[16]) );
  DFFQX1 crc32_r_reg_27_ ( .D(N216), .C(net10623), .Q(crc32_r[27]) );
  DFFQX1 crc32_r_reg_17_ ( .D(N206), .C(net10623), .Q(crc32_r[17]) );
  DFFQX1 crc32_r_reg_11_ ( .D(N200), .C(net10623), .Q(crc32_r[11]) );
  DFFQX1 crc32_r_reg_15_ ( .D(N204), .C(net10623), .Q(crc32_r[15]) );
  DFFQX1 crc32_r_reg_0_ ( .D(N189), .C(net10623), .Q(crc32_r[0]) );
  DFFQX1 crc32_r_reg_4_ ( .D(N193), .C(net10623), .Q(crc32_r[4]) );
  DFFQX1 crc32_r_reg_8_ ( .D(N197), .C(net10623), .Q(crc32_r[8]) );
  DFFQX1 crc32_r_reg_5_ ( .D(N194), .C(net10623), .Q(crc32_r[5]) );
  DFFQX1 crc32_r_reg_1_ ( .D(N190), .C(net10623), .Q(crc32_r[1]) );
  DFFQX1 crc32_r_reg_10_ ( .D(N199), .C(net10623), .Q(crc32_r[10]) );
  DFFQX1 crc32_r_reg_3_ ( .D(N192), .C(net10623), .Q(crc32_r[3]) );
  DFFQX1 crc32_r_reg_6_ ( .D(N195), .C(net10623), .Q(crc32_r[6]) );
  DFFQX1 crc32_r_reg_12_ ( .D(N201), .C(net10623), .Q(crc32_r[12]) );
  DFFQX1 crc32_r_reg_14_ ( .D(N203), .C(net10623), .Q(crc32_r[14]) );
  DFFQX1 crc32_r_reg_18_ ( .D(N207), .C(net10623), .Q(crc32_r[18]) );
  DFFQX1 crc32_r_reg_25_ ( .D(N214), .C(net10623), .Q(crc32_r[25]) );
  DFFQX1 crc32_r_reg_24_ ( .D(N213), .C(net10623), .Q(crc32_r[24]) );
  DFFQX1 crc32_r_reg_9_ ( .D(N198), .C(net10623), .Q(crc32_r[9]) );
  DFFQX1 crc32_r_reg_21_ ( .D(N210), .C(net10623), .Q(crc32_r[21]) );
  DFFQX1 crc32_r_reg_20_ ( .D(N209), .C(net10623), .Q(crc32_r[20]) );
  DFFQX1 crc32_r_reg_7_ ( .D(N196), .C(net10623), .Q(crc32_r[7]) );
  DFFQX1 crc32_r_reg_22_ ( .D(N211), .C(net10623), .Q(crc32_r[22]) );
  DFFQX1 crc32_r_reg_13_ ( .D(N202), .C(net10623), .Q(crc32_r[13]) );
  DFFQX1 crc32_r_reg_2_ ( .D(N191), .C(net10623), .Q(crc32_r[2]) );
  DFFQX1 crc32_r_reg_23_ ( .D(N212), .C(net10623), .Q(crc32_r[23]) );
  DFFQX1 crc32_r_reg_28_ ( .D(N217), .C(net10623), .Q(crc32_r[28]) );
  DFFQX1 crc32_r_reg_29_ ( .D(N218), .C(net10623), .Q(crc32_r[29]) );
  DFFQX1 crc32_r_reg_19_ ( .D(N208), .C(net10623), .Q(crc32_r[19]) );
  DFFQX1 crc32_r_reg_31_ ( .D(N220), .C(net10623), .Q(crc32_r[31]) );
  DFFQX1 crc32_r_reg_30_ ( .D(N219), .C(net10623), .Q(crc32_r[30]) );
  OR2X1 U3 ( .A(n19), .B(i_start), .Y(n1) );
  INVXL U4 ( .A(n1), .Y(n2) );
  INVXL U5 ( .A(n1), .Y(n3) );
  NOR2X1 U6 ( .A(n15), .B(n78), .Y(n4) );
  INVX1 U7 ( .A(n16), .Y(n5) );
  XNOR2XL U8 ( .A(i_shfidat[3]), .B(n117), .Y(n69) );
  INVX1 U9 ( .A(n78), .Y(n6) );
  INVX1 U10 ( .A(n15), .Y(n7) );
  INVX1 U11 ( .A(n75), .Y(n8) );
  XNOR2XL U12 ( .A(i_shfidat[1]), .B(n114), .Y(n48) );
  XNOR2XL U13 ( .A(i_shfidat[2]), .B(n116), .Y(n53) );
  NAND2X1 U14 ( .A(n11), .B(n57), .Y(N188) );
  NAND2X1 U15 ( .A(i_shfo4), .B(n13), .Y(n10) );
  NAND2X1 U16 ( .A(i_shfo4), .B(n11), .Y(n57) );
  INVX1 U17 ( .A(n9), .Y(n11) );
  INVX1 U18 ( .A(n9), .Y(n13) );
  NAND21X1 U19 ( .B(n11), .A(n2), .Y(n43) );
  INVX1 U20 ( .A(n75), .Y(n14) );
  INVX1 U21 ( .A(n9), .Y(n12) );
  NOR2X1 U22 ( .A(n18), .B(i_start), .Y(n65) );
  INVX1 U23 ( .A(i_start), .Y(n15) );
  NOR2X1 U24 ( .A(i_shfi4), .B(n11), .Y(n75) );
  NOR2X1 U25 ( .A(n11), .B(i_start), .Y(n49) );
  OAI21X1 U26 ( .B(n13), .C(n112), .A(n8), .Y(N191) );
  XNOR2XL U27 ( .A(n16), .B(n113), .Y(n112) );
  XNOR2XL U28 ( .A(n17), .B(n18), .Y(n113) );
  OAI21X1 U29 ( .B(n13), .C(n109), .A(n8), .Y(N192) );
  XNOR2XL U30 ( .A(n17), .B(n110), .Y(n109) );
  XNOR2XL U31 ( .A(n18), .B(n6), .Y(n110) );
  NOR2X1 U32 ( .A(n75), .B(n60), .Y(n45) );
  OR2X1 U33 ( .A(i_start), .B(i_shfi4), .Y(n9) );
  OAI21X1 U34 ( .B(n13), .C(n115), .A(n8), .Y(N190) );
  XNOR2XL U35 ( .A(n16), .B(n17), .Y(n115) );
  AOI21X1 U36 ( .B(n17), .C(n7), .A(n75), .Y(n52) );
  AOI21X1 U37 ( .B(n16), .C(n7), .A(n75), .Y(n72) );
  NOR2X1 U38 ( .A(n75), .B(n66), .Y(n47) );
  OAI21X1 U39 ( .B(n13), .C(n16), .A(n8), .Y(N189) );
  INVX1 U40 ( .A(n48), .Y(n18) );
  INVX1 U41 ( .A(n78), .Y(n19) );
  NOR2X1 U42 ( .A(n15), .B(n78), .Y(n60) );
  NOR2X1 U43 ( .A(n15), .B(n48), .Y(n66) );
  INVX1 U44 ( .A(n53), .Y(n17) );
  INVX1 U45 ( .A(n69), .Y(n16) );
  OAI21X1 U46 ( .B(n13), .C(n53), .A(n57), .Y(n54) );
  OAI21X1 U47 ( .B(n13), .C(n48), .A(n57), .Y(n50) );
  OAI21X1 U48 ( .B(n13), .C(n69), .A(n10), .Y(n73) );
  OA21X1 U49 ( .B(n13), .C(n78), .A(n57), .Y(n44) );
  NOR4XL U50 ( .A(n20), .B(n120), .C(n32), .D(n23), .Y(n38) );
  NOR4XL U51 ( .A(n121), .B(n55), .C(n122), .D(n31), .Y(n37) );
  NOR4XL U52 ( .A(n21), .B(n26), .C(n127), .D(n22), .Y(n35) );
  NOR2X1 U53 ( .A(crc32_r[30]), .B(i_start), .Y(n114) );
  XNOR2XL U54 ( .A(i_shfidat[0]), .B(n111), .Y(n78) );
  NOR2X1 U55 ( .A(crc32_r[31]), .B(i_start), .Y(n111) );
  OAI221X1 U56 ( .A(n12), .B(n87), .C(n57), .D(n128), .E(n14), .Y(N200) );
  XNOR2XL U57 ( .A(n88), .B(n69), .Y(n87) );
  XNOR2XL U58 ( .A(n89), .B(n53), .Y(n88) );
  AOI221XL U59 ( .A(crc32_r[7]), .B(n19), .C(n2), .D(n128), .E(n60), .Y(n89)
         );
  OAI221X1 U60 ( .A(n12), .B(n103), .C(n31), .D(n10), .E(n14), .Y(N194) );
  XNOR2XL U61 ( .A(n104), .B(n69), .Y(n103) );
  XNOR2XL U62 ( .A(n105), .B(n53), .Y(n104) );
  AOI221XL U63 ( .A(crc32_r[1]), .B(n19), .C(n2), .D(n31), .E(n4), .Y(n105) );
  OAI221X1 U64 ( .A(n12), .B(n84), .C(n22), .D(n10), .E(n14), .Y(N201) );
  XNOR2XL U65 ( .A(n85), .B(n69), .Y(n84) );
  XNOR2XL U66 ( .A(n86), .B(n53), .Y(n85) );
  AOI221XL U67 ( .A(crc32_r[8]), .B(n18), .C(n65), .D(n22), .E(n66), .Y(n86)
         );
  OAI221X1 U68 ( .A(n12), .B(n95), .C(n21), .D(n57), .E(n14), .Y(N197) );
  XNOR2XL U69 ( .A(n96), .B(n69), .Y(n95) );
  XNOR2XL U70 ( .A(n97), .B(n53), .Y(n96) );
  AOI221XL U71 ( .A(crc32_r[4]), .B(n19), .C(n3), .D(n21), .E(n60), .Y(n97) );
  OAI221X1 U72 ( .A(n12), .B(n98), .C(n125), .D(n10), .E(n14), .Y(N196) );
  XNOR2XL U73 ( .A(n99), .B(n69), .Y(n98) );
  XNOR2XL U74 ( .A(n100), .B(n48), .Y(n99) );
  AOI221XL U75 ( .A(crc32_r[3]), .B(n19), .C(n2), .D(n125), .E(n60), .Y(n100)
         );
  OAI221X1 U76 ( .A(n12), .B(n90), .C(n127), .D(n57), .E(n14), .Y(N199) );
  XNOR2XL U77 ( .A(n91), .B(n69), .Y(n90) );
  XNOR2XL U78 ( .A(n92), .B(n48), .Y(n91) );
  AOI221XL U79 ( .A(crc32_r[6]), .B(n19), .C(n2), .D(n127), .E(n4), .Y(n92) );
  OAI221X1 U80 ( .A(n12), .B(n106), .C(n20), .D(n10), .E(n14), .Y(N193) );
  XNOR2XL U81 ( .A(n107), .B(n69), .Y(n106) );
  XNOR2XL U82 ( .A(n108), .B(n48), .Y(n107) );
  AOI221XL U83 ( .A(crc32_r[0]), .B(n19), .C(n3), .D(n20), .E(n60), .Y(n108)
         );
  OAI221X1 U84 ( .A(n12), .B(n56), .C(n123), .D(n10), .E(n14), .Y(N215) );
  XNOR2XL U85 ( .A(n58), .B(n16), .Y(n56) );
  AOI221XL U86 ( .A(crc32_r[22]), .B(n6), .C(n3), .D(n123), .E(n4), .Y(n58) );
  INVX1 U87 ( .A(crc32_r[22]), .Y(n123) );
  OAI221X1 U88 ( .A(n11), .B(n79), .C(n120), .D(n57), .E(n14), .Y(N203) );
  XNOR2XL U89 ( .A(n80), .B(n18), .Y(n79) );
  AOI221XL U90 ( .A(crc32_r[10]), .B(n19), .C(n3), .D(n120), .E(n4), .Y(n80)
         );
  OAI221X1 U91 ( .A(n12), .B(n93), .C(n26), .D(n10), .E(n14), .Y(N198) );
  XNOR2XL U92 ( .A(n94), .B(n17), .Y(n93) );
  AOI221XL U93 ( .A(crc32_r[5]), .B(n18), .C(n65), .D(n26), .E(n66), .Y(n94)
         );
  OAI221X1 U94 ( .A(n12), .B(n101), .C(n10), .D(n126), .E(n8), .Y(N195) );
  XNOR2XL U95 ( .A(n102), .B(n17), .Y(n101) );
  AOI221XL U96 ( .A(crc32_r[2]), .B(n18), .C(n65), .D(n126), .E(n66), .Y(n102)
         );
  INVX1 U97 ( .A(crc32_r[2]), .Y(n126) );
  OAI221X1 U98 ( .A(n11), .B(n61), .C(n57), .D(n29), .E(n8), .Y(N214) );
  XNOR2XL U99 ( .A(n62), .B(n18), .Y(n61) );
  AOI221XL U100 ( .A(crc32_r[21]), .B(n19), .C(n2), .D(n29), .E(n60), .Y(n62)
         );
  INVX1 U101 ( .A(crc32_r[21]), .Y(n29) );
  OAI221X1 U102 ( .A(n11), .B(n81), .C(n10), .D(n27), .E(n8), .Y(N202) );
  XNOR2XL U103 ( .A(n82), .B(n53), .Y(n81) );
  XNOR2XL U104 ( .A(n83), .B(n48), .Y(n82) );
  AOI221XL U105 ( .A(crc32_r[9]), .B(n19), .C(n3), .D(n27), .E(n4), .Y(n83) );
  OAI221X1 U106 ( .A(n11), .B(n63), .C(n10), .D(n24), .E(n8), .Y(N213) );
  XNOR2XL U107 ( .A(n64), .B(n17), .Y(n63) );
  AOI221XL U108 ( .A(crc32_r[20]), .B(n18), .C(n65), .D(n24), .E(n66), .Y(n64)
         );
  INVX1 U109 ( .A(crc32_r[20]), .Y(n24) );
  NOR2X1 U110 ( .A(crc32_r[28]), .B(i_start), .Y(n117) );
  NOR2X1 U111 ( .A(crc32_r[29]), .B(i_start), .Y(n116) );
  OAI221X1 U112 ( .A(n11), .B(n67), .C(n57), .D(n59), .E(n8), .Y(N212) );
  INVX1 U113 ( .A(crc32_r[19]), .Y(n59) );
  XNOR2XL U114 ( .A(n68), .B(n69), .Y(n67) );
  XNOR2XL U115 ( .A(n70), .B(n53), .Y(n68) );
  NAND2X1 U116 ( .A(n71), .B(n72), .Y(N211) );
  AOI32X1 U117 ( .A(n49), .B(n122), .C(n5), .D(crc32_r[18]), .E(n73), .Y(n71)
         );
  NAND2X1 U118 ( .A(n74), .B(n47), .Y(N207) );
  AOI32X1 U119 ( .A(n48), .B(n121), .C(n49), .D(crc32_r[14]), .E(n50), .Y(n74)
         );
  NAND2X1 U120 ( .A(n51), .B(n52), .Y(N216) );
  AOI32X1 U121 ( .A(n49), .B(n118), .C(n53), .D(crc32_r[23]), .E(n54), .Y(n51)
         );
  INVX1 U122 ( .A(crc32_r[23]), .Y(n118) );
  NAND2X1 U123 ( .A(n76), .B(n52), .Y(N206) );
  AOI32X1 U124 ( .A(n49), .B(n28), .C(n53), .D(crc32_r[13]), .E(n54), .Y(n76)
         );
  INVX1 U125 ( .A(crc32_r[13]), .Y(n28) );
  NAND2X1 U126 ( .A(n46), .B(n47), .Y(N217) );
  AOI32X1 U127 ( .A(n48), .B(n25), .C(n49), .D(crc32_r[24]), .E(n50), .Y(n46)
         );
  INVX1 U128 ( .A(crc32_r[24]), .Y(n25) );
  NAND2X1 U129 ( .A(n77), .B(n72), .Y(N205) );
  AOI32X1 U130 ( .A(n49), .B(n23), .C(n5), .D(crc32_r[12]), .E(n73), .Y(n77)
         );
  OAI221X1 U131 ( .A(crc32_r[15]), .B(n43), .C(n44), .D(n55), .E(n45), .Y(N208) );
  OAI221X1 U132 ( .A(crc32_r[11]), .B(n43), .C(n44), .D(n32), .E(n45), .Y(N204) );
  OAI221X1 U133 ( .A(crc32_r[25]), .B(n43), .C(n44), .D(n30), .E(n45), .Y(N218) );
  INVX1 U134 ( .A(crc32_r[25]), .Y(n30) );
  NOR2X1 U135 ( .A(crc32_r[19]), .B(i_start), .Y(n70) );
  OAI21BBX1 U136 ( .A(N188), .B(crc32_r[26]), .C(n15), .Y(N219) );
  OAI21BBX1 U137 ( .A(N188), .B(crc32_r[27]), .C(n15), .Y(N220) );
  OAI21BBX1 U138 ( .A(N188), .B(crc32_r[17]), .C(n15), .Y(N210) );
  OAI21BBX1 U139 ( .A(N188), .B(crc32_r[16]), .C(n15), .Y(N209) );
  NOR2X1 U140 ( .A(n33), .B(n34), .Y(rx_good) );
  NAND4X1 U141 ( .A(n35), .B(n36), .C(n37), .D(n38), .Y(n34) );
  NAND4X1 U142 ( .A(n39), .B(n40), .C(n41), .D(n42), .Y(n33) );
  NOR43XL U143 ( .B(crc32_r[24]), .C(crc32_r[25]), .D(crc32_r[26]), .A(n125), 
        .Y(n36) );
  NOR4XL U144 ( .A(crc32_r[9]), .B(crc32_r[7]), .C(crc32_r[2]), .D(crc32_r[29]), .Y(n42) );
  NOR4XL U145 ( .A(crc32_r[28]), .B(crc32_r[27]), .C(crc32_r[23]), .D(
        crc32_r[22]), .Y(n41) );
  NOR4XL U146 ( .A(crc32_r[21]), .B(crc32_r[20]), .C(crc32_r[19]), .D(
        crc32_r[17]), .Y(n40) );
  NOR4XL U147 ( .A(crc32_r[16]), .B(crc32_r[13]), .C(crc32_3_0[1]), .D(
        crc32_3_0[0]), .Y(n39) );
  INVX1 U148 ( .A(crc32_r[30]), .Y(crc32_3_0[1]) );
  INVX1 U149 ( .A(crc32_r[31]), .Y(crc32_3_0[0]) );
  INVX1 U150 ( .A(crc32_r[3]), .Y(n125) );
  INVX1 U151 ( .A(crc32_r[6]), .Y(n127) );
  INVX1 U152 ( .A(crc32_r[1]), .Y(n31) );
  INVX1 U153 ( .A(crc32_r[8]), .Y(n22) );
  INVX1 U154 ( .A(crc32_r[10]), .Y(n120) );
  INVX1 U155 ( .A(crc32_r[5]), .Y(n26) );
  INVX1 U156 ( .A(crc32_r[4]), .Y(n21) );
  INVX1 U157 ( .A(crc32_r[0]), .Y(n20) );
  INVX1 U158 ( .A(crc32_r[18]), .Y(n122) );
  INVX1 U159 ( .A(crc32_r[12]), .Y(n23) );
  INVX1 U160 ( .A(crc32_r[14]), .Y(n121) );
  INVX1 U161 ( .A(crc32_r[11]), .Y(n32) );
  INVX1 U162 ( .A(crc32_r[15]), .Y(n55) );
  INVX1 U163 ( .A(crc32_r[28]), .Y(crc32_3_0[3]) );
  INVX1 U164 ( .A(crc32_r[29]), .Y(crc32_3_0[2]) );
  INVX1 U165 ( .A(crc32_r[7]), .Y(n128) );
  INVX1 U166 ( .A(crc32_r[9]), .Y(n27) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phycrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phytx_a0 ( r_txnumk, r_txendk, r_txshrt, r_txauto, prx_cccnt, ptx_txact, 
        ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, i_rdat, i_txreq, i_one, 
        ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4, ptx_crcsidat, ptx_fsm, 
        pcc_crc30, clk, srstz );
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [1:0] prx_cccnt;
  input [7:0] i_rdat;
  output [3:0] ptx_crcsidat;
  output [2:0] ptx_fsm;
  input [3:0] pcc_crc30;
  input r_txendk, r_txshrt, i_txreq, i_one, clk, srstz;
  output ptx_txact, ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, ptx_crcstart,
         ptx_crcshfi4, ptx_crcshfo4;
  wire   n294, hinib, N251, N253, N254, N255, N268, N270, N271, N272, N273,
         N297, N298, N299, net10645, net10651, n237, n238, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293;
  wire   [4:0] bytcnt;
  wire   [3:0] bitcnt;

  SNPS_CLOCK_GATE_HIGH_phytx_a0_0 clk_gate_bitcnt_reg ( .CLK(clk), .EN(N251), 
        .ENCLK(net10645), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phytx_a0_1 clk_gate_bytcnt_reg ( .CLK(clk), .EN(N268), 
        .ENCLK(net10651), .TE(1'b0) );
  DFFQX1 ptx_cc_reg ( .D(n238), .C(clk), .Q(ptx_cc) );
  DFFQX1 bitcnt_reg_1_ ( .D(N253), .C(net10645), .Q(bitcnt[1]) );
  DFFQX1 bitcnt_reg_2_ ( .D(N254), .C(net10645), .Q(bitcnt[2]) );
  DFFQX1 bitcnt_reg_0_ ( .D(n276), .C(net10645), .Q(bitcnt[0]) );
  DFFQX1 bitcnt_reg_3_ ( .D(N255), .C(net10645), .Q(bitcnt[3]) );
  DFFQX1 bytcnt_reg_4_ ( .D(N273), .C(net10651), .Q(bytcnt[4]) );
  DFFQX1 bytcnt_reg_1_ ( .D(N270), .C(net10651), .Q(bytcnt[1]) );
  DFFQX1 cs_txph_reg_0_ ( .D(N297), .C(clk), .Q(ptx_fsm[0]) );
  DFFQX1 cs_txph_reg_2_ ( .D(N299), .C(clk), .Q(ptx_fsm[2]) );
  DFFQX1 cs_txph_reg_1_ ( .D(N298), .C(clk), .Q(ptx_fsm[1]) );
  DFFQX1 hinib_reg ( .D(n237), .C(net10645), .Q(hinib) );
  DFFQX1 bytcnt_reg_0_ ( .D(n275), .C(net10651), .Q(bytcnt[0]) );
  DFFQX1 bytcnt_reg_3_ ( .D(N272), .C(net10651), .Q(bytcnt[3]) );
  DFFQX1 bytcnt_reg_2_ ( .D(N271), .C(net10651), .Q(bytcnt[2]) );
  NAND2X2 U3 ( .A(n11), .B(n27), .Y(n28) );
  NAND2X4 U4 ( .A(n17), .B(n62), .Y(n63) );
  INVX2 U5 ( .A(i_rdat[0]), .Y(n20) );
  INVX2 U6 ( .A(i_rdat[4]), .Y(n226) );
  MUX2X2 U7 ( .D0(n83), .D1(n86), .S(hinib), .Y(n143) );
  NAND2X2 U8 ( .A(n20), .B(n21), .Y(n3) );
  AND3X2 U9 ( .A(n266), .B(n49), .C(n259), .Y(n53) );
  NAND2X2 U10 ( .A(n2), .B(n3), .Y(n157) );
  NAND21X2 U11 ( .B(r_txnumk[1]), .A(bytcnt[1]), .Y(n259) );
  INVX2 U12 ( .A(i_rdat[1]), .Y(n83) );
  INVX3 U13 ( .A(i_rdat[5]), .Y(n86) );
  NAND2X2 U14 ( .A(n170), .B(n157), .Y(n58) );
  MUX2X2 U15 ( .D0(n81), .D1(n66), .S(hinib), .Y(n15) );
  NAND21X2 U16 ( .B(n70), .A(n69), .Y(n126) );
  INVX2 U17 ( .A(r_txnumk[0]), .Y(n47) );
  NOR2X2 U18 ( .A(n133), .B(n269), .Y(n22) );
  INVX3 U19 ( .A(n126), .Y(n133) );
  INVX2 U20 ( .A(i_one), .Y(n73) );
  AND4X2 U21 ( .A(n23), .B(n65), .C(bitcnt[2]), .D(n35), .Y(n136) );
  INVX1 U22 ( .A(ptx_fsm[0]), .Y(n111) );
  NAND21X1 U23 ( .B(n294), .A(prx_cccnt[0]), .Y(n251) );
  INVX1 U24 ( .A(ptx_fsm[2]), .Y(n101) );
  INVX1 U25 ( .A(ptx_fsm[1]), .Y(n90) );
  INVX1 U26 ( .A(bitcnt[3]), .Y(n65) );
  NOR21XL U27 ( .B(bitcnt[3]), .A(n244), .Y(n64) );
  MUX2IX2 U28 ( .D0(n15), .D1(n58), .S(n37), .Y(n59) );
  INVX1 U29 ( .A(i_rdat[3]), .Y(n81) );
  NAND2X1 U30 ( .A(n226), .B(n1), .Y(n2) );
  INVXL U31 ( .A(n21), .Y(n1) );
  NAND2X1 U32 ( .A(i_rdat[6]), .B(n4), .Y(n5) );
  NAND2X1 U33 ( .A(i_rdat[2]), .B(n21), .Y(n6) );
  NAND2X1 U34 ( .A(n5), .B(n6), .Y(n37) );
  INVX1 U35 ( .A(n21), .Y(n4) );
  INVX3 U36 ( .A(n206), .Y(n26) );
  NAND2X1 U37 ( .A(n81), .B(n21), .Y(n12) );
  INVX1 U38 ( .A(n269), .Y(n18) );
  INVX1 U39 ( .A(n143), .Y(ptx_crcsidat[1]) );
  XNOR2XL U40 ( .A(n243), .B(bitcnt[0]), .Y(n7) );
  INVX1 U41 ( .A(n21), .Y(n8) );
  INVX1 U42 ( .A(hinib), .Y(n21) );
  INVX1 U43 ( .A(n267), .Y(n9) );
  BUFXL U44 ( .A(n37), .Y(ptx_crcsidat[2]) );
  NAND21X2 U45 ( .B(n172), .A(n63), .Y(n11) );
  NAND21X2 U46 ( .B(n172), .A(n63), .Y(n206) );
  NAND2X1 U47 ( .A(n66), .B(hinib), .Y(n13) );
  NAND2X1 U48 ( .A(n12), .B(n13), .Y(n170) );
  NAND43XL U49 ( .B(n47), .C(n48), .D(n50), .A(r_txnumk[2]), .Y(n46) );
  INVX1 U50 ( .A(r_txnumk[3]), .Y(n50) );
  INVXL U51 ( .A(n15), .Y(ptx_crcsidat[3]) );
  AND2X1 U52 ( .A(n28), .B(n29), .Y(n23) );
  INVXL U53 ( .A(n77), .Y(n70) );
  NAND31XL U54 ( .C(n79), .A(n226), .B(n86), .Y(n67) );
  XOR2X1 U55 ( .A(n11), .B(n244), .Y(n35) );
  INVXL U56 ( .A(n19), .Y(n75) );
  AND2X2 U57 ( .A(n28), .B(n29), .Y(n14) );
  INVXL U58 ( .A(n17), .Y(n267) );
  OAI22X1 U59 ( .A(bytcnt[2]), .B(n51), .C(bytcnt[3]), .D(n50), .Y(n52) );
  INVXL U60 ( .A(n26), .Y(n16) );
  AND2X2 U61 ( .A(n57), .B(n18), .Y(n17) );
  MUX2XL U62 ( .D0(n147), .D1(n146), .S(n9), .Y(n148) );
  AO21XL U63 ( .B(n194), .C(n17), .A(n193), .Y(n195) );
  NAND21XL U64 ( .B(n17), .A(n145), .Y(n183) );
  NAND21X2 U65 ( .B(n251), .A(n136), .Y(n256) );
  NOR5X2 U66 ( .A(n77), .B(n260), .C(bytcnt[3]), .D(bytcnt[2]), .E(bytcnt[4]), 
        .Y(n19) );
  INVXL U67 ( .A(i_rdat[0]), .Y(n167) );
  INVXL U68 ( .A(n273), .Y(n93) );
  INVXL U69 ( .A(n14), .Y(n203) );
  INVXL U70 ( .A(i_rdat[2]), .Y(n149) );
  NAND2X2 U71 ( .A(n26), .B(bitcnt[1]), .Y(n29) );
  NAND21X2 U72 ( .B(n156), .A(n61), .Y(n62) );
  NAND21X2 U73 ( .B(ptx_crcsidat[1]), .A(n59), .Y(n61) );
  BUFXL U74 ( .A(n81), .Y(n24) );
  NAND21XL U75 ( .B(i_rdat[6]), .A(n66), .Y(n79) );
  OAI221XL U76 ( .A(n183), .B(n213), .C(n227), .D(n149), .E(n148), .Y(n160) );
  NAND32XL U77 ( .B(i_txreq), .C(n126), .A(n125), .Y(n127) );
  NAND21XL U78 ( .B(n256), .A(n158), .Y(n125) );
  INVXL U79 ( .A(n256), .Y(n263) );
  NAND21X1 U80 ( .B(n22), .A(n273), .Y(ptx_fifopop) );
  XNOR2X1 U81 ( .A(n11), .B(bitcnt[2]), .Y(n36) );
  INVXL U82 ( .A(n294), .Y(ptx_txact) );
  NOR2XL U83 ( .A(ptx_fsm[2]), .B(n135), .Y(n294) );
  INVX2 U84 ( .A(i_rdat[7]), .Y(n66) );
  INVXL U85 ( .A(bitcnt[1]), .Y(n27) );
  NAND21X2 U86 ( .B(n251), .A(n134), .Y(n77) );
  NAND21XL U87 ( .B(n156), .A(n67), .Y(n68) );
  NAND6X1 U88 ( .A(n19), .B(n167), .C(n85), .D(n84), .E(i_one), .F(n86), .Y(
        n273) );
  AND4XL U89 ( .A(n149), .B(n83), .C(n82), .D(n24), .Y(n84) );
  AND4XL U90 ( .A(n182), .B(n80), .C(r_txendk), .D(n226), .Y(n82) );
  NAND32XL U91 ( .B(n111), .C(n90), .A(n101), .Y(n228) );
  OAI2B11XL U92 ( .D(n288), .C(n106), .A(i_txreq), .B(n294), .Y(n107) );
  OAI221XL U93 ( .A(n22), .B(n116), .C(n115), .D(n123), .E(n38), .Y(n287) );
  OA21XL U94 ( .B(r_txnumk[0]), .C(n260), .A(n259), .Y(n265) );
  AO21XL U95 ( .B(n112), .C(n103), .A(n101), .Y(n99) );
  AO21XL U96 ( .B(i_rdat[6]), .C(n236), .A(n212), .Y(n242) );
  MUX2XL U97 ( .D0(i_rdat[7]), .D1(i_rdat[5]), .S(n239), .Y(n235) );
  NAND31XL U98 ( .C(n172), .A(n33), .B(n171), .Y(n234) );
  NAND3XL U99 ( .A(r_txauto[6]), .B(n15), .C(n16), .Y(n33) );
  NAND21XL U100 ( .B(r_txauto[6]), .A(n155), .Y(n227) );
  AOI21XL U101 ( .B(n154), .C(n153), .A(n228), .Y(n30) );
  INVXL U102 ( .A(n157), .Y(ptx_crcsidat[0]) );
  NAND32XL U103 ( .B(n101), .C(n90), .A(n111), .Y(n103) );
  NAND21XL U104 ( .B(n72), .A(n121), .Y(n123) );
  OAI22X1 U105 ( .A(bytcnt[1]), .B(n48), .C(bytcnt[0]), .D(n47), .Y(n49) );
  OAI21BBX1 U106 ( .A(bytcnt[4]), .B(n46), .C(r_txnumk[4]), .Y(n55) );
  NAND32X1 U107 ( .B(ptx_fsm[0]), .C(n90), .A(n101), .Y(n269) );
  INVXL U108 ( .A(bitcnt[0]), .Y(n244) );
  OR2X1 U109 ( .A(n113), .B(n31), .Y(n141) );
  OAI22XL U110 ( .A(n112), .B(n111), .C(n289), .D(n110), .Y(n31) );
  MUX4X1 U111 ( .D0(n209), .D1(n208), .D2(n211), .D3(n210), .S0(n239), .S1(n32), .Y(n248) );
  XNOR2XL U112 ( .A(bitcnt[0]), .B(n207), .Y(n32) );
  INVX1 U113 ( .A(n105), .Y(n108) );
  NAND21X1 U114 ( .B(n255), .A(n254), .Y(N251) );
  INVX1 U115 ( .A(n222), .Y(n145) );
  NAND21X1 U116 ( .B(n93), .A(n125), .Y(n105) );
  INVX1 U117 ( .A(n193), .Y(n187) );
  INVX1 U118 ( .A(n183), .Y(n218) );
  INVX1 U119 ( .A(n228), .Y(n182) );
  INVX1 U120 ( .A(n287), .Y(n139) );
  INVX1 U121 ( .A(n128), .Y(n255) );
  NAND21X1 U122 ( .B(n251), .A(n254), .Y(n128) );
  INVX1 U123 ( .A(n127), .Y(n254) );
  AND2X1 U124 ( .A(n270), .B(srstz), .Y(N298) );
  INVX1 U125 ( .A(i_txreq), .Y(n253) );
  NAND21X1 U126 ( .B(n217), .A(n215), .Y(n193) );
  NAND32X1 U127 ( .B(n199), .C(n166), .A(n194), .Y(n197) );
  MUX2BXL U128 ( .D0(n187), .D1(n186), .S(n185), .Y(n188) );
  INVX1 U129 ( .A(n216), .Y(n185) );
  NAND21X1 U130 ( .B(n222), .A(n214), .Y(n186) );
  AO21X1 U131 ( .B(n193), .C(n183), .A(n199), .Y(n169) );
  NAND21X1 U132 ( .B(n199), .A(n187), .Y(n146) );
  INVX1 U133 ( .A(n166), .Y(n215) );
  OAI211X1 U134 ( .C(n198), .D(n197), .A(n196), .B(n195), .Y(n202) );
  INVX1 U135 ( .A(n102), .Y(n96) );
  INVX1 U136 ( .A(n284), .Y(n175) );
  INVX1 U137 ( .A(n144), .Y(n155) );
  INVX1 U138 ( .A(n198), .Y(n214) );
  NAND21XL U139 ( .B(n70), .A(n256), .Y(n258) );
  AND2X1 U140 ( .A(n268), .B(srstz), .Y(N299) );
  INVX1 U141 ( .A(n171), .Y(n212) );
  INVX1 U142 ( .A(n227), .Y(n236) );
  INVX1 U143 ( .A(n234), .Y(n196) );
  AND2X1 U144 ( .A(n257), .B(n258), .Y(ptx_crcshfo4) );
  INVX1 U145 ( .A(n285), .Y(n164) );
  INVX1 U146 ( .A(n282), .Y(n150) );
  INVX1 U147 ( .A(n280), .Y(n219) );
  INVX1 U148 ( .A(n103), .Y(n257) );
  INVX1 U149 ( .A(srstz), .Y(n45) );
  INVX1 U150 ( .A(n268), .Y(n271) );
  INVXL U151 ( .A(n79), .Y(n85) );
  INVX1 U152 ( .A(r_txnumk[1]), .Y(n48) );
  INVX1 U153 ( .A(r_txauto[6]), .Y(n156) );
  INVX1 U154 ( .A(n110), .Y(n172) );
  OAI211X1 U155 ( .C(n91), .D(n90), .A(n89), .B(n88), .Y(n270) );
  OA22XL U156 ( .A(n104), .B(n87), .C(n93), .D(n228), .Y(n88) );
  AOI221XL U157 ( .A(n257), .B(n102), .C(n18), .D(n104), .E(n76), .Y(n91) );
  AOI32XL U158 ( .A(n288), .B(i_txreq), .C(n294), .D(n172), .E(n78), .Y(n89)
         );
  INVX1 U159 ( .A(n141), .Y(n272) );
  INVX1 U160 ( .A(n289), .Y(n106) );
  INVX1 U161 ( .A(n118), .Y(n275) );
  AO21X1 U162 ( .B(n255), .C(n27), .A(n276), .Y(n132) );
  AND2X1 U163 ( .A(n141), .B(srstz), .Y(N297) );
  INVX1 U164 ( .A(n130), .Y(n131) );
  NAND32X1 U165 ( .B(n27), .C(n244), .A(n255), .Y(n130) );
  NAND32X1 U166 ( .B(n100), .C(n105), .A(n99), .Y(n268) );
  INVX1 U167 ( .A(n104), .Y(n100) );
  INVX1 U168 ( .A(n98), .Y(n112) );
  OAI31XL U169 ( .A(n97), .B(n96), .C(n110), .D(n95), .Y(n98) );
  INVX1 U170 ( .A(n94), .Y(n97) );
  INVX1 U171 ( .A(n95), .Y(n76) );
  AND4XL U172 ( .A(n263), .B(n18), .C(n262), .D(n261), .Y(n264) );
  NAND21X1 U173 ( .B(n96), .A(n94), .Y(n78) );
  NAND21X1 U174 ( .B(n221), .A(n145), .Y(n166) );
  NAND32XL U175 ( .B(n73), .C(n269), .A(n126), .Y(n104) );
  NAND21XL U176 ( .B(n80), .A(n19), .Y(n102) );
  MUX3X1 U177 ( .D0(n242), .D1(n241), .D2(n240), .S0(n239), .S1(n7), .Y(n247)
         );
  AO21X1 U178 ( .B(n236), .C(n235), .A(n234), .Y(n240) );
  GEN2XL U179 ( .D(n217), .E(n221), .C(n200), .B(n218), .A(n30), .Y(n201) );
  OA21X1 U180 ( .B(n199), .C(n221), .A(n213), .Y(n200) );
  OA222X1 U181 ( .A(n227), .B(n167), .C(n166), .D(n223), .E(n165), .F(n228), 
        .Y(n168) );
  AOI221XL U182 ( .A(n178), .B(n219), .C(n21), .D(n164), .E(n284), .Y(n165) );
  OA22X1 U183 ( .A(r_txauto[4]), .B(n104), .C(n103), .D(n102), .Y(n109) );
  AO21X1 U184 ( .B(n224), .C(n223), .A(n222), .Y(n225) );
  INVX1 U185 ( .A(n221), .Y(n224) );
  NAND32X1 U186 ( .B(n189), .C(n166), .A(n199), .Y(n147) );
  AND4X1 U187 ( .A(n196), .B(n192), .C(n191), .D(n190), .Y(n209) );
  AOI221XL U188 ( .A(i_rdat[3]), .B(n236), .C(n218), .D(n189), .E(n188), .Y(
        n190) );
  NAND32X1 U189 ( .B(n180), .C(n220), .A(n179), .Y(n181) );
  NOR5X1 U190 ( .A(n160), .B(n159), .C(n30), .D(n158), .E(n212), .Y(n211) );
  INVX1 U191 ( .A(n197), .Y(n159) );
  NAND43X1 U192 ( .B(n233), .C(n232), .D(n231), .A(n230), .Y(n241) );
  AND3X1 U193 ( .A(n215), .B(n214), .C(n213), .Y(n233) );
  AND3X1 U194 ( .A(n218), .B(n217), .C(n216), .Y(n232) );
  OAI221XL U195 ( .A(n229), .B(n228), .C(n227), .D(n226), .E(n225), .Y(n231)
         );
  NAND32XL U196 ( .B(n157), .C(n156), .A(n155), .Y(n171) );
  NAND21X1 U197 ( .B(n194), .A(n184), .Y(n216) );
  INVX1 U198 ( .A(n213), .Y(n194) );
  INVX1 U199 ( .A(n189), .Y(n217) );
  AOI22X1 U200 ( .A(n152), .B(n21), .C(n151), .D(n150), .Y(n154) );
  MUX2BXL U201 ( .D0(n175), .D1(n286), .S(n178), .Y(n153) );
  AOI211X1 U202 ( .C(n260), .D(n281), .A(n220), .B(n219), .Y(n229) );
  INVX1 U203 ( .A(n243), .Y(n207) );
  XNOR2XL U204 ( .A(n245), .B(n34), .Y(n246) );
  AOI21X1 U205 ( .B(n244), .C(n27), .A(n243), .Y(n34) );
  INVX1 U206 ( .A(n184), .Y(n199) );
  INVX1 U207 ( .A(n274), .Y(ptx_goidle) );
  INVX1 U208 ( .A(n92), .Y(n142) );
  INVX1 U209 ( .A(r_txauto[4]), .Y(n87) );
  INVX1 U210 ( .A(n176), .Y(n178) );
  INVX1 U211 ( .A(n192), .Y(n158) );
  AND4X1 U212 ( .A(n272), .B(n271), .C(n270), .D(n269), .Y(ptx_pspyld) );
  INVX1 U213 ( .A(r_txnumk[2]), .Y(n51) );
  AND3X2 U214 ( .A(n14), .B(n64), .C(n36), .Y(n134) );
  INVX1 U215 ( .A(r_txendk), .Y(n56) );
  NAND21X1 U216 ( .B(r_txnumk[2]), .A(bytcnt[2]), .Y(n266) );
  NAND21XL U217 ( .B(r_txnumk[3]), .A(bytcnt[3]), .Y(n261) );
  NAND21X1 U218 ( .B(r_txnumk[4]), .A(bytcnt[4]), .Y(n262) );
  NAND32XL U219 ( .B(ptx_fsm[1]), .C(n111), .A(n101), .Y(n110) );
  NAND21XL U220 ( .B(ptx_fsm[1]), .A(n111), .Y(n135) );
  INVXL U221 ( .A(bytcnt[2]), .Y(n119) );
  INVXL U222 ( .A(bytcnt[1]), .Y(n80) );
  INVXL U223 ( .A(bytcnt[3]), .Y(n72) );
  INVXL U224 ( .A(bytcnt[4]), .Y(n115) );
  OAI211X1 U225 ( .C(r_txauto[5]), .D(n109), .A(n108), .B(n107), .Y(n113) );
  NAND21XL U226 ( .B(bytcnt[0]), .A(n139), .Y(n118) );
  XOR2XL U227 ( .A(ptx_fsm[0]), .B(n272), .Y(n114) );
  OA21XL U228 ( .B(n124), .C(bytcnt[4]), .A(n139), .Y(N273) );
  INVX1 U229 ( .A(n123), .Y(n124) );
  AND2X1 U230 ( .A(n122), .B(n139), .Y(N272) );
  XOR2XL U231 ( .A(bytcnt[3]), .B(n121), .Y(n122) );
  AND2X1 U232 ( .A(n140), .B(n139), .Y(N270) );
  XOR2XL U233 ( .A(bytcnt[1]), .B(bytcnt[0]), .Y(n140) );
  OAI22XL U234 ( .A(n287), .B(n120), .C(n119), .D(n118), .Y(N271) );
  MUX2XL U235 ( .D0(n119), .D1(n117), .S(bytcnt[1]), .Y(n120) );
  NAND21XL U236 ( .B(bytcnt[2]), .A(bytcnt[0]), .Y(n117) );
  AND3X1 U237 ( .A(n39), .B(n40), .C(n114), .Y(n38) );
  XNOR2XL U238 ( .A(n270), .B(ptx_fsm[1]), .Y(n39) );
  AOI21XL U239 ( .B(n268), .C(n101), .A(i_txreq), .Y(n40) );
  INVX1 U240 ( .A(n129), .Y(n276) );
  NAND21XL U241 ( .B(bitcnt[0]), .A(n255), .Y(n129) );
  MUX2IXL U242 ( .D0(n41), .D1(n42), .S(bitcnt[3]), .Y(N255) );
  NAND2XL U243 ( .A(n131), .B(bitcnt[2]), .Y(n41) );
  AOI21X1 U244 ( .B(n255), .C(n245), .A(n132), .Y(n42) );
  MUX2XL U245 ( .D0(n131), .D1(n132), .S(bitcnt[2]), .Y(N254) );
  MUX2AXL U246 ( .D0(n43), .D1(n276), .S(bitcnt[1]), .Y(N253) );
  NAND2XL U247 ( .A(n255), .B(bitcnt[0]), .Y(n43) );
  MUX2IX1 U248 ( .D0(n278), .D1(n277), .S(n44), .Y(n238) );
  NAND3X1 U249 ( .A(srstz), .B(n253), .C(n252), .Y(n44) );
  MUX2XL U250 ( .D0(n138), .D1(n8), .S(n137), .Y(n237) );
  AND3XL U251 ( .A(n133), .B(n263), .C(n253), .Y(n138) );
  AND4XL U252 ( .A(n269), .B(n274), .C(n103), .D(n110), .Y(n74) );
  AND4X1 U253 ( .A(n230), .B(n192), .C(n169), .D(n168), .Y(n210) );
  AOI211XL U254 ( .C(i_rdat[1]), .D(n236), .A(n202), .B(n201), .Y(n208) );
  MUX2XL U255 ( .D0(n251), .D1(n250), .S(prx_cccnt[1]), .Y(n252) );
  NAND21XL U256 ( .B(n249), .A(ptx_txact), .Y(n250) );
  MUX2BXL U257 ( .D0(n248), .D1(n247), .S(n246), .Y(n249) );
  MUX2IXL U258 ( .D0(bitcnt[1]), .D1(n205), .S(n8), .Y(n239) );
  MUX2XL U259 ( .D0(ptx_crcsidat[3]), .D1(pcc_crc30[3]), .S(n257), .Y(n221) );
  MUX2XL U260 ( .D0(ptx_crcsidat[2]), .D1(pcc_crc30[2]), .S(n257), .Y(n189) );
  MUX2BXL U261 ( .D0(n143), .D1(pcc_crc30[1]), .S(n257), .Y(n213) );
  INVX1 U262 ( .A(n163), .Y(n230) );
  GEN2XL U263 ( .D(n8), .E(n281), .C(n180), .B(n182), .A(n212), .Y(n163) );
  OAI221X1 U264 ( .A(n282), .B(n177), .C(n176), .D(n175), .E(n174), .Y(n220)
         );
  MUX2XL U265 ( .D0(bytcnt[0]), .D1(hinib), .S(r_txauto[0]), .Y(n177) );
  MUX2XL U266 ( .D0(n283), .D1(n173), .S(hinib), .Y(n174) );
  NAND21X1 U267 ( .B(n285), .A(n176), .Y(n173) );
  MUX2X1 U268 ( .D0(ptx_crcsidat[0]), .D1(pcc_crc30[0]), .S(n257), .Y(n184) );
  AO21XL U269 ( .B(n281), .C(bytcnt[0]), .A(n164), .Y(n152) );
  OA22XL U270 ( .A(n280), .B(n178), .C(bytcnt[0]), .D(n279), .Y(n179) );
  INVX1 U271 ( .A(n162), .Y(n180) );
  OAI211XL U272 ( .C(n8), .D(bytcnt[0]), .A(n176), .B(n161), .Y(n162) );
  INVX1 U273 ( .A(n283), .Y(n161) );
  NAND43XL U274 ( .B(ptx_cc), .C(n251), .D(n92), .A(ptx_fsm[0]), .Y(n274) );
  MUX2XL U275 ( .D0(bytcnt[0]), .D1(hinib), .S(r_txauto[0]), .Y(n151) );
  NAND21XL U276 ( .B(n260), .A(hinib), .Y(n176) );
  NAND21XL U277 ( .B(ptx_fsm[1]), .A(ptx_fsm[2]), .Y(n92) );
  INVXL U278 ( .A(bytcnt[0]), .Y(n260) );
  NAND21XL U279 ( .B(ptx_fsm[0]), .A(n142), .Y(n192) );
  INVX1 U280 ( .A(n71), .Y(n121) );
  NAND32XL U281 ( .B(n80), .C(n260), .A(bytcnt[2]), .Y(n71) );
  INVXL U282 ( .A(bitcnt[2]), .Y(n245) );
  NAND21XL U283 ( .B(n77), .A(r_txshrt), .Y(n94) );
  AOI31XL U284 ( .A(n110), .B(n228), .C(n103), .D(n77), .Y(n116) );
  AND3XL U285 ( .A(n18), .B(n267), .C(n258), .Y(ptx_crcshfi4) );
  AOI32XL U286 ( .A(n215), .B(n213), .C(n267), .D(n182), .E(n181), .Y(n191) );
  NAND32XL U287 ( .B(n267), .C(n184), .A(n194), .Y(n223) );
  NAND21XL U288 ( .B(n267), .A(n217), .Y(n198) );
  AND4XL U289 ( .A(n267), .B(n266), .C(n265), .D(n264), .Y(ptx_crcstart) );
  NAND32X1 U290 ( .B(n256), .C(n267), .A(n68), .Y(n69) );
  OAI211X1 U291 ( .C(n53), .D(n52), .A(n261), .B(n262), .Y(n54) );
  OAI31XL U292 ( .A(n228), .B(bytcnt[1]), .C(n75), .D(n74), .Y(n95) );
  AOI211XL U293 ( .C(n136), .D(n135), .A(i_txreq), .B(n134), .Y(n137) );
  NAND21XL U294 ( .B(n16), .A(n8), .Y(n243) );
  XOR2XL U295 ( .A(n204), .B(n203), .Y(n205) );
  NAND21XL U296 ( .B(n16), .A(bitcnt[0]), .Y(n204) );
  NAND21XL U297 ( .B(n172), .A(n16), .Y(n144) );
  NAND32XL U298 ( .B(n142), .C(n16), .A(n228), .Y(n222) );
  OAI211X1 U299 ( .C(n73), .D(n56), .A(n54), .B(n55), .Y(n57) );
  NOR2X1 U300 ( .A(n45), .B(n278), .Y(n277) );
  INVX1 U301 ( .A(ptx_cc), .Y(n278) );
  NAND2X1 U302 ( .A(n285), .B(n283), .Y(n286) );
  INVX1 U303 ( .A(n279), .Y(n281) );
  NAND2X1 U304 ( .A(n38), .B(n287), .Y(N268) );
  NOR43XL U305 ( .B(n285), .C(n290), .D(n279), .A(n284), .Y(n289) );
  NOR3XL U306 ( .A(n291), .B(r_txauto[0]), .C(n292), .Y(n284) );
  NAND3X1 U307 ( .A(r_txauto[0]), .B(n292), .C(r_txauto[2]), .Y(n279) );
  AND3X1 U308 ( .A(n282), .B(n280), .C(n283), .Y(n290) );
  NAND3X1 U309 ( .A(n293), .B(n292), .C(r_txauto[2]), .Y(n283) );
  INVX1 U310 ( .A(r_txauto[0]), .Y(n293) );
  NAND3X1 U311 ( .A(n292), .B(n291), .C(r_txauto[0]), .Y(n280) );
  INVX1 U312 ( .A(r_txauto[1]), .Y(n292) );
  NAND2X1 U313 ( .A(r_txauto[1]), .B(n291), .Y(n282) );
  INVX1 U314 ( .A(r_txauto[2]), .Y(n291) );
  NAND3X1 U315 ( .A(r_txauto[2]), .B(r_txauto[0]), .C(r_txauto[1]), .Y(n285)
         );
  INVX1 U316 ( .A(r_txauto[3]), .Y(n288) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyidd_a0 ( i_trans, i_goidle, o_ccidle, o_goidle, o_gobusy, clk, srstz
 );
  input i_trans, i_goidle, clk, srstz;
  output o_ccidle, o_goidle, o_gobusy;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N46, N47, N48, N49, N50, N51,
         N52, N53, N55, N56, N57, N58, N59, N60, N61, N62, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, net10668, net10674, net10679, n29, n30, n31, n32, n33, n34, n35,
         n36, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n53, n54, n55, n56, n57, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n37, n52, n58, n59, n60, n61, n62, n63;
  wire   [7:0] ttranwin;
  wire   [1:0] ntrancnt;
  wire   [7:0] trans0;
  wire   [7:0] ttranwin_minus;
  wire   [7:0] trans1;

  SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 clk_gate_trans1_reg ( .CLK(clk), .EN(N90), 
        .ENCLK(net10668), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 clk_gate_trans0_reg ( .CLK(clk), .EN(N91), 
        .ENCLK(net10674), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 clk_gate_ttranwin_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net10679), .TE(1'b0) );
  phyidd_a0_DW01_sub_0 sub_47 ( .A(trans1), .B(trans0), .CI(1'b0), .DIFF({N53, 
        N52, N51, N50, N49, N48, N47, N46}), .CO() );
  phyidd_a0_DW01_sub_1 sub_24 ( .A({n63, n62, n61, n60, n59, n58, n52, n37}), 
        .B(trans0), .CI(1'b0), .DIFF(ttranwin_minus), .CO() );
  phyidd_a0_DW01_inc_0 add_23 ( .A(ttranwin), .SUM({N18, N17, N16, N15, N14, 
        N13, N12, N11}) );
  DFFQX1 trans1_reg_6_ ( .D(N79), .C(net10668), .Q(trans1[6]) );
  DFFQX1 trans1_reg_7_ ( .D(N80), .C(net10668), .Q(trans1[7]) );
  DFFQX1 trans0_reg_7_ ( .D(N62), .C(net10674), .Q(trans0[7]) );
  DFFQX1 trans1_reg_4_ ( .D(N77), .C(net10668), .Q(trans1[4]) );
  DFFQX1 trans1_reg_5_ ( .D(N78), .C(net10668), .Q(trans1[5]) );
  DFFQX1 trans0_reg_5_ ( .D(N60), .C(net10674), .Q(trans0[5]) );
  DFFQX1 trans0_reg_6_ ( .D(N61), .C(net10674), .Q(trans0[6]) );
  DFFQX1 trans1_reg_3_ ( .D(N76), .C(net10668), .Q(trans1[3]) );
  DFFQX1 trans0_reg_4_ ( .D(N59), .C(net10674), .Q(trans0[4]) );
  DFFQX1 trans1_reg_1_ ( .D(N74), .C(net10668), .Q(trans1[1]) );
  DFFQX1 trans1_reg_2_ ( .D(N75), .C(net10668), .Q(trans1[2]) );
  DFFQX1 ntrancnt_reg_1_ ( .D(n56), .C(clk), .Q(ntrancnt[1]) );
  DFFQX1 trans0_reg_2_ ( .D(N57), .C(net10674), .Q(trans0[2]) );
  DFFQX1 trans0_reg_3_ ( .D(N58), .C(net10674), .Q(trans0[3]) );
  DFFQX1 ntrancnt_reg_0_ ( .D(n57), .C(clk), .Q(ntrancnt[0]) );
  DFFQX1 trans1_reg_0_ ( .D(N73), .C(net10668), .Q(trans1[0]) );
  DFFQX1 trans0_reg_0_ ( .D(N55), .C(net10674), .Q(trans0[0]) );
  DFFQX1 trans0_reg_1_ ( .D(N56), .C(net10674), .Q(trans0[1]) );
  DFFQX1 ttranwin_reg_7_ ( .D(N89), .C(net10679), .Q(ttranwin[7]) );
  DFFQX1 ttranwin_reg_5_ ( .D(N87), .C(net10679), .Q(ttranwin[5]) );
  DFFQX1 ttranwin_reg_1_ ( .D(N83), .C(net10679), .Q(ttranwin[1]) );
  DFFQX1 ttranwin_reg_6_ ( .D(N88), .C(net10679), .Q(ttranwin[6]) );
  DFFQX1 ttranwin_reg_0_ ( .D(N82), .C(net10679), .Q(ttranwin[0]) );
  DFFQX1 ttranwin_reg_4_ ( .D(N86), .C(net10679), .Q(ttranwin[4]) );
  DFFQX1 ttranwin_reg_2_ ( .D(N84), .C(net10679), .Q(ttranwin[2]) );
  DFFQX1 ttranwin_reg_3_ ( .D(N85), .C(net10679), .Q(ttranwin[3]) );
  DFFQX1 ccidle_reg ( .D(n55), .C(clk), .Q(o_ccidle) );
  NAND2X1 U3 ( .A(ntrancnt[0]), .B(n28), .Y(n3) );
  NAND2X1 U4 ( .A(ntrancnt[1]), .B(n26), .Y(n4) );
  INVX1 U5 ( .A(n25), .Y(n50) );
  INVX1 U6 ( .A(n6), .Y(n5) );
  INVX1 U7 ( .A(n14), .Y(o_gobusy) );
  OAI22X1 U8 ( .A(n30), .B(n47), .C(n46), .D(n18), .Y(N88) );
  NAND21X1 U11 ( .B(n13), .A(n12), .Y(n25) );
  NAND2X1 U12 ( .A(n50), .B(n27), .Y(n46) );
  OAI22X1 U13 ( .A(n31), .B(n47), .C(n46), .D(n19), .Y(N87) );
  OAI22X1 U14 ( .A(n32), .B(n47), .C(n46), .D(n20), .Y(N86) );
  OAI22X1 U15 ( .A(n33), .B(n47), .C(n46), .D(n21), .Y(N85) );
  OAI22X1 U16 ( .A(n34), .B(n47), .C(n46), .D(n22), .Y(N84) );
  OAI22X1 U17 ( .A(n35), .B(n47), .C(n46), .D(n23), .Y(N83) );
  INVX1 U18 ( .A(srstz), .Y(n6) );
  NAND21X1 U19 ( .B(n41), .A(n10), .Y(n14) );
  NAND2X1 U20 ( .A(N12), .B(n45), .Y(n35) );
  INVX1 U21 ( .A(n7), .Y(n10) );
  NAND21X1 U22 ( .B(n9), .A(i_trans), .Y(n7) );
  INVX1 U23 ( .A(n36), .Y(n37) );
  OAI22X1 U24 ( .A(n29), .B(n41), .C(n43), .D(n17), .Y(N80) );
  OAI22X1 U25 ( .A(n29), .B(n47), .C(n46), .D(n17), .Y(N89) );
  AO21X1 U26 ( .B(n16), .C(n9), .A(i_goidle), .Y(o_goidle) );
  INVX1 U27 ( .A(ttranwin_minus[6]), .Y(n18) );
  NAND2X1 U28 ( .A(N13), .B(n45), .Y(n34) );
  OAI22X1 U29 ( .A(n30), .B(n4), .C(n43), .D(n18), .Y(N79) );
  NAND31X1 U30 ( .C(N91), .A(n48), .B(n51), .Y(N81) );
  OA21X1 U31 ( .B(n4), .C(n13), .A(n12), .Y(n51) );
  NAND32X1 U32 ( .B(n16), .C(n11), .A(n13), .Y(n48) );
  AND2X1 U33 ( .A(n48), .B(n49), .Y(n47) );
  OAI21BBX1 U34 ( .A(n4), .B(n40), .C(n50), .Y(n49) );
  INVX1 U35 ( .A(ttranwin_minus[5]), .Y(n19) );
  INVX1 U36 ( .A(ttranwin_minus[4]), .Y(n20) );
  NAND2X1 U37 ( .A(N14), .B(n45), .Y(n33) );
  NAND2X1 U38 ( .A(N15), .B(n45), .Y(n32) );
  INVX1 U39 ( .A(n11), .Y(n12) );
  OAI222XL U40 ( .A(n38), .B(n28), .C(n39), .D(n3), .E(n41), .F(n39), .Y(n56)
         );
  OAI21X1 U41 ( .B(n40), .C(n25), .A(n46), .Y(N91) );
  EORX1 U42 ( .A(n39), .B(n42), .C(n39), .D(n43), .Y(n38) );
  INVX1 U43 ( .A(n15), .Y(n42) );
  NAND32X1 U44 ( .B(o_goidle), .C(n44), .A(n14), .Y(n15) );
  OAI21X1 U45 ( .B(n45), .C(i_trans), .A(n5), .Y(n44) );
  OAI22X1 U46 ( .A(n36), .B(n47), .C(n46), .D(n24), .Y(N82) );
  OAI22X1 U47 ( .A(n31), .B(n41), .C(n43), .D(n19), .Y(N78) );
  OAI22X1 U48 ( .A(n32), .B(n4), .C(n43), .D(n20), .Y(N77) );
  NAND2X1 U49 ( .A(n42), .B(i_trans), .Y(n39) );
  INVX1 U50 ( .A(n45), .Y(n16) );
  INVX1 U51 ( .A(ttranwin_minus[3]), .Y(n21) );
  NOR2X1 U52 ( .A(n16), .B(N17), .Y(n30) );
  NAND2X1 U53 ( .A(N16), .B(n45), .Y(n31) );
  INVX1 U54 ( .A(i_trans), .Y(n13) );
  OAI22X1 U55 ( .A(n33), .B(n41), .C(n43), .D(n21), .Y(N76) );
  OAI21X1 U56 ( .B(n41), .C(n25), .A(n46), .Y(N90) );
  ENOX1 U57 ( .A(n30), .B(n3), .C(N52), .D(n27), .Y(N61) );
  ENOX1 U58 ( .A(n31), .B(n40), .C(N51), .D(n27), .Y(N60) );
  INVX1 U59 ( .A(ttranwin_minus[2]), .Y(n22) );
  INVX1 U60 ( .A(ttranwin_minus[1]), .Y(n23) );
  OAI22X1 U61 ( .A(n34), .B(n4), .C(n43), .D(n22), .Y(N75) );
  OAI22X1 U62 ( .A(n35), .B(n41), .C(n43), .D(n23), .Y(N74) );
  ENOX1 U63 ( .A(n32), .B(n3), .C(N50), .D(n27), .Y(N59) );
  OAI211X1 U64 ( .C(o_gobusy), .D(n9), .A(n5), .B(n8), .Y(n55) );
  INVX1 U65 ( .A(o_goidle), .Y(n8) );
  INVX1 U66 ( .A(ttranwin_minus[0]), .Y(n24) );
  OAI22X1 U67 ( .A(n36), .B(n4), .C(n43), .D(n24), .Y(N73) );
  ENOX1 U68 ( .A(n33), .B(n40), .C(N49), .D(n27), .Y(N58) );
  ENOX1 U69 ( .A(n34), .B(n3), .C(N48), .D(n27), .Y(N57) );
  INVX1 U70 ( .A(n43), .Y(n27) );
  ENOX1 U71 ( .A(n35), .B(n40), .C(N47), .D(n27), .Y(N56) );
  INVX1 U72 ( .A(n34), .Y(n58) );
  INVX1 U73 ( .A(n33), .Y(n59) );
  INVX1 U74 ( .A(n32), .Y(n60) );
  INVX1 U75 ( .A(n31), .Y(n61) );
  INVX1 U76 ( .A(n30), .Y(n62) );
  NAND4X1 U77 ( .A(ttranwin[7]), .B(ttranwin[6]), .C(n53), .D(n54), .Y(n45) );
  NOR2X1 U78 ( .A(ttranwin[1]), .B(ttranwin[0]), .Y(n53) );
  NOR4XL U79 ( .A(ttranwin[5]), .B(ttranwin[4]), .C(ttranwin[3]), .D(
        ttranwin[2]), .Y(n54) );
  INVX1 U80 ( .A(n35), .Y(n52) );
  INVX1 U81 ( .A(ttranwin_minus[7]), .Y(n17) );
  INVX1 U82 ( .A(n29), .Y(n63) );
  NAND2X1 U83 ( .A(N11), .B(n45), .Y(n36) );
  AO21X1 U84 ( .B(n10), .C(n26), .A(n6), .Y(n11) );
  OAI22X1 U85 ( .A(n38), .B(n26), .C(ntrancnt[0]), .D(n39), .Y(n57) );
  ENOX1 U86 ( .A(n29), .B(n3), .C(N53), .D(n27), .Y(N62) );
  NOR2X1 U87 ( .A(n16), .B(N18), .Y(n29) );
  NAND2X1 U88 ( .A(ntrancnt[1]), .B(n26), .Y(n41) );
  INVX1 U89 ( .A(o_ccidle), .Y(n9) );
  INVX1 U90 ( .A(ntrancnt[0]), .Y(n26) );
  NAND2X1 U91 ( .A(ntrancnt[0]), .B(ntrancnt[1]), .Y(n43) );
  NAND2X1 U92 ( .A(ntrancnt[0]), .B(n28), .Y(n40) );
  INVX1 U93 ( .A(ntrancnt[1]), .Y(n28) );
  ENOX1 U94 ( .A(n36), .B(n40), .C(N46), .D(n27), .Y(N55) );
endmodule


module phyidd_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module phyidd_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n9), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n7), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n5), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n4), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n3), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U3 ( .A(B[2]), .Y(n5) );
  INVX1 U4 ( .A(B[3]), .Y(n6) );
  INVX1 U5 ( .A(B[4]), .Y(n7) );
  INVX1 U6 ( .A(B[5]), .Y(n8) );
  INVX1 U7 ( .A(B[6]), .Y(n9) );
  INVX1 U8 ( .A(B[1]), .Y(n4) );
  NAND21X1 U9 ( .B(n2), .A(n1), .Y(carry[1]) );
  INVX1 U10 ( .A(B[7]), .Y(n3) );
  INVX1 U11 ( .A(B[0]), .Y(n2) );
endmodule


module phyidd_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n9), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n7), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n5), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n4), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n3), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(B[2]), .Y(n5) );
  INVX1 U2 ( .A(B[3]), .Y(n6) );
  INVX1 U3 ( .A(B[4]), .Y(n7) );
  INVX1 U4 ( .A(B[5]), .Y(n8) );
  INVX1 U5 ( .A(B[6]), .Y(n9) );
  INVX1 U6 ( .A(B[1]), .Y(n4) );
  NAND21X1 U7 ( .B(n2), .A(n1), .Y(carry[1]) );
  INVX1 U8 ( .A(A[0]), .Y(n1) );
  INVX1 U9 ( .A(B[0]), .Y(n2) );
  INVX1 U10 ( .A(B[7]), .Y(n3) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_a0 ( i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, 
        r_rxdb_opt, r_ords_ena, r_pshords, r_rgdcrc, prx_cccnt, prx_rst, 
        prx_setsta, prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, 
        prx_fifopsh, prx_fifowdat, pff_txreq, pid_gobusy, pid_goidle, 
        pid_ccidle, pcc_rxgood, prx_crcstart, prx_crcshfi4, prx_crcsidat, 
        prx_rxcode, prx_adpn, prx_rcvdords, prx_eoprcvd, prx_fsm, clk, srstz
 );
  input [1:0] r_rxdb_opt;
  input [6:0] r_ords_ena;
  output [1:0] prx_cccnt;
  output [1:0] prx_rst;
  output [6:0] prx_setsta;
  output [7:0] prx_fifowdat;
  output [3:0] prx_crcsidat;
  output [4:0] prx_rxcode;
  output [5:0] prx_adpn;
  output [2:0] prx_rcvdords;
  output [3:0] prx_fsm;
  input i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_pshords,
         r_rgdcrc, pff_txreq, pid_gobusy, pid_goidle, pid_ccidle, pcc_rxgood,
         clk, srstz;
  output prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, prx_fifopsh,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd;
  wire   N31, N32, n287, db_gohi, db_golo, k0_det, cctrans, shrtrans, N70, N71,
         N72, N73, N74, N75, N76, N96, N153, N154, N155, N156, N157, N236,
         N238, N239, N246, N247, N248, N249, N250, N251, N275, N276, N277,
         N278, N279, net10696, net10702, net10707, net10712, net10717,
         net10722, net10727, n21, n214, net148177, net148351, net148365,
         net148378, net148388, net148389, net148391, net148392, net148394,
         net148412, net162096, net163489, net167457, net167456, net169093,
         net169136, n1, n2, n3, n4, n6, n7, n9, n10, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n22, n23, n24, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n281, n282,
         n283, n284, n285, n286;
  wire   [5:0] cccnt;
  wire   [2:0] ps_dat5b;
  wire   [2:0] bcnt;
  wire   [7:3] ordsbuf;

  phyrx_db u0_phyrx_db ( .clk(clk), .srstz(n46), .x_cc(i_cc), .ptx_txact(
        ptx_txact), .r_rxdb_opt(r_rxdb_opt), .gohi(db_gohi), .golo(db_golo), 
        .gotrans(prx_trans) );
  phyrx_adp u0_phyrx_adp ( .clk(clk), .srstz(n47), .gohi(db_gohi), .golo(
        db_golo), .gobusy(pid_gobusy), .goidle(pid_goidle), .i_ccidle(
        pid_ccidle), .k0_det(k0_det), .r_adprx_en(r_adprx_en), .r_adp2nd(
        r_adp2nd), .adp_val(prx_adpn), .d_cc(prx_d_cc), .cctrans(cctrans) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 clk_gate_cccnt_reg ( .CLK(clk), .EN(N70), 
        .ENCLK(net10696), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 clk_gate_cs_dat5b_reg ( .CLK(clk), .EN(N153), 
        .ENCLK(net10702), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 clk_gate_bcnt_reg ( .CLK(clk), .EN(N236), 
        .ENCLK(net10707), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 clk_gate_cs_dat4b_reg ( .CLK(clk), .EN(n21), 
        .ENCLK(net10712), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 clk_gate_ordsbuf_reg ( .CLK(clk), .EN(N251), 
        .ENCLK(net10717), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 clk_gate_ordsbuf_reg_0 ( .CLK(clk), .EN(N250), .ENCLK(net10722), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 clk_gate_cs_bmni_reg ( .CLK(clk), .EN(N275), 
        .ENCLK(net10727), .TE(1'b0) );
  DFFQX1 ordsbuf_reg_5_ ( .D(prx_crcsidat[1]), .C(net10717), .Q(ordsbuf[5]) );
  DFFQX1 ordsbuf_reg_6_ ( .D(prx_crcsidat[2]), .C(net10717), .Q(ordsbuf[6]) );
  DFFQX1 ordsbuf_reg_7_ ( .D(prx_fifowdat[7]), .C(net10717), .Q(ordsbuf[7]) );
  DFFQX1 ordsbuf_reg_3_ ( .D(N249), .C(net10722), .Q(ordsbuf[3]) );
  DFFQX1 ordsbuf_reg_4_ ( .D(prx_crcsidat[0]), .C(net10717), .Q(ordsbuf[4]) );
  DFFQX1 cs_dat4b_reg_2_ ( .D(prx_crcsidat[2]), .C(net10712), .Q(
        prx_fifowdat[2]) );
  DFFQX1 cs_dat4b_reg_1_ ( .D(prx_fifowdat[5]), .C(net10712), .Q(
        prx_fifowdat[1]) );
  DFFQX1 cs_dat4b_reg_0_ ( .D(prx_crcsidat[0]), .C(net10712), .Q(
        prx_fifowdat[0]) );
  DFFQX1 cs_dat4b_reg_3_ ( .D(prx_crcsidat[3]), .C(net10712), .Q(prx_rxcode[3]) );
  DFFQX1 cs_dat4b_reg_4_ ( .D(net169093), .C(net10712), .Q(prx_rxcode[4]) );
  DFFQX1 bcnt_reg_1_ ( .D(N238), .C(net10707), .Q(bcnt[1]) );
  DFFQX1 bcnt_reg_2_ ( .D(N239), .C(net10707), .Q(bcnt[2]) );
  DFFQX1 shrtrans_reg ( .D(n214), .C(clk), .Q(shrtrans) );
  DFFQX1 cs_dat5b_reg_0_ ( .D(N154), .C(net10702), .Q(ps_dat5b[0]) );
  DFFQX1 cs_dat5b_reg_2_ ( .D(N156), .C(net10702), .Q(ps_dat5b[2]) );
  DFFQX1 cs_dat5b_reg_1_ ( .D(N155), .C(net10702), .Q(ps_dat5b[1]) );
  DFFQX1 cccnt_reg_1_ ( .D(N72), .C(net10696), .Q(cccnt[1]) );
  DFFQX1 cccnt_reg_2_ ( .D(N73), .C(net10696), .Q(cccnt[2]) );
  DFFQX1 cccnt_reg_4_ ( .D(N75), .C(net10696), .Q(cccnt[4]) );
  DFFQX1 cccnt_reg_3_ ( .D(N74), .C(net10696), .Q(cccnt[3]) );
  DFFQX1 bcnt_reg_0_ ( .D(n281), .C(net10707), .Q(bcnt[0]) );
  DFFQX1 cccnt_reg_0_ ( .D(N71), .C(net10696), .Q(cccnt[0]) );
  DFFQX1 cccnt_reg_5_ ( .D(N76), .C(net10696), .Q(cccnt[5]) );
  DFFQX1 ordsbuf_reg_0_ ( .D(N246), .C(net10722), .Q(prx_rcvdords[0]) );
  DFFQX1 ordsbuf_reg_1_ ( .D(N247), .C(net10722), .Q(prx_rcvdords[1]) );
  DFFQX1 cs_dat5b_reg_3_ ( .D(N157), .C(net10702), .Q(prx_bmc) );
  DFFQX1 cs_bmni_reg_3_ ( .D(N279), .C(net10727), .Q(n287) );
  DFFQX1 ordsbuf_reg_2_ ( .D(N248), .C(net10722), .Q(prx_rcvdords[2]) );
  DFFQX1 cs_bmni_reg_2_ ( .D(N278), .C(net10727), .Q(prx_fsm[2]) );
  DFFQX1 cs_bmni_reg_1_ ( .D(N277), .C(net10727), .Q(prx_fsm[1]) );
  DFFQX1 cs_bmni_reg_0_ ( .D(N276), .C(net10727), .Q(prx_fsm[0]) );
  INVX2 U3 ( .A(n268), .Y(n83) );
  NAND2X2 U4 ( .A(n45), .B(n1), .Y(n2) );
  INVX2 U5 ( .A(net148177), .Y(n1) );
  INVX1 U6 ( .A(cccnt[0]), .Y(net148391) );
  INVX1 U7 ( .A(prx_fsm[1]), .Y(n86) );
  GEN2XL U8 ( .D(shrtrans), .E(net148391), .C(net148392), .B(net162096), .A(
        net148394), .Y(n17) );
  NAND21X1 U9 ( .B(n259), .A(n258), .Y(n263) );
  NAND21X1 U10 ( .B(n257), .A(n256), .Y(n258) );
  INVX1 U11 ( .A(n262), .Y(n35) );
  AO21X1 U12 ( .B(n148), .C(n117), .A(n139), .Y(n118) );
  AO21X1 U13 ( .B(n128), .C(n148), .A(n112), .Y(n113) );
  NAND21X1 U14 ( .B(prx_fsm[2]), .A(prx_fsm[0]), .Y(n87) );
  INVX1 U15 ( .A(n84), .Y(n89) );
  INVX1 U16 ( .A(cccnt[4]), .Y(n277) );
  INVX1 U17 ( .A(n71), .Y(n44) );
  NOR32XL U18 ( .B(ps_dat5b[0]), .C(ps_dat5b[2]), .A(n91), .Y(n71) );
  AOI21X1 U19 ( .B(net148365), .C(n77), .A(n80), .Y(n45) );
  INVX1 U20 ( .A(ps_dat5b[1]), .Y(net148365) );
  AND2X1 U21 ( .A(n22), .B(n28), .Y(n29) );
  INVX1 U22 ( .A(bcnt[2]), .Y(n224) );
  INVX1 U23 ( .A(n188), .Y(n257) );
  AO21X1 U24 ( .B(n54), .C(n56), .A(n48), .Y(N74) );
  AO21X1 U25 ( .B(n52), .C(n56), .A(n48), .Y(N73) );
  AND2X1 U26 ( .A(n47), .B(net148389), .Y(n214) );
  NAND2X1 U27 ( .A(n44), .B(net148177), .Y(n3) );
  NAND2X1 U28 ( .A(n2), .B(n3), .Y(net163489) );
  NAND2X1 U29 ( .A(n227), .B(n72), .Y(n27) );
  INVXL U30 ( .A(prx_crcsidat[1]), .Y(n4) );
  INVXL U31 ( .A(n4), .Y(prx_fifowdat[5]) );
  INVXL U32 ( .A(prx_fifowdat[2]), .Y(n6) );
  INVXL U33 ( .A(prx_fifowdat[6]), .Y(n7) );
  INVXL U34 ( .A(n7), .Y(prx_crcsidat[2]) );
  INVXL U35 ( .A(prx_fifowdat[1]), .Y(n9) );
  INVXL U36 ( .A(prx_crcsidat[0]), .Y(n10) );
  INVXL U37 ( .A(n10), .Y(prx_fifowdat[4]) );
  XNOR2XL U38 ( .A(net167456), .B(ps_dat5b[2]), .Y(n12) );
  XNOR2X1 U39 ( .A(n13), .B(ps_dat5b[2]), .Y(n18) );
  OAI21BBX1 U40 ( .A(n18), .B(net148365), .C(net163489), .Y(N96) );
  NAND43X2 U41 ( .B(n14), .C(n15), .D(n16), .A(cctrans), .Y(n13) );
  INVX3 U42 ( .A(n13), .Y(net148177) );
  INVXL U43 ( .A(n17), .Y(n16) );
  INVXL U44 ( .A(shrtrans), .Y(n15) );
  NAND3XL U45 ( .A(net148388), .B(n17), .C(n15), .Y(n19) );
  INVXL U46 ( .A(net148388), .Y(n14) );
  BUFX1 U47 ( .A(cctrans), .Y(net169136) );
  MUX2BXL U48 ( .D0(shrtrans), .D1(n19), .S(net169136), .Y(net148389) );
  BUFXL U49 ( .A(N96), .Y(net169093) );
  NOR2X2 U50 ( .A(n83), .B(n24), .Y(n23) );
  INVXL U51 ( .A(net169093), .Y(net148351) );
  INVXL U52 ( .A(net148177), .Y(net167456) );
  INVX1 U53 ( .A(net167456), .Y(net167457) );
  BUFXL U54 ( .A(n227), .Y(n20) );
  GEN2X1 U55 ( .D(n61), .E(cccnt[4]), .C(cccnt[5]), .B(net169136), .A(
        net148177), .Y(n268) );
  NAND2X1 U56 ( .A(N96), .B(n269), .Y(n227) );
  NAND2XL U57 ( .A(n20), .B(n72), .Y(n22) );
  AND2X2 U58 ( .A(n27), .B(n23), .Y(prx_fifopsh) );
  AND2X4 U59 ( .A(n263), .B(n35), .Y(n24) );
  AND2XL U60 ( .A(n226), .B(net167457), .Y(N157) );
  INVX1 U61 ( .A(n250), .Y(prx_fsm[3]) );
  INVX1 U62 ( .A(n287), .Y(n250) );
  NAND21X1 U63 ( .B(n287), .A(n89), .Y(n256) );
  NOR32XL U64 ( .B(n261), .C(n287), .A(n260), .Y(n262) );
  MUX2IXL U65 ( .D0(net148412), .D1(n276), .S(ptx_txact), .Y(n30) );
  BUFXL U66 ( .A(prx_rcvdords[2]), .Y(n26) );
  BUFX3 U67 ( .A(prx_fifowdat[1]), .Y(prx_rxcode[1]) );
  BUFX3 U68 ( .A(prx_fifowdat[0]), .Y(prx_rxcode[0]) );
  BUFX3 U69 ( .A(prx_fifowdat[2]), .Y(prx_rxcode[2]) );
  INVXL U70 ( .A(n83), .Y(n28) );
  NAND32X1 U71 ( .B(bcnt[1]), .C(n224), .A(n69), .Y(n72) );
  NAND43X1 U72 ( .B(prx_fsm[0]), .C(prx_fsm[3]), .D(prx_fsm[2]), .A(prx_fsm[1]), .Y(n199) );
  NAND43XL U73 ( .B(cccnt[4]), .C(cccnt[3]), .D(n53), .A(cccnt[5]), .Y(n276)
         );
  INVXL U74 ( .A(prx_fsm[2]), .Y(n261) );
  XNOR2XL U75 ( .A(prx_fsm[0]), .B(prx_fsm[1]), .Y(n260) );
  INVXL U76 ( .A(r_pshords), .Y(n259) );
  NAND21XL U77 ( .B(n251), .A(n257), .Y(n236) );
  NAND21XL U78 ( .B(n269), .A(n230), .Y(n198) );
  NAND32XL U79 ( .B(n269), .C(n190), .A(n189), .Y(n228) );
  AND2XL U80 ( .A(n257), .B(prx_fifowdat[3]), .Y(N249) );
  AOI21XL U81 ( .B(n59), .C(n58), .A(n241), .Y(n31) );
  AOI32XL U82 ( .A(n237), .B(n270), .C(n285), .D(n177), .E(n175), .Y(n176) );
  NAND21XL U83 ( .B(n277), .A(n55), .Y(n58) );
  AND2XL U84 ( .A(cccnt[3]), .B(cccnt[2]), .Y(n61) );
  NAND32X1 U85 ( .B(n287), .C(n87), .A(n86), .Y(n219) );
  NAND2XL U86 ( .A(bcnt[0]), .B(n221), .Y(n40) );
  NAND21XL U87 ( .B(bcnt[0]), .A(n221), .Y(n223) );
  INVX1 U88 ( .A(n240), .Y(n193) );
  NAND21X1 U89 ( .B(n142), .A(n137), .Y(n148) );
  INVX1 U90 ( .A(n208), .Y(n180) );
  INVX1 U91 ( .A(n253), .Y(n254) );
  INVX1 U92 ( .A(N32), .Y(n178) );
  INVX1 U93 ( .A(n249), .Y(n272) );
  NAND2X1 U94 ( .A(n246), .B(n46), .Y(n240) );
  NAND32X1 U95 ( .B(pid_gobusy), .C(n240), .A(n239), .Y(N153) );
  INVX1 U96 ( .A(n232), .Y(n215) );
  INVX1 U97 ( .A(n144), .Y(n137) );
  INVX1 U98 ( .A(n239), .Y(n226) );
  INVX1 U99 ( .A(n141), .Y(n143) );
  NAND21X1 U100 ( .B(N251), .A(n249), .Y(N250) );
  INVX1 U101 ( .A(n106), .Y(n101) );
  INVX1 U102 ( .A(n48), .Y(n47) );
  INVX1 U103 ( .A(n48), .Y(n46) );
  NAND21X1 U104 ( .B(n251), .A(n252), .Y(n246) );
  INVX1 U105 ( .A(n251), .Y(n21) );
  NAND21X1 U106 ( .B(n10), .A(n136), .Y(n142) );
  NAND43X1 U107 ( .B(n165), .C(n171), .D(n167), .A(n166), .Y(n208) );
  AOI221XL U108 ( .A(n127), .B(n126), .C(n125), .D(n153), .E(n124), .Y(n165)
         );
  INVX1 U109 ( .A(n207), .Y(n124) );
  INVX1 U110 ( .A(n121), .Y(n125) );
  OR2X1 U111 ( .A(n202), .B(n183), .Y(n171) );
  NAND21X1 U112 ( .B(n140), .A(n209), .Y(n184) );
  GEN2XL U113 ( .D(n137), .E(n136), .C(n135), .B(n134), .A(n133), .Y(n140) );
  INVX1 U114 ( .A(n128), .Y(n135) );
  AND3X1 U115 ( .A(n141), .B(n10), .C(n132), .Y(n133) );
  AO21X1 U116 ( .B(n204), .C(n203), .A(n202), .Y(n206) );
  INVX1 U117 ( .A(n99), .Y(n136) );
  NAND2X1 U118 ( .A(n248), .B(n272), .Y(n253) );
  AO21X1 U119 ( .B(n179), .C(n171), .A(n168), .Y(N32) );
  NAND21X1 U120 ( .B(n180), .A(n166), .Y(n168) );
  INVX1 U121 ( .A(N31), .Y(n279) );
  INVX1 U122 ( .A(n160), .Y(n157) );
  NAND21X1 U123 ( .B(n251), .A(n237), .Y(n249) );
  NAND21X1 U124 ( .B(n178), .A(n174), .Y(n285) );
  INVX1 U125 ( .A(n174), .Y(n187) );
  OA21X1 U126 ( .B(n198), .C(n197), .A(n215), .Y(N277) );
  OA21X1 U127 ( .B(n177), .C(n197), .A(n215), .Y(N279) );
  NAND43X1 U128 ( .B(pid_goidle), .C(n252), .D(n251), .A(n46), .Y(n232) );
  OR3XL U129 ( .A(n83), .B(n240), .C(pid_gobusy), .Y(n239) );
  AO21X1 U130 ( .B(n134), .C(n131), .A(n137), .Y(n141) );
  NAND21X1 U131 ( .B(r_ordrs4), .A(n102), .Y(n144) );
  INVX1 U132 ( .A(n238), .Y(n221) );
  AO21X1 U133 ( .B(n127), .C(n131), .A(n137), .Y(n106) );
  NAND32X1 U134 ( .B(n21), .C(n48), .A(n238), .Y(N236) );
  INVX1 U135 ( .A(n236), .Y(N251) );
  INVX1 U136 ( .A(srstz), .Y(n48) );
  INVX1 U137 ( .A(n229), .Y(n255) );
  INVX1 U138 ( .A(pid_goidle), .Y(n191) );
  INVX1 U139 ( .A(n234), .Y(n194) );
  INVX1 U140 ( .A(n189), .Y(n177) );
  INVX1 U141 ( .A(n276), .Y(prx_cccnt[0]) );
  NAND32X1 U142 ( .B(n87), .C(n86), .A(n250), .Y(n188) );
  NAND32X1 U143 ( .B(n86), .C(n261), .A(n175), .Y(n84) );
  INVX1 U144 ( .A(n219), .Y(n269) );
  AND4XL U145 ( .A(net167457), .B(net148365), .C(net148378), .D(n77), .Y(n62)
         );
  INVX1 U146 ( .A(n79), .Y(n63) );
  INVX1 U147 ( .A(n119), .Y(prx_fifowdat[3]) );
  OR2X1 U148 ( .A(pff_txreq), .B(n30), .Y(n242) );
  AO21X1 U149 ( .B(n56), .C(net148391), .A(n48), .Y(N71) );
  INVX1 U150 ( .A(n241), .Y(n56) );
  NAND32X1 U151 ( .B(n242), .C(n48), .A(n241), .Y(N70) );
  OR2X1 U152 ( .A(n48), .B(n31), .Y(N76) );
  INVX1 U153 ( .A(n72), .Y(n73) );
  AND3X1 U154 ( .A(prx_eoprcvd), .B(pcc_rxgood), .C(n273), .Y(prx_setsta[3])
         );
  INVX1 U155 ( .A(n247), .Y(prx_eoprcvd) );
  NAND32X1 U156 ( .B(n246), .C(n250), .A(n275), .Y(n247) );
  AO21XL U157 ( .B(n21), .C(n269), .A(prx_setsta[6]), .Y(prx_fiforst) );
  INVX1 U158 ( .A(n264), .Y(prx_setsta[6]) );
  NAND32X1 U159 ( .B(n273), .C(n274), .A(prx_eoprcvd), .Y(n264) );
  INVX1 U160 ( .A(n82), .Y(n252) );
  GEN2XL U161 ( .D(n185), .E(n184), .C(n183), .B(n182), .A(n181), .Y(N31) );
  INVX1 U162 ( .A(n202), .Y(n182) );
  NAND21X1 U163 ( .B(n180), .A(n179), .Y(n181) );
  AO21X1 U164 ( .B(n255), .C(n21), .A(n254), .Y(prx_crcstart) );
  AND2X1 U165 ( .A(prx_crcsidat[1]), .B(prx_fifowdat[7]), .Y(n32) );
  NAND43X1 U166 ( .B(n212), .C(n211), .D(n210), .A(n209), .Y(n248) );
  INVX1 U167 ( .A(n200), .Y(n212) );
  INVX1 U168 ( .A(n201), .Y(n211) );
  OAI211X1 U169 ( .C(n208), .D(n207), .A(n206), .B(n205), .Y(n210) );
  NAND3X1 U170 ( .A(n33), .B(n205), .C(n113), .Y(n202) );
  NAND3X1 U171 ( .A(n106), .B(prx_crcsidat[0]), .C(n132), .Y(n33) );
  NAND21X1 U172 ( .B(prx_crcsidat[2]), .A(n32), .Y(n99) );
  NAND21X1 U173 ( .B(n184), .A(n185), .Y(n167) );
  NAND3X1 U174 ( .A(n34), .B(n204), .C(n118), .Y(n183) );
  NAND4X1 U175 ( .A(n116), .B(prx_crcsidat[0]), .C(n115), .D(n9), .Y(n34) );
  INVX1 U176 ( .A(n100), .Y(n116) );
  NAND32X1 U177 ( .B(n99), .C(n108), .A(prx_fifowdat[3]), .Y(n100) );
  AND2X1 U178 ( .A(n272), .B(n270), .Y(prx_setsta[1]) );
  OAI221X1 U179 ( .A(n120), .B(n121), .C(n161), .D(n142), .E(n152), .Y(n126)
         );
  INVX1 U180 ( .A(n156), .Y(n120) );
  OR2X1 U181 ( .A(n151), .B(n142), .Y(n121) );
  INVX1 U182 ( .A(n105), .Y(n132) );
  NAND21X1 U183 ( .B(n9), .A(n116), .Y(n105) );
  NAND43X1 U184 ( .B(n7), .C(n151), .D(prx_crcsidat[0]), .A(n32), .Y(n160) );
  AND2X1 U185 ( .A(n272), .B(n271), .Y(prx_setsta[2]) );
  AND4X1 U186 ( .A(n153), .B(n10), .C(n32), .D(prx_crcsidat[2]), .Y(n154) );
  INVX1 U187 ( .A(n270), .Y(n271) );
  INVX1 U188 ( .A(n164), .Y(n166) );
  OAI221X1 U189 ( .A(n163), .B(n162), .C(n161), .D(n160), .E(n200), .Y(n164)
         );
  AOI211X1 U190 ( .C(n157), .D(n156), .A(n155), .B(n154), .Y(n163) );
  INVX1 U191 ( .A(n152), .Y(n155) );
  INVX1 U192 ( .A(n75), .Y(n90) );
  OAI31XL U193 ( .A(n172), .B(n171), .C(n170), .D(n169), .Y(n174) );
  INVX1 U194 ( .A(n167), .Y(n172) );
  INVX1 U195 ( .A(n168), .Y(n169) );
  OAI31XL U196 ( .A(n252), .B(n251), .C(n250), .D(n253), .Y(prx_crcshfi4) );
  INVX1 U197 ( .A(n170), .Y(n179) );
  GEN2XL U198 ( .D(n196), .E(n285), .C(n228), .B(n215), .A(n195), .Y(N276) );
  AND4X1 U199 ( .A(n194), .B(n193), .C(n192), .D(n191), .Y(n195) );
  AND2X1 U200 ( .A(n271), .B(n237), .Y(n196) );
  INVX1 U201 ( .A(ptx_txact), .Y(n192) );
  OA21X1 U202 ( .B(n217), .C(n216), .A(n215), .Y(N278) );
  INVX1 U203 ( .A(n199), .Y(n217) );
  AOI211XL U204 ( .C(n248), .D(n270), .A(n213), .B(n256), .Y(n216) );
  INVX1 U205 ( .A(n285), .Y(n213) );
  NAND32X1 U206 ( .B(n255), .C(n190), .A(n176), .Y(n197) );
  AND2X1 U207 ( .A(prx_eoprcvd), .B(n274), .Y(prx_setsta[4]) );
  OAI22XL U208 ( .A(n186), .B(n188), .C(n279), .D(n256), .Y(N246) );
  OAI22XL U209 ( .A(n6), .B(n188), .C(n187), .D(n256), .Y(N248) );
  OAI22XL U210 ( .A(n9), .B(n188), .C(n178), .D(n256), .Y(N247) );
  NAND32X1 U211 ( .B(n139), .C(n123), .A(n122), .Y(n205) );
  NAND21X1 U212 ( .B(n9), .A(n111), .Y(n128) );
  NAND32X1 U213 ( .B(n122), .C(n123), .A(n127), .Y(n204) );
  OAI211X1 U214 ( .C(n220), .D(n219), .A(n265), .B(n218), .Y(n238) );
  INVX1 U215 ( .A(n266), .Y(n220) );
  AND3XL U216 ( .A(n47), .B(n28), .C(n251), .Y(n218) );
  NAND32X1 U217 ( .B(n146), .C(n139), .A(n186), .Y(n209) );
  NAND21X1 U218 ( .B(n286), .A(n98), .Y(n131) );
  OR3XL U219 ( .A(n186), .B(n149), .C(n146), .Y(n203) );
  NAND32X1 U220 ( .B(pid_goidle), .C(n240), .A(n235), .Y(N275) );
  OA22X1 U221 ( .A(ptx_txact), .B(n234), .C(n233), .D(n232), .Y(n235) );
  AND4XL U222 ( .A(n231), .B(n230), .C(n229), .D(n256), .Y(n233) );
  INVX1 U223 ( .A(n228), .Y(n231) );
  INVX1 U224 ( .A(n94), .Y(n111) );
  NAND32X1 U225 ( .B(n144), .C(n108), .A(prx_fifowdat[3]), .Y(n94) );
  INVX1 U226 ( .A(n110), .Y(n159) );
  INVX1 U227 ( .A(n149), .Y(n134) );
  INVX1 U228 ( .A(n98), .Y(n102) );
  INVX1 U229 ( .A(n223), .Y(n281) );
  OR2X1 U230 ( .A(n161), .B(n151), .Y(n152) );
  NAND32X1 U231 ( .B(n162), .C(n123), .A(n122), .Y(n207) );
  AOI21BBXL U232 ( .B(prx_crcsidat[0]), .C(n38), .A(n20), .Y(k0_det) );
  AO21X1 U233 ( .B(n114), .C(n131), .A(n137), .Y(n115) );
  INVX1 U234 ( .A(n139), .Y(n114) );
  INVX1 U235 ( .A(n112), .Y(n127) );
  INVX1 U236 ( .A(n161), .Y(n153) );
  INVX1 U237 ( .A(pcc_rxgood), .Y(n274) );
  NAND5XL U238 ( .A(n127), .B(n159), .C(n102), .D(n6), .E(n186), .Y(n201) );
  NAND21XL U239 ( .B(n250), .A(n89), .Y(n229) );
  INVXL U240 ( .A(n256), .Y(n237) );
  NAND21X1 U241 ( .B(n265), .A(pid_gobusy), .Y(n234) );
  INVX1 U242 ( .A(n88), .Y(n190) );
  NAND32X1 U243 ( .B(n87), .C(n198), .A(n86), .Y(n88) );
  INVX1 U244 ( .A(n85), .Y(n230) );
  NAND21XL U245 ( .B(n257), .A(n199), .Y(n85) );
  NAND32X1 U246 ( .B(n250), .C(n86), .A(n261), .Y(n189) );
  AND4XL U247 ( .A(n269), .B(n28), .C(n267), .D(n266), .Y(prx_setsta[0]) );
  INVX1 U248 ( .A(n265), .Y(prx_idle) );
  INVXL U249 ( .A(cccnt[2]), .Y(net148392) );
  OA21X1 U250 ( .B(n277), .C(n60), .A(n59), .Y(net148394) );
  INVXL U251 ( .A(cccnt[3]), .Y(n60) );
  AOI21X1 U252 ( .B(cccnt[2]), .C(cccnt[1]), .A(cccnt[5]), .Y(net162096) );
  NAND21XL U253 ( .B(n278), .A(cccnt[2]), .Y(n53) );
  NAND21XL U254 ( .B(net148391), .A(cccnt[1]), .Y(n278) );
  NAND21X1 U255 ( .B(net148365), .A(prx_bmc), .Y(n91) );
  NAND31XL U256 ( .C(cccnt[3]), .A(n36), .B(net162096), .Y(net148388) );
  AOI21XL U257 ( .B(cccnt[2]), .C(cccnt[0]), .A(cccnt[4]), .Y(n36) );
  INVXL U258 ( .A(cccnt[5]), .Y(n59) );
  INVXL U259 ( .A(prx_bmc), .Y(n80) );
  INVXL U260 ( .A(ps_dat5b[2]), .Y(net148378) );
  INVXL U261 ( .A(ps_dat5b[0]), .Y(n77) );
  INVX1 U262 ( .A(bcnt[0]), .Y(n69) );
  INVXL U263 ( .A(prx_fsm[0]), .Y(n175) );
  NAND21X1 U264 ( .B(n68), .A(n67), .Y(prx_crcsidat[0]) );
  AO21XL U265 ( .B(n66), .C(n70), .A(n77), .Y(n67) );
  MUX2XL U266 ( .D0(n63), .D1(n62), .S(prx_bmc), .Y(n68) );
  MUX2XL U267 ( .D0(n65), .D1(n75), .S(net167457), .Y(n66) );
  NAND32XL U268 ( .B(net167457), .C(net148378), .A(ps_dat5b[1]), .Y(n79) );
  MUX2IXL U269 ( .D0(prx_rxcode[4]), .D1(prx_rxcode[3]), .S(n287), .Y(n119) );
  NAND21XL U270 ( .B(ps_dat5b[2]), .A(ps_dat5b[1]), .Y(n75) );
  NAND21XL U271 ( .B(n74), .A(prx_bmc), .Y(n65) );
  INVX1 U272 ( .A(n64), .Y(n74) );
  NAND21XL U273 ( .B(ps_dat5b[1]), .A(ps_dat5b[2]), .Y(n64) );
  AO21XL U274 ( .B(n50), .C(cccnt[5]), .A(n242), .Y(n241) );
  INVX1 U275 ( .A(n58), .Y(n50) );
  AO21X1 U276 ( .B(n56), .C(n51), .A(n48), .Y(N72) );
  XOR2XL U277 ( .A(cccnt[1]), .B(cccnt[0]), .Y(n51) );
  AO21X1 U278 ( .B(n57), .C(n56), .A(n48), .Y(N75) );
  XOR2XL U279 ( .A(cccnt[4]), .B(n55), .Y(n57) );
  XNOR2XL U280 ( .A(cccnt[3]), .B(n53), .Y(n54) );
  XNOR2XL U281 ( .A(cccnt[2]), .B(n278), .Y(n52) );
  OR2X1 U282 ( .A(n81), .B(n37), .Y(prx_crcsidat[1]) );
  AOI21XL U283 ( .B(ps_dat5b[0]), .C(n80), .A(n79), .Y(n37) );
  INVX1 U284 ( .A(n93), .Y(prx_crcsidat[3]) );
  GEN2XL U285 ( .D(prx_bmc), .E(ps_dat5b[2]), .C(ps_dat5b[1]), .B(n91), .A(n90), .Y(n92) );
  AND2XL U286 ( .A(n81), .B(prx_bmc), .Y(n38) );
  OAI22X1 U287 ( .A(n78), .B(n80), .C(n77), .D(n79), .Y(prx_fifowdat[6]) );
  MUX2XL U288 ( .D0(ps_dat5b[1]), .D1(n74), .S(net167457), .Y(n76) );
  MUX2X1 U289 ( .D0(n282), .D1(n173), .S(n187), .Y(n270) );
  MUX2X1 U290 ( .D0(n283), .D1(n284), .S(n178), .Y(n173) );
  MUX4X1 U291 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[4]), .D2(r_ords_ena[5]), 
        .D3(r_ords_ena[6]), .S0(N31), .S1(N32), .Y(n282) );
  NOR21XL U292 ( .B(r_ords_ena[0]), .A(n279), .Y(n284) );
  INVX1 U293 ( .A(n150), .Y(n185) );
  OAI211X1 U294 ( .C(n149), .D(n148), .A(n147), .B(n203), .Y(n150) );
  NAND5XL U295 ( .A(prx_fifowdat[1]), .B(prx_fifowdat[2]), .C(prx_fifowdat[3]), 
        .D(n145), .E(n186), .Y(n147) );
  OAI22X1 U296 ( .A(n149), .B(n144), .C(n143), .D(n142), .Y(n145) );
  MUX2X1 U297 ( .D0(r_ords_ena[1]), .D1(r_ords_ena[2]), .S(N31), .Y(n283) );
  OAI211X1 U298 ( .C(n104), .D(n112), .A(n103), .B(n201), .Y(n170) );
  AOI31X1 U299 ( .A(n136), .B(n10), .C(n137), .D(n95), .Y(n104) );
  NAND43X1 U300 ( .B(prx_rxcode[1]), .C(n101), .D(prx_crcsidat[0]), .A(n116), 
        .Y(n103) );
  INVX1 U301 ( .A(n117), .Y(n95) );
  MUX3XL U302 ( .D0(n245), .D1(n244), .D2(n243), .S0(prx_rcvdords[2]), .S1(
        prx_rcvdords[0]), .Y(n275) );
  AND2XL U303 ( .A(r_ords_ena[1]), .B(prx_rcvdords[1]), .Y(n245) );
  MUX2XL U304 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[5]), .S(prx_rcvdords[1]), 
        .Y(n244) );
  MUX4XL U305 ( .D0(r_ords_ena[0]), .D1(r_ords_ena[4]), .D2(r_ords_ena[2]), 
        .D3(r_ords_ena[6]), .S0(prx_rcvdords[2]), .S1(prx_rcvdords[1]), .Y(
        n243) );
  INVX1 U306 ( .A(r_rgdcrc), .Y(n273) );
  NAND43X1 U307 ( .B(ordsbuf[4]), .C(n130), .D(n129), .A(ordsbuf[5]), .Y(n149)
         );
  NAND43X1 U308 ( .B(prx_fifowdat[1]), .C(n119), .D(n6), .A(prx_fifowdat[0]), 
        .Y(n151) );
  NAND21XL U309 ( .B(prx_rcvdords[2]), .A(n39), .Y(n98) );
  NAND32X1 U310 ( .B(n119), .C(r_exist1st), .A(prx_rxcode[1]), .Y(n110) );
  NAND2XL U311 ( .A(ordsbuf[3]), .B(prx_rcvdords[0]), .Y(n109) );
  NOR2XL U312 ( .A(prx_rcvdords[1]), .B(n109), .Y(n39) );
  OR4XL U313 ( .A(prx_rcvdords[2]), .B(n110), .C(n109), .D(n108), .Y(n123) );
  NAND6XL U314 ( .A(prx_rcvdords[2]), .B(prx_rcvdords[1]), .C(ordsbuf[3]), .D(
        n159), .E(n6), .F(n138), .Y(n146) );
  INVXL U315 ( .A(prx_rcvdords[0]), .Y(n138) );
  MUX2AXL U316 ( .D0(n40), .D1(n281), .S(bcnt[1]), .Y(N238) );
  AND2XL U317 ( .A(n226), .B(prx_bmc), .Y(N156) );
  AND2XL U318 ( .A(n226), .B(ps_dat5b[1]), .Y(N154) );
  AND2XL U319 ( .A(n226), .B(ps_dat5b[2]), .Y(N155) );
  OAI22XL U320 ( .A(n225), .B(n238), .C(n224), .D(n223), .Y(N239) );
  MUX2XL U321 ( .D0(n224), .D1(n222), .S(bcnt[1]), .Y(n225) );
  NAND21XL U322 ( .B(bcnt[2]), .A(bcnt[0]), .Y(n222) );
  INVX1 U323 ( .A(ordsbuf[6]), .Y(n129) );
  INVX1 U324 ( .A(ordsbuf[7]), .Y(n130) );
  NAND21X1 U325 ( .B(prx_fifowdat[2]), .A(prx_fifowdat[0]), .Y(n108) );
  NAND43X1 U326 ( .B(ordsbuf[5]), .C(n130), .D(n129), .A(ordsbuf[4]), .Y(n162)
         );
  NAND2X1 U327 ( .A(ordsbuf[5]), .B(n107), .Y(n139) );
  NAND31XL U328 ( .C(r_ordrs4), .A(n26), .B(n39), .Y(n161) );
  NAND21X1 U329 ( .B(ordsbuf[5]), .A(n107), .Y(n112) );
  OAI21BBXL U330 ( .A(n39), .B(prx_rcvdords[2]), .C(r_ordrs4), .Y(n156) );
  NAND21X1 U331 ( .B(prx_rxcode[1]), .A(n111), .Y(n117) );
  NAND6XL U332 ( .A(prx_rxcode[2]), .B(n26), .C(n39), .D(n159), .E(n158), .F(
        n186), .Y(n200) );
  INVX1 U333 ( .A(n162), .Y(n158) );
  NOR5XL U334 ( .A(cccnt[3]), .B(cccnt[2]), .C(cccnt[5]), .D(n278), .E(n277), 
        .Y(prx_cccnt[1]) );
  INVX1 U335 ( .A(n97), .Y(n107) );
  NAND32X1 U336 ( .B(n96), .C(n130), .A(n129), .Y(n97) );
  INVX1 U337 ( .A(ordsbuf[4]), .Y(n96) );
  INVX1 U338 ( .A(prx_fifowdat[0]), .Y(n186) );
  INVXL U339 ( .A(prx_rcvdords[1]), .Y(n122) );
  AND3XL U340 ( .A(pid_goidle), .B(prx_fsm[3]), .C(n275), .Y(prx_setsta[5]) );
  INVX1 U341 ( .A(n49), .Y(n55) );
  NAND21XL U342 ( .B(n53), .A(cccnt[3]), .Y(n49) );
  NAND43X1 U343 ( .B(prx_fsm[0]), .C(prx_fsm[1]), .D(prx_fsm[2]), .A(n250), 
        .Y(n265) );
  OR2XL U344 ( .A(bcnt[2]), .B(bcnt[1]), .Y(n266) );
  MUX2XL U345 ( .D0(net169093), .D1(prx_crcsidat[3]), .S(prx_fsm[3]), .Y(
        prx_fifowdat[7]) );
  NAND32XL U346 ( .B(net167456), .C(net148378), .A(n91), .Y(n70) );
  NAND21XL U347 ( .B(net167456), .A(n92), .Y(n93) );
  OAI31XL U348 ( .A(ps_dat5b[1]), .B(net167456), .C(n77), .D(n70), .Y(n81) );
  XOR2XL U349 ( .A(net167456), .B(prx_bmc), .Y(n267) );
  INVXL U350 ( .A(net169136), .Y(net148412) );
  AOI211XL U351 ( .C(n12), .D(ps_dat5b[0]), .A(n76), .B(n90), .Y(n78) );
  NAND43X1 U352 ( .B(net148351), .C(n7), .D(prx_fifowdat[5]), .A(n10), .Y(n82)
         );
  OAI31XL U353 ( .A(prx_crcsidat[0]), .B(n73), .C(n38), .D(n29), .Y(n251) );
  NOR2X1 U354 ( .A(n279), .B(n285), .Y(prx_rst[0]) );
  NOR2X1 U355 ( .A(N31), .B(n285), .Y(prx_rst[1]) );
  INVX1 U356 ( .A(r_ordrs4), .Y(n286) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_adp ( clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, 
        r_adprx_en, r_adp2nd, adp_val, d_cc, cctrans );
  output [5:0] adp_val;
  input clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, r_adprx_en,
         r_adp2nd;
  output d_cc, cctrans;
  wire   N49, N50, N51, N52, N53, N55, N97, N98, N99, N100, N101, N102, N103,
         N104, N106, N107, N108, N109, N110, N111, N112, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N169, N170, N171, N172, N173, net10744, net10750,
         net10755, net10760, n115, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7;
  wire   [7:0] dcnt_h;
  wire   [5:0] adp_v0;
  wire   [3:0] dcnt_n;
  wire   [5:0] dcnt_e;

  SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 clk_gate_adp_n_reg ( .CLK(clk), .EN(N49), 
        .ENCLK(net10744), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 clk_gate_dcnt_e_reg ( .CLK(clk), .EN(N130), 
        .ENCLK(net10750), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 clk_gate_dcnt_h_reg ( .CLK(clk), .EN(N137), 
        .ENCLK(net10755), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 clk_gate_dcnt_n_reg ( .CLK(clk), .EN(N169), 
        .ENCLK(net10760), .TE(1'b0) );
  phyrx_adp_DW01_inc_0 add_385 ( .A({n8, dcnt_h[6:0]}), .SUM({N104, N103, N102, 
        N101, N100, N99, N98, N97}) );
  phyrx_adp_DW_div_tc_6 div_338 ( .a({dcnt_h[7], n8, dcnt_h[6:0]}), .b({1'b0, 
        1'b1, 1'b1, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, adp_v0}), .remainder({
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7}), .divide_by_0() );
  DFFQX1 adp_n_reg_5_ ( .D(N55), .C(net10744), .Q(adp_val[5]) );
  DFFQX1 dcnt_h_reg_6_ ( .D(N144), .C(net10755), .Q(dcnt_h[6]) );
  DFFQX1 dcnt_h_reg_3_ ( .D(N141), .C(net10755), .Q(dcnt_h[3]) );
  DFFQX1 dcnt_h_reg_4_ ( .D(N142), .C(net10755), .Q(dcnt_h[4]) );
  DFFQX1 dcnt_h_reg_5_ ( .D(N143), .C(net10755), .Q(dcnt_h[5]) );
  DFFQX1 dcnt_h_reg_1_ ( .D(N139), .C(net10755), .Q(dcnt_h[1]) );
  DFFQX1 dcnt_h_reg_2_ ( .D(N140), .C(net10755), .Q(dcnt_h[2]) );
  DFFQX1 dcnt_h_reg_0_ ( .D(N138), .C(net10755), .Q(dcnt_h[0]) );
  DFFQX1 dcnt_h_reg_7_ ( .D(N145), .C(net10755), .Q(dcnt_h[7]) );
  DFFQX1 dcnt_n_reg_2_ ( .D(N172), .C(net10760), .Q(dcnt_n[2]) );
  DFFQX1 dcnt_n_reg_0_ ( .D(N170), .C(net10760), .Q(dcnt_n[0]) );
  DFFQX1 dcnt_e_reg_3_ ( .D(N134), .C(net10750), .Q(dcnt_e[3]) );
  DFFQX1 dcnt_n_reg_1_ ( .D(N171), .C(net10760), .Q(dcnt_n[1]) );
  DFFQX1 adp_n_reg_3_ ( .D(N53), .C(net10744), .Q(adp_val[3]) );
  DFFQX1 adp_n_reg_1_ ( .D(N51), .C(net10744), .Q(adp_val[1]) );
  DFFQX1 adp_n_reg_2_ ( .D(N52), .C(net10744), .Q(adp_val[2]) );
  DFFQX1 adp_n_reg_4_ ( .D(n110), .C(net10744), .Q(adp_val[4]) );
  DFFQX1 adp_n_reg_0_ ( .D(N50), .C(net10744), .Q(adp_val[0]) );
  DFFQX1 cs_d_cc_reg ( .D(n115), .C(clk), .Q(d_cc) );
  DFFQX1 dcnt_e_reg_0_ ( .D(N131), .C(net10750), .Q(dcnt_e[0]) );
  DFFQX1 dcnt_n_reg_3_ ( .D(N173), .C(net10760), .Q(dcnt_n[3]) );
  DFFQX1 dcnt_e_reg_1_ ( .D(N132), .C(net10750), .Q(dcnt_e[1]) );
  DFFQX1 dcnt_e_reg_5_ ( .D(N136), .C(net10750), .Q(dcnt_e[5]) );
  DFFQX1 dcnt_e_reg_2_ ( .D(N133), .C(net10750), .Q(dcnt_e[2]) );
  DFFQX1 dcnt_e_reg_4_ ( .D(N135), .C(net10750), .Q(dcnt_e[4]) );
  AND2X2 U3 ( .A(n1), .B(golo), .Y(n32) );
  OR3X4 U4 ( .A(golo), .B(n5), .C(n89), .Y(n28) );
  INVX1 U5 ( .A(adp_val[2]), .Y(n22) );
  OR2XL U6 ( .A(n104), .B(n106), .Y(n6) );
  NAND42X1 U7 ( .C(adp_val[1]), .D(adp_val[3]), .A(n22), .B(n20), .Y(n21) );
  INVX1 U8 ( .A(adp_val[0]), .Y(n20) );
  INVX1 U9 ( .A(dcnt_e[4]), .Y(n19) );
  NOR3XL U10 ( .A(dcnt_e[4]), .B(n84), .C(dcnt_e[0]), .Y(n14) );
  NAND42X1 U11 ( .C(n25), .D(n24), .A(n9), .B(n23), .Y(n97) );
  AND2X1 U12 ( .A(d_cc), .B(n4), .Y(n1) );
  INVX1 U13 ( .A(adp_val[4]), .Y(n4) );
  INVX1 U14 ( .A(dcnt_e[0]), .Y(n77) );
  INVX1 U15 ( .A(d_cc), .Y(n89) );
  NAND2X1 U16 ( .A(n104), .B(n21), .Y(n62) );
  INVX1 U17 ( .A(n62), .Y(n5) );
  NAND31X2 U18 ( .C(n29), .A(n28), .B(n27), .Y(n30) );
  NOR32X2 U19 ( .B(n89), .C(n62), .A(gohi), .Y(n29) );
  AND3X1 U20 ( .A(gohi), .B(adp_val[4]), .C(n89), .Y(n31) );
  BUFXL U21 ( .A(gohi), .Y(n2) );
  BUFXL U22 ( .A(golo), .Y(n3) );
  AND2X2 U23 ( .A(n107), .B(n6), .Y(cctrans) );
  BUFXL U24 ( .A(n107), .Y(n7) );
  NAND32X1 U25 ( .B(n31), .C(n32), .A(n30), .Y(n107) );
  BUFX3 U26 ( .A(dcnt_h[7]), .Y(n8) );
  NAND31XL U27 ( .C(n71), .A(n97), .B(n63), .Y(n70) );
  XOR2X1 U28 ( .A(dcnt_n[0]), .B(adp_val[0]), .Y(n24) );
  NAND32XL U29 ( .B(n87), .C(n88), .A(n89), .Y(n86) );
  NAND32XL U30 ( .B(n89), .C(n88), .A(n99), .Y(n90) );
  NOR43XL U31 ( .B(dcnt_e[3]), .C(dcnt_e[2]), .D(dcnt_e[4]), .A(n105), .Y(n106) );
  XNOR2XL U32 ( .A(dcnt_n[3]), .B(adp_val[3]), .Y(n9) );
  XOR2X1 U33 ( .A(n19), .B(dcnt_e[5]), .Y(n81) );
  OR4XL U34 ( .A(dcnt_e[3]), .B(n101), .C(n100), .D(n10), .Y(n87) );
  OAI222XL U35 ( .A(dcnt_e[4]), .B(n108), .C(n85), .D(n105), .E(dcnt_e[0]), 
        .F(n84), .Y(n10) );
  NOR21XL U36 ( .B(n98), .A(n11), .Y(N173) );
  XNOR2XL U37 ( .A(n74), .B(n73), .Y(n11) );
  OR2X1 U38 ( .A(n111), .B(n121), .Y(n12) );
  INVX1 U39 ( .A(srstz), .Y(n18) );
  NAND21X1 U40 ( .B(n36), .A(n122), .Y(n40) );
  NAND21X1 U41 ( .B(n61), .A(n126), .Y(n36) );
  NOR21XL U42 ( .B(n40), .A(n39), .Y(n60) );
  MUX2IX1 U43 ( .D0(n38), .D1(n37), .S(n122), .Y(n39) );
  NAND21X1 U44 ( .B(n121), .A(n36), .Y(n38) );
  INVX1 U45 ( .A(n61), .Y(n111) );
  INVX1 U46 ( .A(n37), .Y(n121) );
  INVX1 U47 ( .A(n128), .Y(n88) );
  XOR2X1 U48 ( .A(n41), .B(n123), .Y(n59) );
  NAND21X1 U49 ( .B(n121), .A(n40), .Y(n41) );
  INVX1 U50 ( .A(adp_v0[4]), .Y(n113) );
  NAND32X1 U51 ( .B(n125), .C(adp_v0[0]), .A(n124), .Y(n61) );
  OAI21BX1 U52 ( .C(adp_v0[4]), .B(n125), .A(n124), .Y(n37) );
  INVX1 U53 ( .A(n76), .Y(n50) );
  NAND21X1 U54 ( .B(n18), .A(n5), .Y(n71) );
  INVX1 U55 ( .A(n70), .Y(n98) );
  NAND21X1 U56 ( .B(n14), .A(n81), .Y(n104) );
  NAND21X1 U57 ( .B(n62), .A(n26), .Y(n27) );
  NAND21X1 U58 ( .B(n97), .A(n69), .Y(n26) );
  AND2X1 U59 ( .A(n60), .B(n109), .Y(N52) );
  AND2X1 U60 ( .A(n109), .B(n59), .Y(N53) );
  MUX2BXL U61 ( .D0(n58), .D1(n57), .S(n126), .Y(N51) );
  NAND21X1 U62 ( .B(n111), .A(n110), .Y(n57) );
  AND2X1 U63 ( .A(n109), .B(n12), .Y(n58) );
  INVX1 U64 ( .A(n56), .Y(n110) );
  NAND21X1 U65 ( .B(n121), .A(n109), .Y(n56) );
  AND2X1 U66 ( .A(n109), .B(n61), .Y(N50) );
  AO21X1 U67 ( .B(n78), .C(n112), .A(n88), .Y(n76) );
  AO21X1 U68 ( .B(n80), .C(n79), .A(k0_det), .Y(n101) );
  INVX1 U69 ( .A(n82), .Y(n79) );
  AO21X1 U70 ( .B(n78), .C(n77), .A(n76), .Y(N131) );
  OR2X1 U71 ( .A(n76), .B(n13), .Y(N132) );
  AOI21X1 U72 ( .B(n34), .C(n105), .A(n52), .Y(n13) );
  INVX1 U73 ( .A(n86), .Y(n103) );
  INVX1 U74 ( .A(n87), .Y(n99) );
  INVX1 U75 ( .A(n90), .Y(n102) );
  INVX1 U76 ( .A(n52), .Y(n78) );
  OAI31XL U77 ( .A(n52), .B(n51), .C(n108), .D(n50), .Y(N136) );
  NAND21X1 U78 ( .B(n94), .A(n93), .Y(n129) );
  INVX1 U79 ( .A(n91), .Y(n94) );
  INVX1 U80 ( .A(n92), .Y(n93) );
  INVX1 U81 ( .A(n83), .Y(n100) );
  NAND32X1 U82 ( .B(n84), .C(n82), .A(n81), .Y(n83) );
  NAND42X1 U83 ( .C(n98), .D(n18), .A(n97), .B(n96), .Y(N169) );
  NAND21X1 U84 ( .B(n95), .A(n5), .Y(n96) );
  NAND21X1 U85 ( .B(n109), .A(srstz), .Y(N49) );
  AND2X1 U86 ( .A(n109), .B(n108), .Y(N55) );
  NAND31X1 U87 ( .C(n64), .A(n67), .B(n74), .Y(n63) );
  AND3X1 U88 ( .A(n98), .B(n72), .C(n64), .Y(N171) );
  NAND32X1 U89 ( .B(n77), .C(n19), .A(n54), .Y(n33) );
  INVX1 U90 ( .A(n84), .Y(n54) );
  INVX1 U91 ( .A(n43), .Y(n80) );
  INVX1 U92 ( .A(n46), .Y(n35) );
  INVX1 U93 ( .A(n49), .Y(n47) );
  XOR2X1 U94 ( .A(n22), .B(dcnt_n[2]), .Y(n23) );
  XOR2X1 U95 ( .A(dcnt_n[1]), .B(adp_val[1]), .Y(n25) );
  OR3XL U96 ( .A(dcnt_e[3]), .B(dcnt_e[2]), .C(dcnt_e[1]), .Y(n84) );
  XOR2X1 U97 ( .A(n89), .B(adp_val[4]), .Y(n69) );
  NAND21XL U98 ( .B(n77), .A(dcnt_e[1]), .Y(n105) );
  GEN2XL U99 ( .D(dcnt_e[3]), .E(n46), .C(n47), .B(n78), .A(n45), .Y(N134) );
  OAI31XL U100 ( .A(n44), .B(n43), .C(n92), .D(n50), .Y(n45) );
  AOI211X1 U101 ( .C(n42), .D(n61), .A(n60), .B(n59), .Y(n44) );
  MUX2X1 U102 ( .D0(n12), .D1(n37), .S(n126), .Y(n42) );
  NAND31X1 U103 ( .C(n101), .A(n15), .B(n128), .Y(N137) );
  AOI21XL U104 ( .B(n100), .C(dcnt_e[0]), .A(n99), .Y(n15) );
  AO21X1 U105 ( .B(k0_det), .C(r_adprx_en), .A(n82), .Y(n92) );
  INVXL U106 ( .A(dcnt_e[2]), .Y(n85) );
  OR3XL U107 ( .A(n80), .B(n92), .C(n16), .Y(n52) );
  OAI21X1 U108 ( .B(r_adp2nd), .C(n33), .A(n91), .Y(n16) );
  GEN2XL U109 ( .D(dcnt_e[4]), .E(n49), .C(n51), .B(n78), .A(n76), .Y(N135) );
  GEN2XL U110 ( .D(dcnt_e[2]), .E(n34), .C(n35), .B(n78), .A(n76), .Y(N133) );
  AO22X1 U111 ( .A(N111), .B(n103), .C(N103), .D(n102), .Y(N144) );
  AO22X1 U112 ( .A(N110), .B(n103), .C(N102), .D(n102), .Y(N143) );
  AO22X1 U113 ( .A(N109), .B(n103), .C(N101), .D(n102), .Y(N142) );
  AO22X1 U114 ( .A(N108), .B(n103), .C(N100), .D(n102), .Y(N141) );
  AO22X1 U115 ( .A(N107), .B(n103), .C(N99), .D(n102), .Y(N140) );
  AO22X1 U116 ( .A(N106), .B(n103), .C(N98), .D(n102), .Y(N139) );
  AO22X1 U117 ( .A(N112), .B(n103), .C(N104), .D(n102), .Y(N145) );
  AO22AXL U118 ( .A(N97), .B(n102), .C(n103), .D(dcnt_h[0]), .Y(N138) );
  INVX1 U119 ( .A(n55), .Y(n109) );
  NAND5XL U120 ( .A(dcnt_e[0]), .B(srstz), .C(n54), .D(n81), .E(n53), .Y(n55)
         );
  NAND6XL U121 ( .A(n69), .B(n68), .C(n74), .D(n67), .E(n66), .F(n65), .Y(n95)
         );
  INVXL U122 ( .A(dcnt_n[0]), .Y(n65) );
  AND2X1 U123 ( .A(n75), .B(srstz), .Y(n115) );
  OAI22XL U124 ( .A(n71), .B(n95), .C(dcnt_n[0]), .D(n70), .Y(N170) );
  AND2X1 U125 ( .A(n98), .B(n17), .Y(N172) );
  XNOR2XL U126 ( .A(dcnt_n[2]), .B(n72), .Y(n17) );
  NAND21XL U127 ( .B(n72), .A(dcnt_n[2]), .Y(n73) );
  OR2XL U128 ( .A(dcnt_e[5]), .B(n33), .Y(n43) );
  NAND21XL U129 ( .B(dcnt_e[5]), .A(n14), .Y(n91) );
  NAND21XL U130 ( .B(dcnt_e[1]), .A(n77), .Y(n34) );
  OR2XL U131 ( .A(dcnt_e[2]), .B(n34), .Y(n46) );
  NAND21XL U132 ( .B(dcnt_e[3]), .A(n35), .Y(n49) );
  NAND21XL U133 ( .B(n66), .A(dcnt_n[0]), .Y(n72) );
  NAND21XL U134 ( .B(dcnt_n[0]), .A(n66), .Y(n64) );
  INVXL U135 ( .A(dcnt_n[1]), .Y(n66) );
  INVXL U136 ( .A(dcnt_e[5]), .Y(n108) );
  INVX1 U137 ( .A(n48), .Y(n51) );
  NAND21XL U138 ( .B(dcnt_e[4]), .A(n47), .Y(n48) );
  INVX1 U139 ( .A(r_adprx_en), .Y(n112) );
  INVXL U140 ( .A(dcnt_n[2]), .Y(n67) );
  INVXL U141 ( .A(dcnt_n[3]), .Y(n74) );
  XOR2XL U142 ( .A(n7), .B(d_cc), .Y(n75) );
  NAND21XL U143 ( .B(i_ccidle), .A(n7), .Y(n82) );
  MUX2XL U144 ( .D0(n2), .D1(n3), .S(adp_val[4]), .Y(n68) );
  MUX2XL U145 ( .D0(n2), .D1(n3), .S(d_cc), .Y(n53) );
  OR2X1 U146 ( .A(dcnt_h[1]), .B(dcnt_h[0]), .Y(n114) );
  OAI21BBX1 U147 ( .A(dcnt_h[0]), .B(dcnt_h[1]), .C(n114), .Y(N106) );
  OR2X1 U148 ( .A(n114), .B(dcnt_h[2]), .Y(n116) );
  OAI21BBX1 U149 ( .A(n114), .B(dcnt_h[2]), .C(n116), .Y(N107) );
  OR2X1 U150 ( .A(n116), .B(dcnt_h[3]), .Y(n117) );
  OAI21BBX1 U151 ( .A(n116), .B(dcnt_h[3]), .C(n117), .Y(N108) );
  OR2X1 U152 ( .A(n117), .B(dcnt_h[4]), .Y(n118) );
  OAI21BBX1 U153 ( .A(n117), .B(dcnt_h[4]), .C(n118), .Y(N109) );
  OR2X1 U154 ( .A(n118), .B(dcnt_h[5]), .Y(n119) );
  OAI21BBX1 U155 ( .A(n118), .B(dcnt_h[5]), .C(n119), .Y(N110) );
  XNOR2XL U156 ( .A(n119), .B(dcnt_h[6]), .Y(N111) );
  OR2X1 U157 ( .A(dcnt_h[6]), .B(n119), .Y(n120) );
  XNOR2XL U158 ( .A(n8), .B(n120), .Y(N112) );
  AOI21X1 U159 ( .B(adp_v0[3]), .C(n124), .A(n125), .Y(n123) );
  OAI21X1 U160 ( .B(adp_v0[2]), .C(n125), .A(n124), .Y(n122) );
  OAI21X1 U161 ( .B(adp_v0[1]), .C(n125), .A(n124), .Y(n126) );
  OAI21X1 U162 ( .B(n127), .C(n113), .A(adp_v0[5]), .Y(n124) );
  NOR3XL U163 ( .A(adp_v0[1]), .B(adp_v0[3]), .C(adp_v0[2]), .Y(n127) );
  NOR2X1 U164 ( .A(n113), .B(adp_v0[5]), .Y(n125) );
  OAI2B11X1 U165 ( .D(k0_det), .C(n112), .A(n129), .B(n128), .Y(N130) );
  NOR3XL U166 ( .A(goidle), .B(gobusy), .C(n18), .Y(n128) );
endmodule


module phyrx_adp_DW_div_tc_6 ( a, b, quotient, remainder, divide_by_0 );
  input [8:0] a;
  input [3:0] b;
  output [8:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   u_div_SumTmp_1__0_, u_div_SumTmp_1__2_, u_div_SumTmp_2__0_,
         u_div_SumTmp_3__0_, u_div_SumTmp_4__0_, u_div_SumTmp_5__0_,
         u_div_CryTmp_0__2_, u_div_CryTmp_0__3_, u_div_CryTmp_0__4_,
         u_div_CryTmp_1__2_, u_div_CryTmp_1__4_, u_div_CryTmp_2__4_,
         u_div_CryTmp_3__4_, u_div_CryTmp_4__4_, u_div_CryTmp_5__4_,
         u_div_PartRem_1__2_, u_div_PartRem_1__3_, u_div_PartRem_2__2_,
         u_div_PartRem_2__3_, u_div_PartRem_3__2_, u_div_PartRem_3__3_,
         u_div_PartRem_4__2_, u_div_PartRem_4__3_, u_div_PartRem_5__2_,
         u_div_PartRem_5__3_, u_div_PartRem_7__0_, u_div_PartRem_7__1_, n1, n2,
         n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22;
  wire   [5:1] u_div_QIncCry;
  wire   [5:0] u_div_QInv;
  wire   [6:1] u_div_AIncCry;
  wire   [6:0] u_div_AInv;

  HAD1X1 u_div_u_ha_AInc_6 ( .A(u_div_AInv[6]), .B(u_div_AIncCry[6]), .CO(
        u_div_PartRem_7__1_), .SO(u_div_PartRem_7__0_) );
  HAD1X1 u_div_u_ha_AInc_5 ( .A(u_div_AInv[5]), .B(u_div_AIncCry[5]), .CO(
        u_div_AIncCry[6]), .SO(u_div_SumTmp_5__0_) );
  HAD1X1 u_div_u_ha_AInc_4 ( .A(u_div_AInv[4]), .B(u_div_AIncCry[4]), .CO(
        u_div_AIncCry[5]), .SO(u_div_SumTmp_4__0_) );
  HAD1X1 u_div_u_ha_AInc_3 ( .A(u_div_AInv[3]), .B(u_div_AIncCry[3]), .CO(
        u_div_AIncCry[4]), .SO(u_div_SumTmp_3__0_) );
  HAD1X1 u_div_u_ha_AInc_2 ( .A(u_div_AInv[2]), .B(u_div_AIncCry[2]), .CO(
        u_div_AIncCry[3]), .SO(u_div_SumTmp_2__0_) );
  HAD1X1 u_div_u_ha_AInc_1 ( .A(u_div_AInv[1]), .B(u_div_AIncCry[1]), .CO(
        u_div_AIncCry[2]), .SO(u_div_SumTmp_1__0_) );
  HAD1X1 u_div_u_ha_QInc_4 ( .A(u_div_QInv[4]), .B(u_div_QIncCry[4]), .CO(
        u_div_QIncCry[5]), .SO(quotient[4]) );
  HAD1X1 u_div_u_ha_QInc_3 ( .A(u_div_QInv[3]), .B(u_div_QIncCry[3]), .CO(
        u_div_QIncCry[4]), .SO(quotient[3]) );
  HAD1X1 u_div_u_ha_QInc_2 ( .A(u_div_QInv[2]), .B(u_div_QIncCry[2]), .CO(
        u_div_QIncCry[3]), .SO(quotient[2]) );
  HAD1X1 u_div_u_ha_QInc_1 ( .A(u_div_QInv[1]), .B(u_div_QIncCry[1]), .CO(
        u_div_QIncCry[2]), .SO(quotient[1]) );
  HAD1X1 u_div_u_ha_QInc_0 ( .A(u_div_QInv[0]), .B(a[7]), .CO(u_div_QIncCry[1]), .SO(quotient[0]) );
  AND2X1 u_div_u_ha_AInc_0 ( .A(u_div_AInv[0]), .B(a[8]), .Y(u_div_AIncCry[1])
         );
  XOR2X1 u_div_u_ha_QInc_5 ( .A(u_div_QInv[5]), .B(u_div_QIncCry[5]), .Y(
        quotient[5]) );
  NAND2X1 U1 ( .A(u_div_PartRem_4__2_), .B(n11), .Y(n1) );
  NAND2X1 U2 ( .A(u_div_PartRem_3__2_), .B(n12), .Y(n2) );
  NAND2X1 U3 ( .A(u_div_PartRem_5__2_), .B(n10), .Y(n3) );
  NAND2X1 U4 ( .A(u_div_PartRem_2__2_), .B(u_div_CryTmp_1__2_), .Y(n4) );
  XNOR2XL U5 ( .A(n10), .B(u_div_PartRem_5__2_), .Y(n5) );
  XNOR2XL U6 ( .A(n11), .B(u_div_PartRem_4__2_), .Y(n6) );
  XNOR2XL U7 ( .A(n12), .B(u_div_PartRem_3__2_), .Y(n7) );
  XNOR2XL U8 ( .A(u_div_PartRem_7__0_), .B(u_div_PartRem_7__1_), .Y(n8) );
  NAND21X1 U9 ( .B(u_div_PartRem_4__3_), .A(n1), .Y(u_div_CryTmp_3__4_) );
  MUX2IX1 U10 ( .D0(n17), .D1(n5), .S(u_div_CryTmp_4__4_), .Y(
        u_div_PartRem_4__3_) );
  NAND21X1 U11 ( .B(u_div_PartRem_3__3_), .A(n2), .Y(u_div_CryTmp_2__4_) );
  MUX2IX1 U12 ( .D0(n18), .D1(n6), .S(u_div_CryTmp_3__4_), .Y(
        u_div_PartRem_3__3_) );
  NAND21X1 U13 ( .B(u_div_PartRem_2__3_), .A(n4), .Y(u_div_CryTmp_1__4_) );
  MUX2IX1 U14 ( .D0(n19), .D1(n7), .S(u_div_CryTmp_2__4_), .Y(
        u_div_PartRem_2__3_) );
  INVX1 U15 ( .A(n17), .Y(u_div_PartRem_5__2_) );
  INVX1 U16 ( .A(n18), .Y(u_div_PartRem_4__2_) );
  INVX1 U17 ( .A(n19), .Y(u_div_PartRem_3__2_) );
  INVX1 U18 ( .A(n20), .Y(u_div_PartRem_2__2_) );
  MUX2AXL U19 ( .D0(n20), .D1(u_div_SumTmp_1__2_), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__3_) );
  XOR2X1 U20 ( .A(u_div_CryTmp_1__2_), .B(u_div_PartRem_2__2_), .Y(
        u_div_SumTmp_1__2_) );
  AND2X1 U21 ( .A(u_div_PartRem_7__1_), .B(u_div_PartRem_7__0_), .Y(
        u_div_CryTmp_5__4_) );
  MUX2AXL U22 ( .D0(u_div_PartRem_7__0_), .D1(u_div_PartRem_7__0_), .S(
        u_div_CryTmp_5__4_), .Y(n17) );
  MUX2AXL U23 ( .D0(n10), .D1(n10), .S(u_div_CryTmp_4__4_), .Y(n18) );
  MUX2AXL U24 ( .D0(n12), .D1(n12), .S(u_div_CryTmp_2__4_), .Y(n20) );
  MUX2AXL U25 ( .D0(n11), .D1(n11), .S(u_div_CryTmp_3__4_), .Y(n19) );
  INVX1 U26 ( .A(u_div_CryTmp_0__3_), .Y(n13) );
  NOR21XL U27 ( .B(u_div_CryTmp_0__2_), .A(n14), .Y(u_div_CryTmp_0__3_) );
  INVX1 U28 ( .A(u_div_PartRem_1__2_), .Y(n14) );
  MUX2IX1 U29 ( .D0(n22), .D1(n22), .S(u_div_CryTmp_1__4_), .Y(
        u_div_CryTmp_0__2_) );
  NAND21X1 U30 ( .B(u_div_PartRem_5__3_), .A(n3), .Y(u_div_CryTmp_4__4_) );
  MUX2IX1 U31 ( .D0(n16), .D1(n8), .S(u_div_CryTmp_5__4_), .Y(
        u_div_PartRem_5__3_) );
  MUX2AXL U32 ( .D0(n21), .D1(n21), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__2_) );
  INVX1 U33 ( .A(n21), .Y(u_div_CryTmp_1__2_) );
  XOR2X1 U34 ( .A(a[7]), .B(u_div_CryTmp_4__4_), .Y(u_div_QInv[4]) );
  XOR2X1 U35 ( .A(a[7]), .B(u_div_CryTmp_0__4_), .Y(u_div_QInv[0]) );
  NAND21X1 U36 ( .B(u_div_PartRem_1__3_), .A(n13), .Y(u_div_CryTmp_0__4_) );
  XOR2X1 U37 ( .A(a[7]), .B(u_div_CryTmp_1__4_), .Y(u_div_QInv[1]) );
  XOR2X1 U38 ( .A(a[7]), .B(u_div_CryTmp_2__4_), .Y(u_div_QInv[2]) );
  XOR2X1 U39 ( .A(a[7]), .B(u_div_CryTmp_3__4_), .Y(u_div_QInv[3]) );
  MUX2IX1 U40 ( .D0(u_div_SumTmp_2__0_), .D1(u_div_SumTmp_2__0_), .S(
        u_div_CryTmp_2__4_), .Y(n21) );
  MUX2X1 U41 ( .D0(u_div_SumTmp_5__0_), .D1(u_div_SumTmp_5__0_), .S(
        u_div_CryTmp_5__4_), .Y(n10) );
  XNOR2XL U42 ( .A(a[7]), .B(n15), .Y(u_div_QInv[5]) );
  INVX1 U43 ( .A(u_div_CryTmp_5__4_), .Y(n15) );
  MUX2X1 U44 ( .D0(u_div_SumTmp_4__0_), .D1(u_div_SumTmp_4__0_), .S(
        u_div_CryTmp_4__4_), .Y(n11) );
  MUX2X1 U45 ( .D0(u_div_SumTmp_3__0_), .D1(u_div_SumTmp_3__0_), .S(
        u_div_CryTmp_3__4_), .Y(n12) );
  INVX1 U46 ( .A(u_div_PartRem_7__1_), .Y(n16) );
  INVX1 U47 ( .A(u_div_SumTmp_1__0_), .Y(n22) );
  XOR2X1 U48 ( .A(a[8]), .B(a[6]), .Y(u_div_AInv[6]) );
  XOR2X1 U49 ( .A(a[8]), .B(a[1]), .Y(u_div_AInv[1]) );
  XOR2X1 U50 ( .A(a[8]), .B(a[0]), .Y(u_div_AInv[0]) );
  XOR2X1 U51 ( .A(a[8]), .B(a[2]), .Y(u_div_AInv[2]) );
  XOR2X1 U52 ( .A(a[8]), .B(a[3]), .Y(u_div_AInv[3]) );
  XOR2X1 U53 ( .A(a[8]), .B(a[4]), .Y(u_div_AInv[4]) );
  XOR2X1 U54 ( .A(a[8]), .B(a[5]), .Y(u_div_AInv[5]) );
endmodule


module phyrx_adp_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_db ( clk, srstz, x_cc, ptx_txact, r_rxdb_opt, gohi, golo, gotrans
 );
  input [1:0] r_rxdb_opt;
  input clk, srstz, x_cc, ptx_txact;
  output gohi, golo, gotrans;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, net148062, net148085,
         net148086, net148089, net148090, net148107, net148108, net162175,
         net167897, net168034, net168360, net168382, net168408, net168407,
         net169047, net169046, net169109, net169785, net169885, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;
  wire   [7:1] cc_buf;

  DFFQX1 cc_buf_reg_5_ ( .D(N16), .C(clk), .Q(cc_buf[5]) );
  DFFQX1 cc_buf_reg_4_ ( .D(N15), .C(clk), .Q(cc_buf[4]) );
  DFFQX1 cc_buf_reg_3_ ( .D(N14), .C(clk), .Q(cc_buf[3]) );
  DFFQXX2 cc_buf_reg_2_ ( .D(N13), .C(clk), .Q(net167897), .XQ(n26) );
  DFFQXX2 cc_buf_reg_0_ ( .D(N11), .C(clk), .Q(net168382), .XQ(n23) );
  DFFQX2 cc_buf_reg_1_ ( .D(N12), .C(clk), .Q(cc_buf[1]) );
  DFFQX2 cc_buf_reg_7_ ( .D(N18), .C(clk), .Q(cc_buf[7]) );
  DFFQX1 cc_buf_reg_6_ ( .D(N17), .C(clk), .Q(cc_buf[6]) );
  INVX2 U3 ( .A(n26), .Y(n45) );
  NOR21X2 U4 ( .B(net148086), .A(n49), .Y(n73) );
  INVX2 U5 ( .A(n40), .Y(n49) );
  INVX1 U6 ( .A(net168034), .Y(n5) );
  INVXL U7 ( .A(net168034), .Y(n17) );
  NOR21X2 U8 ( .B(n63), .A(n79), .Y(n62) );
  INVX2 U9 ( .A(net169046), .Y(net169047) );
  NAND21X2 U10 ( .B(cc_buf[7]), .A(n46), .Y(n41) );
  NAND21X2 U11 ( .B(n34), .A(n41), .Y(n35) );
  NAND2XL U12 ( .A(net168034), .B(n33), .Y(n7) );
  INVX3 U13 ( .A(cc_buf[1]), .Y(n33) );
  XNOR2X1 U14 ( .A(n32), .B(n47), .Y(net162175) );
  NAND21X1 U15 ( .B(cc_buf[1]), .A(net168407), .Y(n31) );
  NAND2X1 U16 ( .A(n7), .B(n8), .Y(n46) );
  NAND2X1 U17 ( .A(n5), .B(n6), .Y(n8) );
  INVX1 U18 ( .A(cc_buf[6]), .Y(n34) );
  NOR21XL U19 ( .B(cc_buf[7]), .A(net148090), .Y(n29) );
  INVX1 U20 ( .A(n44), .Y(n27) );
  OAI22X1 U21 ( .A(n70), .B(n69), .C(n68), .D(n67), .Y(n72) );
  INVX1 U22 ( .A(n62), .Y(n57) );
  INVX1 U23 ( .A(n88), .Y(n51) );
  INVX1 U24 ( .A(n83), .Y(n88) );
  INVX1 U25 ( .A(n42), .Y(net148062) );
  NAND21X1 U26 ( .B(net148108), .A(n37), .Y(n42) );
  NOR21XL U27 ( .B(cc_buf[6]), .A(n65), .Y(n66) );
  NAND2X1 U28 ( .A(n68), .B(n2), .Y(n3) );
  NAND2X1 U29 ( .A(n1), .B(cc_buf[3]), .Y(n4) );
  NAND2X1 U30 ( .A(n3), .B(n4), .Y(n78) );
  INVX1 U31 ( .A(n68), .Y(n1) );
  INVXL U32 ( .A(cc_buf[3]), .Y(n2) );
  INVX1 U33 ( .A(n33), .Y(n6) );
  NAND2X1 U34 ( .A(n21), .B(n10), .Y(n11) );
  NAND2X1 U35 ( .A(n9), .B(net162175), .Y(n12) );
  NAND2X1 U36 ( .A(n11), .B(n12), .Y(n79) );
  INVXL U37 ( .A(n21), .Y(n9) );
  INVXL U38 ( .A(net162175), .Y(n10) );
  NAND2X1 U39 ( .A(n32), .B(n47), .Y(n15) );
  NAND2X1 U40 ( .A(n13), .B(n14), .Y(n16) );
  NAND2X1 U41 ( .A(n15), .B(n16), .Y(net169109) );
  INVX1 U42 ( .A(n32), .Y(n13) );
  INVX1 U43 ( .A(n47), .Y(n14) );
  INVX1 U44 ( .A(cc_buf[7]), .Y(n32) );
  BUFX1 U45 ( .A(net168382), .Y(n47) );
  NAND2XL U46 ( .A(net168034), .B(cc_buf[1]), .Y(n19) );
  NAND2X1 U47 ( .A(n17), .B(n18), .Y(n20) );
  NAND2X2 U48 ( .A(n19), .B(n20), .Y(n28) );
  INVXL U49 ( .A(cc_buf[1]), .Y(n18) );
  NAND21X2 U50 ( .B(n32), .A(n28), .Y(net169785) );
  XOR2X1 U51 ( .A(net148107), .B(cc_buf[6]), .Y(n21) );
  NAND2X2 U52 ( .A(n30), .B(n31), .Y(net148107) );
  NOR2X1 U53 ( .A(n23), .B(n33), .Y(n24) );
  NAND4X1 U54 ( .A(n48), .B(n86), .C(cc_buf[3]), .D(n24), .Y(n22) );
  INVX1 U55 ( .A(r_rxdb_opt[0]), .Y(n86) );
  XNOR2XL U56 ( .A(n57), .B(n77), .Y(n56) );
  INVX2 U57 ( .A(net168382), .Y(net168408) );
  INVX1 U58 ( .A(n74), .Y(n25) );
  INVX2 U59 ( .A(n35), .Y(n38) );
  NOR21X1 U60 ( .B(net148086), .A(n49), .Y(n54) );
  NAND21X1 U61 ( .B(n39), .A(net169785), .Y(n36) );
  NAND21X1 U62 ( .B(n23), .A(net168360), .Y(n71) );
  BUFX3 U63 ( .A(net169885), .Y(net168360) );
  NAND2X1 U64 ( .A(n55), .B(n75), .Y(n77) );
  NAND43X1 U65 ( .B(net148089), .C(n24), .D(n34), .A(n41), .Y(n40) );
  NAND21X2 U66 ( .B(net148090), .A(n44), .Y(n37) );
  INVX3 U67 ( .A(n37), .Y(n39) );
  NOR32X2 U68 ( .B(net169785), .C(n37), .A(n38), .Y(net169046) );
  NAND2X2 U69 ( .A(n45), .B(cc_buf[1]), .Y(n30) );
  NAND21X1 U70 ( .B(n45), .A(n33), .Y(n43) );
  NOR21X1 U71 ( .B(n35), .A(n36), .Y(net148085) );
  BUFXL U72 ( .A(net168360), .Y(n48) );
  INVXL U73 ( .A(n24), .Y(n50) );
  NAND31X1 U74 ( .C(n27), .A(n28), .B(n29), .Y(net148086) );
  INVX3 U75 ( .A(n30), .Y(net148090) );
  NAND21X2 U76 ( .B(n23), .A(n43), .Y(n44) );
  NAND21X1 U77 ( .B(n87), .A(n60), .Y(n80) );
  MUX2IX4 U78 ( .D0(n82), .D1(n81), .S(r_rxdb_opt[1]), .Y(golo) );
  INVXL U79 ( .A(net168407), .Y(net169885) );
  NAND3X2 U80 ( .A(n51), .B(n52), .C(r_rxdb_opt[0]), .Y(n53) );
  NAND2X2 U81 ( .A(n53), .B(n85), .Y(gohi) );
  INVX1 U82 ( .A(n56), .Y(n52) );
  XOR2XL U83 ( .A(n23), .B(cc_buf[1]), .Y(n64) );
  INVX3 U84 ( .A(net167897), .Y(net168407) );
  OAI21BBXL U85 ( .A(net169047), .B(n54), .C(n72), .Y(n76) );
  INVX1 U86 ( .A(n61), .Y(n60) );
  AOI21AX1 U87 ( .B(net148062), .C(n25), .A(n22), .Y(n85) );
  OAI21BBX1 U88 ( .A(net169047), .B(n73), .C(n72), .Y(n55) );
  XNOR2X1 U89 ( .A(n77), .B(n57), .Y(n87) );
  NAND2X1 U90 ( .A(net167897), .B(net168382), .Y(n58) );
  NAND2X2 U91 ( .A(net168407), .B(net168408), .Y(n59) );
  NAND2X2 U92 ( .A(n59), .B(n58), .Y(net168034) );
  NAND21X2 U93 ( .B(n83), .A(n80), .Y(n81) );
  OAI21BBX1 U94 ( .A(n62), .B(n75), .C(n76), .Y(n84) );
  INVX1 U95 ( .A(n78), .Y(n63) );
  INVXL U96 ( .A(cc_buf[3]), .Y(n67) );
  AND2X1 U97 ( .A(x_cc), .B(srstz), .Y(N11) );
  XNOR2XL U98 ( .A(n78), .B(n79), .Y(n61) );
  NAND42XL U99 ( .C(cc_buf[3]), .D(n48), .A(n64), .B(n50), .Y(n82) );
  NAND21X1 U100 ( .B(net148090), .A(n71), .Y(net148089) );
  NOR21XL U101 ( .B(net169785), .A(n66), .Y(net148108) );
  XOR2XL U102 ( .A(net169109), .B(net148107), .Y(n65) );
  INVXL U103 ( .A(cc_buf[5]), .Y(n69) );
  XOR2X1 U104 ( .A(n70), .B(cc_buf[5]), .Y(n68) );
  INVX2 U105 ( .A(cc_buf[4]), .Y(n70) );
  INVXL U106 ( .A(n64), .Y(gotrans) );
  AND2XL U107 ( .A(srstz), .B(n48), .Y(N14) );
  AND2XL U108 ( .A(srstz), .B(cc_buf[5]), .Y(N17) );
  AND2XL U109 ( .A(srstz), .B(n47), .Y(N12) );
  AND2XL U110 ( .A(srstz), .B(cc_buf[6]), .Y(N18) );
  AND2XL U111 ( .A(srstz), .B(cc_buf[3]), .Y(N15) );
  AND2XL U112 ( .A(srstz), .B(cc_buf[4]), .Y(N16) );
  NAND21X2 U113 ( .B(net148062), .A(n74), .Y(n83) );
  NAND32X1 U114 ( .B(net148085), .C(n72), .A(n54), .Y(n75) );
  INVX2 U115 ( .A(n84), .Y(n74) );
  NOR32XL U116 ( .B(srstz), .C(cc_buf[1]), .A(ptx_txact), .Y(N13) );
endmodule


module i2cslv_a0 ( i_sda, i_scl, o_sda, i_deva, i_inc, i_fwnak, i_fwack, o_we, 
        o_re, o_r_early, o_idle, o_dec, o_busev, o_ofs, o_lt_ofs, o_wdat, 
        o_lt_buf, o_dbgpo, i_rdat, i_rd_mem, i_clk, i_rstz, i_prefetch );
  input [7:1] i_deva;
  output [3:0] o_busev;
  output [7:0] o_ofs;
  output [7:0] o_lt_ofs;
  output [7:0] o_wdat;
  output [7:0] o_lt_buf;
  output [7:0] o_dbgpo;
  input [7:0] i_rdat;
  input i_sda, i_scl, i_inc, i_fwnak, i_fwack, i_rd_mem, i_clk, i_rstz,
         i_prefetch;
  output o_sda, o_we, o_re, o_r_early, o_idle, o_dec;
  wire   i2c_scl, sdafall, cs_rwb, N74, N75, N76, N77, N78, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, ps_rwbuf_0_, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, net10777, net10783, net10788, net10793,
         net10798, n61, n73, n97, n98, n118, n119, n120, n121, n1, n2, n3, n4,
         n5, n6, n7, n9, n10, n11, n12, n13, n14, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165;
  wire   [1:0] cs_sta;

  i2cdbnc_a0_1 db_scl ( .i_clk(i_clk), .i_rstz(n16), .i_i2c(i_scl), .r_opt({
        1'b1, 1'b0}), .o_i2c(i2c_scl), .rise(o_dbgpo[6]), .fall(o_dbgpo[7]) );
  i2cdbnc_a0_0 db_sda ( .i_clk(i_clk), .i_rstz(n16), .i_i2c(i_sda), .r_opt({
        1'b0, 1'b0}), .o_i2c(ps_rwbuf_0_), .rise(o_dbgpo[5]), .fall(sdafall)
         );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 clk_gate_cs_bit_reg ( .CLK(i_clk), .EN(N74), 
        .ENCLK(net10777), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 clk_gate_adcnt_reg ( .CLK(i_clk), .EN(N114), 
        .ENCLK(net10783), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 clk_gate_rwbuf_reg ( .CLK(i_clk), .EN(N144), 
        .ENCLK(net10788), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 clk_gate_lt_buf_reg ( .CLK(i_clk), .EN(N179), .ENCLK(net10793), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 clk_gate_lt_ofs_reg ( .CLK(i_clk), .EN(
        o_busev[2]), .ENCLK(net10798), .TE(1'b0) );
  DFFQX1 lt_ofs_reg_7_ ( .D(o_wdat[7]), .C(net10798), .Q(o_lt_ofs[7]) );
  DFFQX1 lt_ofs_reg_6_ ( .D(o_wdat[6]), .C(net10798), .Q(o_lt_ofs[6]) );
  DFFQX1 lt_buf_reg_7_ ( .D(N187), .C(net10793), .Q(o_lt_buf[7]) );
  DFFQX1 lt_buf_reg_6_ ( .D(N186), .C(net10793), .Q(o_lt_buf[6]) );
  DFFQX1 lt_ofs_reg_5_ ( .D(o_wdat[5]), .C(net10798), .Q(o_lt_ofs[5]) );
  DFFQX1 lt_ofs_reg_4_ ( .D(o_wdat[4]), .C(net10798), .Q(o_lt_ofs[4]) );
  DFFQX1 lt_buf_reg_5_ ( .D(N185), .C(net10793), .Q(o_lt_buf[5]) );
  DFFQX1 lt_buf_reg_4_ ( .D(N184), .C(net10793), .Q(o_lt_buf[4]) );
  DFFQX1 lt_ofs_reg_3_ ( .D(o_wdat[3]), .C(net10798), .Q(o_lt_ofs[3]) );
  DFFQX1 lt_buf_reg_3_ ( .D(N183), .C(net10793), .Q(o_lt_buf[3]) );
  DFFSQX1 sdat_reg ( .D(n118), .C(i_clk), .XS(n17), .Q(o_sda) );
  DFFQX1 lt_ofs_reg_2_ ( .D(o_wdat[2]), .C(net10798), .Q(o_lt_ofs[2]) );
  DFFQX1 lt_ofs_reg_1_ ( .D(o_wdat[1]), .C(net10798), .Q(o_lt_ofs[1]) );
  DFFQX1 lt_buf_reg_2_ ( .D(N182), .C(net10793), .Q(o_lt_buf[2]) );
  DFFQX1 lt_buf_reg_1_ ( .D(N181), .C(net10793), .Q(o_lt_buf[1]) );
  DFFQX1 lt_ofs_reg_0_ ( .D(o_wdat[0]), .C(net10798), .Q(o_lt_ofs[0]) );
  DFFQX1 lt_buf_reg_0_ ( .D(N180), .C(net10793), .Q(o_lt_buf[0]) );
  DFFRQX1 adcnt_reg_6_ ( .D(N112), .C(net10783), .XR(n19), .Q(o_ofs[6]) );
  DFFRQX1 adcnt_reg_3_ ( .D(N109), .C(net10783), .XR(n18), .Q(o_ofs[3]) );
  DFFRQX1 adcnt_reg_5_ ( .D(N111), .C(net10783), .XR(n18), .Q(o_ofs[5]) );
  DFFRQX1 adcnt_reg_0_ ( .D(N106), .C(net10783), .XR(n18), .Q(o_ofs[0]) );
  DFFRQX1 adcnt_reg_2_ ( .D(N108), .C(net10783), .XR(n18), .Q(o_ofs[2]) );
  DFFRQX1 adcnt_reg_1_ ( .D(N107), .C(net10783), .XR(n18), .Q(o_ofs[1]) );
  DFFSQX1 rwbuf_reg_5_ ( .D(N141), .C(net10788), .XS(n17), .Q(o_wdat[5]) );
  DFFSQX1 rwbuf_reg_7_ ( .D(N143), .C(net10788), .XS(n16), .Q(o_wdat[7]) );
  DFFRQX1 cs_rwb_reg ( .D(n119), .C(i_clk), .XR(n18), .Q(cs_rwb) );
  DFFSQX1 cs_bit_reg_2_ ( .D(N77), .C(net10777), .XS(n17), .Q(o_dbgpo[2]) );
  DFFSQX1 cs_bit_reg_3_ ( .D(N78), .C(net10777), .XS(n17), .Q(o_dbgpo[3]) );
  DFFSQX1 rwbuf_reg_0_ ( .D(N136), .C(net10788), .XS(n16), .Q(o_wdat[0]) );
  DFFSQX1 rwbuf_reg_2_ ( .D(N138), .C(net10788), .XS(n17), .Q(o_wdat[2]) );
  DFFSQX1 rwbuf_reg_6_ ( .D(N142), .C(net10788), .XS(n17), .Q(o_wdat[6]) );
  DFFSQX1 rwbuf_reg_4_ ( .D(N140), .C(net10788), .XS(n17), .Q(o_wdat[4]) );
  DFFRQX1 adcnt_reg_7_ ( .D(N113), .C(net10783), .XR(n18), .Q(o_ofs[7]) );
  DFFSQX1 cs_bit_reg_0_ ( .D(N75), .C(net10777), .XS(n17), .Q(o_dbgpo[0]) );
  DFFSQX1 cs_bit_reg_1_ ( .D(N76), .C(net10777), .XS(n17), .Q(o_dbgpo[1]) );
  DFFSQX1 rwbuf_reg_1_ ( .D(N137), .C(net10788), .XS(n18), .Q(o_wdat[1]) );
  DFFSQX1 rwbuf_reg_3_ ( .D(N139), .C(net10788), .XS(n17), .Q(o_wdat[3]) );
  DFFRQX1 cs_sta_reg_0_ ( .D(n120), .C(i_clk), .XR(n18), .Q(cs_sta[0]) );
  DFFRQX1 cs_sta_reg_1_ ( .D(n121), .C(i_clk), .XR(n19), .Q(cs_sta[1]) );
  DFFRQX1 adcnt_reg_4_ ( .D(N110), .C(net10783), .XR(n18), .Q(o_ofs[4]) );
  INVX1 U3 ( .A(o_dbgpo[7]), .Y(n71) );
  INVX1 U4 ( .A(n27), .Y(o_busev[1]) );
  INVX1 U5 ( .A(cs_sta[0]), .Y(n155) );
  GEN2XL U6 ( .D(o_dbgpo[7]), .E(n161), .C(n65), .B(n131), .A(n56), .Y(n57) );
  INVX1 U7 ( .A(n85), .Y(o_we) );
  INVX1 U8 ( .A(o_wdat[3]), .Y(n100) );
  INVX1 U9 ( .A(o_wdat[4]), .Y(n82) );
  INVX1 U10 ( .A(o_wdat[5]), .Y(n110) );
  NAND21X1 U11 ( .B(n69), .A(o_busev[1]), .Y(n84) );
  INVX1 U12 ( .A(o_wdat[6]), .Y(n83) );
  INVX1 U13 ( .A(n133), .Y(n152) );
  XOR2X1 U14 ( .A(i_deva[1]), .B(o_wdat[0]), .Y(n51) );
  NAND21X1 U15 ( .B(n26), .A(o_dbgpo[0]), .Y(n147) );
  XOR2X1 U16 ( .A(n110), .B(i_deva[5]), .Y(n37) );
  XOR2X1 U17 ( .A(i_deva[2]), .B(o_wdat[1]), .Y(n52) );
  AO21XL U18 ( .B(n138), .C(n93), .A(n152), .Y(n87) );
  NAND21XL U19 ( .B(n79), .A(n85), .Y(N179) );
  NAND42XL U20 ( .C(n146), .D(n133), .A(n132), .B(o_dbgpo[6]), .Y(n135) );
  OA22XL U21 ( .A(n158), .B(n157), .C(n156), .D(n155), .Y(n159) );
  MUX2AXL U22 ( .D0(n1), .D1(n163), .S(o_dbgpo[7]), .Y(n118) );
  AOI22X1 U23 ( .A(n165), .B(i_fwnak), .C(n61), .D(n140), .Y(n1) );
  NAND32XL U24 ( .B(n71), .C(n126), .A(n156), .Y(n68) );
  AOI21XL U25 ( .B(o_dbgpo[7]), .C(n152), .A(n57), .Y(n9) );
  NAND32XL U26 ( .B(n56), .C(n75), .A(n69), .Y(n53) );
  AOI31XL U27 ( .A(n152), .B(n151), .C(n150), .D(n149), .Y(n160) );
  OA21XL U28 ( .B(n147), .C(n146), .A(n145), .Y(n150) );
  NAND32XL U29 ( .B(o_idle), .C(n71), .A(n148), .Y(n97) );
  AO21XL U30 ( .B(n138), .C(n116), .A(n152), .Y(n123) );
  AO21XL U31 ( .B(n138), .C(n106), .A(n152), .Y(n108) );
  AO21XL U32 ( .B(n138), .C(n94), .A(n152), .Y(n96) );
  NAND21X1 U33 ( .B(n142), .A(cs_rwb), .Y(n151) );
  MUX2IX1 U34 ( .D0(n135), .D1(n134), .S(i_prefetch), .Y(o_r_early) );
  OAI32X1 U35 ( .A(i_prefetch), .B(ps_rwbuf_0_), .C(n151), .D(n136), .E(n145), 
        .Y(n137) );
  NAND32X1 U36 ( .B(o_dbgpo[3]), .C(o_dbgpo[2]), .A(n21), .Y(n26) );
  INVX1 U37 ( .A(o_dbgpo[1]), .Y(n21) );
  NAND21XL U38 ( .B(cs_sta[0]), .A(cs_sta[1]), .Y(n127) );
  INVXL U39 ( .A(cs_rwb), .Y(n136) );
  XOR2XL U40 ( .A(i_deva[6]), .B(o_wdat[6]), .Y(n34) );
  INVXL U41 ( .A(ps_rwbuf_0_), .Y(n141) );
  NAND32XL U42 ( .B(n29), .C(o_dbgpo[7]), .A(sdafall), .Y(n73) );
  NAND21XL U43 ( .B(cs_sta[1]), .A(cs_sta[0]), .Y(n126) );
  MUX2BXL U44 ( .D0(n131), .D1(n2), .S(cs_rwb), .Y(n78) );
  AOI21XL U45 ( .B(n156), .C(n77), .A(n76), .Y(n2) );
  MUX2AXL U46 ( .D0(n3), .D1(cs_sta[1]), .S(n9), .Y(n121) );
  AOI21X1 U47 ( .B(n64), .C(n54), .A(n63), .Y(n3) );
  MUX2XL U48 ( .D0(n67), .D1(cs_sta[0]), .S(n9), .Y(n120) );
  AND2XL U49 ( .A(n131), .B(n155), .Y(n66) );
  NAND21XL U50 ( .B(n155), .A(cs_sta[1]), .Y(n148) );
  NAND21XL U51 ( .B(n156), .A(cs_rwb), .Y(n157) );
  NAND2XL U52 ( .A(cs_rwb), .B(n73), .Y(n13) );
  OAI21BBXL U53 ( .A(o_wdat[6]), .B(n122), .C(n4), .Y(N112) );
  MUX2IX1 U54 ( .D0(n117), .D1(n123), .S(o_ofs[6]), .Y(n4) );
  OAI21BBXL U55 ( .A(o_wdat[4]), .B(n122), .C(n5), .Y(N110) );
  MUX2IX1 U56 ( .D0(n107), .D1(n108), .S(o_ofs[4]), .Y(n5) );
  OAI21BBXL U57 ( .A(o_wdat[2]), .B(n122), .C(n6), .Y(N108) );
  MUX2IX1 U58 ( .D0(n95), .D1(n96), .S(o_ofs[2]), .Y(n6) );
  OAI21BBXL U59 ( .A(o_wdat[0]), .B(n122), .C(n7), .Y(N106) );
  MUX2IX1 U60 ( .D0(n86), .D1(n87), .S(o_ofs[0]), .Y(n7) );
  INVXL U61 ( .A(cs_sta[1]), .Y(n161) );
  INVX1 U62 ( .A(n61), .Y(n165) );
  INVX1 U63 ( .A(n20), .Y(n17) );
  INVX1 U64 ( .A(n20), .Y(n18) );
  INVX1 U65 ( .A(n20), .Y(n19) );
  XNOR2XL U66 ( .A(i_fwnak), .B(i_fwack), .Y(n61) );
  INVX1 U67 ( .A(n20), .Y(n16) );
  INVX1 U68 ( .A(i_rstz), .Y(n20) );
  INVX1 U69 ( .A(n84), .Y(n79) );
  INVX1 U70 ( .A(n32), .Y(n74) );
  INVX1 U71 ( .A(n56), .Y(n64) );
  INVX1 U72 ( .A(n55), .Y(n65) );
  NAND21X1 U73 ( .B(o_busev[0]), .A(n98), .Y(n23) );
  INVX1 U74 ( .A(n98), .Y(n62) );
  INVX1 U75 ( .A(n58), .Y(n22) );
  AND2X1 U76 ( .A(n152), .B(n131), .Y(o_dec) );
  NAND32X1 U77 ( .B(n127), .C(n71), .A(n144), .Y(n85) );
  NAND21X1 U78 ( .B(n141), .A(n79), .Y(n134) );
  NAND21X1 U79 ( .B(n147), .A(i_prefetch), .Y(n145) );
  NAND32X1 U80 ( .B(n147), .C(n31), .A(n152), .Y(n27) );
  INVX1 U81 ( .A(o_dbgpo[6]), .Y(n31) );
  INVX1 U82 ( .A(n127), .Y(n138) );
  INVX1 U83 ( .A(n147), .Y(n156) );
  INVX1 U84 ( .A(n26), .Y(n28) );
  INVX1 U85 ( .A(n151), .Y(n132) );
  NOR3XL U86 ( .A(n44), .B(n42), .C(n60), .Y(o_idle) );
  OAI211X1 U87 ( .C(n162), .D(n161), .A(n160), .B(n159), .Y(n163) );
  OA22X1 U88 ( .A(n144), .B(n143), .C(n142), .D(n141), .Y(n162) );
  INVX1 U89 ( .A(i_rd_mem), .Y(n164) );
  NAND32XL U90 ( .B(n31), .C(n72), .A(n142), .Y(n32) );
  OA22X1 U91 ( .A(i_rd_mem), .B(n154), .C(n153), .D(n164), .Y(n158) );
  INVX1 U92 ( .A(i_rdat[7]), .Y(n153) );
  OA21X1 U93 ( .B(n74), .C(n72), .A(n148), .Y(N144) );
  OAI22AX1 U94 ( .D(n72), .C(n153), .A(n83), .B(n32), .Y(N143) );
  INVX1 U95 ( .A(n73), .Y(o_busev[0]) );
  INVX1 U96 ( .A(n68), .Y(o_busev[2]) );
  NAND21X1 U97 ( .B(o_busev[3]), .A(n73), .Y(n56) );
  NAND5XL U98 ( .A(o_dbgpo[6]), .B(n152), .C(n71), .D(n146), .E(n77), .Y(n55)
         );
  INVX1 U99 ( .A(i_prefetch), .Y(n77) );
  INVX1 U100 ( .A(n106), .Y(n113) );
  INVX1 U101 ( .A(n94), .Y(n103) );
  INVX1 U102 ( .A(n53), .Y(n63) );
  INVX1 U103 ( .A(n148), .Y(n149) );
  INVX1 U104 ( .A(i_inc), .Y(n93) );
  NAND21X1 U105 ( .B(o_busev[0]), .A(o_busev[3]), .Y(n98) );
  NAND21X1 U106 ( .B(n97), .A(n142), .Y(n58) );
  OR2X1 U107 ( .A(n62), .B(n10), .Y(N76) );
  AOI21X1 U108 ( .B(n60), .C(n59), .A(n58), .Y(n10) );
  AO21X1 U109 ( .B(n22), .C(n43), .A(n23), .Y(N75) );
  INVX1 U110 ( .A(n142), .Y(n131) );
  INVX1 U111 ( .A(n116), .Y(n124) );
  OAI22XL U112 ( .A(n81), .B(n85), .C(n84), .D(n89), .Y(N182) );
  OAI22XL U113 ( .A(n100), .B(n85), .C(n84), .D(n81), .Y(N183) );
  OAI22XL U114 ( .A(n82), .B(n85), .C(n84), .D(n100), .Y(N184) );
  OAI22XL U115 ( .A(n110), .B(n85), .C(n84), .D(n82), .Y(N185) );
  OAI22XL U116 ( .A(n83), .B(n85), .C(n84), .D(n110), .Y(N186) );
  OAI22XL U117 ( .A(n154), .B(n85), .C(n84), .D(n83), .Y(N187) );
  INVX1 U118 ( .A(n157), .Y(n143) );
  INVX1 U119 ( .A(n25), .Y(n30) );
  NAND3X1 U120 ( .A(n97), .B(n73), .C(n98), .Y(N74) );
  INVX1 U121 ( .A(n126), .Y(n122) );
  BUFX3 U122 ( .A(o_busev[3]), .Y(o_dbgpo[4]) );
  NAND21X1 U123 ( .B(o_dbgpo[0]), .A(n28), .Y(n142) );
  NAND21X1 U124 ( .B(cs_sta[1]), .A(n155), .Y(n133) );
  NAND43X1 U125 ( .B(n52), .C(n51), .D(n50), .A(n49), .Y(n69) );
  AND4X1 U126 ( .A(n48), .B(n47), .C(n46), .D(n45), .Y(n49) );
  NAND43X1 U127 ( .B(n41), .C(n40), .D(n39), .A(n38), .Y(n146) );
  NOR32XL U128 ( .B(n37), .C(n36), .A(n35), .Y(n38) );
  XOR2XL U129 ( .A(i_deva[2]), .B(o_wdat[2]), .Y(n41) );
  XOR2XL U130 ( .A(i_deva[1]), .B(o_wdat[1]), .Y(n40) );
  NAND21X1 U131 ( .B(n34), .A(n33), .Y(n35) );
  XNOR2XL U132 ( .A(i_deva[4]), .B(o_wdat[4]), .Y(n33) );
  XNOR2XL U133 ( .A(i_deva[7]), .B(o_wdat[7]), .Y(n36) );
  XOR2X1 U134 ( .A(n83), .B(i_deva[7]), .Y(n45) );
  XOR2X1 U135 ( .A(n82), .B(i_deva[5]), .Y(n46) );
  XOR2X1 U136 ( .A(n110), .B(i_deva[6]), .Y(n48) );
  XOR2X1 U137 ( .A(n100), .B(i_deva[4]), .Y(n47) );
  XOR2XL U138 ( .A(i_deva[3]), .B(o_wdat[2]), .Y(n50) );
  XOR2XL U139 ( .A(i_deva[3]), .B(o_wdat[3]), .Y(n39) );
  AND3XL U140 ( .A(o_dbgpo[6]), .B(n138), .C(n137), .Y(o_re) );
  INVX1 U141 ( .A(n70), .Y(n144) );
  NAND21X1 U142 ( .B(cs_rwb), .A(n156), .Y(n70) );
  NAND21XL U143 ( .B(n43), .A(o_dbgpo[1]), .Y(n60) );
  INVXL U144 ( .A(o_dbgpo[0]), .Y(n43) );
  INVXL U145 ( .A(o_dbgpo[3]), .Y(n44) );
  INVXL U146 ( .A(o_dbgpo[2]), .Y(n42) );
  NAND6XL U147 ( .A(cs_rwb), .B(o_dbgpo[3]), .C(n30), .D(n148), .E(n29), .F(
        i_rd_mem), .Y(n139) );
  MUX2X1 U148 ( .D0(i_rdat[7]), .D1(o_sda), .S(n139), .Y(n140) );
  NAND2X1 U149 ( .A(n11), .B(n139), .Y(n72) );
  NAND4XL U150 ( .A(n28), .B(cs_rwb), .C(n148), .D(i_rd_mem), .Y(n11) );
  AO22XL U151 ( .A(n74), .B(o_wdat[5]), .C(i_rdat[6]), .D(n72), .Y(N142) );
  AO22XL U152 ( .A(n74), .B(o_wdat[4]), .C(i_rdat[5]), .D(n72), .Y(N141) );
  AO22XL U153 ( .A(n74), .B(o_wdat[3]), .C(i_rdat[4]), .D(n72), .Y(N140) );
  AO22XL U154 ( .A(n74), .B(o_wdat[2]), .C(i_rdat[3]), .D(n72), .Y(N139) );
  AO22XL U155 ( .A(n74), .B(o_wdat[1]), .C(i_rdat[2]), .D(n72), .Y(N138) );
  AO22XL U156 ( .A(n74), .B(o_wdat[0]), .C(i_rdat[1]), .D(n72), .Y(N137) );
  OAI21BBX1 U157 ( .A(i_rdat[0]), .B(n72), .C(n12), .Y(N136) );
  NAND4XL U158 ( .A(o_dbgpo[6]), .B(ps_rwbuf_0_), .C(n142), .D(n136), .Y(n12)
         );
  NOR32XL U159 ( .B(i2c_scl), .C(o_dbgpo[5]), .A(o_dbgpo[7]), .Y(o_busev[3])
         );
  NAND31X1 U160 ( .C(n93), .A(o_ofs[0]), .B(o_ofs[1]), .Y(n94) );
  NAND32X1 U161 ( .B(n115), .C(n114), .A(n113), .Y(n116) );
  INVX1 U162 ( .A(o_ofs[4]), .Y(n115) );
  NAND32X1 U163 ( .B(n105), .C(n104), .A(n103), .Y(n106) );
  INVX1 U164 ( .A(o_ofs[2]), .Y(n105) );
  NAND5XL U165 ( .A(o_dbgpo[1]), .B(i_prefetch), .C(n44), .D(n43), .E(n42), 
        .Y(n75) );
  GEN2XL U166 ( .D(n138), .E(n78), .C(n152), .B(o_dbgpo[7]), .A(o_busev[2]), 
        .Y(N114) );
  INVX1 U167 ( .A(n75), .Y(n76) );
  GEN2XL U168 ( .D(n66), .E(n136), .C(n65), .B(n64), .A(n63), .Y(n67) );
  NAND32XL U169 ( .B(cs_sta[0]), .C(n132), .A(n55), .Y(n54) );
  AND2X1 U170 ( .A(n124), .B(n138), .Y(n117) );
  INVX1 U171 ( .A(i2c_scl), .Y(n29) );
  NAND21XL U172 ( .B(o_dbgpo[1]), .A(n43), .Y(n59) );
  OR2XL U173 ( .A(o_dbgpo[2]), .B(n59), .Y(n25) );
  GEN2XL U174 ( .D(o_dbgpo[3]), .E(n25), .C(n131), .B(n24), .A(n23), .Y(N78)
         );
  INVX1 U175 ( .A(n97), .Y(n24) );
  GEN2XL U176 ( .D(o_dbgpo[2]), .E(n59), .C(n30), .B(n22), .A(n62), .Y(N77) );
  MUX2BXL U177 ( .D0(ps_rwbuf_0_), .D1(n13), .S(n14), .Y(n119) );
  NAND2XL U178 ( .A(o_busev[1]), .B(n73), .Y(n14) );
  AND2X1 U179 ( .A(n113), .B(n138), .Y(n107) );
  AND2X1 U180 ( .A(n103), .B(n138), .Y(n95) );
  AND2X1 U181 ( .A(i_inc), .B(n138), .Y(n86) );
  OAI21BBXL U182 ( .A(o_we), .B(o_wdat[0]), .C(n134), .Y(N180) );
  NAND21XL U183 ( .B(o_ofs[7]), .A(n124), .Y(n125) );
  OAI222XL U184 ( .A(n130), .B(n129), .C(n128), .D(n127), .E(n154), .F(n126), 
        .Y(N113) );
  MUX2X1 U185 ( .D0(n129), .D1(n125), .S(o_ofs[6]), .Y(n128) );
  INVX1 U186 ( .A(n123), .Y(n130) );
  INVXL U187 ( .A(o_ofs[7]), .Y(n129) );
  OAI222XL U188 ( .A(n112), .B(n114), .C(n111), .D(n127), .E(n126), .F(n110), 
        .Y(N111) );
  MUX2X1 U189 ( .D0(n114), .D1(n109), .S(o_ofs[4]), .Y(n111) );
  INVX1 U190 ( .A(n108), .Y(n112) );
  NAND21X1 U191 ( .B(o_ofs[5]), .A(n113), .Y(n109) );
  OAI222XL U192 ( .A(n102), .B(n104), .C(n101), .D(n127), .E(n126), .F(n100), 
        .Y(N109) );
  MUX2X1 U193 ( .D0(n104), .D1(n99), .S(o_ofs[2]), .Y(n101) );
  INVX1 U194 ( .A(n96), .Y(n102) );
  NAND21X1 U195 ( .B(o_ofs[3]), .A(n103), .Y(n99) );
  OAI22XL U196 ( .A(n89), .B(n85), .C(n84), .D(n80), .Y(N181) );
  INVXL U197 ( .A(o_wdat[0]), .Y(n80) );
  INVX1 U198 ( .A(o_ofs[5]), .Y(n114) );
  INVX1 U199 ( .A(o_ofs[3]), .Y(n104) );
  NAND21X1 U200 ( .B(o_ofs[1]), .A(i_inc), .Y(n88) );
  OAI222XL U201 ( .A(n92), .B(n91), .C(n90), .D(n127), .E(n126), .F(n89), .Y(
        N107) );
  MUX2X1 U202 ( .D0(n91), .D1(n88), .S(o_ofs[0]), .Y(n90) );
  INVX1 U203 ( .A(n87), .Y(n92) );
  INVX1 U204 ( .A(o_ofs[1]), .Y(n91) );
  INVXL U205 ( .A(o_wdat[7]), .Y(n154) );
  INVXL U206 ( .A(o_wdat[1]), .Y(n89) );
  INVXL U207 ( .A(o_wdat[2]), .Y(n81) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2cdbnc_a0_0 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n2, n3, n5, n8, n9, n10, n11;

  DFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .C(i_clk), .XS(i_rstz), .Q(N18) );
  DFFSQX1 d_i2c_reg_1_ ( .D(N18), .C(i_clk), .XS(i_rstz), .Q(N19) );
  DFFSQX1 d_i2c_reg_2_ ( .D(N19), .C(i_clk), .XS(i_rstz), .Q(d_i2c_2_) );
  DFFSQXX1 r_i2c_reg ( .D(n9), .C(i_clk), .XS(i_rstz), .Q(o_i2c), .XQ(n11) );
  AND3X1 U3 ( .A(n8), .B(o_i2c), .C(n2), .Y(fall) );
  INVX1 U4 ( .A(n5), .Y(rise) );
  OAI211X1 U5 ( .C(r_opt[0]), .D(d_i2c_2_), .A(n11), .B(n10), .Y(n5) );
  AND2X1 U6 ( .A(N18), .B(N19), .Y(n10) );
  NAND21X1 U7 ( .B(r_opt[1]), .A(d_i2c_2_), .Y(n8) );
  NOR2X1 U8 ( .A(N19), .B(N18), .Y(n2) );
  OR2X1 U9 ( .A(rise), .B(n3), .Y(n9) );
  AOI21X1 U10 ( .B(n8), .C(n2), .A(n11), .Y(n3) );
endmodule


module i2cdbnc_a0_1 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n1, n6, n2, n3, n4, n5;

  DFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .C(i_clk), .XS(i_rstz), .Q(N18) );
  DFFSQX1 d_i2c_reg_1_ ( .D(N18), .C(i_clk), .XS(i_rstz), .Q(N19) );
  DFFSQX1 d_i2c_reg_2_ ( .D(N19), .C(i_clk), .XS(i_rstz), .Q(d_i2c_2_) );
  DFFSQXXL r_i2c_reg ( .D(n6), .C(i_clk), .XS(i_rstz), .Q(o_i2c), .XQ(n1) );
  AND4X1 U3 ( .A(n1), .B(N19), .C(N18), .D(n2), .Y(rise) );
  OR2X1 U4 ( .A(d_i2c_2_), .B(r_opt[0]), .Y(n2) );
  AO21XL U5 ( .B(n5), .C(o_i2c), .A(rise), .Y(n6) );
  INVX1 U6 ( .A(n5), .Y(fall) );
  NAND32XL U7 ( .B(N19), .C(N18), .A(n4), .Y(n5) );
  OA21X1 U8 ( .B(r_opt[1]), .C(n3), .A(o_i2c), .Y(n4) );
  INVXL U9 ( .A(d_i2c_2_), .Y(n3) );
endmodule


module regbank_a0 ( srci, lg_pulse_len, dm_fault, cc1_di, cc2_di, di_rd_det, 
        i_tmrf, i_vcbyval, dnchk_en, r_pwrv_upd, aswkup, lg_dischg, gating_pwr, 
        ps_pwrdn, r_sleep, r_pwrdn, r_ocdrv_enz, r_osc_stop, r_osc_lo, 
        r_osc_gate, r_fw_pwrv, r_cvcwr, r_cvofs, r_otpi_gate, r_pwrctl, 
        r_pwr_i, r_cvctl, r_srcctl, r_dpdmctl, r_ccrx, r_cctrx, r_ccctl, 
        r_fcpwr, r_fcpre, fcp_r_dat, fcp_r_sta, fcp_r_msk, fcp_r_ctl, 
        fcp_r_crc, fcp_r_acc, fcp_r_tui, r_accctl, r_bclk_sel, r_dacwr, 
        r_dac_en, r_sar_en, r_adofs, r_isofs, x_daclsb, r_comp_opt, dac_r_ctl, 
        dac_r_comp, dac_r_cmpsta, dac_r_vs, REVID, atpg_en, sfr_r, sfr_w, 
        set_hold, bkpt_hold, cpurst, sfr_addr, sfr_wdat, sfr_rdat, ff_p0, 
        di_p0, ictlr_idle, ictlr_inc, r_inst_ofs, r_psrd, r_pswr, r_fortxdat, 
        r_fortxrdy, r_fortxen, r_ana_tm, r_gpio_tm, r_gpio_ie, r_gpio_oe, 
        r_gpio_pu, r_gpio_pd, r_gpio_s0, r_gpio_s1, r_gpio_s2, r_gpio_s3, 
        r_regtrm, i_pc, i_goidle, i_gobusy, i_i2c_idle, bus_idle, i2c_stretch, 
        i_i2c_rwbuf, i_i2c_ltbuf, i_i2c_ofs, o_intr, r_auto_gdcrc, r_exist1st, 
        r_ordrs4, r_fifopsh, r_fifopop, r_unlock, r_first, r_last, r_fiforst, 
        r_set_cpmsgid, r_txendk, r_txnumk, r_txshrt, r_auto_discard, 
        r_hold_mcu, r_txauto, r_rxords_ena, r_spec, r_dat_spec, r_dat_portrole, 
        r_dat_datarole, r_discard, r_pshords, r_pg0_sel, r_strtch, r_i2c_attr, 
        r_i2c_ninc, r_hwi2c_en, r_i2c_fwnak, r_i2c_fwack, r_i2c_deva, i2c_ev, 
        prl_c0set, prl_cany0, prl_discard, prl_GCTxDone, prl_cpmsgid, pff_ack, 
        prx_rst, pff_obsd, pff_full, pff_empty, ptx_ack, pff_ptr, prx_adpn, 
        pff_rdat, pff_rxpart, prx_rcvinf, ptx_fsm, prx_fsm, prl_fsm, 
        prx_setsta, clk_1p0m, clk_500, clk, xrstz, xclk, dbgpo, srstz, prstz
 );
  input [5:0] srci;
  input [1:0] lg_pulse_len;
  output [11:0] r_fw_pwrv;
  output [1:0] r_cvcwr;
  input [15:0] r_cvofs;
  output [7:4] r_pwrctl;
  output [7:0] r_pwr_i;
  output [7:0] r_cvctl;
  output [7:0] r_srcctl;
  output [7:0] r_dpdmctl;
  output [7:0] r_ccrx;
  output [7:0] r_cctrx;
  output [7:0] r_ccctl;
  output [6:0] r_fcpwr;
  input [7:0] fcp_r_dat;
  input [7:0] fcp_r_sta;
  input [7:0] fcp_r_msk;
  input [7:0] fcp_r_ctl;
  input [7:0] fcp_r_crc;
  input [7:0] fcp_r_acc;
  input [7:0] fcp_r_tui;
  input [7:0] r_accctl;
  output [14:0] r_dacwr;
  input [7:0] r_dac_en;
  input [7:0] r_sar_en;
  input [7:0] r_adofs;
  input [7:0] r_isofs;
  input [5:0] x_daclsb;
  output [7:0] r_comp_opt;
  input [7:0] dac_r_ctl;
  input [7:0] dac_r_comp;
  input [7:0] dac_r_cmpsta;
  input [63:0] dac_r_vs;
  input [6:0] REVID;
  input [7:0] sfr_addr;
  input [7:0] sfr_wdat;
  output [7:0] sfr_rdat;
  input [7:0] ff_p0;
  input [7:0] di_p0;
  output [14:0] r_inst_ofs;
  output [3:0] r_ana_tm;
  output [1:0] r_gpio_ie;
  output [6:0] r_gpio_oe;
  output [6:0] r_gpio_pu;
  output [6:0] r_gpio_pd;
  output [2:0] r_gpio_s0;
  output [2:0] r_gpio_s1;
  output [2:0] r_gpio_s2;
  output [2:0] r_gpio_s3;
  output [55:0] r_regtrm;
  input [15:0] i_pc;
  input [7:0] i_i2c_rwbuf;
  input [7:0] i_i2c_ltbuf;
  input [7:0] i_i2c_ofs;
  output [4:0] o_intr;
  output [1:0] r_auto_gdcrc;
  output [4:0] r_txnumk;
  output [6:0] r_txauto;
  output [6:0] r_rxords_ena;
  output [1:0] r_spec;
  output [1:0] r_dat_spec;
  output [3:0] r_pg0_sel;
  output [7:1] r_i2c_deva;
  input [7:0] i2c_ev;
  input [2:0] prl_cpmsgid;
  input [1:0] pff_ack;
  input [1:0] prx_rst;
  input [5:0] pff_ptr;
  input [5:0] prx_adpn;
  input [7:0] pff_rdat;
  input [15:0] pff_rxpart;
  input [4:0] prx_rcvinf;
  input [2:0] ptx_fsm;
  input [3:0] prx_fsm;
  input [3:0] prl_fsm;
  input [6:0] prx_setsta;
  output [31:0] dbgpo;
  input dm_fault, cc1_di, cc2_di, di_rd_det, i_tmrf, i_vcbyval, dnchk_en,
         atpg_en, sfr_r, sfr_w, set_hold, bkpt_hold, cpurst, ictlr_idle,
         ictlr_inc, i_goidle, i_gobusy, i_i2c_idle, prl_c0set, prl_cany0,
         prl_discard, prl_GCTxDone, pff_obsd, pff_full, pff_empty, ptx_ack,
         clk_1p0m, clk_500, clk, xrstz, xclk;
  output r_pwrv_upd, aswkup, lg_dischg, gating_pwr, ps_pwrdn, r_sleep, r_pwrdn,
         r_ocdrv_enz, r_osc_stop, r_osc_lo, r_osc_gate, r_otpi_gate, r_fcpre,
         r_bclk_sel, r_psrd, r_pswr, r_fortxdat, r_fortxrdy, r_fortxen,
         r_gpio_tm, bus_idle, i2c_stretch, r_exist1st, r_ordrs4, r_fifopsh,
         r_fifopop, r_unlock, r_first, r_last, r_fiforst, r_set_cpmsgid,
         r_txendk, r_txshrt, r_auto_discard, r_hold_mcu, r_dat_portrole,
         r_dat_datarole, r_discard, r_pshords, r_strtch, r_i2c_attr,
         r_i2c_ninc, r_hwi2c_en, r_i2c_fwnak, r_i2c_fwack, srstz, prstz;
  wire   hit_223, hit_202, hit_197, hit_195, hit_194, hit_151, we_246, we_245,
         we_232, we_231, we_230, we_228, we_227, we_222, we_217, we_215,
         we_214, we_213, we_211, we_209, we_203, we_191, we_187, we_182,
         we_181, we_176, we_175, we_172, we_171, we_148, we_143, regF4_7_,
         regF4_3, regE3_0, regD3_7_, regD3_3, reg25_0_, reg19_7_, reg12_1,
         reg11_7_, reg11_4, regAD_7, N26, N27, N28, N29, N30, N32, N33, N34,
         N35, N36, N37, N38, N39, upd01, phyrst, upd12, upd18, upd19, upd20,
         upd21, lt_reg26_0, i2c_mode_upd, i2c_mode_wdat, upd31, N84, as_p0_chg,
         dmf_wkup, p0_chg_clr, di_rd_det_clr, dm_fault_clr, pwrdn_rstz,
         osc_low_clr, osc_low_rstz, r_pos_gate, m_ovp, m_ovp_sta, setAE_7,
         m_scp, m_scp_sta, s_ovp, s_ovp_sta, s_scp, s_scp_sta, lg_pulse_12m,
         N103, N104, N105, N106, N108, N109, N110, N111, N112, N113, net10815,
         net10821, n1096, n1097, n1121, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1217, n1218, n1219, n1220, n1221, n1222, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151,
         SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153,
         SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155,
         SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157,
         SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159,
         SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161,
         SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163,
         SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165,
         SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167,
         SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169,
         SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171,
         SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173,
         SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175,
         SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177,
         SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179,
         SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181,
         SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183,
         SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185,
         SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187,
         SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189,
         SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191,
         SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193,
         SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195,
         SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197,
         SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199,
         SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201,
         SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203,
         SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205,
         SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207,
         SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209,
         SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211,
         SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213,
         SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215,
         SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217,
         SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219,
         SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221,
         SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223,
         SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225,
         SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227,
         SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229,
         SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231,
         SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233,
         SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235,
         SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237,
         SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239,
         SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241,
         SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243,
         SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245,
         SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247,
         SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249,
         SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251,
         SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253,
         SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255,
         SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257,
         SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259,
         SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261,
         SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263,
         SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265,
         SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267,
         SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269,
         SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271,
         SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273,
         SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275,
         SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277,
         SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279,
         SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281,
         SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283,
         SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285,
         SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287,
         SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289,
         SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291,
         SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293,
         SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295,
         SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297,
         SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299,
         SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301,
         SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303,
         SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305,
         SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307,
         SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309,
         SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311,
         SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313,
         SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315,
         SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317,
         SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319,
         SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321,
         SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323,
         SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325,
         SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327,
         SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329,
         SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331,
         SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333,
         SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335,
         SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337,
         SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339,
         SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341,
         SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343,
         SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345,
         SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347,
         SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349,
         SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351,
         SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353,
         SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355,
         SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357,
         SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359,
         SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361,
         SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363,
         SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365,
         SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367,
         SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369,
         SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371,
         SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373,
         SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375,
         SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377,
         SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379,
         SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381,
         SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383,
         SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385,
         SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387,
         SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389,
         SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391,
         SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393,
         SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395,
         SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397,
         SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399,
         SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401,
         SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403,
         SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405,
         SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407,
         SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409,
         SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411,
         SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413,
         SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415,
         SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417,
         SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419,
         SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421,
         SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423,
         SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425,
         SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427,
         SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429,
         SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431,
         SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433,
         SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435,
         SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437,
         SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439,
         SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441,
         SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443,
         SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445,
         SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447,
         SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449,
         SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451,
         SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453,
         SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455,
         SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457,
         SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459,
         SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461,
         SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463,
         SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465,
         SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467,
         SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469,
         SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471,
         SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473,
         SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475,
         SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477,
         SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479,
         SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481,
         SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483,
         SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485,
         SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487,
         SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489,
         SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491,
         SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493,
         SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495,
         SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497,
         SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499,
         SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501,
         SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503,
         SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505,
         SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507,
         SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509,
         SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511,
         SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513,
         SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515,
         SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517,
         SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519,
         SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521,
         SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523,
         SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525,
         SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527,
         SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529,
         SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531,
         SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533,
         SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535,
         SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537,
         SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539,
         SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541,
         SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543,
         SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545,
         SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547,
         SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549,
         SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551,
         SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553,
         SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555,
         SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557,
         SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559,
         SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561,
         SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563,
         SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565,
         SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567,
         SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569,
         SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571,
         SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573,
         SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575,
         SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577,
         SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579,
         SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581,
         SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583,
         SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585,
         SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587,
         SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589,
         SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591,
         SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593,
         SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595,
         SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597,
         SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599,
         SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601,
         SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603,
         SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605,
         SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607,
         SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609,
         SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611,
         SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613,
         SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615,
         SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617,
         SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619,
         SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621,
         SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623,
         SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625,
         SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627,
         SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629,
         SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631,
         SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633,
         SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635,
         SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637,
         SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639,
         SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641,
         SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643,
         SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645,
         SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647,
         SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649,
         SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651,
         SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653,
         SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655,
         SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657,
         SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659,
         SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661,
         SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663,
         SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665,
         SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667,
         SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669,
         SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671,
         SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673,
         SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675,
         SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677,
         SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679,
         SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681,
         SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683,
         SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685,
         SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687,
         SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689,
         SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691,
         SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693,
         SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695,
         SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697,
         SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699,
         SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701,
         SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703,
         SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705,
         SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707,
         SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709,
         SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711,
         SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713,
         SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715,
         SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717,
         SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719,
         SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721,
         SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723,
         SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725,
         SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727,
         SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729,
         SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731,
         SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733,
         SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735,
         SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737,
         SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739,
         SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741,
         SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743,
         SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745,
         SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747,
         SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749,
         SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751,
         SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753,
         SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755,
         SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757,
         SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759,
         SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761,
         SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763,
         SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765,
         SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767,
         SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769,
         SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771,
         SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773,
         SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775,
         SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777,
         SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779,
         SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781,
         SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783,
         SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785,
         SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787,
         SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789,
         SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791,
         SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793,
         SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795,
         SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797,
         SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799,
         SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801,
         SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803,
         SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805,
         SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807,
         SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809,
         SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811,
         SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813,
         SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815,
         SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817,
         SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819,
         SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821,
         SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823,
         SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825,
         SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827,
         SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829,
         SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831,
         SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833,
         SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835,
         SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837,
         SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839,
         SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841,
         SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843,
         SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845,
         SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847,
         SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849,
         SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851,
         SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853,
         SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855,
         SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857,
         SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859,
         SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861,
         SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863,
         SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865,
         SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867,
         SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869,
         SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871,
         SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873,
         SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875,
         SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877,
         SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879,
         SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881,
         SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883,
         SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885,
         SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887,
         SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889,
         SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891,
         SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893,
         SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895,
         SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897,
         SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899,
         SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901,
         SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903,
         SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905,
         SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907,
         SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909,
         SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911,
         SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913,
         SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915,
         SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917,
         SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919,
         SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921,
         SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923,
         SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925,
         SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927,
         SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929,
         SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931,
         SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933,
         SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935,
         SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937,
         SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939,
         SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941,
         SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943,
         SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945,
         SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947,
         SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949,
         SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951,
         SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953,
         SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955,
         SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957,
         SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959,
         SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961,
         SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963,
         SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965,
         SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967,
         SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969,
         SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971,
         SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973,
         SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975,
         SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977,
         SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979,
         SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981,
         SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983,
         SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985,
         SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987,
         SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989,
         SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991,
         SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993,
         SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995,
         SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997,
         SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999,
         SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001,
         SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003,
         SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005,
         SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007,
         SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009,
         SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011,
         SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013,
         SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015,
         SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017;
  wire   [183:174] hit;
  wire   [167:161] we;
  wire   [3:2] regE3;
  wire   [7:0] regDF;
  wire   [7:0] regDE;
  wire   [7:0] regD4;
  wire   [7:0] reg31;
  wire   [7:0] reg30;
  wire   [7:0] reg28;
  wire   [7:0] reg27;
  wire   [7:1] reg21;
  wire   [4:0] reg20;
  wire   [7:3] reg12;
  wire   [7:0] reg06;
  wire   [7:0] reg05;
  wire   [7:0] regAF;
  wire   [7:0] regAE;
  wire   [5:0] regAD;
  wire   [7:0] regAC;
  wire   [7:0] regAB;
  wire   [7:0] reg94;
  wire   [7:0] irqAE;
  wire   [7:0] irqDF;
  wire   [7:0] irq28;
  wire   [7:0] irq04;
  wire   [7:0] irq03;
  wire   [1:0] drstz;
  wire   [4:0] rstcnt;
  wire   [1:0] r_phyrst;
  wire   [7:0] wd01;
  wire   [7:0] clr03;
  wire   [7:0] set03;
  wire   [7:0] clr04;
  wire   [7:0] set04;
  wire   [7:0] wd12;
  wire   [14:0] inst_ofs_plus;
  wire   [7:0] wd18;
  wire   [7:0] wd19;
  wire   [7:0] wd20;
  wire   [7:0] wd21;
  wire   [7:0] clr28;
  wire   [2:0] oscdwn_shft;
  wire   [3:0] osc_gate_n;
  wire   [7:0] d_p0;
  wire   [7:0] setDF;
  wire   [7:0] clrDF;
  wire   [7:0] clrAE;
  wire   [5:0] setAE;
  wire   [4:0] lg_pulse_cnt;
  wire   [3:0] lt_regE4_3_0;
  wire   [4:2] add_180_carry;

  AND2X1 U0_MASK_0 ( .A(oscdwn_shft[2]), .B(as_p0_chg), .Y(p0_chg_clr) );
  AND2X1 U0_MASK_2 ( .A(regD4[6]), .B(di_rd_det), .Y(di_rd_det_clr) );
  AND2X1 U0_MASK_3 ( .A(regD4[7]), .B(dmf_wkup), .Y(dm_fault_clr) );
  AND2X1 U0_MASK_4 ( .A(regD4[5]), .B(aswkup), .Y(osc_low_clr) );
  glreg_a0_79 u0_reg00 ( .clk(clk), .arstz(n70), .we(we_176), .wdat({n145, 
        n139, n136, n129, n122, sfr_wdat[2], n112, n107}), .rdat({r_txendk, 
        r_txauto}) );
  glreg_a0_78 u0_reg01 ( .clk(clk), .arstz(n62), .we(upd01), .wdat(wd01), 
        .rdat({r_last, r_first, r_unlock, r_txnumk}) );
  glsta_a0_6 u0_reg03 ( .clk(clk), .arstz(n37), .rst0(phyrst), .set2({
        set03[7:4], n1121, set03[2:0]}), .clr1(clr03), .rdat(dbgpo[7:0]), 
        .irq(irq03) );
  glsta_a0_5 u0_reg04 ( .clk(clk), .arstz(n58), .rst0(n17), .set2(set04), 
        .clr1(clr04), .rdat(dbgpo[15:8]), .irq(irq04) );
  glreg_a0_77 u0_reg05 ( .clk(clk), .arstz(n69), .we(we_181), .wdat({n145, 
        n139, n134, n128, n125, n119, n112, n107}), .rdat(reg05) );
  glreg_a0_76 u0_reg06 ( .clk(clk), .arstz(n64), .we(we_182), .wdat({n145, 
        n139, n134, n128, n122, sfr_wdat[2], n112, n107}), .rdat(reg06) );
  glreg_a0_75 u0_reg11 ( .clk(clk), .arstz(n55), .we(we_187), .wdat({n145, 
        n139, n134, n128, n122, sfr_wdat[2], n112, n107}), .rdat({reg11_7_, 
        r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0]}) );
  glreg_a0_74 u0_reg12 ( .clk(clk), .arstz(n67), .we(upd12), .wdat(wd12), 
        .rdat({reg12, r_txshrt, reg12_1, r_pshords}) );
  glreg_WIDTH5_2 u0_reg14 ( .clk(clk), .arstz(n79), .we(r_set_cpmsgid), .wdat(
        {n145, n139, n134, n128, n122}), .rdat({r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1]}) );
  glreg_a0_73 u0_reg15 ( .clk(clk), .arstz(n65), .we(we_191), .wdat({n145, 
        n139, n134, n128, sfr_wdat[3], n117, n112, n107}), .rdat(dbgpo[31:24])
         );
  glreg_a0_72 u0_reg18 ( .clk(clk), .arstz(n60), .we(upd18), .wdat(wd18), 
        .rdat(r_inst_ofs[7:0]) );
  glreg_a0_71 u0_reg19 ( .clk(clk), .arstz(n63), .we(upd19), .wdat(wd19), 
        .rdat({reg19_7_, r_inst_ofs[14:8]}) );
  glreg_a0_70 u0_reg20 ( .clk(clk), .arstz(n59), .we(upd20), .wdat(wd20), 
        .rdat({r_dat_spec, r_dat_datarole, reg20}) );
  glreg_a0_69 u0_reg21 ( .clk(clk), .arstz(n61), .we(upd21), .wdat(wd21), 
        .rdat({reg21, r_dat_portrole}) );
  glreg_6_00000018 u0_reg25 ( .clk(clk), .arstz(n75), .we(n1097), .wdat({n134, 
        n131, n124, sfr_wdat[2], n112, n107}), .rdat({r_i2c_attr, r_pg0_sel, 
        reg25_0_}) );
  glreg_1_1_1 u0_reg26 ( .clk(clk), .arstz(n86), .we(n1096), .wdat(n107), 
        .rdat(lt_reg26_0) );
  glreg_1_1_0 u1_reg26 ( .clk(clk), .arstz(n86), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat(r_hwi2c_en) );
  glreg_7_70 u2_reg26 ( .clk(clk), .arstz(n72), .we(n1096), .wdat({n148, n142, 
        n136, n128, n125, sfr_wdat[2], n112}), .rdat(r_i2c_deva) );
  glreg_a0_68 u0_reg27 ( .clk(clk), .arstz(n56), .we(we_203), .wdat({n145, 
        n139, n134, n128, n125, n117, n114, n109}), .rdat(reg27) );
  glsta_a0_4 u0_reg28 ( .clk(clk), .arstz(n68), .rst0(1'b0), .set2(i2c_ev), 
        .clr1(clr28), .rdat(reg28), .irq(irq28) );
  glreg_a0_67 u0_reg31 ( .clk(clk), .arstz(n57), .we(upd31), .wdat(i_pc[15:8]), 
        .rdat(reg31) );
  glreg_8_00000001 u0_regD1 ( .clk(clk), .arstz(n36), .we(we_209), .wdat({n145, 
        n139, n134, n128, n125, n119, sfr_wdat[1], n109}), .rdat({r_exist1st, 
        r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, r_gpio_oe[6], r_gpio_pu[6], 
        r_gpio_pd[6]}) );
  glreg_8_00000011 u0_regD3 ( .clk(clk), .arstz(n34), .we(we_211), .wdat({n145, 
        n139, n134, n131, n125, n117, sfr_wdat[1], n109}), .rdat({regD3_7_, 
        r_gpio_oe[5], r_gpio_pu[5], r_gpio_pd[5], regD3_3, r_gpio_oe[4], 
        r_gpio_pu[4], r_gpio_pd[4]}) );
  glreg_WIDTH3 u4_regD4 ( .clk(clk), .arstz(n86), .we(n18), .wdat({n146, n140, 
        sfr_wdat[5]}), .rdat(regD4[7:5]) );
  glreg_WIDTH2_2 u3_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n18), .wdat({
        n128, n122}), .rdat(regD4[4:3]) );
  glreg_WIDTH1_5 u2_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n18), .wdat(
        n119), .rdat(regD4[2]) );
  glreg_WIDTH1_4 u1_regD4 ( .clk(clk), .arstz(osc_low_rstz), .we(n18), .wdat(
        n112), .rdat(regD4[1]) );
  glreg_WIDTH1_3 u0_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n18), .wdat(
        n107), .rdat(regD4[0]) );
  glreg_8_000000f0 u0_regD5 ( .clk(clk), .arstz(n30), .we(we_213), .wdat({n148, 
        n142, n136, n131, n125, n117, sfr_wdat[1:0]}), .rdat({r_gpio_pu[3:0], 
        r_gpio_pd[3:0]}) );
  glreg_8_00000098 u0_regD6 ( .clk(clk), .arstz(n32), .we(we_214), .wdat({n148, 
        n140, sfr_wdat[5], n131, n124, n117, sfr_wdat[1:0]}), .rdat({
        r_gpio_oe[1], r_gpio_s1, r_gpio_oe[0], r_gpio_s0}) );
  glreg_8_00000032 u0_regD7 ( .clk(clk), .arstz(n31), .we(we_215), .wdat({n146, 
        n140, n136, n131, n125, n117, n114, sfr_wdat[0]}), .rdat({r_gpio_oe[3], 
        r_gpio_s3, r_gpio_oe[2], r_gpio_s2}) );
  glreg_a0_66 u0_regD9 ( .clk(clk), .arstz(n51), .we(we_217), .wdat({n146, 
        n140, sfr_wdat[5], n129, n125, n117, sfr_wdat[1:0]}), .rdat({r_ana_tm, 
        r_fortxdat, r_fortxrdy, r_fortxen, r_sleep}) );
  glreg_a0_65 u0_regDE ( .clk(clk), .arstz(n53), .we(we_222), .wdat({n146, 
        n140, sfr_wdat[5], n129, n125, n117, n114, sfr_wdat[0]}), .rdat(regDE)
         );
  glsta_a0_3 u0_regDF ( .clk(clk), .arstz(n71), .rst0(1'b0), .set2(setDF), 
        .clr1(clrDF), .rdat(regDF), .irq(irqDF) );
  glreg_a0_64 u0_reg8F ( .clk(clk), .arstz(n49), .we(we_143), .wdat({n146, 
        n140, sfr_wdat[5], n129, n123, n117, n114, sfr_wdat[0]}), .rdat(
        r_dpdmctl) );
  glreg_WIDTH4 u0_reg94 ( .clk(clk), .arstz(n80), .we(we_148), .wdat({n140, 
        sfr_wdat[5], n129, n123}), .rdat(reg94[6:3]) );
  glreg_a0_63 u0_regA1 ( .clk(clk), .arstz(n52), .we(we[161]), .wdat({n146, 
        n140, sfr_wdat[5], n129, n123, n117, n114, n109}), .rdat(r_regtrm[7:0]) );
  glreg_a0_62 u0_regA2 ( .clk(clk), .arstz(n47), .we(we[162]), .wdat({n146, 
        n140, n136, n129, n123, n118, n114, n109}), .rdat(r_regtrm[15:8]) );
  glreg_a0_61 u0_regA3 ( .clk(clk), .arstz(n50), .we(we[163]), .wdat({n146, 
        n141, n136, n129, n123, n118, n113, n109}), .rdat(r_regtrm[23:16]) );
  glreg_a0_60 u0_regA4 ( .clk(clk), .arstz(n54), .we(we[164]), .wdat({n146, 
        n141, n135, n129, n123, n118, n113, n108}), .rdat(r_regtrm[31:24]) );
  glreg_a0_59 u0_regA5 ( .clk(clk), .arstz(n48), .we(we[165]), .wdat({n147, 
        n141, n135, n129, n123, n118, n113, n108}), .rdat(r_regtrm[39:32]) );
  glreg_a0_58 u0_regA6 ( .clk(clk), .arstz(n43), .we(we[166]), .wdat({n147, 
        n141, n135, n130, n123, n118, n113, n108}), .rdat(r_regtrm[47:40]) );
  glreg_a0_57 u0_regA7 ( .clk(clk), .arstz(n46), .we(we[167]), .wdat({n147, 
        n141, n135, n130, n123, n118, n113, n108}), .rdat(r_regtrm[55:48]) );
  glreg_a0_56 u0_regAB ( .clk(clk), .arstz(n41), .we(we_171), .wdat({n147, 
        n141, n135, n130, n123, n118, n113, n108}), .rdat(regAB) );
  glreg_8_00000028 u0_regAC ( .clk(clk), .arstz(n33), .we(we_172), .wdat({n147, 
        n141, n136, n130, n124, n118, n113, n108}), .rdat(regAC) );
  dbnc_WIDTH4_TIMEOUT14_2 u2_ovp_db ( .o_dbc(reg94[2]), .o_chg(), .i_org(
        srci[2]), .clk(clk_500), .rstz(n76) );
  dbnc_WIDTH4_TIMEOUT14_1 u1_ocp_db ( .o_dbc(reg94[1]), .o_chg(), .i_org(
        srci[1]), .clk(clk_500), .rstz(n78) );
  dbnc_WIDTH4_TIMEOUT14_0 u1_uvp_db ( .o_dbc(reg94[0]), .o_chg(), .i_org(
        srci[0]), .clk(clk_500), .rstz(n77) );
  dbnc_WIDTH5_TIMEOUT30 u1_ovp_db ( .o_dbc(m_ovp), .o_chg(m_ovp_sta), .i_org(
        srci[2]), .clk(clk_1p0m), .rstz(n73) );
  dbnc_WIDTH2_4 u0_otpi_db ( .o_dbc(regAD[3]), .o_chg(setAE[3]), .i_org(
        srci[5]), .clk(clk_1p0m), .rstz(n80) );
  dbnc_WIDTH2_3 u0_ocp_db ( .o_dbc(regAD[1]), .o_chg(setAE[1]), .i_org(srci[1]), .clk(clk_1p0m), .rstz(n81) );
  dbnc_WIDTH2_2 u0_uvp_db ( .o_dbc(regAD[0]), .o_chg(setAE[0]), .i_org(srci[0]), .clk(clk_1p0m), .rstz(n85) );
  dbnc_WIDTH2_1 u1_scp_db ( .o_dbc(m_scp), .o_chg(m_scp_sta), .i_org(srci[3]), 
        .clk(clk_1p0m), .rstz(n82) );
  dbnc_WIDTH2_0 u0_dmf_db ( .o_dbc(regAD_7), .o_chg(setAE_7), .i_org(dm_fault), 
        .clk(clk_1p0m), .rstz(n81) );
  dbnc_WIDTH2_TIMEOUT2_14 u0_otps_db ( .o_dbc(reg94[7]), .o_chg(), .i_org(
        srci[5]), .clk(clk), .rstz(n83) );
  dbnc_WIDTH2_TIMEOUT2_13 u0_cc1_db ( .o_dbc(regF4_3), .o_chg(), .i_org(cc1_di), .clk(clk), .rstz(n82) );
  dbnc_WIDTH2_TIMEOUT2_12 u0_cc2_db ( .o_dbc(regF4_7_), .o_chg(), .i_org(
        cc2_di), .clk(clk), .rstz(n84) );
  dbnc_WIDTH2_TIMEOUT2_11 u0_ovp_db ( .o_dbc(s_ovp), .o_chg(s_ovp_sta), 
        .i_org(srci[2]), .clk(clk), .rstz(n83) );
  dbnc_WIDTH2_TIMEOUT2_10 u0_scp_db ( .o_dbc(s_scp), .o_chg(s_scp_sta), 
        .i_org(srci[3]), .clk(clk), .rstz(n85) );
  dbnc_WIDTH2_TIMEOUT2_9 u0_v5oc_db ( .o_dbc(regAD[5]), .o_chg(setAE[5]), 
        .i_org(srci[4]), .clk(clk), .rstz(n84) );
  glsta_a0_2 u0_regAE ( .clk(clk), .arstz(n66), .rst0(1'b0), .set2({setAE_7, 
        1'b0, setAE}), .clr1(clrAE), .rdat(regAE), .irq(irqAE) );
  glreg_a0_55 u0_regAF ( .clk(clk), .arstz(n40), .we(we_175), .wdat({n147, 
        n141, n135, n130, n124, n118, n113, n108}), .rdat(regAF) );
  glreg_WIDTH7_2 u0_regE3 ( .clk(clk), .arstz(n74), .we(we_227), .wdat({n147, 
        n141, n135, n130, n124, n118, n108}), .rdat({r_srcctl[7:4], regE3, 
        regE3_0}) );
  glreg_4_00000004 u1_regE4 ( .clk(clk), .arstz(n79), .we(r_pwrv_upd), .wdat(
        lt_regE4_3_0), .rdat(r_fw_pwrv[3:0]) );
  glreg_8_00000004 u0_regE4 ( .clk(clk), .arstz(n35), .we(we_228), .wdat({n147, 
        n142, n135, n130, n124, n119, n113, n108}), .rdat({r_pwrctl, 
        lt_regE4_3_0}) );
  glreg_8_0000001f u0_regE5 ( .clk(clk), .arstz(n29), .we(r_pwrv_upd), .wdat({
        n147, n142, n136, n131, n125, n119, n114, n109}), .rdat(
        r_fw_pwrv[11:4]) );
  glreg_a0_54 u0_regE6 ( .clk(clk), .arstz(n44), .we(we_230), .wdat({n147, 
        n141, n135, n130, n124, n119, n113, n108}), .rdat(r_ccrx) );
  glreg_a0_53 u0_regE7 ( .clk(clk), .arstz(n39), .we(we_231), .wdat({n148, 
        n142, n136, n130, n124, n119, n114, n109}), .rdat(r_ccctl) );
  glreg_a0_52 u0_regE8 ( .clk(clk), .arstz(n45), .we(we_232), .wdat({n148, 
        n142, n136, n131, n124, n119, n114, n109}), .rdat(r_comp_opt) );
  glreg_a0_51 u0_regF5 ( .clk(clk), .arstz(n38), .we(we_245), .wdat({n148, 
        n142, n135, n130, n124, n119, n114, n109}), .rdat(r_cvctl) );
  glreg_a0_50 u0_regF6 ( .clk(clk), .arstz(n42), .we(we_246), .wdat({n146, 
        n140, n134, n128, n122, sfr_wdat[2], n112, n107}), .rdat(r_cctrx) );
  SNPS_CLOCK_GATE_HIGH_regbank_a0_1 clk_gate_rstcnt_reg ( .CLK(clk), .EN(N26), 
        .ENCLK(net10815), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_regbank_a0_0 clk_gate_lg_pulse_cnt_reg ( .CLK(clk_1p0m), 
        .EN(N108), .ENCLK(net10821), .TE(1'b0) );
  regbank_a0_DW01_add_0 add_526 ( .A(regAC), .B(regAB), .CI(1'b0), .SUM(
        r_pwr_i), .CO() );
  regbank_a0_DW01_inc_0 add_304 ( .A({1'b0, r_inst_ofs}), .SUM({
        SYNOPSYS_UNCONNECTED_1, inst_ofs_plus}) );
  regbank_a0_DW_rightsh_0 srl_133 ( .A({dac_r_vs, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, r_cctrx, r_cvctl, regF4_7_, x_daclsb[5:3], regF4_3, 
        x_daclsb[2:0], r_sar_en, r_dac_en, dac_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_comp_opt, r_ccctl, r_ccrx, r_fw_pwrv[11:4], r_pwrctl, r_fw_pwrv[3:0], 
        r_srcctl[7:4], regE3, r_srcctl[1], regE3_0, dac_r_cmpsta, dac_r_comp, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, regDF, regDE, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_ana_tm, r_fortxdat, 
        r_fortxrdy, r_fortxen, r_sleep, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, r_gpio_oe[3], r_gpio_s3, r_gpio_oe[2], r_gpio_s2, 
        r_gpio_oe[1], r_gpio_s1, r_gpio_oe[0], r_gpio_s0, r_gpio_pu[3:0], 
        r_gpio_pd[3:0], regD4, regD3_7_, r_gpio_oe[5], r_gpio_pu[5], 
        r_gpio_pd[5], regD3_3, r_gpio_oe[4], r_gpio_pu[4], r_gpio_pd[4], 
        i_i2c_rwbuf, r_exist1st, r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, 
        r_gpio_oe[6], r_gpio_pu[6], r_gpio_pd[6], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, reg31, reg30, i_i2c_ltbuf, reg28, reg27, r_i2c_deva, 
        r_hwi2c_en, 1'b0, 1'b0, r_i2c_attr, r_pg0_sel, reg25_0_, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, prx_rcvinf[4], REVID, 
        prx_rcvinf[3], ptx_fsm, prx_fsm, reg21, r_dat_portrole, r_dat_spec, 
        r_dat_datarole, reg20, n11, r_inst_ofs, i_i2c_ofs, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, dbgpo[31:24], r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1], prl_cpmsgid, prl_cany0, 
        prx_rcvinf[2:0], prl_fsm, reg12, r_txshrt, reg12_1, r_pshords, 
        reg11_7_, r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0], 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, pff_empty, 
        pff_full, pff_ptr, reg06, reg05, dbgpo[15:0], pff_rdat, r_last, 
        r_first, r_unlock, r_txnumk, r_txendk, r_txauto, regAF, regAE, regAD_7, 
        1'b0, regAD, regAC, regAB, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_regtrm, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, fcp_r_crc, fcp_r_dat, fcp_r_msk, fcp_r_sta, 
        fcp_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, fcp_r_acc, r_accctl, fcp_r_tui, reg94, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, r_isofs, r_adofs, r_dpdmctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_cvofs, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .DATA_TC(1'b0), .SH({sfr_addr[6:0], 1'b0, 
        1'b0, 1'b0}), .B({SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, 
        SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, 
        SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, 
        SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, 
        SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, 
        SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, 
        SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, 
        SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, 
        SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, 
        SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, 
        SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, 
        SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, 
        SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, 
        SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, 
        SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, 
        SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, 
        SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, 
        SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, 
        SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, 
        SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, 
        SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, 
        SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, 
        SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, 
        SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, 
        SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, 
        SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, 
        SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, 
        SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, 
        SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, 
        SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, 
        SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, 
        SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, 
        SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, 
        SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, 
        SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, 
        SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, 
        SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, 
        SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, 
        SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, 
        SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, 
        SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, 
        SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, 
        SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, 
        SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, 
        SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, 
        SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, 
        SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, 
        SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, 
        SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, 
        SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, 
        SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, 
        SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, 
        SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, 
        SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, 
        SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, 
        SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, 
        SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, 
        SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, 
        SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, 
        SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, 
        SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, 
        SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, 
        SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, 
        SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, 
        SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, 
        SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, 
        SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, 
        SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, 
        SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, 
        SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, 
        SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, 
        SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, 
        SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, 
        SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, 
        SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, 
        SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, 
        SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, 
        SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, 
        SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, 
        SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, 
        SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, 
        SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, 
        SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, 
        SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, 
        SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, 
        SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, 
        SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, 
        SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, 
        SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, 
        SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, 
        SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, 
        SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, 
        SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, 
        SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, 
        SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, 
        SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, 
        SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, 
        SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, 
        SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, 
        SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, 
        SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, 
        SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, 
        SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, 
        SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, 
        SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, 
        SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, 
        SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, 
        SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, 
        SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, 
        SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, 
        SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, 
        SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, 
        SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, 
        SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, 
        SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, 
        SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, 
        SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, 
        SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, 
        SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, 
        SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, 
        SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, 
        SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, 
        SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, 
        SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, 
        SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, 
        SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, 
        SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, 
        SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, 
        SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, 
        SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, 
        SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, 
        SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, 
        SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, 
        SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, 
        SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, 
        SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, 
        SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, 
        SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, 
        SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, 
        SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, 
        SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, 
        SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, 
        SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, 
        SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, 
        SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, 
        SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, 
        SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, 
        SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, 
        SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, 
        SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, 
        SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, 
        SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, 
        SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, 
        SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, 
        SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, 
        SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, 
        SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, 
        SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, 
        SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, 
        SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, 
        SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, 
        SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, 
        SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, 
        SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, 
        SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, 
        SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, 
        SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, 
        SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, 
        SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, 
        SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, 
        SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, 
        SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, 
        SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, 
        SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, 
        SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, 
        SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, 
        SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, 
        SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, 
        SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, 
        SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, 
        SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, 
        SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, 
        SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, 
        SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, 
        SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, 
        SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, 
        SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, 
        SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, 
        SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, 
        SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, 
        SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, 
        SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, 
        SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, 
        SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, 
        SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, 
        SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, 
        SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, 
        SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, 
        SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, 
        SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, 
        SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, 
        SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, 
        SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, 
        SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, 
        SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, 
        SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, 
        SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, 
        SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, 
        SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, 
        SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, 
        SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, 
        SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, 
        SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, 
        SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, 
        SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, 
        SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, 
        SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, 
        SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, 
        SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, 
        SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, 
        SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, 
        SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, 
        SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, 
        SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, 
        SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, 
        SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, 
        SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, 
        SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, 
        SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, 
        SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, 
        SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, 
        SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, 
        SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, 
        SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, 
        SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, 
        SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, 
        SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, 
        SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, 
        SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, 
        SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, 
        SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, 
        SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, 
        SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, 
        SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, 
        SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, 
        SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, 
        SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, 
        SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, 
        SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, 
        SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, 
        SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, 
        SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, 
        SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, 
        SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, 
        SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, 
        SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, 
        SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, 
        SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, 
        SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, 
        SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, 
        SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, 
        SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, 
        SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, 
        SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, 
        SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, 
        SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, 
        SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, 
        SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, 
        SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, 
        SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, 
        SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, 
        SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, 
        SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, 
        SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, 
        SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, 
        SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, 
        SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, 
        SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, 
        SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, 
        SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017, sfr_rdat}) );
  HAD1X1 add_180_U1_1_1 ( .A(N29), .B(N30), .CO(add_180_carry[2]), .SO(N32) );
  HAD1X1 add_180_U1_1_2 ( .A(N28), .B(add_180_carry[2]), .CO(add_180_carry[3]), 
        .SO(N33) );
  HAD1X1 add_180_U1_1_3 ( .A(N27), .B(add_180_carry[3]), .CO(add_180_carry[4]), 
        .SO(N34) );
  DFFRQX1 r_phyrst_reg_0_ ( .D(n1221), .C(clk), .XR(n6), .Q(r_phyrst[0]) );
  DFFRQX1 lg_pulse_cnt_reg_4_ ( .D(N113), .C(net10821), .XR(n87), .Q(
        lg_pulse_cnt[4]) );
  DFFRQX1 lg_pulse_cnt_reg_2_ ( .D(N111), .C(net10821), .XR(n87), .Q(
        lg_pulse_cnt[2]) );
  DFFRQX1 lg_pulse_cnt_reg_3_ ( .D(N112), .C(net10821), .XR(n87), .Q(
        lg_pulse_cnt[3]) );
  DFFRQX1 lg_pulse_cnt_reg_1_ ( .D(N110), .C(net10821), .XR(n87), .Q(
        lg_pulse_cnt[1]) );
  DFFRQX1 rstcnt_reg_0_ ( .D(N39), .C(net10815), .XR(n7), .Q(rstcnt[0]) );
  DFFRQX1 lg_pulse_cnt_reg_0_ ( .D(N109), .C(net10821), .XR(n86), .Q(
        lg_pulse_cnt[0]) );
  DFFRQX1 d_p0_reg_7_ ( .D(ff_p0[7]), .C(clk), .XR(n86), .Q(d_p0[7]) );
  DFFRQX1 d_p0_reg_6_ ( .D(ff_p0[6]), .C(clk), .XR(n86), .Q(d_p0[6]) );
  DFFRQX1 d_p0_reg_5_ ( .D(ff_p0[5]), .C(clk), .XR(n86), .Q(d_p0[5]) );
  DFFRQX1 d_p0_reg_4_ ( .D(ff_p0[4]), .C(clk), .XR(n87), .Q(d_p0[4]) );
  DFFRQX1 d_p0_reg_3_ ( .D(ff_p0[3]), .C(clk), .XR(n86), .Q(d_p0[3]) );
  DFFRQX1 d_p0_reg_2_ ( .D(ff_p0[2]), .C(clk), .XR(n87), .Q(d_p0[2]) );
  DFFRQX1 d_p0_reg_1_ ( .D(ff_p0[1]), .C(clk), .XR(n87), .Q(d_p0[1]) );
  DFFRQX1 d_p0_reg_0_ ( .D(ff_p0[0]), .C(clk), .XR(n87), .Q(d_p0[0]) );
  DFFRQX1 r_phyrst_reg_1_ ( .D(n1220), .C(clk), .XR(n6), .Q(r_phyrst[1]) );
  DFFNRQX1 osc_gate_n_reg_3_ ( .D(osc_gate_n[2]), .XC(xclk), .XR(n6), .Q(
        osc_gate_n[3]) );
  DFFNRQX1 osc_gate_n_reg_0_ ( .D(r_pos_gate), .XC(xclk), .XR(n7), .Q(
        osc_gate_n[0]) );
  DFFNRQX1 osc_gate_n_reg_1_ ( .D(osc_gate_n[0]), .XC(xclk), .XR(n7), .Q(
        osc_gate_n[1]) );
  DFFNRQX1 osc_gate_n_reg_2_ ( .D(osc_gate_n[1]), .XC(xclk), .XR(n6), .Q(
        osc_gate_n[2]) );
  DFFQX1 oscdwn_shft_reg_1_ ( .D(oscdwn_shft[0]), .C(clk), .Q(oscdwn_shft[1])
         );
  DFFQX1 oscdwn_shft_reg_2_ ( .D(n219), .C(clk), .Q(oscdwn_shft[2]) );
  DFFRQX1 rstcnt_reg_1_ ( .D(N38), .C(net10815), .XR(n7), .Q(rstcnt[1]) );
  DFFRQX1 rstcnt_reg_2_ ( .D(N37), .C(net10815), .XR(n6), .Q(rstcnt[2]) );
  DFFRQX1 drstz_reg_1_ ( .D(drstz[0]), .C(clk), .XR(n6), .Q(drstz[1]) );
  DFFRQX1 rstcnt_reg_3_ ( .D(N36), .C(net10815), .XR(n7), .Q(rstcnt[3]) );
  DFFRQX1 rstcnt_reg_4_ ( .D(N35), .C(net10815), .XR(n6), .Q(rstcnt[4]) );
  DFFRQX1 lg_pulse_12m_reg ( .D(n1218), .C(clk), .XR(n87), .Q(lg_pulse_12m) );
  DFFRQX1 lg_pulse_reg ( .D(n1219), .C(clk_1p0m), .XR(n87), .Q(lg_dischg) );
  DFFQX1 oscdwn_shft_reg_0_ ( .D(N84), .C(clk), .Q(oscdwn_shft[0]) );
  DFFRQX1 drstz_reg_0_ ( .D(1'b1), .C(clk), .XR(n7), .Q(drstz[0]) );
  AND2X1 U3 ( .A(n204), .B(n230), .Y(r_dacwr[8]) );
  NOR2X1 U4 ( .A(n239), .B(n184), .Y(n18) );
  INVX1 U5 ( .A(n175), .Y(n4) );
  INVX1 U6 ( .A(sfr_w), .Y(n175) );
  INVX1 U7 ( .A(xrstz), .Y(n5) );
  INVX1 U11 ( .A(n5), .Y(n6) );
  INVX1 U12 ( .A(n5), .Y(n7) );
  BUFXL U13 ( .A(sfr_addr[6]), .Y(n8) );
  BUFXL U14 ( .A(sfr_addr[5]), .Y(n9) );
  INVX1 U15 ( .A(n105), .Y(n10) );
  INVX1 U16 ( .A(n199), .Y(n11) );
  BUFX3 U17 ( .A(n1127), .Y(n12) );
  INVX1 U18 ( .A(n1134), .Y(n13) );
  INVX1 U19 ( .A(n250), .Y(n14) );
  INVX1 U20 ( .A(n186), .Y(n230) );
  BUFX3 U21 ( .A(n244), .Y(n15) );
  AND2X1 U22 ( .A(pff_ack[0]), .B(n15), .Y(set04[4]) );
  BUFX3 U23 ( .A(n1126), .Y(n16) );
  BUFX3 U24 ( .A(phyrst), .Y(n17) );
  BUFXL U25 ( .A(pff_ptr[4]), .Y(dbgpo[20]) );
  BUFXL U26 ( .A(pff_ptr[0]), .Y(dbgpo[16]) );
  BUFXL U27 ( .A(pff_ptr[1]), .Y(dbgpo[17]) );
  BUFXL U28 ( .A(pff_ptr[5]), .Y(dbgpo[21]) );
  BUFXL U29 ( .A(pff_ptr[3]), .Y(dbgpo[19]) );
  BUFXL U30 ( .A(pff_ptr[2]), .Y(dbgpo[18]) );
  INVXL U31 ( .A(n239), .Y(n232) );
  NAND21XL U32 ( .B(n239), .A(n221), .Y(n1189) );
  NAND21XL U33 ( .B(n239), .A(n241), .Y(n1127) );
  NAND21XL U34 ( .B(n175), .A(n224), .Y(n156) );
  NAND21XL U35 ( .B(n175), .A(n227), .Y(n162) );
  NAND21XL U36 ( .B(n175), .A(n238), .Y(n167) );
  NAND21XL U37 ( .B(n175), .A(n240), .Y(n158) );
  NAND21XL U38 ( .B(n175), .A(n237), .Y(n176) );
  NAND21XL U39 ( .B(n186), .A(n226), .Y(n1125) );
  NAND41X1 U40 ( .D(prl_cany0), .A(prx_rcvinf[4]), .B(i_i2c_idle), .C(n1211), 
        .Y(n1185) );
  INVX1 U41 ( .A(n127), .Y(n122) );
  AND2X1 U42 ( .A(n203), .B(n232), .Y(r_dacwr[4]) );
  NAND21X1 U43 ( .B(n191), .A(n112), .Y(n194) );
  NOR2X1 U44 ( .A(n137), .B(n1189), .Y(clr04[5]) );
  NOR2X1 U45 ( .A(n133), .B(n1189), .Y(clr04[4]) );
  NOR2X1 U46 ( .A(n111), .B(n1189), .Y(clr04[0]) );
  NOR3XL U47 ( .A(n1150), .B(n133), .C(n121), .Y(r_discard) );
  NOR2X1 U48 ( .A(n116), .B(n1189), .Y(clr04[1]) );
  NOR2X1 U49 ( .A(n144), .B(n1189), .Y(clr04[6]) );
  NOR2X1 U50 ( .A(n120), .B(n1189), .Y(clr04[2]) );
  NOR2X1 U51 ( .A(n150), .B(n1189), .Y(clr04[7]) );
  NOR2X1 U52 ( .A(n126), .B(n1189), .Y(clr04[3]) );
  INVX1 U53 ( .A(n191), .Y(we_227) );
  AND2X1 U54 ( .A(n205), .B(n232), .Y(we_228) );
  INVX1 U55 ( .A(n143), .Y(n139) );
  INVX1 U56 ( .A(n111), .Y(n107) );
  INVX1 U57 ( .A(n115), .Y(n112) );
  INVX1 U58 ( .A(n150), .Y(n145) );
  INVX1 U59 ( .A(n133), .Y(n128) );
  INVX1 U60 ( .A(n143), .Y(n142) );
  INVX1 U61 ( .A(n150), .Y(n148) );
  INVX1 U62 ( .A(n133), .Y(n130) );
  INVX1 U63 ( .A(n150), .Y(n147) );
  INVX1 U64 ( .A(n111), .Y(n108) );
  INVX1 U65 ( .A(n138), .Y(n135) );
  INVX1 U66 ( .A(n116), .Y(n113) );
  INVX1 U67 ( .A(n144), .Y(n141) );
  INVX1 U68 ( .A(n121), .Y(n118) );
  INVX1 U69 ( .A(n126), .Y(n123) );
  INVX1 U70 ( .A(n143), .Y(n140) );
  INVX1 U71 ( .A(n150), .Y(n146) );
  INVX1 U72 ( .A(n121), .Y(n117) );
  INVX1 U73 ( .A(n138), .Y(n134) );
  INVX1 U74 ( .A(n133), .Y(n129) );
  INVX1 U75 ( .A(n126), .Y(n124) );
  INVX1 U76 ( .A(n138), .Y(n136) );
  INVX1 U77 ( .A(n133), .Y(n131) );
  INVX1 U78 ( .A(n120), .Y(n119) );
  INVX1 U79 ( .A(n111), .Y(n109) );
  INVX1 U80 ( .A(n115), .Y(n114) );
  INVX1 U81 ( .A(n126), .Y(n125) );
  INVX1 U82 ( .A(n88), .Y(n86) );
  INVX1 U83 ( .A(n88), .Y(n87) );
  INVX1 U84 ( .A(n90), .Y(n79) );
  INVX1 U85 ( .A(n89), .Y(n84) );
  INVX1 U86 ( .A(n88), .Y(n85) );
  INVX1 U87 ( .A(n89), .Y(n82) );
  INVX1 U88 ( .A(n90), .Y(n81) );
  INVX1 U89 ( .A(n94), .Y(n66) );
  INVX1 U90 ( .A(n89), .Y(n71) );
  INVX1 U91 ( .A(n100), .Y(n68) );
  INVX1 U92 ( .A(n93), .Y(n58) );
  INVX1 U93 ( .A(n97), .Y(n37) );
  INVX1 U94 ( .A(n96), .Y(n42) );
  INVX1 U95 ( .A(n97), .Y(n38) );
  INVX1 U96 ( .A(n95), .Y(n45) );
  INVX1 U97 ( .A(n97), .Y(n39) );
  INVX1 U98 ( .A(n95), .Y(n44) );
  INVX1 U99 ( .A(n96), .Y(n40) );
  INVX1 U100 ( .A(n89), .Y(n83) );
  INVX1 U101 ( .A(n96), .Y(n41) );
  INVX1 U102 ( .A(n100), .Y(n46) );
  INVX1 U103 ( .A(n95), .Y(n43) );
  INVX1 U104 ( .A(n94), .Y(n48) );
  INVX1 U105 ( .A(n94), .Y(n54) );
  INVX1 U106 ( .A(n97), .Y(n50) );
  INVX1 U107 ( .A(n1222), .Y(n47) );
  INVX1 U108 ( .A(n94), .Y(n52) );
  INVX1 U109 ( .A(n90), .Y(n80) );
  INVX1 U110 ( .A(n96), .Y(n49) );
  INVX1 U111 ( .A(n94), .Y(n53) );
  INVX1 U112 ( .A(n95), .Y(n51) );
  INVX1 U113 ( .A(n96), .Y(n57) );
  INVX1 U114 ( .A(n100), .Y(n56) );
  INVX1 U115 ( .A(n100), .Y(n61) );
  INVX1 U116 ( .A(n93), .Y(n59) );
  INVX1 U117 ( .A(n101), .Y(n63) );
  INVX1 U118 ( .A(n93), .Y(n60) );
  INVX1 U119 ( .A(n93), .Y(n65) );
  INVX1 U120 ( .A(n93), .Y(n67) );
  INVX1 U121 ( .A(n101), .Y(n55) );
  INVX1 U122 ( .A(n89), .Y(n64) );
  INVX1 U123 ( .A(n88), .Y(n69) );
  INVX1 U124 ( .A(n100), .Y(n62) );
  INVX1 U125 ( .A(n98), .Y(n70) );
  INVX1 U126 ( .A(n90), .Y(n72) );
  INVX1 U127 ( .A(n92), .Y(n74) );
  INVX1 U128 ( .A(n92), .Y(n73) );
  INVX1 U129 ( .A(n92), .Y(n75) );
  INVX1 U130 ( .A(n91), .Y(n77) );
  INVX1 U131 ( .A(n91), .Y(n78) );
  INVX1 U132 ( .A(n91), .Y(n76) );
  INVX1 U133 ( .A(atpg_en), .Y(n152) );
  INVX1 U134 ( .A(sfr_wdat[3]), .Y(n127) );
  AND2X1 U135 ( .A(n203), .B(n212), .Y(r_dacwr[7]) );
  AND2X1 U136 ( .A(n203), .B(n217), .Y(r_dacwr[5]) );
  AND2X1 U137 ( .A(n203), .B(n213), .Y(r_dacwr[6]) );
  AND2X1 U138 ( .A(n203), .B(n210), .Y(r_dacwr[3]) );
  AND2X1 U139 ( .A(n203), .B(n206), .Y(r_dacwr[2]) );
  AND2X1 U140 ( .A(n203), .B(n230), .Y(r_dacwr[1]) );
  INVX1 U141 ( .A(n202), .Y(n203) );
  INVX1 U142 ( .A(sfr_wdat[7]), .Y(n149) );
  INVX1 U143 ( .A(sfr_wdat[6]), .Y(n143) );
  INVX1 U144 ( .A(sfr_wdat[0]), .Y(n110) );
  INVX1 U145 ( .A(sfr_wdat[5]), .Y(n137) );
  INVX1 U146 ( .A(sfr_wdat[2]), .Y(n120) );
  INVX1 U147 ( .A(sfr_wdat[1]), .Y(n115) );
  INVX1 U148 ( .A(sfr_wdat[4]), .Y(n132) );
  INVX1 U149 ( .A(sfr_wdat[3]), .Y(n126) );
  NOR2X1 U150 ( .A(n149), .B(n1125), .Y(r_i2c_fwack) );
  NOR2X1 U151 ( .A(n137), .B(n1188), .Y(clr28[5]) );
  NOR2X1 U152 ( .A(n116), .B(n1188), .Y(clr28[1]) );
  NOR2X1 U153 ( .A(n132), .B(n1188), .Y(clr28[4]) );
  NOR2X1 U154 ( .A(n111), .B(n1188), .Y(clr28[0]) );
  NOR2X1 U155 ( .A(n144), .B(n1188), .Y(clr28[6]) );
  NOR2X1 U156 ( .A(n121), .B(n1188), .Y(clr28[2]) );
  NOR2X1 U157 ( .A(n144), .B(n1125), .Y(r_i2c_fwnak) );
  NAND4X1 U158 ( .A(n249), .B(n122), .C(n1180), .D(n139), .Y(n1150) );
  NOR2X1 U159 ( .A(n107), .B(n149), .Y(n1180) );
  AND2X1 U160 ( .A(n206), .B(n205), .Y(r_dacwr[12]) );
  INVX1 U161 ( .A(n1137), .Y(n250) );
  NOR2X1 U162 ( .A(n150), .B(n1188), .Y(clr28[7]) );
  NOR2X1 U163 ( .A(n126), .B(n1188), .Y(clr28[3]) );
  INVX1 U164 ( .A(n164), .Y(r_pwrv_upd) );
  AND2X1 U165 ( .A(n204), .B(n232), .Y(r_dacwr[11]) );
  AND2X1 U166 ( .A(n185), .B(n217), .Y(we_213) );
  AND2X1 U167 ( .A(n185), .B(n210), .Y(we_211) );
  AND2X1 U168 ( .A(n185), .B(n230), .Y(we_209) );
  AND2X1 U169 ( .A(n180), .B(n212), .Y(we[167]) );
  AND2X1 U170 ( .A(n180), .B(n213), .Y(we[166]) );
  AND2X1 U171 ( .A(n180), .B(n217), .Y(we[165]) );
  AND2X1 U172 ( .A(n180), .B(n232), .Y(we[164]) );
  AND2X1 U173 ( .A(n180), .B(n210), .Y(we[163]) );
  AND2X1 U174 ( .A(n180), .B(n206), .Y(we[162]) );
  AND2X1 U175 ( .A(n180), .B(n230), .Y(we[161]) );
  AND2X1 U176 ( .A(n204), .B(n210), .Y(r_dacwr[10]) );
  AND2X1 U177 ( .A(n204), .B(n206), .Y(r_dacwr[9]) );
  AND2X1 U178 ( .A(n204), .B(n213), .Y(we_246) );
  AND2X1 U179 ( .A(n204), .B(n217), .Y(we_245) );
  AND2X1 U180 ( .A(n223), .B(n232), .Y(we_172) );
  AND2X1 U181 ( .A(n213), .B(n221), .Y(we_182) );
  AND2X1 U182 ( .A(n217), .B(n221), .Y(we_181) );
  AND2X1 U183 ( .A(n212), .B(n185), .Y(we_215) );
  AND2X1 U184 ( .A(n213), .B(n185), .Y(we_214) );
  AND2X1 U185 ( .A(n210), .B(n226), .Y(we_203) );
  AND2X1 U186 ( .A(n212), .B(n223), .Y(we_175) );
  AND2X1 U187 ( .A(n210), .B(n223), .Y(we_171) );
  AND2X1 U188 ( .A(n212), .B(n205), .Y(we_231) );
  AND2X1 U189 ( .A(n213), .B(n205), .Y(we_230) );
  AND2X1 U190 ( .A(n212), .B(n188), .Y(we_191) );
  AND2X1 U191 ( .A(n210), .B(n188), .Y(we_187) );
  INVX1 U192 ( .A(n1125), .Y(n1097) );
  INVX1 U193 ( .A(sfr_wdat[0]), .Y(n111) );
  INVX1 U194 ( .A(sfr_wdat[4]), .Y(n133) );
  INVX1 U195 ( .A(sfr_wdat[2]), .Y(n121) );
  INVX1 U196 ( .A(sfr_wdat[6]), .Y(n144) );
  INVX1 U197 ( .A(n168), .Y(n205) );
  INVX1 U198 ( .A(sfr_wdat[5]), .Y(n138) );
  INVX1 U199 ( .A(sfr_wdat[1]), .Y(n116) );
  INVX1 U200 ( .A(sfr_wdat[7]), .Y(n150) );
  INVX1 U201 ( .A(n104), .Y(n102) );
  INVX1 U202 ( .A(n104), .Y(n103) );
  INVX1 U203 ( .A(n101), .Y(n29) );
  INVX1 U204 ( .A(n101), .Y(n30) );
  INVX1 U205 ( .A(n98), .Y(n31) );
  INVX1 U206 ( .A(n98), .Y(n32) );
  INVX1 U207 ( .A(n98), .Y(n33) );
  INVX1 U208 ( .A(n101), .Y(n34) );
  INVX1 U209 ( .A(n91), .Y(n35) );
  INVX1 U210 ( .A(n92), .Y(n36) );
  INVX1 U211 ( .A(n99), .Y(n97) );
  INVX1 U212 ( .A(n243), .Y(n89) );
  INVX1 U213 ( .A(n99), .Y(n91) );
  INVX1 U214 ( .A(n243), .Y(n96) );
  INVX1 U215 ( .A(n99), .Y(n95) );
  INVX1 U216 ( .A(n243), .Y(n94) );
  INVX1 U217 ( .A(n99), .Y(n92) );
  INVX1 U218 ( .A(n243), .Y(n93) );
  INVX1 U219 ( .A(n99), .Y(n90) );
  INVX1 U220 ( .A(n243), .Y(n88) );
  NAND43X1 U221 ( .B(n173), .C(n179), .D(n175), .A(n178), .Y(n239) );
  INVX1 U222 ( .A(n184), .Y(n185) );
  INVX1 U223 ( .A(n153), .Y(n204) );
  INVX1 U224 ( .A(n183), .Y(n200) );
  AND2X1 U225 ( .A(n203), .B(n207), .Y(r_dacwr[0]) );
  INVX1 U226 ( .A(n156), .Y(n213) );
  INVX1 U227 ( .A(n167), .Y(n210) );
  INVX1 U228 ( .A(n158), .Y(n217) );
  INVX1 U229 ( .A(n162), .Y(n212) );
  INVX1 U230 ( .A(n176), .Y(n206) );
  INVX1 U231 ( .A(n166), .Y(n238) );
  NAND21X1 U232 ( .B(n178), .A(n165), .Y(n166) );
  AND2X1 U233 ( .A(n211), .B(n213), .Y(r_fcpwr[3]) );
  INVX1 U234 ( .A(n231), .Y(n221) );
  INVX1 U235 ( .A(prl_c0set), .Y(n254) );
  AND2X1 U236 ( .A(n211), .B(n232), .Y(r_fcpwr[1]) );
  INVX1 U237 ( .A(n229), .Y(hit[178]) );
  INVX1 U238 ( .A(n1148), .Y(n249) );
  AND2X1 U239 ( .A(n217), .B(n228), .Y(r_fcpwr[4]) );
  AND2X1 U240 ( .A(n212), .B(n211), .Y(r_fcpwr[5]) );
  INVX1 U241 ( .A(n1134), .Y(n251) );
  NOR2X1 U242 ( .A(n137), .B(n1187), .Y(clrAE[5]) );
  NOR2X1 U243 ( .A(n116), .B(n1187), .Y(clrAE[1]) );
  NOR2X1 U244 ( .A(n137), .B(n1186), .Y(clrDF[5]) );
  NOR2X1 U245 ( .A(n115), .B(n1186), .Y(clrDF[1]) );
  NOR2X1 U246 ( .A(n137), .B(n1190), .Y(clr03[5]) );
  NOR2X1 U247 ( .A(n116), .B(n1190), .Y(clr03[1]) );
  NOR2X1 U248 ( .A(n133), .B(n1187), .Y(clrAE[4]) );
  NOR2X1 U249 ( .A(n111), .B(n1187), .Y(clrAE[0]) );
  NOR2X1 U250 ( .A(n133), .B(n1186), .Y(clrDF[4]) );
  NOR2X1 U251 ( .A(n111), .B(n1186), .Y(clrDF[0]) );
  NOR2X1 U252 ( .A(n133), .B(n1190), .Y(clr03[4]) );
  NOR2X1 U253 ( .A(n111), .B(n1190), .Y(clr03[0]) );
  NOR2X1 U254 ( .A(n144), .B(n1187), .Y(clrAE[6]) );
  NOR2X1 U255 ( .A(n121), .B(n1187), .Y(clrAE[2]) );
  NOR2X1 U256 ( .A(n144), .B(n1186), .Y(clrDF[6]) );
  NOR2X1 U257 ( .A(n120), .B(n1186), .Y(clrDF[2]) );
  NOR2X1 U258 ( .A(n144), .B(n1190), .Y(clr03[6]) );
  NOR2X1 U259 ( .A(n121), .B(n1190), .Y(clr03[2]) );
  NOR2X1 U260 ( .A(n150), .B(n1187), .Y(clrAE[7]) );
  NOR2X1 U261 ( .A(n126), .B(n1187), .Y(clrAE[3]) );
  NOR2X1 U262 ( .A(n149), .B(n1186), .Y(clrDF[7]) );
  NOR2X1 U263 ( .A(n126), .B(n1186), .Y(clrDF[3]) );
  NOR2X1 U264 ( .A(n150), .B(n1190), .Y(clr03[7]) );
  NOR2X1 U265 ( .A(n126), .B(n1190), .Y(clr03[3]) );
  NAND21X1 U266 ( .B(n1129), .A(n104), .Y(n1128) );
  INVX1 U267 ( .A(n187), .Y(r_set_cpmsgid) );
  INVX1 U268 ( .A(n198), .Y(n242) );
  AND2XL U269 ( .A(n228), .B(n230), .Y(r_dacwr[14]) );
  AND2X1 U270 ( .A(n228), .B(n232), .Y(we_148) );
  AND2X1 U271 ( .A(n211), .B(n217), .Y(r_fcpwr[2]) );
  AND2X1 U272 ( .A(n211), .B(n210), .Y(r_fcpwr[0]) );
  AND2XL U273 ( .A(n225), .B(n230), .Y(we_217) );
  AND2X1 U274 ( .A(n213), .B(n228), .Y(r_fcpwr[6]) );
  AND2X1 U275 ( .A(n213), .B(n225), .Y(we_222) );
  AND2X1 U276 ( .A(n218), .B(n232), .Y(r_cvcwr[0]) );
  AND2X1 U277 ( .A(n218), .B(n217), .Y(r_cvcwr[1]) );
  INVX1 U278 ( .A(n1124), .Y(n1096) );
  INVX1 U279 ( .A(n270), .Y(n208) );
  NOR32XL U280 ( .B(n207), .C(n163), .A(n201), .Y(we_232) );
  AND2X1 U281 ( .A(n207), .B(n228), .Y(r_dacwr[13]) );
  AND2X1 U282 ( .A(n207), .B(n221), .Y(we_176) );
  INVX1 U283 ( .A(n222), .Y(n226) );
  INVX1 U284 ( .A(n234), .Y(n163) );
  INVX1 U285 ( .A(n236), .Y(n241) );
  INVX1 U286 ( .A(n169), .Y(n223) );
  INVX1 U287 ( .A(n170), .Y(n180) );
  INVX1 U288 ( .A(n233), .Y(n188) );
  INVX1 U289 ( .A(ictlr_inc), .Y(n104) );
  INVX1 U290 ( .A(n88), .Y(n99) );
  INVX1 U291 ( .A(n99), .Y(n98) );
  NAND43XL U292 ( .B(n179), .C(n178), .D(n177), .A(sfr_w), .Y(n186) );
  INVX1 U293 ( .A(n177), .Y(n173) );
  INVX1 U294 ( .A(n171), .Y(n178) );
  INVX1 U295 ( .A(n172), .Y(n179) );
  INVX1 U296 ( .A(n214), .Y(n235) );
  INVX1 U297 ( .A(n159), .Y(n207) );
  NAND43XL U298 ( .B(n173), .C(n178), .D(n179), .A(sfr_w), .Y(n159) );
  INVX1 U299 ( .A(n161), .Y(n227) );
  NAND21X1 U300 ( .B(n171), .A(n165), .Y(n161) );
  INVX1 U301 ( .A(n160), .Y(n165) );
  NAND21X1 U302 ( .B(n177), .A(n179), .Y(n160) );
  INVX1 U303 ( .A(n157), .Y(n240) );
  NAND32X1 U304 ( .B(n177), .C(n171), .A(n172), .Y(n157) );
  OAI31XL U305 ( .A(n1147), .B(n1148), .C(n1149), .D(n254), .Y(r_fiforst) );
  NAND2X1 U306 ( .A(n110), .B(n120), .Y(n1149) );
  NAND4X1 U307 ( .A(n126), .B(n132), .C(n143), .D(n149), .Y(n1147) );
  NAND4XL U308 ( .A(hit[183]), .B(sfr_w), .C(n115), .D(n137), .Y(n1148) );
  AND2X1 U309 ( .A(n227), .B(n221), .Y(hit[183]) );
  INVX1 U310 ( .A(n174), .Y(n237) );
  NAND32X1 U311 ( .B(n173), .C(n172), .A(n171), .Y(n174) );
  INVX1 U312 ( .A(n155), .Y(n224) );
  NAND32X1 U313 ( .B(n171), .C(n172), .A(n177), .Y(n155) );
  AND2XL U314 ( .A(hit[178]), .B(sfr_w), .Y(r_fifopsh) );
  AND2X1 U315 ( .A(sfr_r), .B(hit[178]), .Y(r_fifopop) );
  INVX1 U316 ( .A(n1153), .Y(n248) );
  NAND2XL U317 ( .A(hit[174]), .B(sfr_w), .Y(n1187) );
  AND2X1 U318 ( .A(n224), .B(n223), .Y(hit[174]) );
  NAND2XL U319 ( .A(hit_223), .B(sfr_w), .Y(n1186) );
  AND2X1 U320 ( .A(n225), .B(n227), .Y(hit_223) );
  NAND2XL U321 ( .A(hit[179]), .B(sfr_w), .Y(n1190) );
  AND2X1 U322 ( .A(n238), .B(n221), .Y(hit[179]) );
  NAND21X1 U323 ( .B(n19), .A(n220), .Y(N108) );
  NOR2X1 U324 ( .A(n1130), .B(n264), .Y(n1134) );
  NAND4X1 U325 ( .A(n1129), .B(n248), .C(n1142), .D(n104), .Y(upd19) );
  OA21X1 U326 ( .B(prx_rst[0]), .C(prx_rst[1]), .A(set03[1]), .Y(set03[7]) );
  NAND2XL U327 ( .A(hit_197), .B(n4), .Y(n1126) );
  AND2X1 U328 ( .A(n241), .B(n240), .Y(hit_197) );
  NAND2XL U329 ( .A(hit_202), .B(sfr_w), .Y(n1124) );
  AND2X1 U330 ( .A(n226), .B(n237), .Y(hit_202) );
  AND2X1 U331 ( .A(hit_151), .B(sfr_r), .Y(r_fcpre) );
  AND2X1 U332 ( .A(n228), .B(n227), .Y(hit_151) );
  INVX1 U333 ( .A(n189), .Y(n215) );
  NAND2XL U334 ( .A(hit_195), .B(n4), .Y(n1129) );
  AND2X1 U335 ( .A(n238), .B(n241), .Y(hit_195) );
  INVX1 U336 ( .A(n209), .Y(n211) );
  OAI21BBXL U337 ( .A(hit_194), .B(n4), .C(n104), .Y(upd18) );
  AND2X1 U338 ( .A(n237), .B(n241), .Y(hit_194) );
  INVX1 U339 ( .A(n181), .Y(n228) );
  INVX1 U340 ( .A(n182), .Y(n225) );
  INVX1 U341 ( .A(n1141), .Y(n1121) );
  INVX1 U342 ( .A(n216), .Y(n218) );
  INVX1 U343 ( .A(N34), .Y(n265) );
  AND2X1 U344 ( .A(dnchk_en), .B(dm_fault), .Y(dmf_wkup) );
  INVX1 U345 ( .A(n243), .Y(n100) );
  INVX1 U346 ( .A(n243), .Y(n101) );
  BUFX3 U347 ( .A(pff_full), .Y(dbgpo[22]) );
  BUFX3 U348 ( .A(pff_empty), .Y(dbgpo[23]) );
  NAND21XL U349 ( .B(n154), .A(sfr_addr[0]), .Y(n177) );
  NAND21XL U350 ( .B(n154), .A(sfr_addr[4]), .Y(n189) );
  NAND21XL U351 ( .B(n154), .A(sfr_addr[2]), .Y(n171) );
  NAND21XL U352 ( .B(n154), .A(sfr_addr[1]), .Y(n172) );
  NAND21XL U353 ( .B(n154), .A(sfr_addr[3]), .Y(n214) );
  INVX1 U354 ( .A(n20), .Y(srstz) );
  NOR2X1 U355 ( .A(n269), .B(n253), .Y(r_osc_stop) );
  NOR2X1 U356 ( .A(n269), .B(n252), .Y(r_osc_lo) );
  INVX1 U357 ( .A(n1185), .Y(bus_idle) );
  AND2X1 U358 ( .A(pff_ack[1]), .B(n244), .Y(set04[5]) );
  NOR42XL U359 ( .C(n133), .D(n1179), .A(n119), .B(n1150), .Y(n1153) );
  NAND3X1 U360 ( .A(n254), .B(n268), .C(n248), .Y(phyrst) );
  INVX1 U361 ( .A(n195), .Y(n220) );
  NOR2X1 U362 ( .A(n269), .B(n196), .Y(r_pos_gate) );
  AND2X1 U363 ( .A(n193), .B(n220), .Y(n19) );
  NAND3X1 U364 ( .A(n1138), .B(n14), .C(n1135), .Y(upd01) );
  NAND42X1 U365 ( .C(set_hold), .D(cpurst), .A(n1133), .B(n1130), .Y(upd12) );
  AND2X1 U366 ( .A(prx_setsta[1]), .B(n244), .Y(set03[1]) );
  OAI22AX1 U367 ( .D(sfr_wdat[7]), .C(n1128), .A(n104), .B(n199), .Y(wd19[7])
         );
  NAND4X1 U368 ( .A(n249), .B(n1179), .C(n1207), .D(n1208), .Y(n1142) );
  NOR2X1 U369 ( .A(n121), .B(n110), .Y(n1207) );
  NOR4XL U370 ( .A(n145), .B(n122), .C(n143), .D(n132), .Y(n1208) );
  ENOX1 U371 ( .A(n1126), .B(n115), .C(pff_rxpart[9]), .D(n1126), .Y(wd21[1])
         );
  ENOX1 U372 ( .A(n16), .B(n121), .C(pff_rxpart[10]), .D(n1126), .Y(wd21[2])
         );
  ENOX1 U373 ( .A(n16), .B(n127), .C(pff_rxpart[11]), .D(n1126), .Y(wd21[3])
         );
  ENOX1 U374 ( .A(n16), .B(n132), .C(pff_rxpart[12]), .D(n1126), .Y(wd21[4])
         );
  ENOX1 U375 ( .A(n16), .B(n138), .C(pff_rxpart[13]), .D(n1126), .Y(wd21[5])
         );
  ENOX1 U376 ( .A(n16), .B(n144), .C(pff_rxpart[14]), .D(n1126), .Y(wd21[6])
         );
  ENOX1 U377 ( .A(n16), .B(n150), .C(pff_rxpart[15]), .D(n1126), .Y(wd21[7])
         );
  ENOX1 U378 ( .A(n110), .B(n1128), .C(inst_ofs_plus[8]), .D(n103), .Y(wd19[0]) );
  ENOX1 U379 ( .A(n116), .B(n1128), .C(inst_ofs_plus[9]), .D(n103), .Y(wd19[1]) );
  ENOX1 U380 ( .A(n120), .B(n1128), .C(inst_ofs_plus[10]), .D(n103), .Y(
        wd19[2]) );
  ENOX1 U381 ( .A(n127), .B(n1128), .C(inst_ofs_plus[11]), .D(n103), .Y(
        wd19[3]) );
  ENOX1 U382 ( .A(n132), .B(n1128), .C(inst_ofs_plus[12]), .D(n102), .Y(
        wd19[4]) );
  ENOX1 U383 ( .A(n138), .B(n1128), .C(inst_ofs_plus[13]), .D(n103), .Y(
        wd19[5]) );
  ENOX1 U384 ( .A(n110), .B(n1127), .C(pff_rxpart[0]), .D(n1127), .Y(wd20[0])
         );
  ENOX1 U385 ( .A(n116), .B(n12), .C(pff_rxpart[1]), .D(n1127), .Y(wd20[1]) );
  ENOX1 U386 ( .A(n120), .B(n12), .C(pff_rxpart[2]), .D(n1127), .Y(wd20[2]) );
  ENOX1 U387 ( .A(n127), .B(n12), .C(pff_rxpart[3]), .D(n1127), .Y(wd20[3]) );
  ENOX1 U388 ( .A(n132), .B(n12), .C(pff_rxpart[4]), .D(n1127), .Y(wd20[4]) );
  NAND2X1 U389 ( .A(n1140), .B(n12), .Y(upd20) );
  NAND2X1 U390 ( .A(n1140), .B(n16), .Y(upd21) );
  AND2X1 U391 ( .A(prx_setsta[2]), .B(n15), .Y(set03[2]) );
  AND4X1 U392 ( .A(sfr_r), .B(n226), .C(n224), .D(n199), .Y(upd31) );
  AND2X1 U393 ( .A(pff_obsd), .B(n244), .Y(set04[3]) );
  AND2X1 U394 ( .A(prx_setsta[4]), .B(n15), .Y(set03[4]) );
  NAND2X1 U395 ( .A(prx_setsta[3]), .B(n244), .Y(n1141) );
  ENOX1 U396 ( .A(n102), .B(n116), .C(inst_ofs_plus[1]), .D(ictlr_inc), .Y(
        wd18[1]) );
  ENOX1 U397 ( .A(n102), .B(n121), .C(inst_ofs_plus[2]), .D(ictlr_inc), .Y(
        wd18[2]) );
  ENOX1 U398 ( .A(n102), .B(n132), .C(inst_ofs_plus[4]), .D(n103), .Y(wd18[4])
         );
  ENOX1 U399 ( .A(n102), .B(n127), .C(inst_ofs_plus[3]), .D(ictlr_inc), .Y(
        wd18[3]) );
  ENOX1 U400 ( .A(n102), .B(n138), .C(inst_ofs_plus[5]), .D(n103), .Y(wd18[5])
         );
  ENOX1 U401 ( .A(n102), .B(n143), .C(inst_ofs_plus[6]), .D(n103), .Y(wd18[6])
         );
  ENOX1 U402 ( .A(n102), .B(n150), .C(inst_ofs_plus[7]), .D(n103), .Y(wd18[7])
         );
  AND2X1 U403 ( .A(i_gobusy), .B(n15), .Y(set04[2]) );
  AND2X1 U404 ( .A(i_goidle), .B(n244), .Y(set04[1]) );
  AND2X1 U405 ( .A(prl_GCTxDone), .B(n15), .Y(set04[6]) );
  XNOR2XL U406 ( .A(n265), .B(N33), .Y(N37) );
  XNOR2XL U407 ( .A(N35), .B(n265), .Y(N36) );
  XOR2X1 U408 ( .A(N33), .B(N32), .Y(N38) );
  AND2X1 U409 ( .A(prl_discard), .B(n244), .Y(set04[7]) );
  XNOR2XL U410 ( .A(N30), .B(N32), .Y(N39) );
  INVX1 U411 ( .A(n1133), .Y(n264) );
  NAND3X1 U412 ( .A(n252), .B(n196), .C(n253), .Y(N84) );
  XNOR2XL U413 ( .A(di_p0[4]), .B(n258), .Y(n1201) );
  XNOR2XL U414 ( .A(di_p0[6]), .B(n256), .Y(n1203) );
  XNOR2XL U415 ( .A(di_p0[2]), .B(n260), .Y(n1199) );
  XNOR2XL U416 ( .A(di_p0[5]), .B(n257), .Y(n1202) );
  XNOR2XL U417 ( .A(di_p0[7]), .B(n255), .Y(n1204) );
  XNOR2XL U418 ( .A(di_p0[3]), .B(n259), .Y(n1200) );
  NAND2X1 U419 ( .A(n152), .B(aswkup), .Y(pwrdn_rstz) );
  INVX1 U420 ( .A(n1222), .Y(n243) );
  MUX2XL U421 ( .D0(i_pc[1]), .D1(prx_adpn[1]), .S(reg19_7_), .Y(reg30[1]) );
  MUX2XL U422 ( .D0(i_pc[0]), .D1(prx_adpn[0]), .S(reg19_7_), .Y(reg30[0]) );
  MUX2X1 U423 ( .D0(s_ovp), .D1(m_ovp), .S(reg94[4]), .Y(regAD[2]) );
  AND3X1 U424 ( .A(n18), .B(n122), .C(n219), .Y(ps_pwrdn) );
  INVX1 U425 ( .A(n1151), .Y(n219) );
  OR2X1 U426 ( .A(lg_dischg), .B(lg_pulse_12m), .Y(r_srcctl[1]) );
  MUX2XL U427 ( .D0(i_pc[2]), .D1(prx_adpn[2]), .S(reg19_7_), .Y(reg30[2]) );
  NAND42X1 U428 ( .C(bkpt_hold), .D(reg12[3]), .A(n253), .B(n196), .Y(
        r_hold_mcu) );
  NAND3X1 U429 ( .A(n1181), .B(n1182), .C(n1183), .Y(i2c_stretch) );
  AOI22X1 U430 ( .A(reg28[2]), .B(reg27[2]), .C(reg28[3]), .D(reg27[3]), .Y(
        n1181) );
  AOI22X1 U431 ( .A(reg28[0]), .B(reg27[0]), .C(reg28[1]), .D(reg27[1]), .Y(
        n1182) );
  AOI222XL U432 ( .A(reg28[7]), .B(reg27[7]), .C(reg28[4]), .D(reg27[4]), .E(
        reg28[6]), .F(reg27[6]), .Y(n1183) );
  OAI211X1 U433 ( .C(rstcnt[2]), .D(rstcnt[1]), .A(n267), .B(rstcnt[4]), .Y(
        n1192) );
  INVX1 U434 ( .A(regD4[0]), .Y(n253) );
  AOI21X1 U435 ( .B(drstz[1]), .C(n1192), .A(atpg_en), .Y(n20) );
  INVX1 U436 ( .A(rstcnt[3]), .Y(n267) );
  INVX1 U437 ( .A(oscdwn_shft[2]), .Y(n269) );
  INVX1 U438 ( .A(regD4[1]), .Y(n252) );
  NOR4XL U439 ( .A(prl_fsm[3]), .B(prl_fsm[2]), .C(prl_fsm[1]), .D(prl_fsm[0]), 
        .Y(n1211) );
  OAI211X1 U440 ( .C(ictlr_idle), .D(n197), .A(oscdwn_shft[1]), .B(bus_idle), 
        .Y(n1151) );
  AND3X1 U441 ( .A(regD4[1]), .B(n253), .C(n196), .Y(n197) );
  INVX1 U442 ( .A(regD4[2]), .Y(n196) );
  MUX2X1 U443 ( .D0(s_scp), .D1(m_scp), .S(reg94[5]), .Y(regAD[4]) );
  NAND4X1 U444 ( .A(n1166), .B(n1167), .C(n1168), .D(n1169), .Y(o_intr[1]) );
  AOI22X1 U445 ( .A(reg06[6]), .B(irq04[6]), .C(reg06[7]), .D(irq04[7]), .Y(
        n1166) );
  AOI22X1 U446 ( .A(reg06[0]), .B(irq04[0]), .C(reg06[1]), .D(irq04[1]), .Y(
        n1169) );
  AOI22X1 U447 ( .A(reg06[4]), .B(irq04[4]), .C(reg06[5]), .D(irq04[5]), .Y(
        n1167) );
  AND3XL U448 ( .A(n11), .B(sfr_w), .C(n242), .Y(r_pswr) );
  NAND21X1 U449 ( .B(lg_pulse_12m), .A(n194), .Y(n195) );
  OR4X1 U450 ( .A(osc_gate_n[1]), .B(osc_gate_n[0]), .C(osc_gate_n[3]), .D(
        osc_gate_n[2]), .Y(r_osc_gate) );
  NAND31X1 U451 ( .C(n1213), .A(lg_pulse_len[1]), .B(lg_pulse_len[0]), .Y(
        n1212) );
  AND3X1 U452 ( .A(n242), .B(sfr_r), .C(n11), .Y(r_psrd) );
  OAI21AX1 U453 ( .B(lg_pulse_len[0]), .C(lg_pulse_len[1]), .A(n220), .Y(n1213) );
  OAI32X1 U454 ( .A(n1177), .B(i_goidle), .C(n15), .D(r_phyrst[0]), .E(n1178), 
        .Y(n1221) );
  AOI211X1 U455 ( .C(reg11_7_), .D(set03[7]), .A(r_phyrst[1]), .B(n1153), .Y(
        n1178) );
  OAI211X1 U456 ( .C(lg_pulse_len[0]), .D(n1213), .A(n1212), .B(n1214), .Y(
        N112) );
  NAND2X1 U457 ( .A(N105), .B(n19), .Y(n1214) );
  NOR21XL U458 ( .B(regE3_0), .A(gating_pwr), .Y(r_srcctl[0]) );
  AO22X1 U459 ( .A(regAF[4]), .B(regAE[4]), .C(regAF[2]), .D(regAE[2]), .Y(
        gating_pwr) );
  NOR21XL U460 ( .B(n1135), .A(n1136), .Y(wd01[7]) );
  AOI22X1 U461 ( .A(r_last), .B(n1137), .C(n250), .D(n148), .Y(n1136) );
  NOR21XL U462 ( .B(n1138), .A(n1139), .Y(wd01[6]) );
  AOI22X1 U463 ( .A(r_first), .B(n1137), .C(n250), .D(n142), .Y(n1139) );
  AND2X1 U464 ( .A(regE3[3]), .B(n1144), .Y(r_srcctl[3]) );
  AO21X1 U465 ( .B(N103), .C(n19), .A(n195), .Y(N110) );
  AO21X1 U466 ( .B(lg_dischg), .C(n193), .A(n195), .Y(n1219) );
  AO21X1 U467 ( .B(n19), .C(n192), .A(n195), .Y(N109) );
  INVX1 U468 ( .A(lg_pulse_cnt[0]), .Y(n192) );
  OAI21BX1 U469 ( .C(lg_pulse_12m), .B(lg_dischg), .A(n194), .Y(n1218) );
  OAI21X1 U470 ( .B(r_fifopop), .C(r_fifopsh), .A(r_first), .Y(n1138) );
  AOI22X1 U471 ( .A(regAF[5]), .B(regAE[5]), .C(regAD[5]), .D(i_vcbyval), .Y(
        n1144) );
  OAI21X1 U472 ( .B(n132), .C(n1130), .A(n1131), .Y(wd12[4]) );
  AOI21X1 U473 ( .B(reg12[4]), .C(n1130), .A(n264), .Y(n1131) );
  ENOXL U474 ( .A(n110), .B(n251), .C(r_pshords), .D(n251), .Y(wd12[0]) );
  ENOX1 U475 ( .A(n116), .B(n251), .C(reg12_1), .D(n251), .Y(wd12[1]) );
  AO22AXL U476 ( .A(r_txshrt), .B(n251), .C(sfr_wdat[2]), .D(n251), .Y(wd12[2]) );
  ENOX1 U477 ( .A(n138), .B(n251), .C(reg12[5]), .D(n251), .Y(wd12[5]) );
  ENOX1 U478 ( .A(n144), .B(n13), .C(reg12[6]), .D(n251), .Y(wd12[6]) );
  ENOX1 U479 ( .A(n149), .B(n13), .C(reg12[7]), .D(n251), .Y(wd12[7]) );
  OAI21BBX1 U480 ( .A(N106), .B(n19), .C(n1212), .Y(N113) );
  OAI21BBX1 U481 ( .A(n264), .B(reg12[3]), .C(n1132), .Y(wd12[3]) );
  AOI32X1 U482 ( .A(n1133), .B(n1130), .C(set_hold), .D(n1134), .E(n122), .Y(
        n1132) );
  OAI21BBX1 U483 ( .A(N104), .B(n19), .C(n1213), .Y(N111) );
  AND2X1 U484 ( .A(regE3[2]), .B(n1144), .Y(r_srcctl[2]) );
  AOI21X1 U485 ( .B(n1184), .C(n1124), .A(n1185), .Y(i2c_mode_upd) );
  ENOX1 U486 ( .A(n111), .B(n1124), .C(n1124), .D(lt_reg26_0), .Y(
        i2c_mode_wdat) );
  XNOR2XL U487 ( .A(r_hwi2c_en), .B(lt_reg26_0), .Y(n1184) );
  NOR21XL U488 ( .B(regD4[4]), .A(n269), .Y(r_ocdrv_enz) );
  NAND4X1 U489 ( .A(n1170), .B(n1171), .C(n1172), .D(n1173), .Y(o_intr[0]) );
  AOI22X1 U490 ( .A(reg05[4]), .B(irq03[4]), .C(reg05[5]), .D(irq03[5]), .Y(
        n1171) );
  AOI22X1 U491 ( .A(reg05[2]), .B(irq03[2]), .C(reg05[3]), .D(irq03[3]), .Y(
        n1172) );
  NOR21XL U492 ( .B(regD4[3]), .A(n269), .Y(r_pwrdn) );
  AND2X1 U493 ( .A(reg94[7]), .B(reg94[6]), .Y(r_otpi_gate) );
  AOI22X1 U494 ( .A(reg05[6]), .B(irq03[6]), .C(reg05[7]), .D(irq03[7]), .Y(
        n1170) );
  OAI21X1 U495 ( .B(n1206), .C(n1185), .A(n1142), .Y(N26) );
  NOR21XL U496 ( .B(n1143), .A(rstcnt[4]), .Y(n1206) );
  ENOXL U497 ( .A(n111), .B(n1137), .C(r_txnumk[0]), .D(n1137), .Y(wd01[0]) );
  ENOXL U498 ( .A(n116), .B(n14), .C(r_txnumk[1]), .D(n1137), .Y(wd01[1]) );
  ENOXL U499 ( .A(n121), .B(n14), .C(r_txnumk[2]), .D(n1137), .Y(wd01[2]) );
  ENOXL U500 ( .A(n126), .B(n14), .C(r_txnumk[3]), .D(n1137), .Y(wd01[3]) );
  ENOXL U501 ( .A(n132), .B(n14), .C(r_txnumk[4]), .D(n1137), .Y(wd01[4]) );
  ENOX1 U502 ( .A(n138), .B(n14), .C(r_unlock), .D(n1137), .Y(wd01[5]) );
  ENOX1 U503 ( .A(n16), .B(n110), .C(pff_rxpart[8]), .D(n1126), .Y(wd21[0]) );
  ENOX1 U504 ( .A(n144), .B(n1128), .C(inst_ofs_plus[14]), .D(n103), .Y(
        wd19[6]) );
  ENOX1 U505 ( .A(n138), .B(n12), .C(pff_rxpart[5]), .D(n1127), .Y(wd20[5]) );
  ENOX1 U506 ( .A(n143), .B(n12), .C(pff_rxpart[6]), .D(n1127), .Y(wd20[6]) );
  ENOX1 U507 ( .A(n149), .B(n12), .C(pff_rxpart[7]), .D(n1127), .Y(wd20[7]) );
  NAND2X1 U508 ( .A(r_last), .B(r_fifopsh), .Y(n1135) );
  MUX2XL U509 ( .D0(i_pc[3]), .D1(prx_adpn[3]), .S(reg19_7_), .Y(reg30[3]) );
  AOI22X1 U510 ( .A(reg05[0]), .B(irq03[0]), .C(reg05[1]), .D(irq03[1]), .Y(
        n1173) );
  AOI22X1 U511 ( .A(reg06[2]), .B(irq04[2]), .C(reg06[3]), .D(irq04[3]), .Y(
        n1168) );
  MUX2XL U512 ( .D0(i_pc[4]), .D1(prx_adpn[4]), .S(reg19_7_), .Y(reg30[4]) );
  NOR21XL U513 ( .B(prx_setsta[6]), .A(prl_cany0), .Y(set03[6]) );
  MUX2X1 U514 ( .D0(i_pc[5]), .D1(prx_adpn[5]), .S(reg19_7_), .Y(reg30[5]) );
  AO21X1 U515 ( .B(n1145), .C(n1146), .A(reg11_4), .Y(r_rxords_ena[4]) );
  NOR3XL U516 ( .A(r_rxords_ena[0]), .B(r_rxords_ena[2]), .C(r_rxords_ena[1]), 
        .Y(n1145) );
  NOR3XL U517 ( .A(r_rxords_ena[3]), .B(r_rxords_ena[6]), .C(r_rxords_ena[5]), 
        .Y(n1146) );
  ENOX1 U518 ( .A(n102), .B(n110), .C(inst_ofs_plus[0]), .D(n102), .Y(wd18[0])
         );
  AOI21BBXL U519 ( .B(r_auto_gdcrc[1]), .C(n1141), .A(set03[6]), .Y(n1140) );
  AND2X1 U520 ( .A(i_pc[6]), .B(n199), .Y(reg30[6]) );
  AND2X1 U521 ( .A(i_pc[7]), .B(n199), .Y(reg30[7]) );
  INVX1 U522 ( .A(reg19_7_), .Y(n199) );
  OAI31XL U523 ( .A(n263), .B(r_phyrst[1]), .C(n266), .D(n152), .Y(prstz) );
  INVX1 U524 ( .A(drstz[1]), .Y(n263) );
  INVX1 U525 ( .A(n1192), .Y(n266) );
  NAND4X1 U526 ( .A(n1162), .B(n1163), .C(n1164), .D(n1165), .Y(o_intr[2]) );
  AOI22X1 U527 ( .A(reg27[4]), .B(irq28[4]), .C(reg27[5]), .D(irq28[5]), .Y(
        n1163) );
  AOI22X1 U528 ( .A(reg27[0]), .B(irq28[0]), .C(reg27[1]), .D(irq28[1]), .Y(
        n1165) );
  AOI22X1 U529 ( .A(reg27[6]), .B(irq28[6]), .C(reg27[7]), .D(irq28[7]), .Y(
        n1162) );
  AND2X1 U530 ( .A(prx_setsta[5]), .B(n244), .Y(set03[5]) );
  AND2X1 U531 ( .A(ptx_ack), .B(n244), .Y(set04[0]) );
  AOI22X1 U532 ( .A(reg27[2]), .B(irq28[2]), .C(reg27[3]), .D(irq28[3]), .Y(
        n1164) );
  MUX2X1 U533 ( .D0(s_ovp_sta), .D1(m_ovp_sta), .S(reg94[4]), .Y(setAE[2]) );
  MUX2X1 U534 ( .D0(s_scp_sta), .D1(m_scp_sta), .S(reg94[5]), .Y(setAE[4]) );
  XNOR2XL U535 ( .A(d_p0[0]), .B(n262), .Y(setDF[0]) );
  XNOR2XL U536 ( .A(d_p0[1]), .B(n261), .Y(setDF[1]) );
  XNOR2XL U537 ( .A(d_p0[2]), .B(n260), .Y(setDF[2]) );
  XNOR2XL U538 ( .A(d_p0[3]), .B(n259), .Y(setDF[3]) );
  XNOR2XL U539 ( .A(d_p0[4]), .B(n258), .Y(setDF[4]) );
  INVX1 U540 ( .A(prl_cany0), .Y(n244) );
  XNOR2XL U541 ( .A(rstcnt[4]), .B(n267), .Y(N27) );
  XNOR2XL U542 ( .A(n1205), .B(N27), .Y(N29) );
  XNOR2XL U543 ( .A(rstcnt[2]), .B(rstcnt[1]), .Y(n1205) );
  AND2X1 U544 ( .A(prx_setsta[0]), .B(n244), .Y(set03[0]) );
  XOR2X1 U545 ( .A(N29), .B(rstcnt[0]), .Y(N30) );
  XOR2X1 U546 ( .A(rstcnt[2]), .B(N27), .Y(N28) );
  NOR42XL U547 ( .C(n1209), .D(r_inst_ofs[10]), .A(r_inst_ofs[8]), .B(n1210), 
        .Y(n1179) );
  NAND4X1 U548 ( .A(r_inst_ofs[14]), .B(r_inst_ofs[13]), .C(r_inst_ofs[12]), 
        .D(r_inst_ofs[11]), .Y(n1210) );
  NOR2X1 U549 ( .A(n11), .B(r_inst_ofs[9]), .Y(n1209) );
  NAND4X1 U550 ( .A(n1158), .B(n1159), .C(n1160), .D(n1161), .Y(o_intr[3]) );
  AOI22X1 U551 ( .A(regDE[6]), .B(irqDF[6]), .C(regDE[7]), .D(irqDF[7]), .Y(
        n1158) );
  AOI22X1 U552 ( .A(regDE[4]), .B(irqDF[4]), .C(regDE[5]), .D(irqDF[5]), .Y(
        n1159) );
  INVX1 U553 ( .A(reg25_0_), .Y(r_i2c_ninc) );
  NAND4X1 U554 ( .A(n1154), .B(n1155), .C(n1156), .D(n1157), .Y(o_intr[4]) );
  AOI22X1 U555 ( .A(regAF[6]), .B(irqAE[6]), .C(regAF[7]), .D(irqAE[7]), .Y(
        n1154) );
  AOI22X1 U556 ( .A(regAF[0]), .B(irqAE[0]), .C(regAF[1]), .D(irqAE[1]), .Y(
        n1157) );
  AOI22X1 U557 ( .A(regDE[0]), .B(irqDF[0]), .C(regDE[1]), .D(irqDF[1]), .Y(
        n1161) );
  AOI22X1 U558 ( .A(regDE[2]), .B(irqDF[2]), .C(regDE[3]), .D(irqDF[3]), .Y(
        n1160) );
  AOI22X1 U559 ( .A(irqAE[2]), .B(regAF[2]), .C(regAF[3]), .D(irqAE[3]), .Y(
        n1156) );
  AOI22X1 U560 ( .A(irqAE[4]), .B(regAF[4]), .C(irqAE[5]), .D(regAF[5]), .Y(
        n1155) );
  XNOR2XL U561 ( .A(d_p0[6]), .B(n256), .Y(setDF[6]) );
  XNOR2XL U562 ( .A(d_p0[7]), .B(n255), .Y(setDF[7]) );
  XNOR2XL U563 ( .A(d_p0[5]), .B(n257), .Y(setDF[5]) );
  OAI22X1 U564 ( .A(r_phyrst[0]), .B(n268), .C(n1176), .D(n1177), .Y(n1220) );
  NOR2X1 U565 ( .A(i_goidle), .B(n15), .Y(n1176) );
  INVX1 U566 ( .A(ff_p0[5]), .Y(n257) );
  INVX1 U567 ( .A(ff_p0[7]), .Y(n255) );
  INVX1 U568 ( .A(ff_p0[1]), .Y(n261) );
  INVX1 U569 ( .A(ff_p0[2]), .Y(n260) );
  INVX1 U570 ( .A(ff_p0[3]), .Y(n259) );
  INVX1 U571 ( .A(ff_p0[4]), .Y(n258) );
  INVX1 U572 ( .A(ff_p0[6]), .Y(n256) );
  INVX1 U573 ( .A(ff_p0[0]), .Y(n262) );
  NAND2X1 U574 ( .A(rstcnt[4]), .B(n1143), .Y(n1133) );
  NOR4XL U575 ( .A(rstcnt[0]), .B(rstcnt[1]), .C(rstcnt[2]), .D(rstcnt[3]), 
        .Y(n1143) );
  NAND32X1 U576 ( .B(lg_pulse_cnt[1]), .C(lg_pulse_cnt[0]), .A(n1217), .Y(n193) );
  NOR3XL U577 ( .A(lg_pulse_cnt[2]), .B(lg_pulse_cnt[4]), .C(lg_pulse_cnt[3]), 
        .Y(n1217) );
  INVX1 U578 ( .A(r_phyrst[1]), .Y(n268) );
  NAND2X1 U579 ( .A(r_phyrst[0]), .B(n268), .Y(n1177) );
  NAND21X1 U580 ( .B(n20), .A(n7), .Y(n1222) );
  NAND32X1 U581 ( .B(di_rd_det_clr), .C(n1222), .A(n1191), .Y(aswkup) );
  NOR3XL U582 ( .A(dm_fault_clr), .B(p0_chg_clr), .C(i_tmrf), .Y(n1191) );
  INVX1 U583 ( .A(regD3_3), .Y(r_gpio_ie[0]) );
  OAI21X1 U584 ( .B(osc_low_clr), .C(n1222), .A(n152), .Y(osc_low_rstz) );
  AOI22X1 U585 ( .A(regDE[0]), .B(n1197), .C(regDE[1]), .D(n1198), .Y(n1196)
         );
  XNOR2XL U586 ( .A(di_p0[1]), .B(n261), .Y(n1198) );
  XNOR2XL U587 ( .A(di_p0[0]), .B(n262), .Y(n1197) );
  INVX1 U588 ( .A(regD3_7_), .Y(r_gpio_ie[1]) );
  NAND4X1 U589 ( .A(n1193), .B(n1194), .C(n1195), .D(n1196), .Y(as_p0_chg) );
  AOI22X1 U590 ( .A(regDE[6]), .B(n1203), .C(regDE[7]), .D(n1204), .Y(n1193)
         );
  AOI22X1 U591 ( .A(regDE[4]), .B(n1201), .C(regDE[5]), .D(n1202), .Y(n1194)
         );
  AOI22X1 U592 ( .A(regDE[2]), .B(n1199), .C(regDE[3]), .D(n1200), .Y(n1195)
         );
  INVX1 U593 ( .A(sfr_addr[7]), .Y(n154) );
  NAND32XL U594 ( .B(n235), .C(n183), .A(n105), .Y(n184) );
  NAND21X1 U595 ( .B(n233), .A(n232), .Y(n1130) );
  NAND21X1 U596 ( .B(n233), .A(n213), .Y(n187) );
  INVXL U597 ( .A(n8), .Y(n106) );
  NAND32XL U598 ( .B(n190), .C(n189), .A(n106), .Y(n231) );
  NAND32XL U599 ( .B(n215), .C(n190), .A(n106), .Y(n170) );
  NAND21X1 U600 ( .B(n190), .A(n163), .Y(n168) );
  NAND21X1 U601 ( .B(n190), .A(n200), .Y(n153) );
  AND4XL U602 ( .A(n212), .B(n270), .C(n235), .D(n189), .Y(we_143) );
  NAND32X1 U603 ( .B(n235), .C(n234), .A(n105), .Y(n236) );
  NAND32X1 U604 ( .B(n234), .C(n214), .A(n105), .Y(n222) );
  NAND32XL U605 ( .B(n214), .C(n183), .A(n105), .Y(n182) );
  NAND21X1 U606 ( .B(n105), .A(n235), .Y(n201) );
  NAND21X1 U607 ( .B(n231), .A(n230), .Y(n1137) );
  NAND21X1 U608 ( .B(n231), .A(n237), .Y(n229) );
  NAND21X1 U609 ( .B(n168), .A(n210), .Y(n191) );
  NAND21X1 U610 ( .B(n168), .A(n217), .Y(n164) );
  NAND32XL U611 ( .B(n214), .C(n208), .A(n215), .Y(n209) );
  NAND32XL U612 ( .B(n189), .C(n208), .A(n214), .Y(n181) );
  NAND21X1 U613 ( .B(n222), .A(n232), .Y(n1188) );
  NAND21X1 U614 ( .B(n222), .A(n227), .Y(n198) );
  NAND21X1 U615 ( .B(n201), .A(n200), .Y(n202) );
  NAND32XL U616 ( .B(n189), .C(n201), .A(n106), .Y(n233) );
  NAND32XL U617 ( .B(n215), .C(n201), .A(n106), .Y(n169) );
  NOR2XL U618 ( .A(n8), .B(n10), .Y(n270) );
  INVXL U619 ( .A(n9), .Y(n105) );
  NAND21XL U620 ( .B(n235), .A(n10), .Y(n190) );
  NAND43X1 U621 ( .B(n8), .C(n10), .D(n215), .A(n214), .Y(n216) );
  NAND21XL U622 ( .B(n215), .A(n8), .Y(n234) );
  NAND21XL U623 ( .B(n189), .A(n8), .Y(n183) );
  XOR2X1 U624 ( .A(add_180_carry[4]), .B(rstcnt[4]), .Y(N35) );
  OR2X1 U625 ( .A(lg_pulse_cnt[1]), .B(lg_pulse_cnt[0]), .Y(n245) );
  OAI21BBX1 U626 ( .A(lg_pulse_cnt[0]), .B(lg_pulse_cnt[1]), .C(n245), .Y(N103) );
  OR2X1 U627 ( .A(n245), .B(lg_pulse_cnt[2]), .Y(n246) );
  OAI21BBX1 U628 ( .A(n245), .B(lg_pulse_cnt[2]), .C(n246), .Y(N104) );
  XNOR2XL U629 ( .A(lg_pulse_cnt[3]), .B(n246), .Y(N105) );
  OR2X1 U630 ( .A(lg_pulse_cnt[3]), .B(n246), .Y(n247) );
  XNOR2XL U631 ( .A(lg_pulse_cnt[4]), .B(n247), .Y(N106) );
endmodule


module regbank_a0_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394;

  INVX4 U2565 ( .A(n3650), .Y(n3762) );
  OR2XL U2566 ( .A(A[314]), .B(n3650), .Y(n3642) );
  OR2XL U2567 ( .A(A[306]), .B(n3650), .Y(n3640) );
  INVX4 U2568 ( .A(n3650), .Y(n3775) );
  MUX2IX2 U2569 ( .D0(A[128]), .D1(A[384]), .S(n3775), .Y(n4359) );
  INVX4 U2570 ( .A(n3781), .Y(n3700) );
  INVX3 U2571 ( .A(n3834), .Y(n3668) );
  BUFX3 U2572 ( .A(n3749), .Y(n3602) );
  INVXL U2573 ( .A(n3751), .Y(n3749) );
  MUX2IX1 U2574 ( .D0(n3652), .D1(n3653), .S(n3740), .Y(n4334) );
  INVX2 U2575 ( .A(n3742), .Y(n3740) );
  NOR2X2 U2576 ( .A(n3775), .B(A[608]), .Y(n4373) );
  NOR2X2 U2577 ( .A(n3808), .B(A[624]), .Y(n4366) );
  INVX6 U2578 ( .A(n3781), .Y(n3808) );
  INVX2 U2579 ( .A(n3829), .Y(n3823) );
  BUFX3 U2580 ( .A(n3821), .Y(n3603) );
  INVXL U2581 ( .A(n3706), .Y(n3821) );
  INVX12 U2582 ( .A(n3670), .Y(n3830) );
  BUFX3 U2583 ( .A(n3747), .Y(n3604) );
  INVXL U2584 ( .A(n3752), .Y(n3747) );
  INVX2 U2585 ( .A(n3808), .Y(n3786) );
  INVX2 U2586 ( .A(n3808), .Y(n3785) );
  INVX2 U2587 ( .A(n3771), .Y(n3615) );
  INVXL U2588 ( .A(n3655), .Y(n3766) );
  MUX4X1 U2589 ( .D0(A[241]), .D1(A[753]), .D2(A[497]), .D3(A[1009]), .S0(
        n3817), .S1(n3768), .Y(n4271) );
  MUX4X1 U2590 ( .D0(A[249]), .D1(A[761]), .D2(A[505]), .D3(A[1017]), .S0(
        n3817), .S1(n3768), .Y(n4272) );
  MUX4XL U2591 ( .D0(n4292), .D1(n4293), .D2(n4294), .D3(n4295), .S0(n3817), 
        .S1(n3740), .Y(n4291) );
  MUX4XL U2592 ( .D0(A[181]), .D1(A[693]), .D2(A[437]), .D3(A[949]), .S0(n3817), .S1(n3805), .Y(n4001) );
  MUX4XL U2593 ( .D0(A[141]), .D1(A[653]), .D2(A[397]), .D3(A[909]), .S0(n3817), .S1(n3626), .Y(n4013) );
  INVX6 U2594 ( .A(n3828), .Y(n3817) );
  BUFX3 U2595 ( .A(n3735), .Y(n3605) );
  BUFX4 U2596 ( .A(n3735), .Y(n3606) );
  INVXL U2597 ( .A(n3743), .Y(n3735) );
  INVX3 U2598 ( .A(n3744), .Y(n3733) );
  INVXL U2599 ( .A(SH[3]), .Y(n3744) );
  INVX2 U2600 ( .A(n3742), .Y(n3741) );
  BUFX4 U2601 ( .A(SH[3]), .Y(n3732) );
  MUX2IXL U2602 ( .D0(A[233]), .D1(A[489]), .S(n3760), .Y(n4274) );
  MUX2X2 U2603 ( .D0(A[570]), .D1(A[826]), .S(n3760), .Y(n3641) );
  BUFX3 U2604 ( .A(n3760), .Y(n3614) );
  INVX2 U2605 ( .A(n3760), .Y(n3644) );
  MUX2IX1 U2606 ( .D0(A[218]), .D1(A[474]), .S(n3760), .Y(n4216) );
  INVX8 U2607 ( .A(n3781), .Y(n3760) );
  INVX8 U2608 ( .A(n3812), .Y(n3708) );
  INVX8 U2609 ( .A(SH[8]), .Y(n3812) );
  INVX6 U2610 ( .A(n3708), .Y(n3781) );
  BUFX3 U2611 ( .A(SH[8]), .Y(n3620) );
  INVX1 U2612 ( .A(SH[3]), .Y(n3742) );
  INVX1 U2613 ( .A(A[216]), .Y(n3687) );
  INVX1 U2614 ( .A(A[626]), .Y(n3647) );
  NOR2X1 U2615 ( .A(n3759), .B(A[634]), .Y(n4239) );
  INVX1 U2616 ( .A(A[282]), .Y(n3651) );
  INVX1 U2617 ( .A(A[794]), .Y(n3675) );
  INVX1 U2618 ( .A(A[538]), .Y(n3674) );
  INVX1 U2619 ( .A(A[674]), .Y(n3657) );
  INVX1 U2620 ( .A(A[162]), .Y(n3656) );
  INVX1 U2621 ( .A(A[930]), .Y(n3659) );
  INVX1 U2622 ( .A(A[418]), .Y(n3658) );
  INVX1 U2623 ( .A(n3780), .Y(n3801) );
  INVX2 U2624 ( .A(n3834), .Y(n3707) );
  INVX1 U2625 ( .A(n3729), .Y(n3827) );
  INVX2 U2626 ( .A(n3827), .Y(n3728) );
  INVX1 U2627 ( .A(SH[3]), .Y(n3743) );
  INVX1 U2628 ( .A(A[240]), .Y(n3701) );
  INVX1 U2629 ( .A(A[752]), .Y(n3702) );
  INVX1 U2630 ( .A(A[496]), .Y(n3703) );
  INVX1 U2631 ( .A(A[504]), .Y(n3715) );
  INVX1 U2632 ( .A(A[760]), .Y(n3714) );
  INVX1 U2633 ( .A(A[248]), .Y(n3713) );
  INVX1 U2634 ( .A(A[688]), .Y(n3722) );
  INVX1 U2635 ( .A(A[176]), .Y(n3721) );
  INVX1 U2636 ( .A(A[432]), .Y(n3723) );
  INVX1 U2637 ( .A(A[944]), .Y(n3724) );
  INVX1 U2638 ( .A(A[168]), .Y(n3683) );
  INVX1 U2639 ( .A(A[680]), .Y(n3682) );
  INVX1 U2640 ( .A(A[424]), .Y(n3685) );
  INVX1 U2641 ( .A(A[936]), .Y(n3684) );
  INVX1 U2642 ( .A(A[472]), .Y(n3686) );
  INVX1 U2643 ( .A(A[352]), .Y(n3691) );
  INVX1 U2644 ( .A(A[360]), .Y(n3667) );
  AND3X1 U2645 ( .A(n3726), .B(n3788), .C(n3643), .Y(n4377) );
  INVX1 U2646 ( .A(A[584]), .Y(n3643) );
  INVX1 U2647 ( .A(A[304]), .Y(n3673) );
  MUX2IX1 U2648 ( .D0(A[520]), .D1(A[776]), .S(n3762), .Y(n4394) );
  INVX1 U2649 ( .A(A[689]), .Y(n3636) );
  INVX1 U2650 ( .A(A[177]), .Y(n3635) );
  INVX1 U2651 ( .A(A[433]), .Y(n3637) );
  INVX1 U2652 ( .A(A[945]), .Y(n3638) );
  INVX1 U2653 ( .A(n3699), .Y(n3725) );
  NOR2X1 U2654 ( .A(n3773), .B(A[609]), .Y(n4314) );
  INVX2 U2655 ( .A(n3830), .Y(n3822) );
  INVX1 U2656 ( .A(n3830), .Y(n3824) );
  MUX4IX1 U2657 ( .D0(n3635), .D1(n3636), .D2(n3637), .D3(n3638), .S0(n3619), 
        .S1(n3711), .Y(n4285) );
  OR2X1 U2658 ( .A(n3745), .B(n4329), .Y(n3665) );
  INVX1 U2659 ( .A(n3758), .Y(n3757) );
  MUX2IX1 U2660 ( .D0(n3612), .D1(n3613), .S(n3810), .Y(n3692) );
  NAND2X1 U2661 ( .A(n4199), .B(n3607), .Y(n3608) );
  NAND2X1 U2662 ( .A(n4198), .B(n3660), .Y(n3609) );
  NAND2X1 U2663 ( .A(n3608), .B(n3609), .Y(B[2]) );
  INVX1 U2664 ( .A(n3660), .Y(n3607) );
  NOR2X1 U2665 ( .A(n3830), .B(A[832]), .Y(n3610) );
  NOR2X1 U2666 ( .A(n3799), .B(n3611), .Y(n4376) );
  INVX1 U2667 ( .A(n3610), .Y(n3611) );
  INVX1 U2668 ( .A(n3801), .Y(n3799) );
  MUX2IX1 U2669 ( .D0(n3717), .D1(n3718), .S(n3668), .Y(n3612) );
  MUX2IX1 U2670 ( .D0(n3719), .D1(n3720), .S(n3668), .Y(n3613) );
  INVX1 U2671 ( .A(A[160]), .Y(n3717) );
  INVX1 U2672 ( .A(A[672]), .Y(n3718) );
  INVX1 U2673 ( .A(A[416]), .Y(n3719) );
  INVX1 U2674 ( .A(A[928]), .Y(n3720) );
  INVX2 U2675 ( .A(n3813), .Y(n3810) );
  INVX6 U2676 ( .A(n3834), .Y(n3670) );
  MUX2IX1 U2677 ( .D0(A[657]), .D1(A[913]), .S(n3760), .Y(n4293) );
  MUX2IX1 U2678 ( .D0(A[232]), .D1(A[488]), .S(n3708), .Y(n4339) );
  INVX2 U2679 ( .A(n3810), .Y(n3795) );
  INVX1 U2680 ( .A(n3706), .Y(n3833) );
  BUFX1 U2681 ( .A(n3670), .Y(n3690) );
  INVXL U2682 ( .A(SH[4]), .Y(n3751) );
  INVX1 U2683 ( .A(n3758), .Y(n3756) );
  INVX1 U2684 ( .A(SH[6]), .Y(n3758) );
  INVX1 U2685 ( .A(n3751), .Y(n3748) );
  INVX1 U2686 ( .A(SH[7]), .Y(n3660) );
  INVX1 U2687 ( .A(n3742), .Y(n3739) );
  INVX2 U2688 ( .A(n3743), .Y(n3734) );
  INVX1 U2689 ( .A(n3778), .Y(n3772) );
  INVX3 U2690 ( .A(n3779), .Y(n3769) );
  INVX1 U2691 ( .A(n3615), .Y(n3616) );
  INVX1 U2692 ( .A(n3615), .Y(n3617) );
  INVX2 U2693 ( .A(n3828), .Y(n3618) );
  INVX3 U2694 ( .A(n3828), .Y(n3619) );
  MUX2IX1 U2695 ( .D0(n4313), .D1(n4314), .S(n3619), .Y(n3680) );
  INVX2 U2696 ( .A(n3828), .Y(n3818) );
  BUFX4 U2697 ( .A(SH[8]), .Y(n3621) );
  BUFX1 U2698 ( .A(SH[8]), .Y(n3688) );
  INVX1 U2699 ( .A(n3707), .Y(n3832) );
  INVXL U2700 ( .A(n3826), .Y(n3622) );
  INVXL U2701 ( .A(n3826), .Y(n3623) );
  MUX2IX1 U2702 ( .D0(A[656]), .D1(A[912]), .S(n3688), .Y(n4354) );
  INVXL U2703 ( .A(n3766), .Y(n3624) );
  INVXL U2704 ( .A(n3624), .Y(n3625) );
  INVXL U2705 ( .A(n3624), .Y(n3626) );
  INVXL U2706 ( .A(n3624), .Y(n3627) );
  INVX1 U2707 ( .A(n3602), .Y(n3661) );
  MUX2IX1 U2708 ( .D0(A[473]), .D1(A[217]), .S(n3777), .Y(n4281) );
  INVX4 U2709 ( .A(n3780), .Y(n3711) );
  INVX1 U2710 ( .A(n3809), .Y(n3777) );
  MUX2IX1 U2711 ( .D0(n4337), .D1(n4336), .S(n3751), .Y(n4335) );
  MUX2IX1 U2712 ( .D0(A[440]), .D1(A[184]), .S(n3812), .Y(n4349) );
  MUX2X2 U2713 ( .D0(n3696), .D1(n3697), .S(n3734), .Y(n4337) );
  MUX4X1 U2714 ( .D0(n3682), .D1(n3683), .D2(n3684), .D3(n3685), .S0(n3834), 
        .S1(n3620), .Y(n3694) );
  INVX3 U2715 ( .A(n3825), .Y(n3819) );
  MUX2IX1 U2716 ( .D0(n4351), .D1(n4352), .S(n3604), .Y(n4332) );
  MUX2IX1 U2717 ( .D0(n4358), .D1(n4357), .S(n3744), .Y(n4351) );
  MUX4XL U2718 ( .D0(n3899), .D1(n3900), .D2(n3901), .D3(n3902), .S0(n3819), 
        .S1(n3740), .Y(n3893) );
  MUX4XL U2719 ( .D0(n3885), .D1(n3886), .D2(n3887), .D3(n3888), .S0(n3819), 
        .S1(n3740), .Y(n3874) );
  MUX4XL U2720 ( .D0(A[246]), .D1(A[758]), .D2(A[502]), .D3(A[1014]), .S0(
        n3819), .S1(n3768), .Y(n3916) );
  MUX4XL U2721 ( .D0(A[143]), .D1(A[655]), .D2(A[399]), .D3(A[911]), .S0(n3819), .S1(n3767), .Y(n3869) );
  MUX4X1 U2722 ( .D0(n3722), .D1(n3721), .D2(n3724), .D3(n3723), .S0(n3834), 
        .S1(n3621), .Y(n3693) );
  NAND2X1 U2723 ( .A(n4349), .B(n3628), .Y(n3629) );
  NAND2XL U2724 ( .A(n4350), .B(n3729), .Y(n3630) );
  NAND2X1 U2725 ( .A(n3630), .B(n3629), .Y(n3695) );
  INVXL U2726 ( .A(n3729), .Y(n3628) );
  NOR2XL U2727 ( .A(A[284]), .B(n3795), .Y(n4118) );
  NOR2XL U2728 ( .A(A[276]), .B(n3795), .Y(n4116) );
  NOR2XL U2729 ( .A(A[308]), .B(n3795), .Y(n4112) );
  INVX3 U2730 ( .A(n3812), .Y(n3809) );
  BUFX12 U2731 ( .A(n3812), .Y(n3650) );
  MUX2X1 U2732 ( .D0(n3686), .D1(n3687), .S(n3812), .Y(n4346) );
  INVX2 U2733 ( .A(n3809), .Y(n3784) );
  MUX4XL U2734 ( .D0(n3849), .D1(n3850), .D2(n3851), .D3(n3852), .S0(n3746), 
        .S1(n3739), .Y(n3839) );
  MUX4XL U2735 ( .D0(n3856), .D1(n3857), .D2(n3858), .D3(n3859), .S0(n3746), 
        .S1(n3740), .Y(n3838) );
  MUX4XL U2736 ( .D0(n4073), .D1(n4074), .D2(n4075), .D3(n4076), .S0(n3746), 
        .S1(n3737), .Y(n4055) );
  MUX4XL U2737 ( .D0(n3922), .D1(n3923), .D2(n3924), .D3(n3925), .S0(n3746), 
        .S1(n3739), .Y(n3912) );
  MUX4XL U2738 ( .D0(n3929), .D1(n3930), .D2(n3931), .D3(n3932), .S0(n3746), 
        .S1(n3739), .Y(n3911) );
  MUX4XL U2739 ( .D0(n3993), .D1(n3994), .D2(n3995), .D3(n3996), .S0(n3746), 
        .S1(n3738), .Y(n3983) );
  MUX4XL U2740 ( .D0(n4066), .D1(n4067), .D2(n4068), .D3(n4069), .S0(n3746), 
        .S1(n3737), .Y(n4056) );
  MUX4XL U2741 ( .D0(n4000), .D1(n4001), .D2(n4002), .D3(n4003), .S0(n3746), 
        .S1(n3738), .Y(n3982) );
  NOR2XL U2742 ( .A(A[305]), .B(n3785), .Y(n4319) );
  MUX2IX1 U2743 ( .D0(A[224]), .D1(A[480]), .S(n3621), .Y(n4338) );
  MUX4X1 U2744 ( .D0(n4273), .D1(n4274), .D2(n4275), .D3(n4276), .S0(n3732), 
        .S1(n3822), .Y(n4269) );
  MUX4IX1 U2745 ( .D0(n4324), .D1(n4323), .D2(n4326), .D3(n4325), .S0(n3832), 
        .S1(n3740), .Y(n3663) );
  MUX2IX1 U2746 ( .D0(n4291), .D1(n4290), .S(n3661), .Y(n4265) );
  INVXL U2747 ( .A(n3699), .Y(n3726) );
  INVX1 U2748 ( .A(n3707), .Y(n3645) );
  INVXL U2749 ( .A(n3807), .Y(n3790) );
  INVX3 U2750 ( .A(n3810), .Y(n3778) );
  INVXL U2751 ( .A(n3810), .Y(n3789) );
  INVX3 U2752 ( .A(n3778), .Y(n3771) );
  MUX2IX1 U2753 ( .D0(n4353), .D1(n4354), .S(n3819), .Y(n3631) );
  MUX2IX1 U2754 ( .D0(n4355), .D1(n4356), .S(n3819), .Y(n3632) );
  MUX2IX1 U2755 ( .D0(n3631), .D1(n3632), .S(n3732), .Y(n4352) );
  NOR2X1 U2756 ( .A(A[408]), .B(n3784), .Y(n4355) );
  INVX2 U2757 ( .A(n3781), .Y(n3761) );
  MUX2IX1 U2758 ( .D0(n4300), .D1(n4299), .S(n3758), .Y(n4263) );
  INVX1 U2759 ( .A(n3668), .Y(n3706) );
  MUX2IX1 U2760 ( .D0(n4394), .D1(n4393), .S(n3830), .Y(n4392) );
  MUX2IXL U2761 ( .D0(A[32]), .D1(A[544]), .S(n3729), .Y(n3633) );
  MUX2IXL U2762 ( .D0(A[288]), .D1(A[800]), .S(n3729), .Y(n3634) );
  MUX2IXL U2763 ( .D0(n3633), .D1(n3634), .S(n3762), .Y(n4390) );
  MUX2IX1 U2764 ( .D0(A[121]), .D1(A[377]), .S(n3807), .Y(n4306) );
  MUX4X1 U2765 ( .D0(n3703), .D1(n3704), .D2(n3701), .D3(n3702), .S0(n3729), 
        .S1(n3780), .Y(n3696) );
  MUX4IX1 U2766 ( .D0(n3639), .D1(n3640), .D2(n3641), .D3(n3642), .S0(n3646), 
        .S1(n3739), .Y(n4253) );
  MUX2X2 U2767 ( .D0(A[818]), .D1(A[562]), .S(n3778), .Y(n3639) );
  NOR21X1 U2768 ( .B(n3813), .A(A[696]), .Y(n4350) );
  INVXL U2769 ( .A(n3780), .Y(n3767) );
  AND2X1 U2770 ( .A(n3673), .B(n3621), .Y(n4382) );
  AND2X1 U2771 ( .A(n3691), .B(n3620), .Y(n4372) );
  NOR2XL U2772 ( .A(A[1000]), .B(n3784), .Y(n4341) );
  NOR2XL U2773 ( .A(A[274]), .B(n3650), .Y(n4254) );
  INVX1 U2774 ( .A(n3777), .Y(n3776) );
  MUX2IXL U2775 ( .D0(A[378]), .D1(A[122]), .S(n3655), .Y(n4237) );
  INVXL U2776 ( .A(n3726), .Y(n3646) );
  AND2XL U2777 ( .A(n3777), .B(n3647), .Y(n4238) );
  MUX4X1 U2778 ( .D0(n4208), .D1(n4209), .D2(n4210), .D3(n4211), .S0(n3733), 
        .S1(n3603), .Y(n4204) );
  MUX2IX1 U2779 ( .D0(n4369), .D1(n4368), .S(n3745), .Y(n4362) );
  INVX1 U2780 ( .A(A[1016]), .Y(n3716) );
  INVX1 U2781 ( .A(A[1008]), .Y(n3704) );
  INVX1 U2782 ( .A(A[992]), .Y(n3672) );
  INVX1 U2783 ( .A(A[984]), .Y(n3712) );
  MUX2IXL U2784 ( .D0(A[712]), .D1(A[968]), .S(n3620), .Y(n4348) );
  NAND2X1 U2785 ( .A(n4376), .B(n3745), .Y(n3648) );
  NAND2XL U2786 ( .A(n4377), .B(n3741), .Y(n3649) );
  NAND2X1 U2787 ( .A(n3648), .B(n3649), .Y(n4360) );
  MUX4IX1 U2788 ( .D0(n4361), .D1(n4360), .D2(n4363), .D3(n4362), .S0(n3755), 
        .S1(n3602), .Y(n3710) );
  MUX4IX1 U2789 ( .D0(n4333), .D1(n4332), .D2(n4335), .D3(n4334), .S0(n3755), 
        .S1(n3757), .Y(n3731) );
  MUX2IX1 U2790 ( .D0(A[536]), .D1(A[792]), .S(n3620), .Y(n4389) );
  MUX4IX1 U2791 ( .D0(n4379), .D1(n4378), .D2(n4381), .D3(n4380), .S0(n3755), 
        .S1(n3602), .Y(n3709) );
  INVXL U2792 ( .A(n3812), .Y(n3811) );
  MUX2IX1 U2793 ( .D0(A[664]), .D1(A[920]), .S(n3688), .Y(n4356) );
  INVX8 U2794 ( .A(SH[9]), .Y(n3834) );
  NOR21XL U2795 ( .B(n3651), .A(n3788), .Y(n4256) );
  MUX4X1 U2796 ( .D0(A[434]), .D1(A[946]), .D2(A[178]), .D3(A[690]), .S0(n3707), .S1(n3644), .Y(n4220) );
  MUX2IXL U2797 ( .D0(A[521]), .D1(A[777]), .S(n3768), .Y(n4331) );
  INVX3 U2798 ( .A(n3780), .Y(n3768) );
  MUX4X1 U2799 ( .D0(A[161]), .D1(A[673]), .D2(A[417]), .D3(A[929]), .S0(n3818), .S1(n3711), .Y(n4284) );
  MUX4X1 U2800 ( .D0(A[137]), .D1(A[649]), .D2(A[393]), .D3(A[905]), .S0(n3618), .S1(n3711), .Y(n4297) );
  MUX2IX1 U2801 ( .D0(n4315), .D1(n4316), .S(n3618), .Y(n3681) );
  MUX4X1 U2802 ( .D0(n4383), .D1(n4382), .D2(n4385), .D3(n4384), .S0(n3706), 
        .S1(n3741), .Y(n4381) );
  MUX2IX1 U2803 ( .D0(n4342), .D1(n4343), .S(n3654), .Y(n3652) );
  MUX2IX1 U2804 ( .D0(n4344), .D1(n4345), .S(n3654), .Y(n3653) );
  NAND31XL U2805 ( .C(A[960]), .A(n3769), .B(n3725), .Y(n4342) );
  NAND31XL U2806 ( .C(A[976]), .A(n3769), .B(n3707), .Y(n4343) );
  NAND2XL U2807 ( .A(n4348), .B(n3817), .Y(n4344) );
  INVXL U2808 ( .A(n3752), .Y(n3654) );
  MUX4X1 U2809 ( .D0(A[136]), .D1(A[648]), .D2(A[392]), .D3(A[904]), .S0(SH[9]), .S1(n3621), .Y(n4358) );
  NAND31XL U2810 ( .C(A[962]), .A(n3770), .B(n3823), .Y(n4212) );
  INVXL U2811 ( .A(n3708), .Y(n3787) );
  INVXL U2812 ( .A(n3708), .Y(n3788) );
  INVXL U2813 ( .A(n3809), .Y(n3655) );
  NOR2XL U2814 ( .A(n3771), .B(A[633]), .Y(n4308) );
  MUX2IXL U2815 ( .D0(A[825]), .D1(A[569]), .S(n3780), .Y(n4322) );
  INVX6 U2816 ( .A(n3708), .Y(n3780) );
  MUX4X1 U2817 ( .D0(n4373), .D1(n4372), .D2(n4375), .D3(n4374), .S0(n3645), 
        .S1(n3741), .Y(n4361) );
  MUX2IXL U2818 ( .D0(A[561]), .D1(A[817]), .S(n3811), .Y(n4320) );
  MUX2IXL U2819 ( .D0(A[185]), .D1(A[441]), .S(n3769), .Y(n4288) );
  MUX4IX1 U2820 ( .D0(n3693), .D1(n3692), .D2(n3695), .D3(n3694), .S0(n3751), 
        .S1(n3741), .Y(n4333) );
  INVXL U2821 ( .A(n3825), .Y(n3689) );
  INVXL U2822 ( .A(n3781), .Y(n3759) );
  MUX4XL U2823 ( .D0(A[39]), .D1(A[551]), .D2(A[295]), .D3(A[807]), .S0(n3819), 
        .S1(n3700), .Y(n3903) );
  NAND31XL U2824 ( .C(A[965]), .A(n3700), .B(n3823), .Y(n3993) );
  NAND31XL U2825 ( .C(A[963]), .A(n3700), .B(n3823), .Y(n4139) );
  MUX4X1 U2826 ( .D0(n4305), .D1(n4306), .D2(n4307), .D3(n4308), .S0(n3732), 
        .S1(n3603), .Y(n4304) );
  MUX4XL U2827 ( .D0(A[174]), .D1(A[686]), .D2(A[430]), .D3(A[942]), .S0(n3819), .S1(n3767), .Y(n3931) );
  MUX4XL U2828 ( .D0(A[166]), .D1(A[678]), .D2(A[422]), .D3(A[934]), .S0(n3819), .S1(n3765), .Y(n3929) );
  MUX4XL U2829 ( .D0(A[35]), .D1(A[547]), .D2(A[291]), .D3(A[803]), .S0(n3815), 
        .S1(n3666), .Y(n4193) );
  MUX4XL U2830 ( .D0(A[43]), .D1(A[555]), .D2(A[299]), .D3(A[811]), .S0(n3815), 
        .S1(n3764), .Y(n4194) );
  MUX4XL U2831 ( .D0(A[242]), .D1(A[754]), .D2(A[498]), .D3(A[1010]), .S0(
        n3707), .S1(n3711), .Y(n4206) );
  MUX4X1 U2832 ( .D0(n4251), .D1(n4250), .D2(n4253), .D3(n4252), .S0(n3755), 
        .S1(n3602), .Y(n4234) );
  MUX4IX1 U2833 ( .D0(n3656), .D1(n3657), .D2(n3658), .D3(n3659), .S0(n3707), 
        .S1(n3768), .Y(n4219) );
  MUX2X2 U2834 ( .D0(n4264), .D1(n4263), .S(n3660), .Y(B[1]) );
  MUX4IX1 U2835 ( .D0(n3662), .D1(n3663), .D2(n3664), .D3(n3665), .S0(n3755), 
        .S1(n3661), .Y(n4299) );
  MUX4IX1 U2836 ( .D0(n4319), .D1(n4320), .D2(n4321), .D3(n4322), .S0(n3619), 
        .S1(n3740), .Y(n3662) );
  MUX2X1 U2837 ( .D0(n4327), .D1(n4328), .S(n3733), .Y(n3664) );
  MUX2IX1 U2838 ( .D0(n3680), .D1(n3681), .S(n3740), .Y(n4302) );
  MUX4X1 U2839 ( .D0(A[41]), .D1(A[553]), .D2(A[297]), .D3(A[809]), .S0(n3725), 
        .S1(n3711), .Y(n4328) );
  NOR2XL U2840 ( .A(A[368]), .B(n3783), .Y(n4364) );
  INVXL U2841 ( .A(n3785), .Y(n3666) );
  NOR21XL U2842 ( .B(n3667), .A(n3783), .Y(n4374) );
  MUX2IX1 U2843 ( .D0(A[528]), .D1(A[784]), .S(n3621), .Y(n4387) );
  MUX2IX1 U2844 ( .D0(A[120]), .D1(A[376]), .S(n3620), .Y(n4365) );
  MUX4IX1 U2845 ( .D0(n4238), .D1(n4239), .D2(n4236), .D3(n4237), .S0(n3733), 
        .S1(n3832), .Y(n3676) );
  INVXL U2846 ( .A(n3791), .Y(n3669) );
  INVX1 U2847 ( .A(n3806), .Y(n3791) );
  INVX3 U2848 ( .A(n3670), .Y(n3825) );
  MUX2IX1 U2849 ( .D0(n4347), .D1(n4346), .S(n3830), .Y(n4345) );
  INVXL U2850 ( .A(n3617), .Y(n3671) );
  NOR21XL U2851 ( .B(n3672), .A(n3784), .Y(n4340) );
  INVXL U2852 ( .A(SH[9]), .Y(n3699) );
  MUX2XL U2853 ( .D0(n3675), .D1(n3674), .S(n3813), .Y(n4257) );
  MUX4IX1 U2854 ( .D0(n3676), .D1(n3677), .D2(n3678), .D3(n3679), .S0(n3755), 
        .S1(n3661), .Y(n4235) );
  MUX2X1 U2855 ( .D0(n4240), .D1(n4241), .S(n3734), .Y(n3677) );
  MUX4IX1 U2856 ( .D0(n4244), .D1(n4245), .D2(n4246), .D3(n4247), .S0(n3690), 
        .S1(n3739), .Y(n3678) );
  MUX2IX1 U2857 ( .D0(n4248), .D1(n4249), .S(n3741), .Y(n3679) );
  INVX2 U2858 ( .A(n3755), .Y(n3754) );
  NOR2XL U2859 ( .A(A[361]), .B(n3785), .Y(n4315) );
  NOR2XL U2860 ( .A(n3773), .B(A[617]), .Y(n4316) );
  MUX4X1 U2861 ( .D0(n4257), .D1(n4256), .D2(n4255), .D3(n4254), .S0(n3829), 
        .S1(n3745), .Y(n4252) );
  NOR2XL U2862 ( .A(A[369]), .B(n3786), .Y(n4305) );
  NOR2XL U2863 ( .A(A[345]), .B(n3786), .Y(n4311) );
  NOR2XL U2864 ( .A(A[401]), .B(n3786), .Y(n4292) );
  NOR2XL U2865 ( .A(A[409]), .B(n3786), .Y(n4294) );
  NOR2XL U2866 ( .A(A[273]), .B(n3777), .Y(n4323) );
  NOR2XL U2867 ( .A(A[281]), .B(n3777), .Y(n4325) );
  INVX2 U2868 ( .A(SH[8]), .Y(n3813) );
  NOR2XL U2869 ( .A(n3744), .B(n3905), .Y(n3891) );
  MUX2IXL U2870 ( .D0(n3843), .D1(n3844), .S(n3733), .Y(n3842) );
  MUX4XL U2871 ( .D0(n4021), .D1(n4022), .D2(n4023), .D3(n4024), .S0(n3733), 
        .S1(n3822), .Y(n4020) );
  MUX4XL U2872 ( .D0(n3989), .D1(n3990), .D2(n3991), .D3(n3992), .S0(n3733), 
        .S1(n3823), .Y(n3985) );
  MUX4XL U2873 ( .D0(n4062), .D1(n4063), .D2(n4064), .D3(n4065), .S0(n3733), 
        .S1(n3822), .Y(n4058) );
  NOR2XL U2874 ( .A(A[353]), .B(n3785), .Y(n4313) );
  INVX3 U2875 ( .A(n3668), .Y(n3828) );
  NOR2XL U2876 ( .A(A[272]), .B(n3782), .Y(n4386) );
  NOR2XL U2877 ( .A(n3772), .B(A[606]), .Y(n3957) );
  NOR2XL U2878 ( .A(n3772), .B(A[630]), .Y(n3952) );
  NOR2XL U2879 ( .A(n3772), .B(A[638]), .Y(n3953) );
  NOR2XL U2880 ( .A(n3772), .B(A[615]), .Y(n3886) );
  NOR2XL U2881 ( .A(n3773), .B(A[631]), .Y(n3879) );
  NOR2XL U2882 ( .A(n3772), .B(A[605]), .Y(n4028) );
  INVX2 U2883 ( .A(n3834), .Y(n3729) );
  MUX4XL U2884 ( .D0(n3950), .D1(n3951), .D2(n3952), .D3(n3953), .S0(n3734), 
        .S1(n3822), .Y(n3949) );
  MUX4XL U2885 ( .D0(n3918), .D1(n3919), .D2(n3920), .D3(n3921), .S0(n3739), 
        .S1(n3822), .Y(n3914) );
  MUX4XL U2886 ( .D0(n3877), .D1(n3878), .D2(n3879), .D3(n3880), .S0(n3733), 
        .S1(n3823), .Y(n3876) );
  MUX4XL U2887 ( .D0(n3845), .D1(n3846), .D2(n3847), .D3(n3848), .S0(n3732), 
        .S1(n3822), .Y(n3841) );
  MUX4XL U2888 ( .D0(n4167), .D1(n4168), .D2(n4169), .D3(n4170), .S0(n3732), 
        .S1(n3822), .Y(n4166) );
  MUX4XL U2889 ( .D0(n4135), .D1(n4136), .D2(n4137), .D3(n4138), .S0(n3732), 
        .S1(n3822), .Y(n4131) );
  INVX2 U2890 ( .A(n3778), .Y(n3773) );
  MUX4X1 U2891 ( .D0(n4386), .D1(n4387), .D2(n4388), .D3(n4389), .S0(n3689), 
        .S1(n3741), .Y(n4380) );
  INVX1 U2892 ( .A(n3752), .Y(n3746) );
  MUX2IX1 U2893 ( .D0(A[530]), .D1(A[786]), .S(n3762), .Y(n4255) );
  MUX4X1 U2894 ( .D0(n4268), .D1(n4267), .D2(n4266), .D3(n4265), .S0(n3755), 
        .S1(n3758), .Y(n4264) );
  MUX2IX1 U2895 ( .D0(A[824]), .D1(A[568]), .S(n3650), .Y(n4385) );
  MUX4X1 U2896 ( .D0(n3714), .D1(n3713), .D2(n3716), .D3(n3715), .S0(n3825), 
        .S1(n3806), .Y(n3697) );
  MUX4XL U2897 ( .D0(n4094), .D1(n4095), .D2(n4096), .D3(n4097), .S0(n3733), 
        .S1(n3603), .Y(n4093) );
  MUX4X1 U2898 ( .D0(n4301), .D1(n4302), .D2(n4303), .D3(n4304), .S0(n3754), 
        .S1(n3602), .Y(n4300) );
  MUX2IX1 U2899 ( .D0(n3730), .D1(n3731), .S(SH[7]), .Y(B[0]) );
  INVXL U2900 ( .A(n3670), .Y(n3829) );
  MUX4XL U2901 ( .D0(n3970), .D1(n3971), .D2(n3972), .D3(n3973), .S0(n3817), 
        .S1(n3738), .Y(n3964) );
  MUX4XL U2902 ( .D0(A[245]), .D1(A[757]), .D2(A[501]), .D3(A[1013]), .S0(
        n3618), .S1(n3705), .Y(n3987) );
  MUX4XL U2903 ( .D0(A[253]), .D1(A[765]), .D2(A[509]), .D3(A[1021]), .S0(
        n3619), .S1(n3627), .Y(n3988) );
  MUX4XL U2904 ( .D0(n4189), .D1(n4190), .D2(n4191), .D3(n4192), .S0(n3618), 
        .S1(n3738), .Y(n4183) );
  AND2X1 U2905 ( .A(n3712), .B(n3811), .Y(n4347) );
  MUX2IX1 U2906 ( .D0(n3709), .D1(n3710), .S(n3756), .Y(n3730) );
  MUX4X1 U2907 ( .D0(n4341), .D1(n4340), .D2(n4339), .D3(n4338), .S0(n3743), 
        .S1(n3831), .Y(n4336) );
  INVXL U2908 ( .A(n3729), .Y(n3831) );
  MUX4XL U2909 ( .D0(A[38]), .D1(A[550]), .D2(A[294]), .D3(A[806]), .S0(n3619), 
        .S1(n3773), .Y(n3974) );
  INVXL U2910 ( .A(n3813), .Y(n3807) );
  INVX1 U2911 ( .A(n3825), .Y(n3727) );
  INVXL U2912 ( .A(n3759), .Y(n3698) );
  INVX3 U2913 ( .A(n3708), .Y(n3779) );
  NAND31XL U2914 ( .C(A[978]), .A(n3770), .B(n3707), .Y(n4213) );
  NAND31XL U2915 ( .C(A[977]), .A(n3700), .B(n3726), .Y(n4278) );
  NAND31XL U2916 ( .C(A[981]), .A(n3770), .B(n3622), .Y(n3994) );
  MUX2IXL U2917 ( .D0(n4004), .D1(n4005), .S(n3603), .Y(n4003) );
  MUX2IXL U2918 ( .D0(n3997), .D1(n3998), .S(n3603), .Y(n3996) );
  MUX2IXL U2919 ( .D0(n3956), .D1(n3957), .S(n3603), .Y(n3955) );
  MUX2IXL U2920 ( .D0(n3933), .D1(n3934), .S(n3603), .Y(n3932) );
  MUX2IXL U2921 ( .D0(n3906), .D1(n3907), .S(n3603), .Y(n3905) );
  MUX2IXL U2922 ( .D0(n3883), .D1(n3884), .S(n3603), .Y(n3882) );
  MUX2IXL U2923 ( .D0(n3853), .D1(n3854), .S(n3603), .Y(n3852) );
  INVXL U2924 ( .A(n3800), .Y(n3705) );
  INVX1 U2925 ( .A(n3779), .Y(n3770) );
  MUX2IX1 U2926 ( .D0(A[560]), .D1(A[816]), .S(n3708), .Y(n4383) );
  NOR2XL U2927 ( .A(A[400]), .B(n3813), .Y(n4353) );
  NOR2XL U2928 ( .A(A[1007]), .B(n3671), .Y(n3848) );
  MUX4XL U2929 ( .D0(n3864), .D1(n3865), .D2(n3866), .D3(n3867), .S0(n3727), 
        .S1(n3732), .Y(n3863) );
  MUX4XL U2930 ( .D0(n4043), .D1(n4044), .D2(n4045), .D3(n4046), .S0(n3816), 
        .S1(n3737), .Y(n4037) );
  MUX4XL U2931 ( .D0(A[37]), .D1(A[549]), .D2(A[293]), .D3(A[805]), .S0(n3816), 
        .S1(n3768), .Y(n4047) );
  MUX4XL U2932 ( .D0(A[45]), .D1(A[557]), .D2(A[301]), .D3(A[813]), .S0(n3816), 
        .S1(n3669), .Y(n4048) );
  MUX4XL U2933 ( .D0(A[244]), .D1(A[756]), .D2(A[500]), .D3(A[1012]), .S0(
        n3816), .S1(n3763), .Y(n4060) );
  MUX4XL U2934 ( .D0(A[252]), .D1(A[764]), .D2(A[508]), .D3(A[1020]), .S0(
        n3816), .S1(n3768), .Y(n4061) );
  MUX2IXL U2935 ( .D0(n4311), .D1(n4312), .S(n3725), .Y(n4310) );
  MUX4XL U2936 ( .D0(n4277), .D1(n4278), .D2(n4279), .D3(n4280), .S0(n3604), 
        .S1(n3740), .Y(n4267) );
  NOR2XL U2937 ( .A(n3774), .B(A[614]), .Y(n3959) );
  NOR2XL U2938 ( .A(n3774), .B(n3830), .Y(n3890) );
  NOR2XL U2939 ( .A(n3774), .B(A[622]), .Y(n3960) );
  NOR2XL U2940 ( .A(n3774), .B(A[629]), .Y(n4023) );
  NOR2XL U2941 ( .A(n3774), .B(A[703]), .Y(n3861) );
  NOR2XL U2942 ( .A(n3774), .B(A[636]), .Y(n4097) );
  NOR2XL U2943 ( .A(n3774), .B(A[700]), .Y(n4078) );
  NOR2XL U2944 ( .A(n3774), .B(A[699]), .Y(n4151) );
  MUX4XL U2945 ( .D0(n3966), .D1(n3967), .D2(n3968), .D3(n3969), .S0(n3623), 
        .S1(n3738), .Y(n3965) );
  MUX4XL U2946 ( .D0(n3937), .D1(n3938), .D2(n3939), .D3(n3940), .S0(n3623), 
        .S1(n3739), .Y(n3936) );
  MUX4XL U2947 ( .D0(A[46]), .D1(A[558]), .D2(A[302]), .D3(A[814]), .S0(n3622), 
        .S1(n3626), .Y(n3975) );
  MUX4XL U2948 ( .D0(A[142]), .D1(A[654]), .D2(A[398]), .D3(A[910]), .S0(n3623), .S1(n3765), .Y(n3942) );
  MUX4XL U2949 ( .D0(A[182]), .D1(A[694]), .D2(A[438]), .D3(A[950]), .S0(n3622), .S1(n3803), .Y(n3930) );
  MUX4XL U2950 ( .D0(A[33]), .D1(A[545]), .D2(A[289]), .D3(A[801]), .S0(n3725), 
        .S1(n3711), .Y(n4327) );
  NAND32XL U2951 ( .B(A[598]), .C(n3666), .A(n3824), .Y(n3954) );
  NAND32XL U2952 ( .B(A[599]), .C(n3805), .A(n3824), .Y(n3881) );
  NAND32XL U2953 ( .B(A[597]), .C(n3765), .A(n3824), .Y(n4025) );
  NAND32XL U2954 ( .B(A[596]), .C(n3767), .A(n3824), .Y(n4098) );
  NAND31XL U2955 ( .C(A[964]), .A(n3802), .B(n3823), .Y(n4066) );
  NAND31XL U2956 ( .C(A[980]), .A(n3770), .B(n3729), .Y(n4067) );
  NAND32XL U2957 ( .B(A[595]), .C(n3770), .A(n3824), .Y(n4171) );
  NAND32XL U2958 ( .B(A[593]), .C(n3700), .A(n3824), .Y(n4309) );
  NAND32XL U2959 ( .B(A[594]), .C(n3769), .A(n3824), .Y(n4240) );
  MUX4XL U2960 ( .D0(n3958), .D1(n3666), .D2(n3959), .D3(n3960), .S0(n3733), 
        .S1(n3822), .Y(n3947) );
  NOR2XL U2961 ( .A(n3666), .B(A[637]), .Y(n4024) );
  NOR2XL U2962 ( .A(n3666), .B(A[604]), .Y(n4101) );
  NOR2XL U2963 ( .A(n3666), .B(A[628]), .Y(n4096) );
  NOR2XL U2964 ( .A(n3666), .B(A[620]), .Y(n4105) );
  NOR2XL U2965 ( .A(n3666), .B(A[612]), .Y(n4103) );
  NOR2XL U2966 ( .A(n3775), .B(A[600]), .Y(n4371) );
  NOR2XL U2967 ( .A(n3775), .B(A[632]), .Y(n4367) );
  NOR2XL U2968 ( .A(n3775), .B(A[616]), .Y(n4375) );
  INVX1 U2969 ( .A(n3671), .Y(n3774) );
  MUX2IXL U2970 ( .D0(A[563]), .D1(A[819]), .S(n3761), .Y(n4186) );
  MUX2IXL U2971 ( .D0(A[131]), .D1(A[387]), .S(n3761), .Y(n4160) );
  MUX2IXL U2972 ( .D0(A[130]), .D1(A[386]), .S(n3614), .Y(n4233) );
  MUX2IXL U2973 ( .D0(A[134]), .D1(A[390]), .S(n3802), .Y(n3943) );
  MUX2IXL U2974 ( .D0(A[659]), .D1(A[915]), .S(n3761), .Y(n4155) );
  INVXL U2975 ( .A(n3742), .Y(n3738) );
  INVXL U2976 ( .A(n3826), .Y(n3816) );
  INVXL U2977 ( .A(n3646), .Y(n3820) );
  INVXL U2978 ( .A(n3745), .Y(n3737) );
  INVXL U2979 ( .A(n3751), .Y(n3750) );
  INVXL U2980 ( .A(n3755), .Y(n3753) );
  MUX4XL U2981 ( .D0(A[250]), .D1(A[762]), .D2(A[506]), .D3(A[1018]), .S0(
        n3726), .S1(n3711), .Y(n4207) );
  MUX2IXL U2982 ( .D0(A[713]), .D1(A[969]), .S(n3769), .Y(n4283) );
  MUX2IXL U2983 ( .D0(A[714]), .D1(A[970]), .S(n3760), .Y(n4218) );
  MUX2IXL U2984 ( .D0(A[219]), .D1(A[475]), .S(n3763), .Y(n4143) );
  MUX4XL U2985 ( .D0(A[251]), .D1(A[763]), .D2(A[507]), .D3(A[1019]), .S0(
        n3816), .S1(n3802), .Y(n4134) );
  MUX2IXL U2986 ( .D0(A[715]), .D1(A[971]), .S(n3626), .Y(n4145) );
  MUX4XL U2987 ( .D0(n4054), .D1(n4055), .D2(n4056), .D3(n4057), .S0(n3753), 
        .S1(n3756), .Y(n4053) );
  MUX4XL U2988 ( .D0(n3981), .D1(n3982), .D2(n3983), .D3(n3984), .S0(n3753), 
        .S1(n3756), .Y(n3980) );
  MUX4XL U2989 ( .D0(n3837), .D1(n3838), .D2(n3839), .D3(n3840), .S0(n3753), 
        .S1(n3757), .Y(n3836) );
  MUX2IXL U2990 ( .D0(A[221]), .D1(A[477]), .S(n3763), .Y(n3997) );
  MUX4XL U2991 ( .D0(A[254]), .D1(A[766]), .D2(A[510]), .D3(A[1022]), .S0(
        n3819), .S1(n3764), .Y(n3917) );
  INVX1 U2992 ( .A(n3827), .Y(n3815) );
  INVXL U2993 ( .A(n3655), .Y(n3763) );
  INVXL U2994 ( .A(n3655), .Y(n3764) );
  INVX1 U2995 ( .A(n3698), .Y(n3765) );
  INVX1 U2996 ( .A(n3743), .Y(n3736) );
  INVX1 U2997 ( .A(SH[4]), .Y(n3752) );
  INVX1 U2998 ( .A(SH[5]), .Y(n3755) );
  INVXL U2999 ( .A(SH[3]), .Y(n3745) );
  INVXL U3000 ( .A(n3833), .Y(n3826) );
  INVX1 U3001 ( .A(n3814), .Y(n3804) );
  INVX1 U3002 ( .A(n3814), .Y(n3803) );
  INVX1 U3003 ( .A(n3814), .Y(n3802) );
  INVXL U3004 ( .A(n3813), .Y(n3806) );
  INVXL U3005 ( .A(n3698), .Y(n3805) );
  INVXL U3006 ( .A(n3669), .Y(n3792) );
  INVXL U3007 ( .A(n3669), .Y(n3794) );
  INVXL U3008 ( .A(n3669), .Y(n3793) );
  INVX1 U3009 ( .A(n3765), .Y(n3797) );
  INVX1 U3010 ( .A(n3805), .Y(n3796) );
  INVXL U3011 ( .A(n3801), .Y(n3800) );
  INVX1 U3012 ( .A(n3801), .Y(n3798) );
  INVX1 U3013 ( .A(n3809), .Y(n3783) );
  INVX1 U3014 ( .A(n3809), .Y(n3782) );
  INVXL U3015 ( .A(n3770), .Y(n3814) );
  MUX2IXL U3016 ( .D0(A[235]), .D1(A[491]), .S(n3625), .Y(n4136) );
  MUX4XL U3017 ( .D0(n3895), .D1(n3896), .D2(n3897), .D3(n3898), .S0(n3622), 
        .S1(n3740), .Y(n3894) );
  MUX4XL U3018 ( .D0(A[47]), .D1(A[559]), .D2(A[303]), .D3(A[815]), .S0(n3622), 
        .S1(n3768), .Y(n3904) );
  MUX4XL U3019 ( .D0(A[175]), .D1(A[687]), .D2(A[431]), .D3(A[943]), .S0(n3623), .S1(n3765), .Y(n3858) );
  MUX4XL U3020 ( .D0(A[167]), .D1(A[679]), .D2(A[423]), .D3(A[935]), .S0(n3622), .S1(n3765), .Y(n3856) );
  MUX4XL U3021 ( .D0(A[40]), .D1(A[552]), .D2(A[296]), .D3(A[808]), .S0(n3670), 
        .S1(n3762), .Y(n4391) );
  MUX2X1 U3022 ( .D0(n3835), .D1(n3836), .S(SH[7]), .Y(B[7]) );
  MUX2IX1 U3023 ( .D0(n3841), .D1(n3842), .S(n3604), .Y(n3840) );
  MUX4X1 U3024 ( .D0(A[255]), .D1(A[767]), .D2(A[511]), .D3(A[1023]), .S0(
        n3815), .S1(n3767), .Y(n3844) );
  MUX4X1 U3025 ( .D0(A[247]), .D1(A[759]), .D2(A[503]), .D3(A[1015]), .S0(
        n3623), .S1(n3705), .Y(n3843) );
  NOR2X1 U3026 ( .A(A[999]), .B(n3796), .Y(n3847) );
  MUX2IX1 U3027 ( .D0(A[239]), .D1(A[495]), .S(n3626), .Y(n3846) );
  MUX2IX1 U3028 ( .D0(A[231]), .D1(A[487]), .S(n3627), .Y(n3845) );
  NOR2X1 U3029 ( .A(A[991]), .B(n3798), .Y(n3854) );
  MUX2IX1 U3030 ( .D0(A[223]), .D1(A[479]), .S(n3805), .Y(n3853) );
  NAND2X1 U3031 ( .A(n3855), .B(n3622), .Y(n3851) );
  MUX2IX1 U3032 ( .D0(A[719]), .D1(A[975]), .S(n3767), .Y(n3855) );
  NAND31X1 U3033 ( .C(A[983]), .A(n3802), .B(n3623), .Y(n3850) );
  NAND31X1 U3034 ( .C(A[967]), .A(n3770), .B(n3622), .Y(n3849) );
  MUX2IX1 U3035 ( .D0(n3860), .D1(n3861), .S(n3820), .Y(n3859) );
  MUX2IX1 U3036 ( .D0(A[191]), .D1(A[447]), .S(n3802), .Y(n3860) );
  MUX4X1 U3037 ( .D0(A[183]), .D1(A[695]), .D2(A[439]), .D3(A[951]), .S0(n3623), .S1(n3804), .Y(n3857) );
  MUX2IX1 U3038 ( .D0(n3862), .D1(n3863), .S(n3748), .Y(n3837) );
  MUX2IX1 U3039 ( .D0(A[671]), .D1(A[927]), .S(n3805), .Y(n3867) );
  NOR2X1 U3040 ( .A(A[415]), .B(n3796), .Y(n3866) );
  MUX2IX1 U3041 ( .D0(A[663]), .D1(A[919]), .S(n3802), .Y(n3865) );
  NOR2X1 U3042 ( .A(A[407]), .B(n3798), .Y(n3864) );
  MUX2IX1 U3043 ( .D0(n3868), .D1(n3869), .S(n3736), .Y(n3862) );
  NAND2X1 U3044 ( .A(n3870), .B(n3827), .Y(n3868) );
  MUX2IX1 U3045 ( .D0(A[135]), .D1(A[391]), .S(n3765), .Y(n3870) );
  MUX2IX1 U3046 ( .D0(n3871), .D1(n3872), .S(n3756), .Y(n3835) );
  MUX4X1 U3047 ( .D0(n3873), .D1(n3874), .D2(n3875), .D3(n3876), .S0(n3753), 
        .S1(n3602), .Y(n3872) );
  NOR2X1 U3048 ( .A(n3772), .B(A[639]), .Y(n3880) );
  MUX2IX1 U3049 ( .D0(A[127]), .D1(A[383]), .S(n3764), .Y(n3878) );
  NOR2X1 U3050 ( .A(A[375]), .B(n3796), .Y(n3877) );
  MUX2IX1 U3051 ( .D0(n3881), .D1(n3882), .S(n3736), .Y(n3875) );
  NOR2X1 U3052 ( .A(n3772), .B(A[607]), .Y(n3884) );
  NOR2X1 U3053 ( .A(A[351]), .B(n3793), .Y(n3883) );
  NOR2X1 U3054 ( .A(n3772), .B(A[623]), .Y(n3888) );
  NOR2X1 U3055 ( .A(A[367]), .B(n3792), .Y(n3887) );
  NOR2X1 U3056 ( .A(A[359]), .B(n3794), .Y(n3885) );
  MUX2X1 U3057 ( .D0(n3889), .D1(n3890), .S(n3741), .Y(n3873) );
  NOR3XL U3058 ( .A(n3826), .B(A[839]), .C(n3799), .Y(n3889) );
  MUX4X1 U3059 ( .D0(n3891), .D1(n3892), .D2(n3893), .D3(n3894), .S0(n3753), 
        .S1(n3750), .Y(n3871) );
  MUX2IX1 U3060 ( .D0(A[575]), .D1(A[831]), .S(n3767), .Y(n3898) );
  NOR2X1 U3061 ( .A(A[319]), .B(n3800), .Y(n3897) );
  MUX2IX1 U3062 ( .D0(A[567]), .D1(A[823]), .S(n3763), .Y(n3896) );
  NOR2X1 U3063 ( .A(A[311]), .B(n3796), .Y(n3895) );
  MUX2IX1 U3064 ( .D0(A[543]), .D1(A[799]), .S(n3774), .Y(n3902) );
  NOR2X1 U3065 ( .A(A[287]), .B(n3800), .Y(n3901) );
  MUX2IX1 U3066 ( .D0(A[535]), .D1(A[791]), .S(n3805), .Y(n3900) );
  NOR2X1 U3067 ( .A(A[279]), .B(n3793), .Y(n3899) );
  MUX2IX1 U3068 ( .D0(n3903), .D1(n3904), .S(n3736), .Y(n3892) );
  MUX2IX1 U3069 ( .D0(A[527]), .D1(A[783]), .S(n3805), .Y(n3907) );
  NOR2X1 U3070 ( .A(A[271]), .B(n3792), .Y(n3906) );
  MUX2X1 U3071 ( .D0(n3908), .D1(n3909), .S(SH[7]), .Y(B[6]) );
  MUX4X1 U3072 ( .D0(n3910), .D1(n3911), .D2(n3912), .D3(n3913), .S0(n3753), 
        .S1(n3757), .Y(n3909) );
  MUX2IX1 U3073 ( .D0(n3914), .D1(n3915), .S(n3604), .Y(n3913) );
  MUX2IX1 U3074 ( .D0(n3916), .D1(n3917), .S(n3736), .Y(n3915) );
  NOR2X1 U3075 ( .A(A[1006]), .B(n3797), .Y(n3921) );
  NOR2X1 U3076 ( .A(A[998]), .B(n3800), .Y(n3920) );
  MUX2IX1 U3077 ( .D0(A[238]), .D1(A[494]), .S(n3805), .Y(n3919) );
  MUX2IX1 U3078 ( .D0(A[230]), .D1(A[486]), .S(n3767), .Y(n3918) );
  MUX2IX1 U3079 ( .D0(n3926), .D1(n3927), .S(n3820), .Y(n3925) );
  NOR2X1 U3080 ( .A(A[990]), .B(n3793), .Y(n3927) );
  MUX2IX1 U3081 ( .D0(A[222]), .D1(A[478]), .S(n3805), .Y(n3926) );
  NAND2X1 U3082 ( .A(n3928), .B(n3622), .Y(n3924) );
  MUX2IX1 U3083 ( .D0(A[718]), .D1(A[974]), .S(n3804), .Y(n3928) );
  NAND31X1 U3084 ( .C(A[982]), .A(n3666), .B(n3622), .Y(n3923) );
  NAND31X1 U3085 ( .C(A[966]), .A(n3666), .B(n3623), .Y(n3922) );
  NOR2X1 U3086 ( .A(n3617), .B(A[702]), .Y(n3934) );
  MUX2IX1 U3087 ( .D0(A[190]), .D1(A[446]), .S(n3763), .Y(n3933) );
  MUX2IX1 U3088 ( .D0(n3935), .D1(n3936), .S(n3748), .Y(n3910) );
  MUX2IX1 U3089 ( .D0(A[670]), .D1(A[926]), .S(n3765), .Y(n3940) );
  NOR2X1 U3090 ( .A(A[414]), .B(n3792), .Y(n3939) );
  MUX2IX1 U3091 ( .D0(A[662]), .D1(A[918]), .S(n3803), .Y(n3938) );
  NOR2X1 U3092 ( .A(A[406]), .B(n3792), .Y(n3937) );
  MUX2IX1 U3093 ( .D0(n3941), .D1(n3942), .S(n3736), .Y(n3935) );
  NAND2X1 U3094 ( .A(n3943), .B(n3827), .Y(n3941) );
  MUX2IX1 U3095 ( .D0(n3944), .D1(n3945), .S(n3756), .Y(n3908) );
  MUX4X1 U3096 ( .D0(n3946), .D1(n3947), .D2(n3948), .D3(n3949), .S0(n3753), 
        .S1(n3750), .Y(n3945) );
  MUX2IX1 U3097 ( .D0(A[126]), .D1(A[382]), .S(n3764), .Y(n3951) );
  NOR2X1 U3098 ( .A(A[374]), .B(n3793), .Y(n3950) );
  MUX2IX1 U3099 ( .D0(n3954), .D1(n3955), .S(n3736), .Y(n3948) );
  NOR2X1 U3100 ( .A(A[350]), .B(n3792), .Y(n3956) );
  NOR2X1 U3101 ( .A(A[358]), .B(n3698), .Y(n3958) );
  MUX2X1 U3102 ( .D0(n3961), .D1(n3890), .S(n3741), .Y(n3946) );
  NOR3XL U3103 ( .A(n3826), .B(A[838]), .C(n3800), .Y(n3961) );
  MUX4X1 U3104 ( .D0(n3962), .D1(n3963), .D2(n3964), .D3(n3965), .S0(n3753), 
        .S1(n3750), .Y(n3944) );
  MUX2IX1 U3105 ( .D0(A[574]), .D1(A[830]), .S(n3804), .Y(n3969) );
  NOR2X1 U3106 ( .A(A[318]), .B(n3800), .Y(n3968) );
  MUX2IX1 U3107 ( .D0(A[566]), .D1(A[822]), .S(n3802), .Y(n3967) );
  NOR2X1 U3108 ( .A(A[310]), .B(n3794), .Y(n3966) );
  MUX2IX1 U3109 ( .D0(A[542]), .D1(A[798]), .S(n3765), .Y(n3973) );
  NOR2X1 U3110 ( .A(A[286]), .B(n3794), .Y(n3972) );
  MUX2IX1 U3111 ( .D0(A[534]), .D1(A[790]), .S(n3805), .Y(n3971) );
  NOR2X1 U3112 ( .A(A[278]), .B(n3793), .Y(n3970) );
  MUX2IX1 U3113 ( .D0(n3974), .D1(n3975), .S(n3736), .Y(n3963) );
  NOR2X1 U3114 ( .A(n3742), .B(n3976), .Y(n3962) );
  MUX2IX1 U3115 ( .D0(n3977), .D1(n3978), .S(n3727), .Y(n3976) );
  MUX2IX1 U3116 ( .D0(A[526]), .D1(A[782]), .S(n3802), .Y(n3978) );
  NOR2X1 U3117 ( .A(A[270]), .B(n3800), .Y(n3977) );
  MUX2X1 U3118 ( .D0(n3979), .D1(n3980), .S(SH[7]), .Y(B[5]) );
  MUX2IX1 U3119 ( .D0(n3985), .D1(n3986), .S(n3604), .Y(n3984) );
  MUX2IX1 U3120 ( .D0(n3987), .D1(n3988), .S(n3606), .Y(n3986) );
  NOR2X1 U3121 ( .A(A[1005]), .B(n3698), .Y(n3992) );
  NOR2X1 U3122 ( .A(A[997]), .B(n3800), .Y(n3991) );
  MUX2IX1 U3123 ( .D0(A[237]), .D1(A[493]), .S(n3764), .Y(n3990) );
  MUX2IX1 U3124 ( .D0(A[229]), .D1(A[485]), .S(n3625), .Y(n3989) );
  NOR2X1 U3125 ( .A(A[989]), .B(n3797), .Y(n3998) );
  NAND2X1 U3126 ( .A(n3999), .B(n3623), .Y(n3995) );
  MUX2IX1 U3127 ( .D0(A[717]), .D1(A[973]), .S(n3803), .Y(n3999) );
  NOR2X1 U3128 ( .A(n3617), .B(A[701]), .Y(n4005) );
  MUX2IX1 U3129 ( .D0(A[189]), .D1(A[445]), .S(n3767), .Y(n4004) );
  MUX4X1 U3130 ( .D0(A[173]), .D1(A[685]), .D2(A[429]), .D3(A[941]), .S0(n3618), .S1(n3768), .Y(n4002) );
  MUX4X1 U3131 ( .D0(A[165]), .D1(A[677]), .D2(A[421]), .D3(A[933]), .S0(n3619), .S1(n3705), .Y(n4000) );
  MUX2IX1 U3132 ( .D0(n4006), .D1(n4007), .S(n3748), .Y(n3981) );
  MUX4X1 U3133 ( .D0(n4008), .D1(n4009), .D2(n4010), .D3(n4011), .S0(n3619), 
        .S1(n3737), .Y(n4007) );
  MUX2IX1 U3134 ( .D0(A[669]), .D1(A[925]), .S(n3764), .Y(n4011) );
  NOR2X1 U3135 ( .A(A[413]), .B(n3800), .Y(n4010) );
  MUX2IX1 U3136 ( .D0(A[661]), .D1(A[917]), .S(n3627), .Y(n4009) );
  NOR2X1 U3137 ( .A(A[405]), .B(n3797), .Y(n4008) );
  MUX2IX1 U3138 ( .D0(n4012), .D1(n4013), .S(n3736), .Y(n4006) );
  NAND2X1 U3139 ( .A(n4014), .B(n3826), .Y(n4012) );
  MUX2IX1 U3140 ( .D0(A[133]), .D1(A[389]), .S(n3764), .Y(n4014) );
  MUX2IX1 U3141 ( .D0(n4015), .D1(n4016), .S(n3756), .Y(n3979) );
  MUX4X1 U3142 ( .D0(n4017), .D1(n4018), .D2(n4019), .D3(n4020), .S0(n3753), 
        .S1(n3750), .Y(n4016) );
  MUX2IX1 U3143 ( .D0(A[125]), .D1(A[381]), .S(n3625), .Y(n4022) );
  NOR2X1 U3144 ( .A(A[373]), .B(n3796), .Y(n4021) );
  MUX2IX1 U3145 ( .D0(n4025), .D1(n4026), .S(n3736), .Y(n4019) );
  MUX2IX1 U3146 ( .D0(n4027), .D1(n4028), .S(n3820), .Y(n4026) );
  NOR2X1 U3147 ( .A(A[349]), .B(n3797), .Y(n4027) );
  MUX4X1 U3148 ( .D0(n4029), .D1(n4030), .D2(n4031), .D3(n4032), .S0(n3817), 
        .S1(n3737), .Y(n4018) );
  NOR2X1 U3149 ( .A(n3773), .B(A[621]), .Y(n4032) );
  NOR2X1 U3150 ( .A(A[365]), .B(n3797), .Y(n4031) );
  NOR2X1 U3151 ( .A(n3763), .B(A[613]), .Y(n4030) );
  NOR2X1 U3152 ( .A(A[357]), .B(n3793), .Y(n4029) );
  MUX2X1 U3153 ( .D0(n4033), .D1(n4034), .S(n3732), .Y(n4017) );
  NOR3XL U3154 ( .A(n3826), .B(n3776), .C(A[589]), .Y(n4034) );
  NOR3XL U3155 ( .A(n3831), .B(A[837]), .C(n3799), .Y(n4033) );
  MUX4X1 U3156 ( .D0(n4035), .D1(n4036), .D2(n4037), .D3(n4038), .S0(n3753), 
        .S1(n3750), .Y(n4015) );
  MUX4X1 U3157 ( .D0(n4039), .D1(n4040), .D2(n4041), .D3(n4042), .S0(n3618), 
        .S1(n3736), .Y(n4038) );
  MUX2IX1 U3158 ( .D0(A[573]), .D1(A[829]), .S(n3763), .Y(n4042) );
  NOR2X1 U3159 ( .A(A[317]), .B(n3794), .Y(n4041) );
  MUX2IX1 U3160 ( .D0(A[565]), .D1(A[821]), .S(n3625), .Y(n4040) );
  NOR2X1 U3161 ( .A(A[309]), .B(n3792), .Y(n4039) );
  MUX2IX1 U3162 ( .D0(A[541]), .D1(A[797]), .S(n3627), .Y(n4046) );
  NOR2X1 U3163 ( .A(A[285]), .B(n3796), .Y(n4045) );
  MUX2IX1 U3164 ( .D0(A[533]), .D1(A[789]), .S(n3626), .Y(n4044) );
  NOR2X1 U3165 ( .A(A[277]), .B(n3797), .Y(n4043) );
  MUX2IX1 U3166 ( .D0(n4047), .D1(n4048), .S(n3606), .Y(n4036) );
  NOR2X1 U3167 ( .A(n3745), .B(n4049), .Y(n4035) );
  MUX2IX1 U3168 ( .D0(n4050), .D1(n4051), .S(n3820), .Y(n4049) );
  MUX2IX1 U3169 ( .D0(A[525]), .D1(A[781]), .S(n3625), .Y(n4051) );
  NOR2X1 U3170 ( .A(A[269]), .B(n3796), .Y(n4050) );
  MUX2X1 U3171 ( .D0(n4052), .D1(n4053), .S(SH[7]), .Y(B[4]) );
  MUX2IX1 U3172 ( .D0(n4058), .D1(n4059), .S(n3748), .Y(n4057) );
  MUX2IX1 U3173 ( .D0(n4060), .D1(n4061), .S(n3606), .Y(n4059) );
  NOR2X1 U3174 ( .A(A[1004]), .B(n3797), .Y(n4065) );
  NOR2X1 U3175 ( .A(A[996]), .B(n3797), .Y(n4064) );
  MUX2IX1 U3176 ( .D0(A[236]), .D1(A[492]), .S(n3626), .Y(n4063) );
  MUX2IX1 U3177 ( .D0(A[228]), .D1(A[484]), .S(n3625), .Y(n4062) );
  MUX2IX1 U3178 ( .D0(n4070), .D1(n4071), .S(n3820), .Y(n4069) );
  NOR2X1 U3179 ( .A(A[988]), .B(n3796), .Y(n4071) );
  MUX2IX1 U3180 ( .D0(A[220]), .D1(A[476]), .S(n3625), .Y(n4070) );
  NAND2X1 U3181 ( .A(n4072), .B(n3623), .Y(n4068) );
  MUX2IX1 U3182 ( .D0(A[716]), .D1(A[972]), .S(n3763), .Y(n4072) );
  MUX2IX1 U3183 ( .D0(n4077), .D1(n4078), .S(n3820), .Y(n4076) );
  MUX2IX1 U3184 ( .D0(A[188]), .D1(A[444]), .S(n3764), .Y(n4077) );
  MUX4X1 U3185 ( .D0(A[172]), .D1(A[684]), .D2(A[428]), .D3(A[940]), .S0(n3728), .S1(n3627), .Y(n4075) );
  MUX4X1 U3186 ( .D0(A[180]), .D1(A[692]), .D2(A[436]), .D3(A[948]), .S0(n3728), .S1(n3764), .Y(n4074) );
  MUX4X1 U3187 ( .D0(A[164]), .D1(A[676]), .D2(A[420]), .D3(A[932]), .S0(n3728), .S1(n3626), .Y(n4073) );
  MUX2IX1 U3188 ( .D0(n4079), .D1(n4080), .S(n3748), .Y(n4054) );
  MUX4X1 U3189 ( .D0(n4081), .D1(n4082), .D2(n4083), .D3(n4084), .S0(n3728), 
        .S1(n3738), .Y(n4080) );
  MUX2IX1 U3190 ( .D0(A[668]), .D1(A[924]), .S(n3625), .Y(n4084) );
  NOR2X1 U3191 ( .A(A[412]), .B(n3797), .Y(n4083) );
  MUX2IX1 U3192 ( .D0(A[660]), .D1(A[916]), .S(n3626), .Y(n4082) );
  NOR2X1 U3193 ( .A(A[404]), .B(n3796), .Y(n4081) );
  MUX2IX1 U3194 ( .D0(n4085), .D1(n4086), .S(n3606), .Y(n4079) );
  MUX4X1 U3195 ( .D0(A[140]), .D1(A[652]), .D2(A[396]), .D3(A[908]), .S0(n3728), .S1(n3626), .Y(n4086) );
  NAND2X1 U3196 ( .A(n4087), .B(n3826), .Y(n4085) );
  MUX2IX1 U3197 ( .D0(A[132]), .D1(A[388]), .S(n3763), .Y(n4087) );
  MUX2IX1 U3198 ( .D0(n4088), .D1(n4089), .S(n3756), .Y(n4052) );
  MUX4X1 U3199 ( .D0(n4090), .D1(n4091), .D2(n4092), .D3(n4093), .S0(n3754), 
        .S1(n3750), .Y(n4089) );
  MUX2IX1 U3200 ( .D0(A[124]), .D1(A[380]), .S(n3627), .Y(n4095) );
  NOR2X1 U3201 ( .A(A[372]), .B(n3797), .Y(n4094) );
  MUX2IX1 U3202 ( .D0(n4098), .D1(n4099), .S(n3606), .Y(n4092) );
  MUX2IX1 U3203 ( .D0(n4100), .D1(n4101), .S(n3820), .Y(n4099) );
  NOR2X1 U3204 ( .A(A[348]), .B(n3796), .Y(n4100) );
  MUX4X1 U3205 ( .D0(n4102), .D1(n4103), .D2(n4104), .D3(n4105), .S0(n3728), 
        .S1(n3737), .Y(n4091) );
  NOR2X1 U3206 ( .A(A[364]), .B(n3698), .Y(n4104) );
  NOR2X1 U3207 ( .A(A[356]), .B(n3698), .Y(n4102) );
  MUX2X1 U3208 ( .D0(n4106), .D1(n4107), .S(n3732), .Y(n4090) );
  NOR3XL U3209 ( .A(n3826), .B(n3776), .C(A[588]), .Y(n4107) );
  NOR3XL U3210 ( .A(n3831), .B(A[836]), .C(n3799), .Y(n4106) );
  MUX4X1 U3211 ( .D0(n4108), .D1(n4109), .D2(n4110), .D3(n4111), .S0(n3754), 
        .S1(n3750), .Y(n4088) );
  MUX4X1 U3212 ( .D0(n4112), .D1(n4113), .D2(n4114), .D3(n4115), .S0(n3728), 
        .S1(n3737), .Y(n4111) );
  MUX2IX1 U3213 ( .D0(A[572]), .D1(A[828]), .S(n3764), .Y(n4115) );
  NOR2X1 U3214 ( .A(A[316]), .B(n3698), .Y(n4114) );
  MUX2IX1 U3215 ( .D0(A[564]), .D1(A[820]), .S(n3627), .Y(n4113) );
  MUX4X1 U3216 ( .D0(n4116), .D1(n4117), .D2(n4118), .D3(n4119), .S0(n3816), 
        .S1(n3737), .Y(n4110) );
  MUX2IX1 U3217 ( .D0(A[540]), .D1(A[796]), .S(n3627), .Y(n4119) );
  MUX2IX1 U3218 ( .D0(A[532]), .D1(A[788]), .S(n3625), .Y(n4117) );
  MUX2IX1 U3219 ( .D0(n4120), .D1(n4121), .S(n3606), .Y(n4109) );
  MUX4X1 U3220 ( .D0(A[44]), .D1(A[556]), .D2(A[300]), .D3(A[812]), .S0(n3816), 
        .S1(n3705), .Y(n4121) );
  MUX4X1 U3221 ( .D0(A[36]), .D1(A[548]), .D2(A[292]), .D3(A[804]), .S0(n3816), 
        .S1(n3765), .Y(n4120) );
  NOR2X1 U3222 ( .A(n3745), .B(n4122), .Y(n4108) );
  MUX2IX1 U3223 ( .D0(n4123), .D1(n4124), .S(n3820), .Y(n4122) );
  MUX2IX1 U3224 ( .D0(A[524]), .D1(A[780]), .S(n3626), .Y(n4124) );
  NOR2X1 U3225 ( .A(A[268]), .B(n3794), .Y(n4123) );
  MUX2X1 U3226 ( .D0(n4125), .D1(n4126), .S(SH[7]), .Y(B[3]) );
  MUX4X1 U3227 ( .D0(n4127), .D1(n4128), .D2(n4129), .D3(n4130), .S0(n3754), 
        .S1(n3757), .Y(n4126) );
  MUX2IX1 U3228 ( .D0(n4131), .D1(n4132), .S(n3748), .Y(n4130) );
  MUX2IX1 U3229 ( .D0(n4133), .D1(n4134), .S(n3606), .Y(n4132) );
  MUX4X1 U3230 ( .D0(A[243]), .D1(A[755]), .D2(A[499]), .D3(A[1011]), .S0(
        n3816), .S1(n3705), .Y(n4133) );
  NOR2X1 U3231 ( .A(A[1003]), .B(n3794), .Y(n4138) );
  NOR2X1 U3232 ( .A(A[995]), .B(n3794), .Y(n4137) );
  MUX2IX1 U3233 ( .D0(A[227]), .D1(A[483]), .S(n3625), .Y(n4135) );
  MUX4X1 U3234 ( .D0(n4139), .D1(n4140), .D2(n4141), .D3(n4142), .S0(n3604), 
        .S1(n3737), .Y(n4129) );
  MUX2IX1 U3235 ( .D0(n4143), .D1(n4144), .S(n3820), .Y(n4142) );
  NOR2X1 U3236 ( .A(A[987]), .B(n3794), .Y(n4144) );
  NAND2X1 U3237 ( .A(n4145), .B(n3824), .Y(n4141) );
  NAND31X1 U3238 ( .C(A[979]), .A(n3770), .B(n3823), .Y(n4140) );
  MUX4X1 U3239 ( .D0(n4146), .D1(n4147), .D2(n4148), .D3(n4149), .S0(n3604), 
        .S1(n3738), .Y(n4128) );
  MUX2IX1 U3240 ( .D0(n4150), .D1(n4151), .S(n3820), .Y(n4149) );
  MUX2IX1 U3241 ( .D0(A[187]), .D1(A[443]), .S(n3627), .Y(n4150) );
  MUX4X1 U3242 ( .D0(A[171]), .D1(A[683]), .D2(A[427]), .D3(A[939]), .S0(n3815), .S1(n3803), .Y(n4148) );
  MUX4X1 U3243 ( .D0(A[179]), .D1(A[691]), .D2(A[435]), .D3(A[947]), .S0(n3815), .S1(n3804), .Y(n4147) );
  MUX4X1 U3244 ( .D0(A[163]), .D1(A[675]), .D2(A[419]), .D3(A[931]), .S0(n3815), .S1(n3767), .Y(n4146) );
  MUX2IX1 U3245 ( .D0(n4152), .D1(n4153), .S(n3748), .Y(n4127) );
  MUX4X1 U3246 ( .D0(n4154), .D1(n4155), .D2(n4156), .D3(n4157), .S0(n3815), 
        .S1(n3737), .Y(n4153) );
  MUX2IX1 U3247 ( .D0(A[667]), .D1(A[923]), .S(n3761), .Y(n4157) );
  NOR2X1 U3248 ( .A(A[411]), .B(n3793), .Y(n4156) );
  NOR2X1 U3249 ( .A(A[403]), .B(n3793), .Y(n4154) );
  MUX2IX1 U3250 ( .D0(n4158), .D1(n4159), .S(n3606), .Y(n4152) );
  MUX4X1 U3251 ( .D0(A[139]), .D1(A[651]), .D2(A[395]), .D3(A[907]), .S0(n3815), .S1(n3767), .Y(n4159) );
  NAND2X1 U3252 ( .A(n4160), .B(n3826), .Y(n4158) );
  MUX2IX1 U3253 ( .D0(n4161), .D1(n4162), .S(n3756), .Y(n4125) );
  MUX4X1 U3254 ( .D0(n4163), .D1(n4164), .D2(n4165), .D3(n4166), .S0(n3754), 
        .S1(n3750), .Y(n4162) );
  NOR2X1 U3255 ( .A(n3772), .B(A[635]), .Y(n4170) );
  NOR2X1 U3256 ( .A(n3772), .B(A[627]), .Y(n4169) );
  MUX2IX1 U3257 ( .D0(A[123]), .D1(A[379]), .S(n3761), .Y(n4168) );
  NOR2X1 U3258 ( .A(A[371]), .B(n3793), .Y(n4167) );
  MUX2IX1 U3259 ( .D0(n4171), .D1(n4172), .S(n3734), .Y(n4165) );
  MUX2IX1 U3260 ( .D0(n4173), .D1(n4174), .S(n3727), .Y(n4172) );
  NOR2X1 U3261 ( .A(n3773), .B(A[603]), .Y(n4174) );
  NOR2X1 U3262 ( .A(A[347]), .B(n3793), .Y(n4173) );
  MUX4X1 U3263 ( .D0(n4175), .D1(n4176), .D2(n4177), .D3(n4178), .S0(n3815), 
        .S1(n3738), .Y(n4164) );
  NOR2X1 U3264 ( .A(n3705), .B(A[619]), .Y(n4178) );
  NOR2X1 U3265 ( .A(A[363]), .B(n3792), .Y(n4177) );
  NOR2X1 U3266 ( .A(n3773), .B(A[611]), .Y(n4176) );
  NOR2X1 U3267 ( .A(A[355]), .B(n3792), .Y(n4175) );
  MUX2X1 U3268 ( .D0(n4179), .D1(n4180), .S(n3741), .Y(n4163) );
  NOR3XL U3269 ( .A(n3832), .B(n3776), .C(A[587]), .Y(n4180) );
  NOR3XL U3270 ( .A(n3831), .B(A[835]), .C(n3798), .Y(n4179) );
  MUX4X1 U3271 ( .D0(n4181), .D1(n4182), .D2(n4183), .D3(n4184), .S0(n3754), 
        .S1(n3602), .Y(n4161) );
  MUX4X1 U3272 ( .D0(n4185), .D1(n4186), .D2(n4187), .D3(n4188), .S0(n3815), 
        .S1(n3738), .Y(n4184) );
  MUX2IX1 U3273 ( .D0(A[571]), .D1(A[827]), .S(n3761), .Y(n4188) );
  NOR2X1 U3274 ( .A(A[315]), .B(n3792), .Y(n4187) );
  NOR2X1 U3275 ( .A(A[307]), .B(n3792), .Y(n4185) );
  MUX2IX1 U3276 ( .D0(A[539]), .D1(A[795]), .S(n3761), .Y(n4192) );
  NOR2X1 U3277 ( .A(A[283]), .B(n3791), .Y(n4191) );
  MUX2IX1 U3278 ( .D0(A[531]), .D1(A[787]), .S(n3761), .Y(n4190) );
  NOR2X1 U3279 ( .A(A[275]), .B(n3791), .Y(n4189) );
  MUX2IX1 U3280 ( .D0(n4193), .D1(n4194), .S(n3734), .Y(n4182) );
  NOR2X1 U3281 ( .A(n3745), .B(n4195), .Y(n4181) );
  MUX2IX1 U3282 ( .D0(n4196), .D1(n4197), .S(n3727), .Y(n4195) );
  MUX2IX1 U3283 ( .D0(A[523]), .D1(A[779]), .S(n3761), .Y(n4197) );
  NOR2X1 U3284 ( .A(A[267]), .B(n3791), .Y(n4196) );
  MUX4X1 U3285 ( .D0(n4200), .D1(n4201), .D2(n4202), .D3(n4203), .S0(n3754), 
        .S1(n3757), .Y(n4199) );
  MUX2IX1 U3286 ( .D0(n4204), .D1(n4205), .S(n3602), .Y(n4203) );
  MUX2IX1 U3287 ( .D0(n4206), .D1(n4207), .S(n3606), .Y(n4205) );
  NOR2X1 U3288 ( .A(A[1002]), .B(n3791), .Y(n4211) );
  NOR2X1 U3289 ( .A(A[994]), .B(n3790), .Y(n4210) );
  MUX2IX1 U3290 ( .D0(A[234]), .D1(A[490]), .S(n3761), .Y(n4209) );
  MUX2IX1 U3291 ( .D0(A[226]), .D1(A[482]), .S(n3760), .Y(n4208) );
  MUX4X1 U3292 ( .D0(n4212), .D1(n4213), .D2(n4214), .D3(n4215), .S0(n3604), 
        .S1(n3739), .Y(n4202) );
  MUX2IX1 U3293 ( .D0(n4216), .D1(n4217), .S(n3707), .Y(n4215) );
  NOR2X1 U3294 ( .A(A[986]), .B(n3790), .Y(n4217) );
  NAND2X1 U3295 ( .A(n4218), .B(n3824), .Y(n4214) );
  MUX4X1 U3296 ( .D0(n4219), .D1(n4220), .D2(n4221), .D3(n4222), .S0(n3604), 
        .S1(n3738), .Y(n4201) );
  MUX2IX1 U3297 ( .D0(n4223), .D1(n4224), .S(n3727), .Y(n4222) );
  NOR2X1 U3298 ( .A(n3617), .B(A[698]), .Y(n4224) );
  MUX2IX1 U3299 ( .D0(A[186]), .D1(A[442]), .S(n3760), .Y(n4223) );
  MUX4X1 U3300 ( .D0(A[170]), .D1(A[682]), .D2(A[426]), .D3(A[938]), .S0(n3707), .S1(n3768), .Y(n4221) );
  MUX2IX1 U3301 ( .D0(n4225), .D1(n4226), .S(n3602), .Y(n4200) );
  MUX4X1 U3302 ( .D0(n4227), .D1(n4228), .D2(n4229), .D3(n4230), .S0(n3728), 
        .S1(n3739), .Y(n4226) );
  MUX2IX1 U3303 ( .D0(A[666]), .D1(A[922]), .S(n3614), .Y(n4230) );
  NOR2X1 U3304 ( .A(A[410]), .B(n3790), .Y(n4229) );
  MUX2IX1 U3305 ( .D0(A[658]), .D1(A[914]), .S(n3760), .Y(n4228) );
  NOR2X1 U3306 ( .A(A[402]), .B(n3790), .Y(n4227) );
  MUX2IX1 U3307 ( .D0(n4231), .D1(n4232), .S(n3734), .Y(n4225) );
  MUX4X1 U3308 ( .D0(A[138]), .D1(A[650]), .D2(A[394]), .D3(A[906]), .S0(n3728), .S1(n3769), .Y(n4232) );
  NAND2X1 U3309 ( .A(n4233), .B(n3825), .Y(n4231) );
  MUX2IX1 U3310 ( .D0(n4234), .D1(n4235), .S(n3756), .Y(n4198) );
  NOR2X1 U3311 ( .A(A[370]), .B(n3789), .Y(n4236) );
  MUX2IX1 U3312 ( .D0(n4242), .D1(n4243), .S(n3690), .Y(n4241) );
  NOR2X1 U3313 ( .A(n3766), .B(A[602]), .Y(n4243) );
  NOR2X1 U3314 ( .A(A[346]), .B(n3789), .Y(n4242) );
  NOR2X1 U3315 ( .A(n3617), .B(A[618]), .Y(n4247) );
  NOR2X1 U3316 ( .A(A[362]), .B(n3789), .Y(n4246) );
  NOR2X1 U3317 ( .A(n3616), .B(A[610]), .Y(n4245) );
  NOR2X1 U3318 ( .A(A[354]), .B(n3789), .Y(n4244) );
  NOR3XL U3319 ( .A(n3831), .B(n3776), .C(A[586]), .Y(n4249) );
  NOR3XL U3320 ( .A(n3832), .B(A[834]), .C(n3798), .Y(n4248) );
  MUX2IX1 U3321 ( .D0(n4258), .D1(n4259), .S(n3734), .Y(n4251) );
  MUX4X1 U3322 ( .D0(A[42]), .D1(A[554]), .D2(A[298]), .D3(A[810]), .S0(n3690), 
        .S1(n3770), .Y(n4259) );
  MUX4X1 U3323 ( .D0(A[34]), .D1(A[546]), .D2(A[290]), .D3(A[802]), .S0(n3690), 
        .S1(n3770), .Y(n4258) );
  NOR2X1 U3324 ( .A(n3745), .B(n4260), .Y(n4250) );
  MUX2IX1 U3325 ( .D0(n4261), .D1(n4262), .S(n3727), .Y(n4260) );
  MUX2IX1 U3326 ( .D0(A[522]), .D1(A[778]), .S(n3759), .Y(n4262) );
  NOR2X1 U3327 ( .A(A[266]), .B(n3787), .Y(n4261) );
  MUX2IX1 U3328 ( .D0(n4269), .D1(n4270), .S(n3748), .Y(n4268) );
  MUX2IX1 U3329 ( .D0(n4271), .D1(n4272), .S(n3734), .Y(n4270) );
  NOR2X1 U3330 ( .A(A[1001]), .B(n3787), .Y(n4276) );
  NOR2X1 U3331 ( .A(A[993]), .B(n3787), .Y(n4275) );
  MUX2IX1 U3332 ( .D0(A[225]), .D1(A[481]), .S(n3769), .Y(n4273) );
  MUX2IX1 U3333 ( .D0(n4281), .D1(n4282), .S(n3822), .Y(n4280) );
  NOR2X1 U3334 ( .A(A[985]), .B(n3787), .Y(n4282) );
  NAND2X1 U3335 ( .A(n4283), .B(n3833), .Y(n4279) );
  NAND31X1 U3336 ( .C(A[961]), .A(n3769), .B(n3823), .Y(n4277) );
  MUX4X1 U3337 ( .D0(n4284), .D1(n4285), .D2(n4286), .D3(n4287), .S0(n3746), 
        .S1(n3739), .Y(n4266) );
  MUX2IX1 U3338 ( .D0(n4288), .D1(n4289), .S(n3833), .Y(n4287) );
  NOR2X1 U3339 ( .A(n3616), .B(A[697]), .Y(n4289) );
  MUX4X1 U3340 ( .D0(A[169]), .D1(A[681]), .D2(A[425]), .D3(A[937]), .S0(n3818), .S1(n3711), .Y(n4286) );
  MUX2IX1 U3341 ( .D0(A[665]), .D1(A[921]), .S(n3769), .Y(n4295) );
  MUX2IX1 U3342 ( .D0(n4296), .D1(n4297), .S(n3734), .Y(n4290) );
  NAND2X1 U3343 ( .A(n4298), .B(n3825), .Y(n4296) );
  MUX2IX1 U3344 ( .D0(A[129]), .D1(A[385]), .S(n3711), .Y(n4298) );
  NOR2X1 U3345 ( .A(n3771), .B(A[625]), .Y(n4307) );
  MUX2IX1 U3346 ( .D0(n4309), .D1(n4310), .S(n3734), .Y(n4303) );
  NOR2X1 U3347 ( .A(n3773), .B(A[601]), .Y(n4312) );
  MUX2X1 U3348 ( .D0(n4317), .D1(n4318), .S(n3741), .Y(n4301) );
  NOR3XL U3349 ( .A(n3832), .B(n3776), .C(A[585]), .Y(n4318) );
  NOR3XL U3350 ( .A(n3832), .B(A[833]), .C(n3799), .Y(n4317) );
  NOR2X1 U3351 ( .A(A[313]), .B(n3785), .Y(n4321) );
  MUX2IX1 U3352 ( .D0(A[537]), .D1(A[793]), .S(n3700), .Y(n4326) );
  MUX2IX1 U3353 ( .D0(A[529]), .D1(A[785]), .S(n3762), .Y(n4324) );
  MUX2IX1 U3354 ( .D0(n4330), .D1(n4331), .S(n3727), .Y(n4329) );
  NOR2X1 U3355 ( .A(A[265]), .B(n3791), .Y(n4330) );
  NAND2X1 U3356 ( .A(n4359), .B(n3825), .Y(n4357) );
  MUX4X1 U3357 ( .D0(n4364), .D1(n4365), .D2(n4366), .D3(n4367), .S0(n3732), 
        .S1(n3823), .Y(n4363) );
  MUX2IX1 U3358 ( .D0(n4370), .D1(n4371), .S(n3833), .Y(n4369) );
  NOR2X1 U3359 ( .A(A[344]), .B(n3783), .Y(n4370) );
  NAND32X1 U3360 ( .B(A[592]), .C(n3769), .A(n3824), .Y(n4368) );
  NOR2X1 U3361 ( .A(A[312]), .B(n3782), .Y(n4384) );
  NOR2X1 U3362 ( .A(A[280]), .B(n3782), .Y(n4388) );
  MUX2IX1 U3363 ( .D0(n4390), .D1(n4391), .S(n3605), .Y(n4379) );
  NOR2X1 U3364 ( .A(n3745), .B(n4392), .Y(n4378) );
  NOR2X1 U3365 ( .A(A[264]), .B(n3795), .Y(n4393) );
endmodule


module regbank_a0_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module regbank_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regbank_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regbank_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_50 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10838;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_50 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10838), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10838), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10838), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10838), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10838), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10838), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10838), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10838), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10838), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_51 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10856;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_51 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10856), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10856), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10856), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10856), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10856), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10856), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10856), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10856), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10856), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_52 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10874;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_52 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10874), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10874), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10874), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10874), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10874), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10874), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10874), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10874), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10874), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_53 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10892;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_53 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10892), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10892), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10892), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10892), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10892), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10892), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10892), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10892), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10892), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_54 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10910;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_54 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10910), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10910), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10910), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10910), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10910), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10910), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10910), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10910), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10910), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_0000001f ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10928;

  SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10928), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10928), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10928), .XR(arstz), .Q(rdat[6]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10928), .XS(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10928), .XR(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10928), .XS(arstz), .Q(rdat[3]) );
  DFFSQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10928), .XS(arstz), .Q(rdat[2]) );
  DFFSQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10928), .XS(arstz), .Q(rdat[1]) );
  DFFSQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10928), .XS(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000004 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10946;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10946), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10946), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10946), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10946), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10946), .XR(arstz), .Q(rdat[4]) );
  DFFSQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10946), .XS(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10946), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10946), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10946), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_4_00000004 ( clk, arstz, we, wdat, rdat );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we;
  wire   net10964;

  SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10964), .TE(1'b0) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10964), .XR(arstz), .Q(rdat[3]) );
  DFFSQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10964), .XS(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10964), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10964), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH7_2 ( clk, arstz, we, wdat, rdat );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we;
  wire   net10982;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10982), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10982), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10982), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10982), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10982), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10982), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10982), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10982), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_55 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11000;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_55 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11000), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11000), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11000), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11000), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11000), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11000), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11000), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11000), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11000), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_55 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_2 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_2 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[2]), .Y(n1) );
  INVX1 U4 ( .A(set2[4]), .Y(n2) );
  INVX1 U5 ( .A(set2[7]), .Y(n6) );
  INVX1 U6 ( .A(set2[5]), .Y(n3) );
  INVX1 U7 ( .A(set2[0]), .Y(n5) );
  INVX1 U8 ( .A(set2[1]), .Y(n4) );
  INVX1 U9 ( .A(set2[3]), .Y(n15) );
  NAND3X1 U10 ( .A(n16), .B(n6), .C(n3), .Y(n21) );
  NAND4X1 U11 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U12 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U13 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U14 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U15 ( .C(n5), .D(n14), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U16 ( .A(rdat[0]), .Y(n14) );
  AOI211X1 U17 ( .C(n4), .D(n13), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U18 ( .A(rdat[1]), .Y(n13) );
  AOI211X1 U19 ( .C(n1), .D(n12), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U20 ( .A(rdat[2]), .Y(n12) );
  AOI211X1 U21 ( .C(n15), .D(n11), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U22 ( .A(rdat[3]), .Y(n11) );
  AOI211X1 U23 ( .C(n2), .D(n10), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U24 ( .A(rdat[4]), .Y(n10) );
  AOI211X1 U25 ( .C(n3), .D(n9), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U26 ( .A(rdat[5]), .Y(n9) );
  AOI211X1 U27 ( .C(n16), .D(n8), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U28 ( .A(rdat[6]), .Y(n8) );
  AOI211X1 U29 ( .C(n6), .D(n7), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U30 ( .A(rdat[7]), .Y(n7) );
  NOR2X1 U31 ( .A(rdat[3]), .B(n15), .Y(irq[3]) );
  NOR2X1 U32 ( .A(rdat[2]), .B(n1), .Y(irq[2]) );
  NOR2X1 U33 ( .A(rdat[5]), .B(n3), .Y(irq[5]) );
  NOR2X1 U34 ( .A(rdat[4]), .B(n2), .Y(irq[4]) );
  NOR2X1 U35 ( .A(rdat[0]), .B(n5), .Y(irq[0]) );
  NOR2X1 U36 ( .A(rdat[1]), .B(n4), .Y(irq[1]) );
  NOR2X1 U37 ( .A(rdat[7]), .B(n6), .Y(irq[7]) );
  NOR2X1 U38 ( .A(rdat[6]), .B(n16), .Y(irq[6]) );
  INVX1 U39 ( .A(set2[6]), .Y(n16) );
endmodule


module glreg_WIDTH8_2 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11018;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11018), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11018), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11018), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11018), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11018), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11018), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11018), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11018), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11018), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_9 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n2, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n10), .C(clk), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n7), .A(n2), .Y(n11) );
  NOR3XL U4 ( .A(n7), .B(n2), .C(db_cnt[0]), .Y(o_chg) );
  XNOR2XL U5 ( .A(d_org_0_), .B(o_dbc), .Y(n7) );
  INVX1 U6 ( .A(db_cnt[1]), .Y(n2) );
  MUX2X1 U7 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n10) );
  NOR2X1 U8 ( .A(db_cnt[0]), .B(n11), .Y(n8) );
  NOR21XL U9 ( .B(db_cnt[0]), .A(n11), .Y(n9) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_10 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n2, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n10), .C(clk), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n7), .A(n2), .Y(n11) );
  NOR3XL U4 ( .A(n7), .B(n2), .C(db_cnt[0]), .Y(o_chg) );
  INVX1 U5 ( .A(db_cnt[1]), .Y(n2) );
  XNOR2XL U6 ( .A(d_org_0_), .B(o_dbc), .Y(n7) );
  MUX2X1 U7 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n10) );
  NOR2X1 U8 ( .A(db_cnt[0]), .B(n11), .Y(n8) );
  NOR21XL U9 ( .B(db_cnt[0]), .A(n11), .Y(n9) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_11 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n2, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n10), .C(clk), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n7), .A(n2), .Y(n11) );
  XNOR2XL U4 ( .A(d_org_0_), .B(o_dbc), .Y(n7) );
  NOR3XL U5 ( .A(n7), .B(n2), .C(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(db_cnt[1]), .Y(n2) );
  MUX2X1 U7 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n10) );
  NOR2X1 U8 ( .A(db_cnt[0]), .B(n11), .Y(n8) );
  NOR21XL U9 ( .B(db_cnt[0]), .A(n11), .Y(n9) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_12 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n2, n7, n8, n9, n10, n11, n12;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n10), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n9), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n11), .C(clk), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n8), .A(n7), .Y(n12) );
  MUX2X1 U4 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n11) );
  INVX1 U5 ( .A(n2), .Y(o_chg) );
  NAND32X1 U6 ( .B(n8), .C(n7), .A(n1), .Y(n2) );
  INVX1 U7 ( .A(db_cnt[0]), .Y(n1) );
  NOR2X1 U8 ( .A(db_cnt[0]), .B(n12), .Y(n9) );
  XNOR2XL U9 ( .A(d_org_0_), .B(o_dbc), .Y(n8) );
  NOR21XL U10 ( .B(db_cnt[0]), .A(n12), .Y(n10) );
  INVX1 U11 ( .A(db_cnt[1]), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_13 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n2, n7, n8, n9, n10, n11, n12;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n10), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n9), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n11), .C(clk), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n8), .A(n7), .Y(n12) );
  MUX2X1 U4 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n11) );
  INVX1 U5 ( .A(n2), .Y(o_chg) );
  NAND32X1 U6 ( .B(n8), .C(n7), .A(n1), .Y(n2) );
  INVX1 U7 ( .A(db_cnt[0]), .Y(n1) );
  NOR2X1 U8 ( .A(db_cnt[0]), .B(n12), .Y(n9) );
  XNOR2XL U9 ( .A(d_org_0_), .B(o_dbc), .Y(n8) );
  NOR21XL U10 ( .B(db_cnt[0]), .A(n12), .Y(n10) );
  INVX1 U11 ( .A(db_cnt[1]), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_14 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n3, n4, n5, n6, n1, n2, n7, n8;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n5), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n6), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n4), .C(clk), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n8), .A(n7), .Y(n3) );
  MUX2X1 U4 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n4) );
  INVX1 U5 ( .A(n2), .Y(o_chg) );
  NAND32X1 U6 ( .B(n8), .C(n7), .A(n1), .Y(n2) );
  INVX1 U7 ( .A(db_cnt[0]), .Y(n1) );
  NOR2X1 U8 ( .A(db_cnt[0]), .B(n3), .Y(n6) );
  XNOR2XL U9 ( .A(d_org_0_), .B(o_dbc), .Y(n8) );
  NOR21XL U10 ( .B(db_cnt[0]), .A(n3), .Y(n5) );
  INVX1 U11 ( .A(db_cnt[1]), .Y(n7) );
endmodule


module dbnc_WIDTH2_0 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n3, n4, n7, n8, n9;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(d_org_0_), .B(o_dbc), .Y(n1) );
  AND3X1 U4 ( .A(db_cnt[0]), .B(db_cnt[1]), .C(n1), .Y(o_chg) );
  INVX1 U5 ( .A(n3), .Y(n7) );
  NAND21X1 U6 ( .B(db_cnt[0]), .A(n1), .Y(n3) );
  MUX2X1 U7 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n9) );
  MUX2X1 U8 ( .D0(n4), .D1(n7), .S(db_cnt[1]), .Y(n8) );
  AND2X1 U9 ( .A(db_cnt[0]), .B(n1), .Y(n4) );
endmodule


module dbnc_WIDTH2_1 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n3, n4, n7, n8, n9;
  wire   [1:0] db_cnt;

  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(d_org_0_), .B(o_dbc), .Y(n1) );
  AND3X1 U4 ( .A(db_cnt[0]), .B(db_cnt[1]), .C(n1), .Y(o_chg) );
  INVX1 U5 ( .A(n3), .Y(n7) );
  NAND21X1 U6 ( .B(db_cnt[0]), .A(n1), .Y(n3) );
  MUX2X1 U7 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n9) );
  MUX2X1 U8 ( .D0(n4), .D1(n7), .S(db_cnt[1]), .Y(n8) );
  AND2X1 U9 ( .A(db_cnt[0]), .B(n1), .Y(n4) );
endmodule


module dbnc_WIDTH2_2 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n3, n4, n7, n8, n9;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(d_org_0_), .B(o_dbc), .Y(n1) );
  AND3X1 U4 ( .A(db_cnt[0]), .B(db_cnt[1]), .C(n1), .Y(o_chg) );
  INVX1 U5 ( .A(n3), .Y(n7) );
  NAND21X1 U6 ( .B(db_cnt[0]), .A(n1), .Y(n3) );
  MUX2X1 U7 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n9) );
  MUX2X1 U8 ( .D0(n4), .D1(n7), .S(db_cnt[1]), .Y(n8) );
  AND2X1 U9 ( .A(db_cnt[0]), .B(n1), .Y(n4) );
endmodule


module dbnc_WIDTH2_3 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n3, n4, n7, n8, n9;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(d_org_0_), .B(o_dbc), .Y(n1) );
  AND3X1 U4 ( .A(db_cnt[0]), .B(db_cnt[1]), .C(n1), .Y(o_chg) );
  INVX1 U5 ( .A(n3), .Y(n7) );
  NAND21X1 U6 ( .B(db_cnt[0]), .A(n1), .Y(n3) );
  MUX2X1 U7 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n9) );
  MUX2X1 U8 ( .D0(n4), .D1(n7), .S(db_cnt[1]), .Y(n8) );
  AND2X1 U9 ( .A(db_cnt[0]), .B(n1), .Y(n4) );
endmodule


module dbnc_WIDTH2_4 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n5, n6, n1, n3, n4, n7;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n6), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n5), .C(clk), .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(d_org_0_), .B(o_dbc), .Y(n1) );
  AND3X1 U4 ( .A(db_cnt[0]), .B(db_cnt[1]), .C(n1), .Y(o_chg) );
  INVX1 U5 ( .A(n3), .Y(n7) );
  NAND21X1 U6 ( .B(db_cnt[0]), .A(n1), .Y(n3) );
  MUX2X1 U7 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n5) );
  MUX2X1 U8 ( .D0(n4), .D1(n7), .S(db_cnt[1]), .Y(n6) );
  AND2X1 U9 ( .A(db_cnt[0]), .B(n1), .Y(n4) );
endmodule


module dbnc_WIDTH5_TIMEOUT30 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N7, N8, N9, N10, N11, N17, N18, N19, N20, N21, N22,
         net11036, n1, n3, n4, n5, n6, n2, n7, n8, n9;
  wire   [4:0] db_cnt;
  wire   [4:2] add_165_carry;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH5_TIMEOUT30 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N17), .ENCLK(net11036), .TE(1'b0) );
  HAD1X1 add_165_U1_1_1 ( .A(db_cnt[1]), .B(db_cnt[0]), .CO(add_165_carry[2]), 
        .SO(N8) );
  HAD1X1 add_165_U1_1_2 ( .A(db_cnt[2]), .B(add_165_carry[2]), .CO(
        add_165_carry[3]), .SO(N9) );
  HAD1X1 add_165_U1_1_3 ( .A(db_cnt[3]), .B(add_165_carry[3]), .CO(
        add_165_carry[4]), .SO(N10) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N19), .C(net11036), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_4_ ( .D(N22), .C(net11036), .XR(rstz), .Q(db_cnt[4]) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N21), .C(net11036), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N20), .C(net11036), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N18), .C(net11036), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n6), .C(net11036), .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n7) );
  INVX1 U4 ( .A(n2), .Y(o_chg) );
  NAND21X1 U5 ( .B(n1), .A(n7), .Y(n2) );
  AND2X1 U6 ( .A(N10), .B(n3), .Y(N21) );
  AND2X1 U7 ( .A(N9), .B(n3), .Y(N20) );
  AND2X1 U8 ( .A(N8), .B(n3), .Y(N19) );
  INVX1 U9 ( .A(n9), .Y(n3) );
  NAND21X1 U10 ( .B(n8), .A(n1), .Y(n9) );
  XNOR2XL U11 ( .A(d_org_0_), .B(o_dbc), .Y(n8) );
  NAND4X1 U12 ( .A(db_cnt[4]), .B(db_cnt[3]), .C(n4), .D(db_cnt[2]), .Y(n1) );
  NOR21XL U13 ( .B(db_cnt[1]), .A(db_cnt[0]), .Y(n4) );
  NAND43X1 U14 ( .B(db_cnt[0]), .C(db_cnt[1]), .D(n7), .A(n5), .Y(N17) );
  NOR3XL U15 ( .A(db_cnt[2]), .B(db_cnt[4]), .C(db_cnt[3]), .Y(n5) );
  MUX2X1 U16 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n6) );
  AND2X1 U17 ( .A(N11), .B(n3), .Y(N22) );
  AND2X1 U18 ( .A(N7), .B(n3), .Y(N18) );
  INVX1 U19 ( .A(db_cnt[0]), .Y(N7) );
  XOR2X1 U20 ( .A(add_165_carry[4]), .B(db_cnt[4]), .Y(N11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH5_TIMEOUT30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_0 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N15, N16, N17, N18, N19, net11054, n4, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n2, n3, n5, n14, n15;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11054), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N19), .C(net11054), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N16), .C(net11054), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N17), .C(net11054), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N18), .C(net11054), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 d_org_reg_1_ ( .D(n13), .C(net11054), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n3), .A(n4), .Y(n7) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  XNOR2XL U5 ( .A(d_org_0_), .B(o_dbc), .Y(n3) );
  AOI21BBXL U6 ( .B(db_cnt[1]), .C(n7), .A(N16), .Y(n9) );
  OAI32X1 U7 ( .A(n6), .B(n7), .C(n5), .D(n8), .E(n15), .Y(N19) );
  NAND3X1 U8 ( .A(db_cnt[1]), .B(n15), .C(db_cnt[2]), .Y(n6) );
  OA21X1 U9 ( .B(n7), .C(db_cnt[2]), .A(n9), .Y(n8) );
  INVX1 U10 ( .A(db_cnt[3]), .Y(n15) );
  NOR2X1 U11 ( .A(n7), .B(db_cnt[0]), .Y(N16) );
  NAND4X1 U12 ( .A(db_cnt[3]), .B(db_cnt[2]), .C(db_cnt[1]), .D(n5), .Y(n4) );
  MUX2X1 U13 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n13) );
  INVX1 U14 ( .A(n1), .Y(o_chg) );
  NAND21X1 U15 ( .B(n4), .A(n2), .Y(n1) );
  NAND32X1 U16 ( .B(db_cnt[0]), .C(n2), .A(n12), .Y(N15) );
  NOR3XL U17 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n12) );
  OAI21X1 U18 ( .B(n9), .C(n14), .A(n10), .Y(N18) );
  NAND42X1 U19 ( .C(n7), .D(n5), .A(db_cnt[1]), .B(n14), .Y(n10) );
  INVX1 U20 ( .A(db_cnt[2]), .Y(n14) );
  INVX1 U21 ( .A(db_cnt[0]), .Y(n5) );
  NOR2X1 U22 ( .A(n11), .B(n7), .Y(N17) );
  XNOR2XL U23 ( .A(db_cnt[1]), .B(db_cnt[0]), .Y(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_1 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N15, N16, N17, N18, N19, net11072, n4, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n2, n3, n5, n14, n15;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11072), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N19), .C(net11072), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N16), .C(net11072), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N17), .C(net11072), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N18), .C(net11072), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 d_org_reg_1_ ( .D(n13), .C(net11072), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n3), .A(n4), .Y(n7) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  XNOR2XL U5 ( .A(d_org_0_), .B(o_dbc), .Y(n3) );
  AOI21BBXL U6 ( .B(db_cnt[1]), .C(n7), .A(N16), .Y(n9) );
  OAI32X1 U7 ( .A(n6), .B(n7), .C(n5), .D(n8), .E(n15), .Y(N19) );
  NAND3X1 U8 ( .A(db_cnt[1]), .B(n15), .C(db_cnt[2]), .Y(n6) );
  OA21X1 U9 ( .B(n7), .C(db_cnt[2]), .A(n9), .Y(n8) );
  INVX1 U10 ( .A(db_cnt[3]), .Y(n15) );
  NOR2X1 U11 ( .A(n7), .B(db_cnt[0]), .Y(N16) );
  NAND4X1 U12 ( .A(db_cnt[3]), .B(db_cnt[2]), .C(db_cnt[1]), .D(n5), .Y(n4) );
  MUX2X1 U13 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n13) );
  INVX1 U14 ( .A(n1), .Y(o_chg) );
  NAND21X1 U15 ( .B(n4), .A(n2), .Y(n1) );
  NAND32X1 U16 ( .B(db_cnt[0]), .C(n2), .A(n12), .Y(N15) );
  NOR3XL U17 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n12) );
  OAI21X1 U18 ( .B(n9), .C(n14), .A(n10), .Y(N18) );
  NAND42X1 U19 ( .C(n7), .D(n5), .A(db_cnt[1]), .B(n14), .Y(n10) );
  INVX1 U20 ( .A(db_cnt[2]), .Y(n14) );
  INVX1 U21 ( .A(db_cnt[0]), .Y(n5) );
  NOR2X1 U22 ( .A(n11), .B(n7), .Y(N17) );
  XNOR2XL U23 ( .A(db_cnt[1]), .B(db_cnt[0]), .Y(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_2 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N15, N16, N17, N18, N19, net11090, n4, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n2, n3, n5, n14, n15;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11090), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N19), .C(net11090), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N16), .C(net11090), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N17), .C(net11090), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N18), .C(net11090), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 d_org_reg_1_ ( .D(n13), .C(net11090), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n3), .A(n4), .Y(n7) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  XNOR2XL U5 ( .A(d_org_0_), .B(o_dbc), .Y(n3) );
  AOI21BBXL U6 ( .B(db_cnt[1]), .C(n7), .A(N16), .Y(n9) );
  OAI32X1 U7 ( .A(n6), .B(n7), .C(n5), .D(n8), .E(n15), .Y(N19) );
  NAND3X1 U8 ( .A(db_cnt[1]), .B(n15), .C(db_cnt[2]), .Y(n6) );
  OA21X1 U9 ( .B(n7), .C(db_cnt[2]), .A(n9), .Y(n8) );
  INVX1 U10 ( .A(db_cnt[3]), .Y(n15) );
  NOR2X1 U11 ( .A(n7), .B(db_cnt[0]), .Y(N16) );
  NAND4X1 U12 ( .A(db_cnt[3]), .B(db_cnt[2]), .C(db_cnt[1]), .D(n5), .Y(n4) );
  MUX2X1 U13 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n13) );
  INVX1 U14 ( .A(n1), .Y(o_chg) );
  NAND21X1 U15 ( .B(n4), .A(n2), .Y(n1) );
  NAND32X1 U16 ( .B(db_cnt[0]), .C(n2), .A(n12), .Y(N15) );
  NOR3XL U17 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n12) );
  OAI21X1 U18 ( .B(n9), .C(n14), .A(n10), .Y(N18) );
  NAND42X1 U19 ( .C(n7), .D(n5), .A(db_cnt[1]), .B(n14), .Y(n10) );
  INVX1 U20 ( .A(db_cnt[2]), .Y(n14) );
  INVX1 U21 ( .A(db_cnt[0]), .Y(n5) );
  NOR2X1 U22 ( .A(n11), .B(n7), .Y(N17) );
  XNOR2XL U23 ( .A(db_cnt[1]), .B(db_cnt[0]), .Y(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000028 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11108;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11108), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11108), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11108), .XR(arstz), .Q(rdat[6]) );
  DFFSQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11108), .XS(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11108), .XS(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11108), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11108), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11108), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11108), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_56 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11126;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_56 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11126), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11126), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11126), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11126), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11126), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11126), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11126), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11126), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11126), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_56 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_57 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11144;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_57 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11144), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11144), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11144), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11144), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11144), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11144), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11144), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11144), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11144), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_57 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_58 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11162;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_58 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11162), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11162), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11162), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11162), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11162), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11162), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11162), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11162), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11162), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_58 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_59 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11180;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_59 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11180), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11180), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11180), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11180), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11180), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11180), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11180), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11180), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11180), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_59 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_60 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11198;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_60 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11198), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11198), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11198), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11198), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11198), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11198), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11198), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11198), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11198), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_60 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_61 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11216;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_61 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11216), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11216), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11216), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11216), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11216), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11216), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11216), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11216), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11216), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_61 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_62 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11234;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_62 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11234), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11234), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11234), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11234), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11234), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11234), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11234), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11234), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11234), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_62 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_63 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11252;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_63 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11252), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11252), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11252), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11252), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11252), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11252), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11252), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11252), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11252), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_63 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH4 ( clk, arstz, we, wdat, rdat );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we;
  wire   net11270;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11270), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11270), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11270), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11270), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11270), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_64 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11288;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_64 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11288), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11288), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11288), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11288), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11288), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11288), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11288), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11288), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11288), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_64 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_3 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_3 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[0]), .Y(n16) );
  INVX1 U4 ( .A(set2[1]), .Y(n15) );
  INVX1 U5 ( .A(set2[2]), .Y(n14) );
  INVX1 U6 ( .A(set2[3]), .Y(n13) );
  INVX1 U7 ( .A(set2[4]), .Y(n12) );
  NAND3X1 U8 ( .A(n10), .B(n9), .C(n11), .Y(n21) );
  NAND4X1 U9 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U10 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U11 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U12 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U13 ( .C(n16), .D(n8), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U14 ( .A(rdat[0]), .Y(n8) );
  AOI211X1 U15 ( .C(n15), .D(n7), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U16 ( .A(rdat[1]), .Y(n7) );
  AOI211X1 U17 ( .C(n14), .D(n6), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U18 ( .A(rdat[2]), .Y(n6) );
  AOI211X1 U19 ( .C(n13), .D(n5), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U20 ( .A(rdat[3]), .Y(n5) );
  AOI211X1 U21 ( .C(n12), .D(n4), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U22 ( .A(rdat[4]), .Y(n4) );
  AOI211X1 U23 ( .C(n11), .D(n3), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U24 ( .A(rdat[5]), .Y(n3) );
  AOI211X1 U25 ( .C(n10), .D(n2), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U26 ( .A(rdat[6]), .Y(n2) );
  AOI211X1 U27 ( .C(n9), .D(n1), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U28 ( .A(rdat[7]), .Y(n1) );
  NOR2X1 U29 ( .A(rdat[0]), .B(n16), .Y(irq[0]) );
  NOR2X1 U30 ( .A(rdat[1]), .B(n15), .Y(irq[1]) );
  NOR2X1 U31 ( .A(rdat[2]), .B(n14), .Y(irq[2]) );
  NOR2X1 U32 ( .A(rdat[3]), .B(n13), .Y(irq[3]) );
  INVX1 U33 ( .A(set2[6]), .Y(n10) );
  INVX1 U34 ( .A(set2[7]), .Y(n9) );
  INVX1 U35 ( .A(set2[5]), .Y(n11) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n12), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n10), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[5]), .B(n11), .Y(irq[5]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n9), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_3 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11306;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11306), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11306), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11306), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11306), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11306), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11306), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11306), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11306), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11306), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_65 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11324;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_65 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11324), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11324), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11324), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11324), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11324), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11324), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11324), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11324), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11324), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_65 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_66 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11342;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_66 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11342), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11342), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11342), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11342), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11342), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11342), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11342), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11342), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11342), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_66 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000032 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11360;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11360), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11360), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11360), .XR(arstz), .Q(rdat[3]) );
  DFFSQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11360), .XS(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11360), .XR(arstz), .Q(rdat[6]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11360), .XS(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11360), .XR(arstz), .Q(rdat[2]) );
  DFFSQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11360), .XS(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11360), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000098 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11378;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11378), .TE(1'b0) );
  DFFSQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11378), .XS(arstz), .Q(rdat[7]) );
  DFFSQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11378), .XS(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11378), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11378), .XR(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11378), .XS(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11378), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11378), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11378), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_000000f0 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11396;

  SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11396), .TE(1'b0) );
  DFFSQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11396), .XS(arstz), .Q(rdat[7]) );
  DFFSQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11396), .XS(arstz), .Q(rdat[6]) );
  DFFSQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11396), .XS(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11396), .XS(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11396), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11396), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11396), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11396), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_3 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  MUX2XL U2 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n2) );
endmodule


module glreg_WIDTH1_4 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  MUX2XL U2 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n2) );
endmodule


module glreg_WIDTH1_5 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n1;

  DFFRQX1 mem_reg_0_ ( .D(n1), .C(clk), .XR(arstz), .Q(rdat[0]) );
  MUX2XL U2 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n1) );
endmodule


module glreg_WIDTH2_2 ( clk, arstz, we, wdat, rdat );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we;
  wire   n2, n3;

  DFFRQX1 mem_reg_1_ ( .D(n3), .C(clk), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  MUX2XL U2 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n2) );
  MUX2XL U3 ( .D0(rdat[1]), .D1(wdat[1]), .S(we), .Y(n3) );
endmodule


module glreg_WIDTH3 ( clk, arstz, we, wdat, rdat );
  input [2:0] wdat;
  output [2:0] rdat;
  input clk, arstz, we;
  wire   net11414;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11414), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11414), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11414), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11414), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000011 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11432;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11432), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11432), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11432), .XR(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11432), .XS(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11432), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11432), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11432), .XR(arstz), .Q(rdat[2]) );
  DFFSQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11432), .XS(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11432), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000001 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11450;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11450), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11450), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11450), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11450), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11450), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11450), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11450), .XR(arstz), .Q(rdat[2]) );
  DFFSQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11450), .XS(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11450), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_67 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11468;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_67 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11468), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11468), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11468), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11468), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11468), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11468), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11468), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11468), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11468), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_67 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_4 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_4 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  INVXL U2 ( .A(set2[7]), .Y(n4) );
  NOR4XL U3 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U4 ( .A(set2[3]), .Y(n14) );
  INVX1 U5 ( .A(set2[0]), .Y(n1) );
  NAND3X1 U6 ( .A(n3), .B(n4), .C(n2), .Y(n21) );
  INVX1 U7 ( .A(set2[1]), .Y(n16) );
  INVX1 U8 ( .A(set2[4]), .Y(n13) );
  INVX1 U9 ( .A(set2[6]), .Y(n3) );
  INVX1 U10 ( .A(set2[2]), .Y(n15) );
  INVX1 U11 ( .A(set2[5]), .Y(n2) );
  NAND4X1 U12 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U13 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U14 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U15 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U16 ( .C(n1), .D(n12), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U17 ( .A(rdat[0]), .Y(n12) );
  AOI211X1 U18 ( .C(n16), .D(n11), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U19 ( .A(rdat[1]), .Y(n11) );
  AOI211X1 U20 ( .C(n15), .D(n10), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U21 ( .A(rdat[2]), .Y(n10) );
  AOI211X1 U22 ( .C(n14), .D(n9), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U23 ( .A(rdat[3]), .Y(n9) );
  AOI211X1 U24 ( .C(n13), .D(n8), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U25 ( .A(rdat[4]), .Y(n8) );
  AOI211X1 U26 ( .C(n2), .D(n7), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U27 ( .A(rdat[5]), .Y(n7) );
  AOI211X1 U28 ( .C(n3), .D(n6), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U29 ( .A(rdat[6]), .Y(n6) );
  AOI211X1 U30 ( .C(n4), .D(n5), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U31 ( .A(rdat[7]), .Y(n5) );
  NOR2X1 U32 ( .A(rdat[7]), .B(n4), .Y(irq[7]) );
  NOR2X1 U33 ( .A(rdat[6]), .B(n3), .Y(irq[6]) );
  NOR2X1 U34 ( .A(rdat[3]), .B(n14), .Y(irq[3]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n15), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n1), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[4]), .B(n13), .Y(irq[4]) );
  NOR2X1 U38 ( .A(rdat[5]), .B(n2), .Y(irq[5]) );
  NOR2X1 U39 ( .A(rdat[1]), .B(n16), .Y(irq[1]) );
endmodule


module glreg_WIDTH8_4 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11486;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11486), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11486), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11486), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11486), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11486), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11486), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11486), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11486), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11486), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_68 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11504;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_68 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11504), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11504), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11504), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11504), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11504), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11504), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11504), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11504), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11504), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_68 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_7_70 ( clk, arstz, we, wdat, rdat );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we;
  wire   net11522;

  SNPS_CLOCK_GATE_HIGH_glreg_7_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11522), .TE(1'b0) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11522), .XS(arstz), .Q(rdat[4]) );
  DFFSQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11522), .XS(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11522), .XS(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11522), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11522), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11522), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11522), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_7_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_1_1_0 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFSQX1 mem_reg_0_ ( .D(n2), .C(clk), .XS(arstz), .Q(rdat[0]) );
  MUX2X1 U2 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n2) );
endmodule


module glreg_1_1_1 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n1;

  DFFSQX1 mem_reg_0_ ( .D(n1), .C(clk), .XS(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n1) );
endmodule


module glreg_6_00000018 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net11540;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11540), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11540), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11540), .XR(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11540), .XS(arstz), .Q(rdat[4]) );
  DFFSQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11540), .XS(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11540), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11540), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_69 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11558;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_69 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11558), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11558), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11558), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11558), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11558), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11558), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11558), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11558), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11558), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_69 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_70 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11576;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11576), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11576), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11576), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11576), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11576), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11576), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11576), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11576), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11576), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_71 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11594;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_71 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11594), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11594), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11594), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11594), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11594), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11594), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11594), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11594), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11594), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_71 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_72 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11612;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_72 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11612), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11612), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11612), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11612), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11612), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11612), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11612), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11612), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11612), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_72 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_73 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11630;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_73 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11630), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11630), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11630), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11630), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11630), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11630), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11630), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11630), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11630), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_73 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_2 ( clk, arstz, we, wdat, rdat );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we;
  wire   net11648;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11648), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11648), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11648), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11648), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11648), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11648), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_74 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11666;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_74 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11666), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11666), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11666), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11666), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11666), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11666), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11666), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11666), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11666), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_74 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_75 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11684;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_75 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11684), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11684), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11684), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11684), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11684), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11684), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11684), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11684), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11684), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_75 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_76 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11702;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_76 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11702), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11702), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11702), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11702), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11702), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11702), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11702), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11702), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11702), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_76 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_77 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11720;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_77 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11720), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11720), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11720), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11720), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11720), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11720), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11720), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11720), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11720), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_77 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_5 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_5 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR3XL U2 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NAND3X1 U3 ( .A(n14), .B(n3), .C(n2), .Y(n21) );
  INVX1 U4 ( .A(set2[4]), .Y(n1) );
  INVX1 U5 ( .A(set2[3]), .Y(n4) );
  INVX1 U6 ( .A(set2[2]), .Y(n5) );
  INVX1 U7 ( .A(set2[1]), .Y(n15) );
  INVX1 U8 ( .A(set2[5]), .Y(n2) );
  NAND4X1 U9 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U10 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U11 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  NOR4XL U12 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  INVX1 U13 ( .A(set2[6]), .Y(n14) );
  INVX1 U14 ( .A(set2[0]), .Y(n16) );
  INVX1 U15 ( .A(set2[7]), .Y(n3) );
  NOR2X1 U16 ( .A(rdat[4]), .B(n1), .Y(irq[4]) );
  NOR2X1 U17 ( .A(rdat[5]), .B(n2), .Y(irq[5]) );
  AOI211X1 U18 ( .C(n2), .D(n8), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U19 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U20 ( .C(n1), .D(n9), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U21 ( .A(rdat[4]), .Y(n9) );
  AOI211X1 U22 ( .C(n16), .D(n13), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U23 ( .A(rdat[0]), .Y(n13) );
  AOI211X1 U24 ( .C(n15), .D(n12), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U25 ( .A(rdat[1]), .Y(n12) );
  AOI211X1 U26 ( .C(n5), .D(n11), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U27 ( .A(rdat[2]), .Y(n11) );
  AOI211X1 U28 ( .C(n4), .D(n10), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U29 ( .A(rdat[3]), .Y(n10) );
  AOI211X1 U30 ( .C(n14), .D(n7), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U31 ( .A(rdat[6]), .Y(n7) );
  AOI211X1 U32 ( .C(n3), .D(n6), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U33 ( .A(rdat[7]), .Y(n6) );
  NOR2X1 U34 ( .A(rdat[2]), .B(n5), .Y(irq[2]) );
  NOR2X1 U35 ( .A(rdat[3]), .B(n4), .Y(irq[3]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n16), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n14), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[1]), .B(n15), .Y(irq[1]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n3), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_5 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11738;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11738), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11738), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11738), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11738), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11738), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11738), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11738), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11738), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11738), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_6 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_6 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  INVX1 U2 ( .A(set2[7]), .Y(n2) );
  INVX1 U3 ( .A(set2[3]), .Y(n5) );
  NAND4X1 U4 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR3XL U5 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U6 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U7 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U8 ( .A(set2[1]), .Y(n1) );
  INVX1 U9 ( .A(set2[2]), .Y(n3) );
  INVX1 U10 ( .A(set2[4]), .Y(n6) );
  NOR4XL U11 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NAND3X1 U12 ( .A(n4), .B(n2), .C(n15), .Y(n21) );
  INVX1 U13 ( .A(set2[6]), .Y(n4) );
  INVX1 U14 ( .A(set2[0]), .Y(n16) );
  AOI211X1 U15 ( .C(n16), .D(n14), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U16 ( .A(rdat[0]), .Y(n14) );
  AOI211X1 U17 ( .C(n1), .D(n13), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U18 ( .A(rdat[1]), .Y(n13) );
  AOI211X1 U19 ( .C(n3), .D(n12), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U20 ( .A(rdat[2]), .Y(n12) );
  AOI211X1 U21 ( .C(n5), .D(n11), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U22 ( .A(rdat[3]), .Y(n11) );
  AOI211X1 U23 ( .C(n6), .D(n10), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U24 ( .A(rdat[4]), .Y(n10) );
  AOI211X1 U25 ( .C(n15), .D(n9), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U26 ( .A(rdat[5]), .Y(n9) );
  AOI211X1 U27 ( .C(n4), .D(n8), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U28 ( .A(rdat[6]), .Y(n8) );
  AOI211X1 U29 ( .C(n2), .D(n7), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U30 ( .A(rdat[7]), .Y(n7) );
  NOR2X1 U31 ( .A(rdat[6]), .B(n4), .Y(irq[6]) );
  NOR2X1 U32 ( .A(rdat[7]), .B(n2), .Y(irq[7]) );
  NOR2X1 U33 ( .A(rdat[2]), .B(n3), .Y(irq[2]) );
  NOR2X1 U34 ( .A(rdat[0]), .B(n16), .Y(irq[0]) );
  NOR2X1 U35 ( .A(rdat[1]), .B(n1), .Y(irq[1]) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n6), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[3]), .B(n5), .Y(irq[3]) );
  INVX1 U38 ( .A(set2[5]), .Y(n15) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n15), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_6 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11756;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11756), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11756), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11756), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11756), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11756), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11756), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11756), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11756), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11756), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_78 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11774;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_78 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11774), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11774), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11774), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11774), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11774), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11774), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11774), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11774), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11774), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_78 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_79 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11792;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_79 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11792), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11792), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11792), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11792), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11792), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11792), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11792), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11792), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11792), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_79 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ictlr_a0 ( bkpt_ena, bkpt_pc, memaddr_c, memaddr, mcu_psr_c, mcu_psw, 
        hit_ps_c, hit_ps, mempsack, memdatao, o_set_hold, o_bkp_hold, 
        o_ofs_inc, o_inst, d_inst, sfr_psrack, sfr_psofs, sfr_psr, sfr_psw, 
        dw_rst, dw_ena, sfr_wdat, pmem_pgm, pmem_re, pmem_csb, pmem_clk, 
        pmem_a, pmem_q0, pmem_q1, pmem_twlb, wd_twlb, we_twlb, pwrdn_rst, 
        r_pwdn_en, r_multi, r_hold_mcu, clk, srst );
  input [14:0] bkpt_pc;
  input [14:0] memaddr_c;
  input [14:0] memaddr;
  input [7:0] memdatao;
  output [7:0] o_inst;
  output [7:0] d_inst;
  input [14:0] sfr_psofs;
  input [7:0] sfr_wdat;
  output [1:0] pmem_clk;
  output [15:0] pmem_a;
  input [7:0] pmem_q0;
  input [7:0] pmem_q1;
  output [1:0] pmem_twlb;
  input [1:0] wd_twlb;
  input bkpt_ena, mcu_psr_c, mcu_psw, hit_ps_c, hit_ps, sfr_psr, sfr_psw,
         dw_rst, dw_ena, we_twlb, pwrdn_rst, r_pwdn_en, r_multi, r_hold_mcu,
         clk, srst;
  output mempsack, o_set_hold, o_bkp_hold, o_ofs_inc, sfr_psrack, pmem_pgm,
         pmem_re, pmem_csb;
  wire   N152, N153, N154, c_buf_22__7_, c_buf_22__6_, c_buf_22__5_,
         c_buf_22__4_, c_buf_22__3_, c_buf_22__2_, c_buf_22__1_, c_buf_22__0_,
         c_buf_21__7_, c_buf_21__6_, c_buf_21__5_, c_buf_21__4_, c_buf_21__3_,
         c_buf_21__2_, c_buf_21__1_, c_buf_21__0_, c_buf_20__7_, c_buf_20__6_,
         c_buf_20__5_, c_buf_20__4_, c_buf_20__3_, c_buf_20__2_, c_buf_20__1_,
         c_buf_20__0_, c_buf_19__7_, c_buf_19__6_, c_buf_19__5_, c_buf_19__4_,
         c_buf_19__3_, c_buf_19__2_, c_buf_19__1_, c_buf_19__0_, c_buf_18__7_,
         c_buf_18__6_, c_buf_18__5_, c_buf_18__4_, c_buf_18__3_, c_buf_18__2_,
         c_buf_18__1_, c_buf_18__0_, c_buf_17__7_, c_buf_17__6_, c_buf_17__5_,
         c_buf_17__4_, c_buf_17__3_, c_buf_17__2_, c_buf_17__1_, c_buf_17__0_,
         c_buf_16__7_, c_buf_16__6_, c_buf_16__5_, c_buf_16__4_, c_buf_16__3_,
         c_buf_16__2_, c_buf_16__1_, c_buf_16__0_, d_psrd, r_rdy, N353, N354,
         N355, N356, N357, N358, N359, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N479, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491,
         N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502,
         N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634,
         N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645,
         N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656,
         N657, N658, N659, N660, N661, N662, N757, N758, N759, N786, N787,
         N788, N789, N790, N791, N792, N793, N795, N796, N797, N798, N799,
         N800, N801, N820, N821, N822, N823, N824, N825, N826, N827, N828,
         N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839,
         N840, N842, N843, N844, N845, N846, N853, N854, N855, N856, N857,
         N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868,
         N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895,
         N896, N897, N898, N899, cs_n, un_hold, N974, net11818, net11824,
         net11829, net11834, net11839, net11844, net11849, net11854, net11859,
         net11864, net11869, net11874, net11879, net11884, net11889, net11894,
         net11899, net11904, net11909, net11914, net11919, net11924, net11929,
         net11934, net11939, net11944, net11949, net11954, net11959, net11964,
         n93, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923;
  wire   [3:0] d_hold;
  wire   [1:0] dummy;
  wire   [3:0] cs_ft;
  wire   [4:0] c_ptr;
  wire   [14:0] c_adr;
  wire   [14:13] adr_p;
  wire   [7:0] rd_buf;
  wire   [7:0] dbg_01;
  wire   [7:0] dbg_02;
  wire   [7:0] dbg_03;
  wire   [7:0] dbg_04;
  wire   [7:0] dbg_05;
  wire   [7:0] dbg_06;
  wire   [7:0] dbg_07;
  wire   [7:0] dbg_08;
  wire   [7:0] dbg_09;
  wire   [7:0] dbg_0a;
  wire   [7:0] dbg_0b;
  wire   [7:0] dbg_0c;
  wire   [7:0] dbg_0d;
  wire   [7:0] dbg_0e;
  wire   [7:0] dbg_0f;
  wire   [7:0] wr_buf;
  wire   [14:0] pre_1_adr;
  wire   [6:0] wspp_cnt;

  SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 clk_gate_wspp_cnt_reg ( .CLK(clk), .EN(N899), 
        .ENCLK(net11818), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 clk_gate_a_bit_reg ( .CLK(clk), .EN(N898), 
        .ENCLK(net11824), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 clk_gate_adr_p_reg ( .CLK(clk), .EN(N853), 
        .ENCLK(net11829), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 clk_gate_c_buf_reg_23_ ( .CLK(clk), .EN(
        N897), .ENCLK(net11834), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 clk_gate_c_buf_reg_22_ ( .CLK(clk), .EN(
        N896), .ENCLK(net11839), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 clk_gate_c_buf_reg_21_ ( .CLK(clk), .EN(
        N895), .ENCLK(net11844), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 clk_gate_c_buf_reg_20_ ( .CLK(clk), .EN(
        N894), .ENCLK(net11849), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 clk_gate_c_buf_reg_19_ ( .CLK(clk), .EN(
        N893), .ENCLK(net11854), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 clk_gate_c_buf_reg_18_ ( .CLK(clk), .EN(
        N892), .ENCLK(net11859), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 clk_gate_c_buf_reg_17_ ( .CLK(clk), .EN(
        N891), .ENCLK(net11864), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 clk_gate_c_buf_reg_16_ ( .CLK(clk), .EN(
        N890), .ENCLK(net11869), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 clk_gate_c_buf_reg_15_ ( .CLK(clk), .EN(
        N889), .ENCLK(net11874), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 clk_gate_c_buf_reg_14_ ( .CLK(clk), .EN(
        N888), .ENCLK(net11879), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 clk_gate_c_buf_reg_13_ ( .CLK(clk), .EN(
        N887), .ENCLK(net11884), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 clk_gate_c_buf_reg_12_ ( .CLK(clk), .EN(
        N886), .ENCLK(net11889), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 clk_gate_c_buf_reg_11_ ( .CLK(clk), .EN(
        N885), .ENCLK(net11894), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 clk_gate_c_buf_reg_10_ ( .CLK(clk), .EN(
        N884), .ENCLK(net11899), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 clk_gate_c_buf_reg_9_ ( .CLK(clk), .EN(N883), .ENCLK(net11904), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 clk_gate_c_buf_reg_8_ ( .CLK(clk), .EN(N882), .ENCLK(net11909), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 clk_gate_c_buf_reg_7_ ( .CLK(clk), .EN(N881), .ENCLK(net11914), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 clk_gate_c_buf_reg_6_ ( .CLK(clk), .EN(N880), .ENCLK(net11919), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 clk_gate_c_buf_reg_5_ ( .CLK(clk), .EN(N879), 
        .ENCLK(net11924), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 clk_gate_c_buf_reg_4_ ( .CLK(clk), .EN(N878), 
        .ENCLK(net11929), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 clk_gate_c_buf_reg_3_ ( .CLK(clk), .EN(N877), 
        .ENCLK(net11934), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 clk_gate_c_buf_reg_2_ ( .CLK(clk), .EN(N876), 
        .ENCLK(net11939), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 clk_gate_c_buf_reg_1_ ( .CLK(clk), .EN(N875), 
        .ENCLK(net11944), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 clk_gate_c_buf_reg_0_ ( .CLK(clk), .EN(N874), 
        .ENCLK(net11949), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 clk_gate_c_ptr_reg ( .CLK(clk), .EN(n93), 
        .ENCLK(net11954), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 clk_gate_c_adr_reg ( .CLK(clk), .EN(N825), 
        .ENCLK(net11959), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 clk_gate_cs_ft_reg ( .CLK(clk), .EN(N820), 
        .ENCLK(net11964), .TE(1'b0) );
  ictlr_a0_DW01_inc_1 add_242 ( .A(c_adr), .SUM({N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431}) );
  ictlr_a0_DW01_inc_2 r492 ( .A({adr_p, pmem_a[15:9], pmem_a[5:0]}), .SUM(
        pre_1_adr) );
  DFFNQXL ck_n_reg_1_ ( .D(n642), .XC(clk), .Q(pmem_clk[1]) );
  DFFNQXL ck_n_reg_0_ ( .D(n641), .XC(clk), .Q(pmem_clk[0]) );
  DFFQX1 wspp_cnt_reg_1_ ( .D(N796), .C(net11818), .Q(wspp_cnt[1]) );
  DFFQX1 wspp_cnt_reg_2_ ( .D(N797), .C(net11818), .Q(wspp_cnt[2]) );
  DFFQX1 wspp_cnt_reg_0_ ( .D(N795), .C(net11818), .Q(wspp_cnt[0]) );
  DFFQX1 dummy_reg_1_ ( .D(n650), .C(clk), .Q(dummy[1]) );
  DFFQX1 dummy_reg_0_ ( .D(n651), .C(clk), .Q(dummy[0]) );
  DFFQX1 d_hold_reg_0_ ( .D(n923), .C(clk), .Q(d_hold[0]) );
  DFFQX1 d_hold_reg_3_ ( .D(N154), .C(clk), .Q(d_hold[3]) );
  DFFQX1 d_hold_reg_1_ ( .D(N152), .C(clk), .Q(d_hold[1]) );
  DFFQX1 d_hold_reg_2_ ( .D(N153), .C(clk), .Q(d_hold[2]) );
  DFFQX1 d_psrd_reg ( .D(n649), .C(net11964), .Q(d_psrd) );
  DFFQX1 c_adr_reg_12_ ( .D(N838), .C(net11959), .Q(c_adr[12]) );
  DFFQX1 c_adr_reg_14_ ( .D(N840), .C(net11959), .Q(c_adr[14]) );
  DFFQX1 c_adr_reg_13_ ( .D(N839), .C(net11959), .Q(c_adr[13]) );
  DFFQX1 c_adr_reg_11_ ( .D(N837), .C(net11959), .Q(c_adr[11]) );
  DFFQX1 c_adr_reg_10_ ( .D(N836), .C(net11959), .Q(c_adr[10]) );
  DFFQX1 c_adr_reg_9_ ( .D(N835), .C(net11959), .Q(c_adr[9]) );
  DFFQX1 c_adr_reg_8_ ( .D(N834), .C(net11959), .Q(c_adr[8]) );
  DFFQX1 c_adr_reg_7_ ( .D(N833), .C(net11959), .Q(c_adr[7]) );
  DFFQX1 c_adr_reg_6_ ( .D(N832), .C(net11959), .Q(c_adr[6]) );
  DFFQX1 c_adr_reg_5_ ( .D(N831), .C(net11959), .Q(c_adr[5]) );
  DFFQX1 c_ptr_reg_4_ ( .D(N846), .C(net11954), .Q(c_ptr[4]) );
  DFFQX1 c_ptr_reg_3_ ( .D(N845), .C(net11954), .Q(c_ptr[3]) );
  DFFQX1 c_ptr_reg_2_ ( .D(N844), .C(net11954), .Q(c_ptr[2]) );
  DFFQX1 c_ptr_reg_0_ ( .D(N842), .C(net11954), .Q(c_ptr[0]) );
  DFFQX1 c_ptr_reg_1_ ( .D(N843), .C(net11954), .Q(c_ptr[1]) );
  DFFQX1 adr_p_reg_14_ ( .D(N868), .C(net11829), .Q(adr_p[14]) );
  DFFQX1 wspp_cnt_reg_5_ ( .D(N800), .C(net11818), .Q(wspp_cnt[5]) );
  DFFQX1 wspp_cnt_reg_3_ ( .D(N798), .C(net11818), .Q(wspp_cnt[3]) );
  DFFQX1 wspp_cnt_reg_4_ ( .D(N799), .C(net11818), .Q(wspp_cnt[4]) );
  DFFQX1 wspp_cnt_reg_6_ ( .D(N801), .C(net11818), .Q(wspp_cnt[6]) );
  DFFQX1 adr_p_reg_13_ ( .D(N867), .C(net11829), .Q(adr_p[13]) );
  DFFNQXL cs_n_reg ( .D(n643), .XC(clk), .Q(cs_n) );
  DFFQX1 re_p_reg ( .D(n647), .C(clk), .Q(pmem_re) );
  DFFQX1 pgm_p_reg ( .D(n644), .C(net11964), .Q(pmem_pgm) );
  DFFQX1 un_hold_reg ( .D(N974), .C(clk), .Q(un_hold) );
  DFFQX1 c_buf_reg_20__2_ ( .D(N641), .C(net11849), .Q(c_buf_20__2_) );
  DFFQX1 c_buf_reg_23__2_ ( .D(N788), .C(net11834), .Q(wr_buf[2]) );
  DFFQX1 c_buf_reg_22__6_ ( .D(N661), .C(net11839), .Q(c_buf_22__6_) );
  DFFQX1 c_buf_reg_22__5_ ( .D(N660), .C(net11839), .Q(c_buf_22__5_) );
  DFFQX1 c_buf_reg_22__4_ ( .D(N659), .C(net11839), .Q(c_buf_22__4_) );
  DFFQX1 c_buf_reg_22__3_ ( .D(N658), .C(net11839), .Q(c_buf_22__3_) );
  DFFQX1 c_buf_reg_22__2_ ( .D(N657), .C(net11839), .Q(c_buf_22__2_) );
  DFFQX1 c_buf_reg_22__1_ ( .D(N656), .C(net11839), .Q(c_buf_22__1_) );
  DFFQX1 c_buf_reg_22__0_ ( .D(N655), .C(net11839), .Q(c_buf_22__0_) );
  DFFQX1 c_buf_reg_21__6_ ( .D(N653), .C(net11844), .Q(c_buf_21__6_) );
  DFFQX1 c_buf_reg_21__5_ ( .D(N652), .C(net11844), .Q(c_buf_21__5_) );
  DFFQX1 c_buf_reg_21__4_ ( .D(N651), .C(net11844), .Q(c_buf_21__4_) );
  DFFQX1 c_buf_reg_21__3_ ( .D(N650), .C(net11844), .Q(c_buf_21__3_) );
  DFFQX1 c_buf_reg_21__2_ ( .D(N649), .C(net11844), .Q(c_buf_21__2_) );
  DFFQX1 c_buf_reg_21__1_ ( .D(N648), .C(net11844), .Q(c_buf_21__1_) );
  DFFQX1 c_buf_reg_21__0_ ( .D(N647), .C(net11844), .Q(c_buf_21__0_) );
  DFFQX1 c_buf_reg_20__6_ ( .D(N645), .C(net11849), .Q(c_buf_20__6_) );
  DFFQX1 c_buf_reg_20__5_ ( .D(N644), .C(net11849), .Q(c_buf_20__5_) );
  DFFQX1 c_buf_reg_20__4_ ( .D(N643), .C(net11849), .Q(c_buf_20__4_) );
  DFFQX1 c_buf_reg_20__3_ ( .D(N642), .C(net11849), .Q(c_buf_20__3_) );
  DFFQX1 c_buf_reg_20__1_ ( .D(N640), .C(net11849), .Q(c_buf_20__1_) );
  DFFQX1 c_buf_reg_20__0_ ( .D(N639), .C(net11849), .Q(c_buf_20__0_) );
  DFFQX1 c_buf_reg_19__6_ ( .D(N637), .C(net11854), .Q(c_buf_19__6_) );
  DFFQX1 c_buf_reg_19__5_ ( .D(N636), .C(net11854), .Q(c_buf_19__5_) );
  DFFQX1 c_buf_reg_19__4_ ( .D(N635), .C(net11854), .Q(c_buf_19__4_) );
  DFFQX1 c_buf_reg_19__3_ ( .D(N634), .C(net11854), .Q(c_buf_19__3_) );
  DFFQX1 c_buf_reg_19__2_ ( .D(N633), .C(net11854), .Q(c_buf_19__2_) );
  DFFQX1 c_buf_reg_19__1_ ( .D(N632), .C(net11854), .Q(c_buf_19__1_) );
  DFFQX1 c_buf_reg_19__0_ ( .D(N631), .C(net11854), .Q(c_buf_19__0_) );
  DFFQX1 c_buf_reg_18__6_ ( .D(N629), .C(net11859), .Q(c_buf_18__6_) );
  DFFQX1 c_buf_reg_18__5_ ( .D(N628), .C(net11859), .Q(c_buf_18__5_) );
  DFFQX1 c_buf_reg_18__4_ ( .D(N627), .C(net11859), .Q(c_buf_18__4_) );
  DFFQX1 c_buf_reg_18__3_ ( .D(N626), .C(net11859), .Q(c_buf_18__3_) );
  DFFQX1 c_buf_reg_18__2_ ( .D(N625), .C(net11859), .Q(c_buf_18__2_) );
  DFFQX1 c_buf_reg_18__1_ ( .D(N624), .C(net11859), .Q(c_buf_18__1_) );
  DFFQX1 c_buf_reg_18__0_ ( .D(N623), .C(net11859), .Q(c_buf_18__0_) );
  DFFQX1 c_buf_reg_17__6_ ( .D(N621), .C(net11864), .Q(c_buf_17__6_) );
  DFFQX1 c_buf_reg_17__5_ ( .D(N620), .C(net11864), .Q(c_buf_17__5_) );
  DFFQX1 c_buf_reg_17__4_ ( .D(N619), .C(net11864), .Q(c_buf_17__4_) );
  DFFQX1 c_buf_reg_17__3_ ( .D(N618), .C(net11864), .Q(c_buf_17__3_) );
  DFFQX1 c_buf_reg_17__2_ ( .D(N617), .C(net11864), .Q(c_buf_17__2_) );
  DFFQX1 c_buf_reg_17__1_ ( .D(N616), .C(net11864), .Q(c_buf_17__1_) );
  DFFQX1 c_buf_reg_17__0_ ( .D(N615), .C(net11864), .Q(c_buf_17__0_) );
  DFFQX1 c_buf_reg_16__6_ ( .D(N613), .C(net11869), .Q(c_buf_16__6_) );
  DFFQX1 c_buf_reg_16__5_ ( .D(N612), .C(net11869), .Q(c_buf_16__5_) );
  DFFQX1 c_buf_reg_16__4_ ( .D(N611), .C(net11869), .Q(c_buf_16__4_) );
  DFFQX1 c_buf_reg_16__2_ ( .D(N609), .C(net11869), .Q(c_buf_16__2_) );
  DFFQX1 c_buf_reg_16__1_ ( .D(N608), .C(net11869), .Q(c_buf_16__1_) );
  DFFQX1 c_buf_reg_16__0_ ( .D(N607), .C(net11869), .Q(c_buf_16__0_) );
  DFFQX1 c_buf_reg_15__5_ ( .D(N604), .C(net11874), .Q(dbg_0f[5]) );
  DFFQX1 c_buf_reg_15__4_ ( .D(N603), .C(net11874), .Q(dbg_0f[4]) );
  DFFQX1 c_buf_reg_15__2_ ( .D(N601), .C(net11874), .Q(dbg_0f[2]) );
  DFFQX1 c_buf_reg_15__1_ ( .D(N600), .C(net11874), .Q(dbg_0f[1]) );
  DFFQX1 c_buf_reg_15__0_ ( .D(N599), .C(net11874), .Q(dbg_0f[0]) );
  DFFQX1 c_buf_reg_14__6_ ( .D(N597), .C(net11879), .Q(dbg_0e[6]) );
  DFFQX1 c_buf_reg_14__5_ ( .D(N596), .C(net11879), .Q(dbg_0e[5]) );
  DFFQX1 c_buf_reg_14__4_ ( .D(N595), .C(net11879), .Q(dbg_0e[4]) );
  DFFQX1 c_buf_reg_14__3_ ( .D(N594), .C(net11879), .Q(dbg_0e[3]) );
  DFFQX1 c_buf_reg_14__2_ ( .D(N593), .C(net11879), .Q(dbg_0e[2]) );
  DFFQX1 c_buf_reg_14__1_ ( .D(N592), .C(net11879), .Q(dbg_0e[1]) );
  DFFQX1 c_buf_reg_14__0_ ( .D(N591), .C(net11879), .Q(dbg_0e[0]) );
  DFFQX1 c_buf_reg_13__5_ ( .D(N588), .C(net11884), .Q(dbg_0d[5]) );
  DFFQX1 c_buf_reg_13__4_ ( .D(N587), .C(net11884), .Q(dbg_0d[4]) );
  DFFQX1 c_buf_reg_13__2_ ( .D(N585), .C(net11884), .Q(dbg_0d[2]) );
  DFFQX1 c_buf_reg_13__1_ ( .D(N584), .C(net11884), .Q(dbg_0d[1]) );
  DFFQX1 c_buf_reg_13__0_ ( .D(N583), .C(net11884), .Q(dbg_0d[0]) );
  DFFQX1 c_buf_reg_12__5_ ( .D(N580), .C(net11889), .Q(dbg_0c[5]) );
  DFFQX1 c_buf_reg_12__4_ ( .D(N579), .C(net11889), .Q(dbg_0c[4]) );
  DFFQX1 c_buf_reg_12__2_ ( .D(N577), .C(net11889), .Q(dbg_0c[2]) );
  DFFQX1 c_buf_reg_12__1_ ( .D(N576), .C(net11889), .Q(dbg_0c[1]) );
  DFFQX1 c_buf_reg_12__0_ ( .D(N575), .C(net11889), .Q(dbg_0c[0]) );
  DFFQX1 c_buf_reg_11__2_ ( .D(N569), .C(net11894), .Q(dbg_0b[2]) );
  DFFQX1 c_buf_reg_11__1_ ( .D(N568), .C(net11894), .Q(dbg_0b[1]) );
  DFFQX1 c_buf_reg_10__2_ ( .D(N561), .C(net11899), .Q(dbg_0a[2]) );
  DFFQX1 c_buf_reg_10__1_ ( .D(N560), .C(net11899), .Q(dbg_0a[1]) );
  DFFQX1 c_buf_reg_9__4_ ( .D(N555), .C(net11904), .Q(dbg_09[4]) );
  DFFQX1 c_buf_reg_9__2_ ( .D(N553), .C(net11904), .Q(dbg_09[2]) );
  DFFQX1 c_buf_reg_9__1_ ( .D(N552), .C(net11904), .Q(dbg_09[1]) );
  DFFQX1 c_buf_reg_9__0_ ( .D(N551), .C(net11904), .Q(dbg_09[0]) );
  DFFQX1 c_buf_reg_8__2_ ( .D(N545), .C(net11909), .Q(dbg_08[2]) );
  DFFQX1 c_buf_reg_8__1_ ( .D(N544), .C(net11909), .Q(dbg_08[1]) );
  DFFQX1 c_buf_reg_7__2_ ( .D(N537), .C(net11914), .Q(dbg_07[2]) );
  DFFQX1 c_buf_reg_7__1_ ( .D(N536), .C(net11914), .Q(dbg_07[1]) );
  DFFQX1 c_buf_reg_6__4_ ( .D(N531), .C(net11919), .Q(dbg_06[4]) );
  DFFQX1 c_buf_reg_6__2_ ( .D(N529), .C(net11919), .Q(dbg_06[2]) );
  DFFQX1 c_buf_reg_5__2_ ( .D(N521), .C(net11924), .Q(dbg_05[2]) );
  DFFQX1 c_buf_reg_4__2_ ( .D(N513), .C(net11929), .Q(dbg_04[2]) );
  DFFQX1 c_buf_reg_3__2_ ( .D(N505), .C(net11934), .Q(dbg_03[2]) );
  DFFQX1 c_buf_reg_2__2_ ( .D(N497), .C(net11939), .Q(dbg_02[2]) );
  DFFQX1 c_buf_reg_1__2_ ( .D(N489), .C(net11944), .Q(dbg_01[2]) );
  DFFQX1 c_buf_reg_6__1_ ( .D(N528), .C(net11919), .Q(dbg_06[1]) );
  DFFQX1 c_buf_reg_5__1_ ( .D(N520), .C(net11924), .Q(dbg_05[1]) );
  DFFQX1 c_buf_reg_4__1_ ( .D(N512), .C(net11929), .Q(dbg_04[1]) );
  DFFQX1 c_buf_reg_3__1_ ( .D(N504), .C(net11934), .Q(dbg_03[1]) );
  DFFQX1 c_buf_reg_2__1_ ( .D(N496), .C(net11939), .Q(dbg_02[1]) );
  DFFQX1 c_buf_reg_1__1_ ( .D(N488), .C(net11944), .Q(dbg_01[1]) );
  DFFQX1 c_buf_reg_6__0_ ( .D(N527), .C(net11919), .Q(dbg_06[0]) );
  DFFQX1 c_buf_reg_0__2_ ( .D(N481), .C(net11949), .Q(rd_buf[2]) );
  DFFQX1 c_buf_reg_0__1_ ( .D(N480), .C(net11949), .Q(rd_buf[1]) );
  DFFQX1 c_buf_reg_23__4_ ( .D(N790), .C(net11834), .Q(wr_buf[4]) );
  DFFQX1 c_buf_reg_23__6_ ( .D(N792), .C(net11834), .Q(wr_buf[6]) );
  DFFQX1 c_buf_reg_23__3_ ( .D(N789), .C(net11834), .Q(wr_buf[3]) );
  DFFQX1 c_buf_reg_23__5_ ( .D(N791), .C(net11834), .Q(wr_buf[5]) );
  DFFQX1 c_buf_reg_23__1_ ( .D(N787), .C(net11834), .Q(wr_buf[1]) );
  DFFQX1 c_buf_reg_23__0_ ( .D(N786), .C(net11834), .Q(wr_buf[0]) );
  DFFQX1 r_twlb_reg_1_ ( .D(n645), .C(clk), .Q(pmem_twlb[1]) );
  DFFQX1 r_twlb_reg_0_ ( .D(n646), .C(clk), .Q(pmem_twlb[0]) );
  DFFQX1 c_buf_reg_16__3_ ( .D(N610), .C(net11869), .Q(c_buf_16__3_) );
  DFFQX1 c_buf_reg_15__6_ ( .D(N605), .C(net11874), .Q(dbg_0f[6]) );
  DFFQX1 c_buf_reg_15__3_ ( .D(N602), .C(net11874), .Q(dbg_0f[3]) );
  DFFQX1 c_buf_reg_13__6_ ( .D(N589), .C(net11884), .Q(dbg_0d[6]) );
  DFFQX1 c_buf_reg_13__3_ ( .D(N586), .C(net11884), .Q(dbg_0d[3]) );
  DFFQX1 c_buf_reg_12__6_ ( .D(N581), .C(net11889), .Q(dbg_0c[6]) );
  DFFQX1 c_buf_reg_12__3_ ( .D(N578), .C(net11889), .Q(dbg_0c[3]) );
  DFFQX1 c_buf_reg_11__6_ ( .D(N573), .C(net11894), .Q(dbg_0b[6]) );
  DFFQX1 c_buf_reg_11__5_ ( .D(N572), .C(net11894), .Q(dbg_0b[5]) );
  DFFQX1 c_buf_reg_11__4_ ( .D(N571), .C(net11894), .Q(dbg_0b[4]) );
  DFFQX1 c_buf_reg_11__3_ ( .D(N570), .C(net11894), .Q(dbg_0b[3]) );
  DFFQX1 c_buf_reg_11__0_ ( .D(N567), .C(net11894), .Q(dbg_0b[0]) );
  DFFQX1 c_buf_reg_10__6_ ( .D(N565), .C(net11899), .Q(dbg_0a[6]) );
  DFFQX1 c_buf_reg_10__5_ ( .D(N564), .C(net11899), .Q(dbg_0a[5]) );
  DFFQX1 c_buf_reg_10__4_ ( .D(N563), .C(net11899), .Q(dbg_0a[4]) );
  DFFQX1 c_buf_reg_10__3_ ( .D(N562), .C(net11899), .Q(dbg_0a[3]) );
  DFFQX1 c_buf_reg_10__0_ ( .D(N559), .C(net11899), .Q(dbg_0a[0]) );
  DFFQX1 c_buf_reg_9__6_ ( .D(N557), .C(net11904), .Q(dbg_09[6]) );
  DFFQX1 c_buf_reg_9__5_ ( .D(N556), .C(net11904), .Q(dbg_09[5]) );
  DFFQX1 c_buf_reg_9__3_ ( .D(N554), .C(net11904), .Q(dbg_09[3]) );
  DFFQX1 c_buf_reg_8__6_ ( .D(N549), .C(net11909), .Q(dbg_08[6]) );
  DFFQX1 c_buf_reg_8__5_ ( .D(N548), .C(net11909), .Q(dbg_08[5]) );
  DFFQX1 c_buf_reg_8__4_ ( .D(N547), .C(net11909), .Q(dbg_08[4]) );
  DFFQX1 c_buf_reg_8__3_ ( .D(N546), .C(net11909), .Q(dbg_08[3]) );
  DFFQX1 c_buf_reg_8__0_ ( .D(N543), .C(net11909), .Q(dbg_08[0]) );
  DFFQX1 c_buf_reg_7__6_ ( .D(N541), .C(net11914), .Q(dbg_07[6]) );
  DFFQX1 c_buf_reg_7__5_ ( .D(N540), .C(net11914), .Q(dbg_07[5]) );
  DFFQX1 c_buf_reg_7__4_ ( .D(N539), .C(net11914), .Q(dbg_07[4]) );
  DFFQX1 c_buf_reg_7__3_ ( .D(N538), .C(net11914), .Q(dbg_07[3]) );
  DFFQX1 c_buf_reg_7__0_ ( .D(N535), .C(net11914), .Q(dbg_07[0]) );
  DFFQX1 c_buf_reg_6__6_ ( .D(N533), .C(net11919), .Q(dbg_06[6]) );
  DFFQX1 c_buf_reg_5__6_ ( .D(N525), .C(net11924), .Q(dbg_05[6]) );
  DFFQX1 c_buf_reg_4__6_ ( .D(N517), .C(net11929), .Q(dbg_04[6]) );
  DFFQX1 c_buf_reg_3__6_ ( .D(N509), .C(net11934), .Q(dbg_03[6]) );
  DFFQX1 c_buf_reg_2__6_ ( .D(N501), .C(net11939), .Q(dbg_02[6]) );
  DFFQX1 c_buf_reg_1__6_ ( .D(N493), .C(net11944), .Q(dbg_01[6]) );
  DFFQX1 c_buf_reg_6__5_ ( .D(N532), .C(net11919), .Q(dbg_06[5]) );
  DFFQX1 c_buf_reg_5__5_ ( .D(N524), .C(net11924), .Q(dbg_05[5]) );
  DFFQX1 c_buf_reg_4__5_ ( .D(N516), .C(net11929), .Q(dbg_04[5]) );
  DFFQX1 c_buf_reg_3__5_ ( .D(N508), .C(net11934), .Q(dbg_03[5]) );
  DFFQX1 c_buf_reg_2__5_ ( .D(N500), .C(net11939), .Q(dbg_02[5]) );
  DFFQX1 c_buf_reg_1__5_ ( .D(N492), .C(net11944), .Q(dbg_01[5]) );
  DFFQX1 c_buf_reg_5__4_ ( .D(N523), .C(net11924), .Q(dbg_05[4]) );
  DFFQX1 c_buf_reg_4__4_ ( .D(N515), .C(net11929), .Q(dbg_04[4]) );
  DFFQX1 c_buf_reg_3__4_ ( .D(N507), .C(net11934), .Q(dbg_03[4]) );
  DFFQX1 c_buf_reg_2__4_ ( .D(N499), .C(net11939), .Q(dbg_02[4]) );
  DFFQX1 c_buf_reg_1__4_ ( .D(N491), .C(net11944), .Q(dbg_01[4]) );
  DFFQX1 c_buf_reg_6__3_ ( .D(N530), .C(net11919), .Q(dbg_06[3]) );
  DFFQX1 c_buf_reg_5__3_ ( .D(N522), .C(net11924), .Q(dbg_05[3]) );
  DFFQX1 c_buf_reg_4__3_ ( .D(N514), .C(net11929), .Q(dbg_04[3]) );
  DFFQX1 c_buf_reg_3__3_ ( .D(N506), .C(net11934), .Q(dbg_03[3]) );
  DFFQX1 c_buf_reg_2__3_ ( .D(N498), .C(net11939), .Q(dbg_02[3]) );
  DFFQX1 c_buf_reg_1__3_ ( .D(N490), .C(net11944), .Q(dbg_01[3]) );
  DFFQX1 c_buf_reg_5__0_ ( .D(N519), .C(net11924), .Q(dbg_05[0]) );
  DFFQX1 c_buf_reg_4__0_ ( .D(N511), .C(net11929), .Q(dbg_04[0]) );
  DFFQX1 c_buf_reg_3__0_ ( .D(N503), .C(net11934), .Q(dbg_03[0]) );
  DFFQX1 c_buf_reg_2__0_ ( .D(N495), .C(net11939), .Q(dbg_02[0]) );
  DFFQX1 c_buf_reg_1__0_ ( .D(N487), .C(net11944), .Q(dbg_01[0]) );
  DFFQX1 c_buf_reg_0__6_ ( .D(N485), .C(net11949), .Q(rd_buf[6]) );
  DFFQX1 c_buf_reg_0__5_ ( .D(N484), .C(net11949), .Q(rd_buf[5]) );
  DFFQX1 c_buf_reg_0__3_ ( .D(N482), .C(net11949), .Q(rd_buf[3]) );
  DFFQX1 c_buf_reg_0__4_ ( .D(N483), .C(net11949), .Q(rd_buf[4]) );
  DFFQX1 c_buf_reg_0__0_ ( .D(N479), .C(net11949), .Q(rd_buf[0]) );
  DFFQX1 cs_ft_reg_3_ ( .D(N824), .C(net11964), .Q(cs_ft[3]) );
  DFFQX1 r_rdy_reg ( .D(n648), .C(clk), .Q(r_rdy) );
  DFFQX1 cs_ft_reg_1_ ( .D(N822), .C(net11964), .Q(cs_ft[1]) );
  DFFQX1 cs_ft_reg_2_ ( .D(N823), .C(net11964), .Q(cs_ft[2]) );
  DFFQX1 c_buf_reg_22__7_ ( .D(N662), .C(net11839), .Q(c_buf_22__7_) );
  DFFQX1 c_buf_reg_21__7_ ( .D(N654), .C(net11844), .Q(c_buf_21__7_) );
  DFFQX1 c_buf_reg_20__7_ ( .D(N646), .C(net11849), .Q(c_buf_20__7_) );
  DFFQX1 c_buf_reg_19__7_ ( .D(N638), .C(net11854), .Q(c_buf_19__7_) );
  DFFQX1 c_buf_reg_18__7_ ( .D(N630), .C(net11859), .Q(c_buf_18__7_) );
  DFFQX1 c_buf_reg_17__7_ ( .D(N622), .C(net11864), .Q(c_buf_17__7_) );
  DFFQX1 c_buf_reg_16__7_ ( .D(N614), .C(net11869), .Q(c_buf_16__7_) );
  DFFQX1 c_buf_reg_15__7_ ( .D(N606), .C(net11874), .Q(dbg_0f[7]) );
  DFFQX1 c_buf_reg_14__7_ ( .D(N598), .C(net11879), .Q(dbg_0e[7]) );
  DFFQX1 c_buf_reg_13__7_ ( .D(N590), .C(net11884), .Q(dbg_0d[7]) );
  DFFQX1 c_buf_reg_12__7_ ( .D(N582), .C(net11889), .Q(dbg_0c[7]) );
  DFFQX1 c_buf_reg_11__7_ ( .D(N574), .C(net11894), .Q(dbg_0b[7]) );
  DFFQX1 c_buf_reg_10__7_ ( .D(N566), .C(net11899), .Q(dbg_0a[7]) );
  DFFQX1 c_buf_reg_9__7_ ( .D(N558), .C(net11904), .Q(dbg_09[7]) );
  DFFQX1 c_buf_reg_8__7_ ( .D(N550), .C(net11909), .Q(dbg_08[7]) );
  DFFQX1 c_buf_reg_7__7_ ( .D(N542), .C(net11914), .Q(dbg_07[7]) );
  DFFQX1 c_buf_reg_6__7_ ( .D(N534), .C(net11919), .Q(dbg_06[7]) );
  DFFQX1 c_buf_reg_5__7_ ( .D(N526), .C(net11924), .Q(dbg_05[7]) );
  DFFQX1 c_buf_reg_4__7_ ( .D(N518), .C(net11929), .Q(dbg_04[7]) );
  DFFQX1 c_buf_reg_3__7_ ( .D(N510), .C(net11934), .Q(dbg_03[7]) );
  DFFQX1 c_buf_reg_2__7_ ( .D(N502), .C(net11939), .Q(dbg_02[7]) );
  DFFQX1 c_buf_reg_1__7_ ( .D(N494), .C(net11944), .Q(dbg_01[7]) );
  DFFQX1 c_buf_reg_0__7_ ( .D(N486), .C(net11949), .Q(rd_buf[7]) );
  DFFQX1 c_buf_reg_23__7_ ( .D(N793), .C(net11834), .Q(wr_buf[7]) );
  DFFQX1 cs_ft_reg_0_ ( .D(N821), .C(net11964), .Q(cs_ft[0]) );
  DFFQX1 c_adr_reg_4_ ( .D(N830), .C(net11959), .Q(c_adr[4]) );
  DFFQX1 c_adr_reg_3_ ( .D(N829), .C(net11959), .Q(c_adr[3]) );
  DFFQX4 adr_p_reg_6_ ( .D(N860), .C(net11829), .Q(pmem_a[9]) );
  DFFQX4 a_bit_reg_0_ ( .D(N757), .C(net11824), .Q(pmem_a[6]) );
  DFFQX4 adr_p_reg_8_ ( .D(N862), .C(net11829), .Q(pmem_a[11]) );
  DFFQX4 adr_p_reg_9_ ( .D(N863), .C(net11829), .Q(pmem_a[12]) );
  DFFQX4 adr_p_reg_7_ ( .D(N861), .C(net11829), .Q(pmem_a[10]) );
  DFFQX4 adr_p_reg_12_ ( .D(N866), .C(net11829), .Q(pmem_a[15]) );
  DFFQX4 adr_p_reg_11_ ( .D(N865), .C(net11829), .Q(pmem_a[14]) );
  DFFQX4 adr_p_reg_10_ ( .D(N864), .C(net11829), .Q(pmem_a[13]) );
  DFFQX4 adr_p_reg_0_ ( .D(N854), .C(net11829), .Q(pmem_a[0]) );
  DFFQX4 a_bit_reg_1_ ( .D(N758), .C(net11824), .Q(pmem_a[7]) );
  DFFQX4 adr_p_reg_4_ ( .D(N858), .C(net11829), .Q(pmem_a[4]) );
  DFFQX4 adr_p_reg_3_ ( .D(N857), .C(net11829), .Q(pmem_a[3]) );
  DFFQX4 adr_p_reg_2_ ( .D(N856), .C(net11829), .Q(pmem_a[2]) );
  DFFQX4 adr_p_reg_5_ ( .D(N859), .C(net11829), .Q(pmem_a[5]) );
  DFFQX4 adr_p_reg_1_ ( .D(N855), .C(net11829), .Q(pmem_a[1]) );
  DFFQX4 a_bit_reg_2_ ( .D(N759), .C(net11824), .Q(pmem_a[8]) );
  DFFQX1 c_adr_reg_2_ ( .D(N828), .C(net11959), .Q(c_adr[2]) );
  DFFQX1 c_adr_reg_1_ ( .D(N827), .C(net11959), .Q(c_adr[1]) );
  DFFQX1 c_adr_reg_0_ ( .D(N826), .C(net11959), .Q(c_adr[0]) );
  INVX1 U3 ( .A(c_adr[2]), .Y(n360) );
  INVX1 U4 ( .A(c_adr[1]), .Y(n359) );
  OA222X1 U5 ( .A(memaddr_c[4]), .B(n163), .C(n162), .D(n161), .E(memaddr_c[5]), .F(n160), .Y(n167) );
  XNOR3X1 U6 ( .A(memaddr[4]), .B(c_adr[4]), .C(n30), .Y(n396) );
  NAND5XL U7 ( .A(n575), .B(n574), .C(n573), .D(n572), .E(n571), .Y(o_inst[3])
         );
  AND3X1 U8 ( .A(n128), .B(n130), .C(n127), .Y(n129) );
  NAND5XL U9 ( .A(n419), .B(n418), .C(n417), .D(n416), .E(n415), .Y(o_inst[7])
         );
  INVX1 U10 ( .A(n835), .Y(n83) );
  NAND21X1 U11 ( .B(pwrdn_rst), .A(n85), .Y(n835) );
  XNOR2XL U12 ( .A(n137), .B(c_adr[14]), .Y(n1) );
  INVXL U13 ( .A(n344), .Y(n2) );
  INVXL U14 ( .A(n2), .Y(n3) );
  NAND3XL U15 ( .A(pmem_a[6]), .B(n918), .C(pmem_a[7]), .Y(n916) );
  INVX1 U16 ( .A(n357), .Y(n4) );
  INVX1 U17 ( .A(n357), .Y(n5) );
  INVX1 U18 ( .A(n340), .Y(n6) );
  INVX1 U19 ( .A(n426), .Y(n7) );
  INVX1 U20 ( .A(n426), .Y(n8) );
  INVX1 U21 ( .A(n341), .Y(n9) );
  INVX1 U22 ( .A(n465), .Y(n10) );
  INVX1 U23 ( .A(n465), .Y(n11) );
  INVX1 U24 ( .A(n503), .Y(n12) );
  INVX1 U25 ( .A(n503), .Y(n13) );
  INVX1 U26 ( .A(n339), .Y(n14) );
  INVX1 U27 ( .A(n542), .Y(n15) );
  INVX1 U28 ( .A(n542), .Y(n16) );
  INVX1 U29 ( .A(n746), .Y(n17) );
  INVX1 U30 ( .A(n581), .Y(n18) );
  INVX1 U31 ( .A(n581), .Y(n19) );
  INVX1 U32 ( .A(n894), .Y(n20) );
  INVX1 U33 ( .A(n784), .Y(n21) );
  INVX1 U34 ( .A(n621), .Y(n22) );
  INVX1 U35 ( .A(n621), .Y(n23) );
  BUFX3 U36 ( .A(n292), .Y(n24) );
  INVX1 U37 ( .A(n848), .Y(n25) );
  INVX1 U38 ( .A(n782), .Y(n26) );
  INVX1 U39 ( .A(n782), .Y(n27) );
  INVX1 U40 ( .A(n674), .Y(n28) );
  INVX1 U41 ( .A(n674), .Y(n29) );
  NAND21XL U42 ( .B(n152), .A(memaddr_c[2]), .Y(n214) );
  XOR2XL U43 ( .A(memaddr_c[2]), .B(n232), .Y(n233) );
  NAND2XL U44 ( .A(n165), .B(memaddr_c[6]), .Y(n208) );
  OR2X1 U45 ( .A(n370), .B(n407), .Y(n678) );
  NAND21X1 U46 ( .B(n376), .A(n375), .Y(n691) );
  INVX1 U47 ( .A(n376), .Y(n374) );
  NAND21XL U48 ( .B(n81), .A(n746), .Y(n757) );
  AO21XL U49 ( .B(n354), .C(n327), .A(n840), .Y(n823) );
  AND4XL U50 ( .A(o_inst[4]), .B(o_inst[3]), .C(o_inst[2]), .D(o_inst[1]), .Y(
        n734) );
  NAND5XL U51 ( .A(n498), .B(n497), .C(n496), .D(n495), .E(n494), .Y(o_inst[5]) );
  NAND5XL U52 ( .A(n459), .B(n458), .C(n457), .D(n456), .E(n455), .Y(o_inst[6]) );
  INVXL U53 ( .A(n835), .Y(n84) );
  INVX1 U54 ( .A(n386), .Y(n392) );
  OAI21BBX1 U55 ( .A(n158), .B(n157), .C(n205), .Y(n161) );
  NAND21XL U56 ( .B(n153), .A(memaddr_c[1]), .Y(n197) );
  OAI22XL U57 ( .A(memaddr_c[2]), .B(n360), .C(memaddr_c[3]), .D(n362), .Y(n47) );
  NAND21XL U58 ( .B(n164), .A(memaddr_c[5]), .Y(n204) );
  XOR2XL U59 ( .A(memaddr_c[1]), .B(n238), .Y(n251) );
  AND3X1 U60 ( .A(pmem_clk[0]), .B(n33), .C(n830), .Y(n828) );
  XNOR3XL U61 ( .A(memaddr[3]), .B(c_adr[3]), .C(n377), .Y(n53) );
  XOR3XL U62 ( .A(memaddr[2]), .B(c_adr[2]), .C(n363), .Y(n390) );
  AOI21X1 U63 ( .B(memaddr[3]), .C(n362), .A(n361), .Y(n30) );
  AOI21AXL U64 ( .B(memaddr[0]), .C(n364), .A(n365), .Y(n31) );
  NOR43XL U65 ( .B(n84), .C(r_rdy), .D(n751), .A(n334), .Y(n330) );
  XOR2XL U66 ( .A(n765), .B(c_adr[3]), .Y(n246) );
  NAND21XL U67 ( .B(c_adr[3]), .A(n765), .Y(n221) );
  NAND21XL U68 ( .B(n765), .A(c_adr[3]), .Y(n133) );
  INVX1 U69 ( .A(n782), .Y(n777) );
  INVX1 U70 ( .A(n757), .Y(n766) );
  NAND21X1 U71 ( .B(n336), .A(n782), .Y(n344) );
  NAND21X1 U72 ( .B(n757), .A(n62), .Y(n782) );
  NAND32X1 U73 ( .B(n786), .C(n785), .A(n784), .Y(N853) );
  AOI21X1 U74 ( .B(n810), .C(we_twlb), .A(N853), .Y(n32) );
  INVX1 U75 ( .A(n784), .Y(n749) );
  INVX1 U76 ( .A(n320), .Y(n819) );
  AO21X1 U77 ( .B(n786), .C(n755), .A(n785), .Y(n93) );
  INVX1 U78 ( .A(n308), .Y(n74) );
  INVX1 U79 ( .A(n308), .Y(n67) );
  INVX1 U80 ( .A(n308), .Y(n76) );
  INVX1 U81 ( .A(n80), .Y(n69) );
  INVX1 U82 ( .A(n80), .Y(n63) );
  INVX1 U83 ( .A(n80), .Y(n78) );
  INVX1 U84 ( .A(n308), .Y(n71) );
  INVX1 U85 ( .A(n308), .Y(n64) );
  INVX1 U86 ( .A(n80), .Y(n73) );
  INVX1 U87 ( .A(n80), .Y(n66) );
  INVX1 U88 ( .A(n80), .Y(n77) );
  INVX1 U89 ( .A(n308), .Y(n75) );
  INVX1 U90 ( .A(n80), .Y(n72) );
  INVX1 U91 ( .A(n80), .Y(n70) );
  INVX1 U92 ( .A(n308), .Y(n68) );
  INVX1 U93 ( .A(n80), .Y(n65) );
  INVX1 U94 ( .A(n308), .Y(n79) );
  INVX1 U95 ( .A(n740), .Y(n754) );
  NAND21X1 U96 ( .B(n794), .A(n810), .Y(n740) );
  INVX1 U97 ( .A(n823), .Y(n818) );
  INVX1 U98 ( .A(n800), .Y(n790) );
  INVX1 U99 ( .A(n318), .Y(n789) );
  NAND21X1 U100 ( .B(n813), .A(n844), .Y(n318) );
  INVX1 U101 ( .A(n83), .Y(n81) );
  NOR3XL U102 ( .A(n827), .B(n81), .C(n826), .Y(n33) );
  NAND2X1 U103 ( .A(n857), .B(n84), .Y(n840) );
  INVX1 U104 ( .A(n83), .Y(n82) );
  NAND21X1 U105 ( .B(n405), .A(n400), .Y(n711) );
  NAND21X1 U106 ( .B(n407), .A(n374), .Y(n693) );
  NAND21X1 U107 ( .B(n399), .A(n406), .Y(n717) );
  NAND21X1 U108 ( .B(n404), .A(n406), .Y(n723) );
  NAND21X1 U109 ( .B(n370), .A(n375), .Y(n687) );
  OR2X1 U110 ( .A(n370), .B(n399), .Y(n681) );
  NAND21X1 U111 ( .B(n405), .A(n406), .Y(n721) );
  NAND21X1 U112 ( .B(n399), .A(n374), .Y(n685) );
  NAND21X1 U113 ( .B(n407), .A(n400), .Y(n715) );
  OR2X1 U114 ( .A(n370), .B(n405), .Y(n680) );
  NAND21X1 U115 ( .B(n405), .A(n374), .Y(n683) );
  NAND21X1 U116 ( .B(n399), .A(n400), .Y(n707) );
  NAND21X1 U117 ( .B(n407), .A(n406), .Y(n719) );
  NAND21X1 U118 ( .B(n404), .A(n400), .Y(n713) );
  NAND21X1 U119 ( .B(n405), .A(n382), .Y(n699) );
  NAND21X1 U120 ( .B(n407), .A(n392), .Y(n705) );
  NAND21X1 U121 ( .B(n407), .A(n382), .Y(n697) );
  NAND21X1 U122 ( .B(n399), .A(n392), .Y(n703) );
  NAND21X1 U123 ( .B(n404), .A(n392), .Y(n709) );
  NAND21X1 U124 ( .B(n405), .A(n392), .Y(n701) );
  NAND21X1 U125 ( .B(n399), .A(n382), .Y(n689) );
  NAND21X1 U126 ( .B(n404), .A(n382), .Y(n695) );
  INVX1 U127 ( .A(n404), .Y(n375) );
  NAND21X1 U128 ( .B(n751), .A(n62), .Y(n784) );
  NAND6XL U129 ( .A(n215), .B(n214), .C(n213), .D(n212), .E(n211), .F(n210), 
        .Y(n755) );
  OA21X1 U130 ( .B(n224), .C(n198), .A(n197), .Y(n213) );
  AND4X1 U131 ( .A(n209), .B(n208), .C(n207), .D(n206), .Y(n210) );
  AND4X1 U132 ( .A(n49), .B(n205), .C(n204), .D(n203), .Y(n211) );
  OAI211X1 U133 ( .C(n291), .D(n329), .A(n321), .B(n849), .Y(n322) );
  AND4X1 U134 ( .A(n202), .B(n201), .C(n200), .D(n199), .Y(n212) );
  INVX1 U135 ( .A(n80), .Y(n62) );
  INVX1 U136 ( .A(n676), .Y(n80) );
  NAND21X1 U137 ( .B(n332), .A(n849), .Y(n320) );
  INVX1 U138 ( .A(n279), .Y(n336) );
  NAND21X1 U139 ( .B(n757), .A(n750), .Y(n279) );
  NAND42X1 U140 ( .C(n754), .D(n753), .A(n752), .B(n801), .Y(n785) );
  NAND21X1 U141 ( .B(n751), .A(n750), .Y(n752) );
  AO21X1 U142 ( .B(n780), .C(n775), .A(n777), .Y(N894) );
  AO21X1 U143 ( .B(n48), .C(n775), .A(n26), .Y(N886) );
  AO21X1 U144 ( .B(n763), .C(n775), .A(n27), .Y(N882) );
  AO21X1 U145 ( .B(n761), .C(n775), .A(n777), .Y(N878) );
  NAND2X1 U146 ( .A(n747), .B(n84), .Y(n753) );
  INVX1 U147 ( .A(n214), .Y(n154) );
  NAND21X1 U148 ( .B(n301), .A(n747), .Y(n292) );
  INVX1 U149 ( .A(n208), .Y(n168) );
  INVX1 U150 ( .A(n105), .Y(n107) );
  INVX1 U151 ( .A(n111), .Y(n109) );
  INVX1 U152 ( .A(n302), .Y(n786) );
  NAND21X1 U153 ( .B(n332), .A(n301), .Y(n302) );
  INVX1 U154 ( .A(n204), .Y(n166) );
  NAND32X1 U155 ( .B(n327), .C(n795), .A(n806), .Y(n800) );
  INVX1 U156 ( .A(n327), .Y(n813) );
  INVX1 U157 ( .A(n841), .Y(n810) );
  INVX1 U158 ( .A(n741), .Y(n743) );
  INVX1 U159 ( .A(n795), .Y(n844) );
  INVX1 U160 ( .A(n796), .Y(n816) );
  NAND21X1 U161 ( .B(n795), .A(n794), .Y(n796) );
  INVX1 U162 ( .A(n341), .Y(n342) );
  INVX1 U163 ( .A(n340), .Y(n343) );
  INVX1 U164 ( .A(srst), .Y(n85) );
  INVX1 U165 ( .A(n788), .Y(n827) );
  INVX1 U166 ( .A(n825), .Y(n832) );
  INVX1 U167 ( .A(n806), .Y(n794) );
  INVX1 U168 ( .A(n159), .Y(n139) );
  INVX1 U169 ( .A(n143), .Y(n147) );
  INVX1 U170 ( .A(n152), .Y(n146) );
  INVX1 U171 ( .A(n252), .Y(n253) );
  INVX1 U172 ( .A(n265), .Y(n266) );
  INVX1 U173 ( .A(n255), .Y(n256) );
  INVX1 U174 ( .A(n751), .Y(n746) );
  INVX1 U175 ( .A(n742), .Y(n301) );
  INVX1 U176 ( .A(n352), .Y(n616) );
  NAND21X1 U177 ( .B(n833), .A(n667), .Y(n352) );
  INVX1 U178 ( .A(n421), .Y(n846) );
  INVX1 U179 ( .A(n305), .Y(n283) );
  OAI31XL U180 ( .A(n839), .B(pmem_csb), .C(n840), .D(n838), .Y(n643) );
  AO21X1 U181 ( .B(n837), .C(n836), .A(n82), .Y(n838) );
  NAND21X1 U182 ( .B(n396), .A(n390), .Y(n376) );
  INVX1 U183 ( .A(n391), .Y(n400) );
  NAND32X1 U184 ( .B(n390), .C(n53), .A(n396), .Y(n391) );
  INVX1 U185 ( .A(n398), .Y(n406) );
  NAND32X1 U186 ( .B(n397), .C(n53), .A(n396), .Y(n398) );
  NAND21X1 U187 ( .B(n396), .A(n397), .Y(n370) );
  AND4X1 U188 ( .A(n414), .B(n413), .C(n412), .D(n411), .Y(n415) );
  OA222X1 U189 ( .A(n705), .B(n389), .C(n703), .D(n388), .E(n701), .F(n387), 
        .Y(n414) );
  OA222X1 U190 ( .A(n711), .B(n395), .C(n709), .D(n394), .E(n707), .F(n393), 
        .Y(n413) );
  OA222X1 U191 ( .A(n717), .B(n403), .C(n715), .D(n402), .E(n713), .F(n401), 
        .Y(n412) );
  OA222X1 U192 ( .A(n699), .B(n385), .C(n697), .D(n384), .E(n695), .F(n383), 
        .Y(n416) );
  OA222X1 U193 ( .A(n681), .B(n422), .C(n680), .D(n368), .E(n678), .F(n367), 
        .Y(n419) );
  OA222X1 U194 ( .A(n687), .B(n373), .C(n685), .D(n372), .E(n683), .F(n371), 
        .Y(n418) );
  NAND21X1 U195 ( .B(n366), .A(n31), .Y(n405) );
  NAND21X1 U196 ( .B(n31), .A(n366), .Y(n407) );
  NAND21X1 U197 ( .B(n31), .A(n369), .Y(n399) );
  NAND21X1 U198 ( .B(n369), .A(n31), .Y(n404) );
  INVX1 U199 ( .A(n390), .Y(n397) );
  INVX1 U200 ( .A(n366), .Y(n369) );
  AND4X1 U201 ( .A(n570), .B(n569), .C(n568), .D(n567), .Y(n571) );
  OA222X1 U202 ( .A(n705), .B(n557), .C(n703), .D(n556), .E(n701), .F(n555), 
        .Y(n570) );
  OA222X1 U203 ( .A(n711), .B(n560), .C(n709), .D(n559), .E(n707), .F(n558), 
        .Y(n569) );
  OA222X1 U204 ( .A(n717), .B(n563), .C(n715), .D(n562), .E(n713), .F(n561), 
        .Y(n568) );
  AND4X1 U205 ( .A(n454), .B(n453), .C(n452), .D(n451), .Y(n455) );
  OA222X1 U206 ( .A(n705), .B(n441), .C(n703), .D(n440), .E(n701), .F(n439), 
        .Y(n454) );
  OA222X1 U207 ( .A(n711), .B(n444), .C(n709), .D(n443), .E(n707), .F(n442), 
        .Y(n453) );
  OA222X1 U208 ( .A(n717), .B(n447), .C(n715), .D(n446), .E(n713), .F(n445), 
        .Y(n452) );
  AND4X1 U209 ( .A(n531), .B(n530), .C(n529), .D(n528), .Y(n532) );
  OA222X1 U210 ( .A(n705), .B(n518), .C(n703), .D(n517), .E(n701), .F(n516), 
        .Y(n531) );
  OA222X1 U211 ( .A(n711), .B(n521), .C(n709), .D(n520), .E(n707), .F(n519), 
        .Y(n530) );
  OA222X1 U212 ( .A(n717), .B(n524), .C(n715), .D(n523), .E(n713), .F(n522), 
        .Y(n529) );
  AND4X1 U213 ( .A(n727), .B(n726), .C(n725), .D(n724), .Y(n728) );
  OA222X1 U214 ( .A(n705), .B(n704), .C(n703), .D(n702), .E(n701), .F(n700), 
        .Y(n727) );
  OA222X1 U215 ( .A(n711), .B(n710), .C(n709), .D(n708), .E(n707), .F(n706), 
        .Y(n726) );
  OA222X1 U216 ( .A(n717), .B(n716), .C(n715), .D(n714), .E(n713), .F(n712), 
        .Y(n725) );
  AND4X1 U217 ( .A(n493), .B(n492), .C(n491), .D(n490), .Y(n494) );
  OA222X1 U218 ( .A(n705), .B(n480), .C(n703), .D(n479), .E(n701), .F(n478), 
        .Y(n493) );
  OA222X1 U219 ( .A(n711), .B(n483), .C(n709), .D(n482), .E(n707), .F(n481), 
        .Y(n492) );
  OA222X1 U220 ( .A(n717), .B(n486), .C(n715), .D(n485), .E(n713), .F(n484), 
        .Y(n491) );
  AND4X1 U221 ( .A(n609), .B(n608), .C(n607), .D(n606), .Y(n610) );
  OA222X1 U222 ( .A(n705), .B(n596), .C(n703), .D(n595), .E(n701), .F(n594), 
        .Y(n609) );
  OA222X1 U223 ( .A(n711), .B(n599), .C(n709), .D(n598), .E(n707), .F(n597), 
        .Y(n608) );
  OA222X1 U224 ( .A(n717), .B(n602), .C(n715), .D(n601), .E(n713), .F(n600), 
        .Y(n607) );
  AND4X1 U225 ( .A(n660), .B(n659), .C(n658), .D(n657), .Y(n661) );
  OA222X1 U226 ( .A(n705), .B(n636), .C(n703), .D(n635), .E(n701), .F(n634), 
        .Y(n660) );
  OA222X1 U227 ( .A(n711), .B(n639), .C(n709), .D(n638), .E(n707), .F(n637), 
        .Y(n659) );
  OA222X1 U228 ( .A(n717), .B(n653), .C(n715), .D(n652), .E(n713), .F(n640), 
        .Y(n658) );
  INVX1 U229 ( .A(n378), .Y(n382) );
  NAND21X1 U230 ( .B(n390), .A(n53), .Y(n378) );
  NAND21X1 U231 ( .B(n397), .A(n53), .Y(n386) );
  OA222X1 U232 ( .A(n699), .B(n477), .C(n697), .D(n476), .E(n695), .F(n475), 
        .Y(n495) );
  OA222X1 U233 ( .A(n687), .B(n471), .C(n685), .D(n470), .E(n683), .F(n469), 
        .Y(n497) );
  OA222X1 U234 ( .A(n681), .B(n499), .C(n680), .D(n468), .E(n678), .F(n467), 
        .Y(n498) );
  OA222X1 U235 ( .A(n699), .B(n438), .C(n697), .D(n437), .E(n695), .F(n436), 
        .Y(n456) );
  OA222X1 U236 ( .A(n687), .B(n432), .C(n685), .D(n431), .E(n683), .F(n430), 
        .Y(n458) );
  OA222X1 U237 ( .A(n681), .B(n461), .C(n680), .D(n429), .E(n678), .F(n428), 
        .Y(n459) );
  NAND5XL U238 ( .A(n665), .B(n664), .C(n663), .D(n662), .E(n661), .Y(
        o_inst[1]) );
  OA222X1 U239 ( .A(n699), .B(n633), .C(n697), .D(n632), .E(n695), .F(n631), 
        .Y(n662) );
  OA222X1 U240 ( .A(n687), .B(n627), .C(n685), .D(n626), .E(n683), .F(n625), 
        .Y(n664) );
  OA222X1 U241 ( .A(n681), .B(n668), .C(n680), .D(n624), .E(n678), .F(n623), 
        .Y(n665) );
  NAND5XL U242 ( .A(n614), .B(n613), .C(n612), .D(n611), .E(n610), .Y(
        o_inst[2]) );
  OA222X1 U243 ( .A(n699), .B(n593), .C(n697), .D(n592), .E(n695), .F(n591), 
        .Y(n611) );
  OA222X1 U244 ( .A(n687), .B(n587), .C(n685), .D(n586), .E(n683), .F(n585), 
        .Y(n613) );
  OA222X1 U245 ( .A(n681), .B(n617), .C(n680), .D(n584), .E(n678), .F(n583), 
        .Y(n614) );
  NAND5XL U246 ( .A(n536), .B(n535), .C(n534), .D(n533), .E(n532), .Y(
        o_inst[4]) );
  OA222X1 U247 ( .A(n699), .B(n515), .C(n697), .D(n514), .E(n695), .F(n513), 
        .Y(n533) );
  OA222X1 U248 ( .A(n687), .B(n509), .C(n685), .D(n508), .E(n683), .F(n507), 
        .Y(n535) );
  OA222X1 U249 ( .A(n681), .B(n538), .C(n680), .D(n506), .E(n678), .F(n505), 
        .Y(n536) );
  NAND5XL U250 ( .A(n732), .B(n731), .C(n730), .D(n729), .E(n728), .Y(
        o_inst[0]) );
  OA222X1 U251 ( .A(n699), .B(n698), .C(n697), .D(n696), .E(n695), .F(n694), 
        .Y(n729) );
  OA222X1 U252 ( .A(n687), .B(n686), .C(n685), .D(n684), .E(n683), .F(n682), 
        .Y(n731) );
  OA222X1 U253 ( .A(n681), .B(n791), .C(n680), .D(n679), .E(n678), .F(n677), 
        .Y(n732) );
  OA222X1 U254 ( .A(n699), .B(n554), .C(n697), .D(n553), .E(n695), .F(n552), 
        .Y(n572) );
  OA222X1 U255 ( .A(n687), .B(n548), .C(n685), .D(n547), .E(n683), .F(n546), 
        .Y(n574) );
  OA222X1 U256 ( .A(n681), .B(n577), .C(n680), .D(n545), .E(n678), .F(n544), 
        .Y(n575) );
  NAND32X1 U257 ( .B(n287), .C(n298), .A(n300), .Y(n857) );
  INVX1 U258 ( .A(n156), .Y(n163) );
  INVX1 U259 ( .A(n164), .Y(n160) );
  INVX1 U260 ( .A(n203), .Y(n162) );
  INVX1 U261 ( .A(n153), .Y(n151) );
  OA222X1 U262 ( .A(memaddr_c[11]), .B(n184), .C(n183), .D(n182), .E(
        memaddr_c[10]), .F(n181), .Y(n187) );
  INVX1 U263 ( .A(n201), .Y(n183) );
  AO21X1 U264 ( .B(n180), .C(n179), .A(n178), .Y(n182) );
  INVX1 U265 ( .A(n207), .Y(n178) );
  NAND21X1 U266 ( .B(n192), .A(n49), .Y(n200) );
  OA222X1 U267 ( .A(memaddr_c[13]), .B(n191), .C(n190), .D(n189), .E(
        memaddr_c[12]), .F(n188), .Y(n192) );
  INVX1 U268 ( .A(n199), .Y(n190) );
  NAND21X1 U269 ( .B(n187), .A(n202), .Y(n189) );
  NAND32X1 U270 ( .B(n155), .C(n154), .A(n197), .Y(n157) );
  INVX1 U271 ( .A(n308), .Y(n676) );
  AOI32X1 U272 ( .A(n209), .B(n175), .C(n206), .D(n174), .E(n173), .Y(n180) );
  INVX1 U273 ( .A(memaddr_c[8]), .Y(n173) );
  AO21X1 U274 ( .B(n60), .C(n170), .A(n169), .Y(n175) );
  INVX1 U275 ( .A(n288), .Y(n329) );
  NAND32X1 U276 ( .B(n830), .C(n755), .A(n300), .Y(n288) );
  OAI21BBX1 U277 ( .A(N432), .B(n21), .C(n34), .Y(N827) );
  AOI21XL U278 ( .B(memaddr_c[1]), .C(n24), .A(n82), .Y(n34) );
  OAI21BBX1 U279 ( .A(N433), .B(n21), .C(n35), .Y(N828) );
  AOI21XL U280 ( .B(memaddr_c[2]), .C(n24), .A(n82), .Y(n35) );
  OAI21BBX1 U281 ( .A(N436), .B(n749), .C(n36), .Y(N831) );
  AOI21XL U282 ( .B(memaddr_c[5]), .C(n292), .A(n82), .Y(n36) );
  OAI21BBX1 U283 ( .A(N438), .B(n749), .C(n37), .Y(N833) );
  AOI21XL U284 ( .B(memaddr_c[7]), .C(n292), .A(n82), .Y(n37) );
  OAI21BBX1 U285 ( .A(N439), .B(n749), .C(n38), .Y(N834) );
  AOI21XL U286 ( .B(memaddr_c[8]), .C(n292), .A(n82), .Y(n38) );
  OAI21BBX1 U287 ( .A(N440), .B(n749), .C(n39), .Y(N835) );
  AOI21X1 U288 ( .B(memaddr_c[9]), .C(n292), .A(n835), .Y(n39) );
  OAI21BBX1 U289 ( .A(N441), .B(n21), .C(n40), .Y(N836) );
  AOI21X1 U290 ( .B(memaddr_c[10]), .C(n292), .A(n835), .Y(n40) );
  OAI21BBX1 U291 ( .A(N442), .B(n749), .C(n41), .Y(N837) );
  AOI21X1 U292 ( .B(memaddr_c[11]), .C(n292), .A(n835), .Y(n41) );
  OAI21BBX1 U293 ( .A(N443), .B(n749), .C(n42), .Y(N838) );
  AOI21X1 U294 ( .B(memaddr_c[12]), .C(n292), .A(n835), .Y(n42) );
  OAI21BBX1 U295 ( .A(N444), .B(n749), .C(n43), .Y(N839) );
  AOI21XL U296 ( .B(memaddr_c[13]), .C(n292), .A(n81), .Y(n43) );
  OAI21BBX1 U297 ( .A(N434), .B(n749), .C(n44), .Y(N829) );
  AOI21XL U298 ( .B(memaddr_c[3]), .C(n292), .A(n82), .Y(n44) );
  OAI21BBX1 U299 ( .A(N435), .B(n21), .C(n45), .Y(N830) );
  AOI21XL U300 ( .B(memaddr_c[4]), .C(n24), .A(n82), .Y(n45) );
  OAI21BBX1 U301 ( .A(N437), .B(n21), .C(n46), .Y(N832) );
  AOI21XL U302 ( .B(memaddr_c[6]), .C(n24), .A(n82), .Y(n46) );
  AO21X1 U303 ( .B(n778), .C(n780), .A(n26), .Y(N896) );
  AO21X1 U304 ( .B(n776), .C(n780), .A(n27), .Y(N895) );
  AO21X1 U305 ( .B(n771), .C(n781), .A(n777), .Y(N893) );
  AO21X1 U306 ( .B(n771), .C(n778), .A(n26), .Y(N892) );
  AO21X1 U307 ( .B(n771), .C(n776), .A(n27), .Y(N891) );
  AO21X1 U308 ( .B(n771), .C(n775), .A(n777), .Y(N890) );
  AO21X1 U309 ( .B(n48), .C(n781), .A(n26), .Y(N889) );
  AO21X1 U310 ( .B(n48), .C(n778), .A(n27), .Y(N888) );
  AO21X1 U311 ( .B(n48), .C(n776), .A(n777), .Y(N887) );
  AO21X1 U312 ( .B(n763), .C(n781), .A(n26), .Y(N885) );
  AO21X1 U313 ( .B(n763), .C(n778), .A(n27), .Y(N884) );
  AO21X1 U314 ( .B(n763), .C(n776), .A(n777), .Y(N883) );
  AO21X1 U315 ( .B(n761), .C(n781), .A(n26), .Y(N881) );
  AO21X1 U316 ( .B(n761), .C(n778), .A(n27), .Y(N880) );
  AO21X1 U317 ( .B(n761), .C(n776), .A(n777), .Y(N879) );
  AO21X1 U318 ( .B(n759), .C(n781), .A(n26), .Y(N877) );
  AO21X1 U319 ( .B(n759), .C(n778), .A(n27), .Y(N876) );
  AO21X1 U320 ( .B(n759), .C(n776), .A(n777), .Y(N875) );
  AO21X1 U321 ( .B(n759), .C(n775), .A(n26), .Y(N874) );
  NAND32X1 U322 ( .B(n790), .C(n783), .A(n782), .Y(N897) );
  AO21X1 U323 ( .B(n781), .C(n780), .A(n779), .Y(n783) );
  INVX1 U324 ( .A(n787), .Y(n779) );
  INVX1 U325 ( .A(n756), .Y(n768) );
  INVX1 U326 ( .A(n304), .Y(n750) );
  OR2X1 U327 ( .A(n751), .B(n335), .Y(n747) );
  INVX1 U328 ( .A(n306), .Y(n332) );
  INVX1 U329 ( .A(n774), .Y(n780) );
  NAND21X1 U330 ( .B(n773), .A(n772), .Y(n774) );
  NAND2X1 U331 ( .A(n47), .B(n102), .Y(n111) );
  NAND2X1 U332 ( .A(n184), .B(memaddr_c[11]), .Y(n199) );
  INVX1 U333 ( .A(n674), .Y(n675) );
  NAND21X1 U334 ( .B(n768), .A(n673), .Y(n674) );
  INVX1 U335 ( .A(n621), .Y(n622) );
  NAND21X1 U336 ( .B(n768), .A(n620), .Y(n621) );
  INVX1 U337 ( .A(n581), .Y(n582) );
  NAND21X1 U338 ( .B(n768), .A(n580), .Y(n581) );
  INVX1 U339 ( .A(n542), .Y(n543) );
  NAND21X1 U340 ( .B(n768), .A(n541), .Y(n542) );
  INVX1 U341 ( .A(n503), .Y(n504) );
  NAND21X1 U342 ( .B(n768), .A(n502), .Y(n503) );
  INVX1 U343 ( .A(n465), .Y(n466) );
  NAND21X1 U344 ( .B(n768), .A(n464), .Y(n465) );
  INVX1 U345 ( .A(n426), .Y(n427) );
  NAND21X1 U346 ( .B(n768), .A(n425), .Y(n426) );
  INVX1 U347 ( .A(n357), .Y(n358) );
  NAND21X1 U348 ( .B(n768), .A(n356), .Y(n357) );
  NAND2X1 U349 ( .A(n188), .B(memaddr_c[12]), .Y(n202) );
  OAI211X1 U350 ( .C(n892), .D(n320), .A(n825), .B(n837), .Y(n741) );
  INVX1 U351 ( .A(memaddr_c[14]), .Y(n798) );
  NOR3XL U352 ( .A(n765), .B(n773), .C(n764), .Y(n48) );
  INVX1 U353 ( .A(n762), .Y(n763) );
  NAND32X1 U354 ( .B(n765), .C(n764), .A(n773), .Y(n762) );
  INVX1 U355 ( .A(n760), .Y(n761) );
  NAND32X1 U356 ( .B(n773), .C(n764), .A(n765), .Y(n760) );
  INVX1 U357 ( .A(n286), .Y(n291) );
  EORX1 U358 ( .A(n191), .B(memaddr_c[13]), .C(n1), .D(n798), .Y(n49) );
  AO21X1 U359 ( .B(sfr_psr), .C(n88), .A(n849), .Y(n327) );
  INVX1 U360 ( .A(n910), .Y(n88) );
  NAND21X1 U361 ( .B(n739), .A(n813), .Y(n841) );
  INVX1 U362 ( .A(n102), .Y(n101) );
  NAND21X1 U363 ( .B(n174), .A(memaddr_c[8]), .Y(n206) );
  NAND21X1 U364 ( .B(n60), .A(memaddr_c[7]), .Y(n209) );
  NAND43X1 U365 ( .B(n746), .C(n754), .D(n745), .A(n744), .Y(N820) );
  AO21X1 U366 ( .B(n904), .C(n847), .A(n909), .Y(n745) );
  AND4X1 U367 ( .A(n846), .B(n818), .C(n743), .D(n742), .Y(n744) );
  NAND21X1 U368 ( .B(memaddr_c[14]), .A(n1), .Y(n215) );
  NAND21X1 U369 ( .B(memaddr_c[9]), .A(n59), .Y(n179) );
  OA21X1 U370 ( .B(n778), .C(n776), .A(n336), .Y(N843) );
  INVX1 U371 ( .A(memaddr_c[7]), .Y(n170) );
  INVX1 U372 ( .A(memaddr_c[11]), .Y(n126) );
  AND2X1 U373 ( .A(n336), .B(n293), .Y(N842) );
  AND2X1 U374 ( .A(n285), .B(n336), .Y(N846) );
  XOR2X1 U375 ( .A(n767), .B(n284), .Y(n285) );
  NAND21X1 U376 ( .B(n765), .A(n283), .Y(n284) );
  INVX1 U377 ( .A(n128), .Y(n92) );
  INVX1 U378 ( .A(n87), .Y(n849) );
  NAND21X1 U379 ( .B(n59), .A(memaddr_c[9]), .Y(n201) );
  NAND2X1 U380 ( .A(n181), .B(memaddr_c[10]), .Y(n207) );
  INVX1 U381 ( .A(memaddr_c[10]), .Y(n120) );
  NAND21X1 U382 ( .B(n739), .A(n84), .Y(n795) );
  NAND21X1 U383 ( .B(n850), .A(n844), .Y(n340) );
  AND4X1 U384 ( .A(n251), .B(n250), .C(n249), .D(n248), .Y(n274) );
  OR3XL U385 ( .A(n790), .B(n789), .C(n50), .Y(N898) );
  AOI21X1 U386 ( .B(n788), .C(n906), .A(n787), .Y(n50) );
  INVX1 U387 ( .A(n799), .Y(n804) );
  MUX2BXL U388 ( .D0(n231), .D1(n229), .S(n230), .Y(n232) );
  AO21XL U389 ( .B(n672), .C(n801), .A(n81), .Y(n341) );
  NAND21X1 U390 ( .B(n908), .A(n84), .Y(n787) );
  NAND21X1 U391 ( .B(n847), .A(n893), .Y(n826) );
  INVX1 U392 ( .A(n894), .Y(n847) );
  INVX1 U393 ( .A(n666), .Y(n833) );
  AOI21XL U394 ( .B(n793), .C(n792), .A(n81), .Y(N899) );
  AO21X1 U395 ( .B(n850), .C(n791), .A(n846), .Y(n792) );
  NAND21X1 U396 ( .B(n904), .A(n847), .Y(n793) );
  NAND21X1 U397 ( .B(n299), .A(n315), .Y(n788) );
  NAND32X1 U398 ( .B(n300), .C(n299), .A(n298), .Y(n825) );
  INVX1 U399 ( .A(n892), .Y(n839) );
  OAI31XL U400 ( .A(n886), .B(n910), .C(n326), .D(n911), .Y(n806) );
  INVX1 U401 ( .A(sfr_psw), .Y(n326) );
  MUX2AXL U402 ( .D0(n857), .D1(sfr_psr), .S(n848), .Y(sfr_psrack) );
  MUX2AXL U403 ( .D0(n242), .D1(n240), .S(n141), .Y(n156) );
  AO21X1 U404 ( .B(n141), .C(n223), .A(n222), .Y(n159) );
  AO21X1 U405 ( .B(n142), .C(n221), .A(n220), .Y(n141) );
  AO21X1 U406 ( .B(n150), .C(n217), .A(n216), .Y(n145) );
  AO21X1 U407 ( .B(n219), .C(n145), .A(n218), .Y(n142) );
  INVX1 U408 ( .A(n149), .Y(n216) );
  MUX2AXL U409 ( .D0(n246), .D1(n244), .S(n142), .Y(n143) );
  INVX1 U410 ( .A(n144), .Y(n218) );
  MUX2AXL U411 ( .D0(n237), .D1(n235), .S(n150), .Y(n153) );
  NAND2X1 U412 ( .A(n219), .B(n144), .Y(n229) );
  NAND21X1 U413 ( .B(n220), .A(n221), .Y(n244) );
  NAND21X1 U414 ( .B(n222), .A(n223), .Y(n240) );
  NAND2X1 U415 ( .A(n217), .B(n149), .Y(n235) );
  OR2X1 U416 ( .A(n171), .B(n225), .Y(n176) );
  NAND21X1 U417 ( .B(n139), .A(n61), .Y(n171) );
  MUX2AXL U418 ( .D0(n231), .D1(n229), .S(n145), .Y(n152) );
  OR2X1 U419 ( .A(n176), .B(n226), .Y(n185) );
  OR2X1 U420 ( .A(n185), .B(n227), .Y(n138) );
  NAND21X1 U421 ( .B(n226), .A(n253), .Y(n265) );
  NAND21X1 U422 ( .B(n227), .A(n266), .Y(n263) );
  NAND21X1 U423 ( .B(n225), .A(n256), .Y(n252) );
  NAND21X1 U424 ( .B(n51), .A(n61), .Y(n255) );
  AO21X1 U425 ( .B(n245), .C(n221), .A(n220), .Y(n241) );
  AO21X1 U426 ( .B(n230), .C(n219), .A(n218), .Y(n245) );
  AO21X1 U427 ( .B(n236), .C(n217), .A(n216), .Y(n230) );
  OR2X1 U428 ( .A(n228), .B(n263), .Y(n264) );
  AOI21X1 U429 ( .B(n241), .C(n223), .A(n222), .Y(n51) );
  MUX2BXL U430 ( .D0(n246), .D1(n244), .S(n245), .Y(n247) );
  MUX2BXL U431 ( .D0(n242), .D1(n240), .S(n241), .Y(n243) );
  MUX2BXL U432 ( .D0(n237), .D1(n235), .S(n236), .Y(n238) );
  INVX1 U433 ( .A(n196), .Y(n224) );
  AND4X1 U434 ( .A(n775), .B(n767), .C(n773), .D(n765), .Y(n193) );
  INVX1 U435 ( .A(n278), .Y(n775) );
  AO21X1 U436 ( .B(n299), .C(n287), .A(n294), .Y(n751) );
  INVX1 U437 ( .A(n289), .Y(n321) );
  OR2X1 U438 ( .A(n300), .B(n830), .Y(n742) );
  NAND21X1 U439 ( .B(n848), .A(n301), .Y(n801) );
  INVX1 U440 ( .A(n829), .Y(n667) );
  NAND2X1 U441 ( .A(n836), .B(n788), .Y(n421) );
  NAND21X1 U442 ( .B(n839), .A(n893), .Y(n334) );
  INVX1 U443 ( .A(n906), .Y(n851) );
  INVX1 U444 ( .A(n739), .Y(n354) );
  INVX1 U445 ( .A(n908), .Y(n316) );
  NAND21X1 U446 ( .B(n773), .A(n781), .Y(n305) );
  NAND21X1 U447 ( .B(n850), .A(n354), .Y(n671) );
  GEN2XL U448 ( .D(n834), .E(n833), .C(n832), .B(n84), .A(n831), .Y(n642) );
  AND3X1 U449 ( .A(pmem_clk[1]), .B(n33), .C(n830), .Y(n831) );
  GEN2XL U450 ( .D(n834), .E(n829), .C(n832), .B(n83), .A(n828), .Y(n641) );
  OA21X1 U451 ( .B(memaddr[3]), .C(n362), .A(n377), .Y(n361) );
  NAND21X1 U452 ( .B(memaddr[0]), .A(c_adr[0]), .Y(n365) );
  OA222X1 U453 ( .A(n693), .B(n381), .C(n691), .D(n380), .E(n689), .F(n379), 
        .Y(n417) );
  INVX1 U454 ( .A(c_buf_17__7_), .Y(n381) );
  INVX1 U455 ( .A(c_buf_16__7_), .Y(n380) );
  INVX1 U456 ( .A(dbg_0f[7]), .Y(n379) );
  OA222X1 U457 ( .A(n723), .B(n410), .C(n721), .D(n409), .E(n719), .F(n408), 
        .Y(n411) );
  INVX1 U458 ( .A(rd_buf[7]), .Y(n410) );
  INVX1 U459 ( .A(dbg_02[7]), .Y(n409) );
  INVX1 U460 ( .A(dbg_01[7]), .Y(n408) );
  OAI21BBX1 U461 ( .A(memaddr[2]), .B(n360), .C(n52), .Y(n377) );
  OAI21X1 U462 ( .B(memaddr[2]), .C(n360), .A(n363), .Y(n52) );
  OAI21BX1 U463 ( .C(memaddr[1]), .B(c_adr[1]), .A(n54), .Y(n363) );
  OAI21X1 U464 ( .B(memaddr[1]), .C(n359), .A(n365), .Y(n54) );
  XOR3XL U465 ( .A(memaddr[1]), .B(c_adr[1]), .C(n365), .Y(n366) );
  OA222X1 U466 ( .A(n693), .B(n435), .C(n691), .D(n434), .E(n689), .F(n433), 
        .Y(n457) );
  INVX1 U467 ( .A(c_buf_17__6_), .Y(n435) );
  INVX1 U468 ( .A(c_buf_16__6_), .Y(n434) );
  INVX1 U469 ( .A(dbg_0f[6]), .Y(n433) );
  OA222X1 U470 ( .A(n693), .B(n551), .C(n691), .D(n550), .E(n689), .F(n549), 
        .Y(n573) );
  INVX1 U471 ( .A(c_buf_17__3_), .Y(n551) );
  INVX1 U472 ( .A(c_buf_16__3_), .Y(n550) );
  INVX1 U473 ( .A(dbg_0f[3]), .Y(n549) );
  OA222X1 U474 ( .A(n693), .B(n474), .C(n691), .D(n473), .E(n689), .F(n472), 
        .Y(n496) );
  INVX1 U475 ( .A(c_buf_17__5_), .Y(n474) );
  INVX1 U476 ( .A(c_buf_16__5_), .Y(n473) );
  INVX1 U477 ( .A(dbg_0f[5]), .Y(n472) );
  OA222X1 U478 ( .A(n693), .B(n590), .C(n691), .D(n589), .E(n689), .F(n588), 
        .Y(n612) );
  INVX1 U479 ( .A(c_buf_17__2_), .Y(n590) );
  INVX1 U480 ( .A(c_buf_16__2_), .Y(n589) );
  INVX1 U481 ( .A(dbg_0f[2]), .Y(n588) );
  OA222X1 U482 ( .A(n693), .B(n630), .C(n691), .D(n629), .E(n689), .F(n628), 
        .Y(n663) );
  INVX1 U483 ( .A(c_buf_17__1_), .Y(n630) );
  INVX1 U484 ( .A(c_buf_16__1_), .Y(n629) );
  INVX1 U485 ( .A(dbg_0f[1]), .Y(n628) );
  OA222X1 U486 ( .A(n693), .B(n512), .C(n691), .D(n511), .E(n689), .F(n510), 
        .Y(n534) );
  INVX1 U487 ( .A(c_buf_17__4_), .Y(n512) );
  INVX1 U488 ( .A(c_buf_16__4_), .Y(n511) );
  INVX1 U489 ( .A(dbg_0f[4]), .Y(n510) );
  OA222X1 U490 ( .A(n693), .B(n692), .C(n691), .D(n690), .E(n689), .F(n688), 
        .Y(n730) );
  INVX1 U491 ( .A(c_buf_17__0_), .Y(n692) );
  INVX1 U492 ( .A(c_buf_16__0_), .Y(n690) );
  INVX1 U493 ( .A(dbg_0f[0]), .Y(n688) );
  OA222X1 U494 ( .A(n723), .B(n566), .C(n721), .D(n565), .E(n719), .F(n564), 
        .Y(n567) );
  INVX1 U495 ( .A(rd_buf[3]), .Y(n566) );
  INVX1 U496 ( .A(dbg_02[3]), .Y(n565) );
  INVX1 U497 ( .A(dbg_01[3]), .Y(n564) );
  OA222X1 U498 ( .A(n723), .B(n450), .C(n721), .D(n449), .E(n719), .F(n448), 
        .Y(n451) );
  INVX1 U499 ( .A(rd_buf[6]), .Y(n450) );
  INVX1 U500 ( .A(dbg_02[6]), .Y(n449) );
  INVX1 U501 ( .A(dbg_01[6]), .Y(n448) );
  OA222X1 U502 ( .A(n723), .B(n527), .C(n721), .D(n526), .E(n719), .F(n525), 
        .Y(n528) );
  INVX1 U503 ( .A(rd_buf[4]), .Y(n527) );
  INVX1 U504 ( .A(dbg_02[4]), .Y(n526) );
  INVX1 U505 ( .A(dbg_01[4]), .Y(n525) );
  OA222X1 U506 ( .A(n723), .B(n722), .C(n721), .D(n720), .E(n719), .F(n718), 
        .Y(n724) );
  INVX1 U507 ( .A(rd_buf[0]), .Y(n722) );
  INVX1 U508 ( .A(dbg_02[0]), .Y(n720) );
  INVX1 U509 ( .A(dbg_01[0]), .Y(n718) );
  OA222X1 U510 ( .A(n723), .B(n489), .C(n721), .D(n488), .E(n719), .F(n487), 
        .Y(n490) );
  INVX1 U511 ( .A(rd_buf[5]), .Y(n489) );
  INVX1 U512 ( .A(dbg_02[5]), .Y(n488) );
  INVX1 U513 ( .A(dbg_01[5]), .Y(n487) );
  OA222X1 U514 ( .A(n723), .B(n605), .C(n721), .D(n604), .E(n719), .F(n603), 
        .Y(n606) );
  INVX1 U515 ( .A(rd_buf[2]), .Y(n605) );
  INVX1 U516 ( .A(dbg_02[2]), .Y(n604) );
  INVX1 U517 ( .A(dbg_01[2]), .Y(n603) );
  OA222X1 U518 ( .A(n723), .B(n656), .C(n721), .D(n655), .E(n719), .F(n654), 
        .Y(n657) );
  INVX1 U519 ( .A(rd_buf[1]), .Y(n656) );
  INVX1 U520 ( .A(dbg_02[1]), .Y(n655) );
  INVX1 U521 ( .A(dbg_01[1]), .Y(n654) );
  INVXL U522 ( .A(c_adr[0]), .Y(n364) );
  INVX1 U523 ( .A(c_adr[3]), .Y(n362) );
  NAND21X1 U524 ( .B(cs_ft[0]), .A(cs_ft[1]), .Y(n287) );
  INVX1 U525 ( .A(wr_buf[7]), .Y(n422) );
  INVX1 U526 ( .A(dbg_04[7]), .Y(n401) );
  INVX1 U527 ( .A(dbg_07[7]), .Y(n393) );
  INVX1 U528 ( .A(dbg_0a[7]), .Y(n387) );
  INVX1 U529 ( .A(c_buf_18__7_), .Y(n371) );
  INVX1 U530 ( .A(c_buf_21__7_), .Y(n367) );
  INVX1 U531 ( .A(dbg_0c[7]), .Y(n383) );
  INVX1 U532 ( .A(dbg_05[7]), .Y(n402) );
  INVX1 U533 ( .A(dbg_08[7]), .Y(n394) );
  INVX1 U534 ( .A(dbg_0b[7]), .Y(n388) );
  INVX1 U535 ( .A(c_buf_19__7_), .Y(n372) );
  INVX1 U536 ( .A(c_buf_22__7_), .Y(n368) );
  INVX1 U537 ( .A(dbg_0d[7]), .Y(n384) );
  INVX1 U538 ( .A(dbg_03[7]), .Y(n403) );
  INVX1 U539 ( .A(dbg_06[7]), .Y(n395) );
  INVX1 U540 ( .A(dbg_09[7]), .Y(n389) );
  INVX1 U541 ( .A(c_buf_20__7_), .Y(n373) );
  INVX1 U542 ( .A(dbg_0e[7]), .Y(n385) );
  INVX1 U543 ( .A(cs_ft[2]), .Y(n300) );
  INVX1 U544 ( .A(cs_ft[3]), .Y(n298) );
  INVX1 U545 ( .A(mcu_psw), .Y(n850) );
  INVX1 U546 ( .A(r_rdy), .Y(n845) );
  INVX1 U547 ( .A(dbg_04[3]), .Y(n561) );
  INVX1 U548 ( .A(dbg_07[3]), .Y(n558) );
  INVX1 U549 ( .A(dbg_0a[3]), .Y(n555) );
  INVX1 U550 ( .A(dbg_04[4]), .Y(n522) );
  INVX1 U551 ( .A(dbg_07[4]), .Y(n519) );
  INVX1 U552 ( .A(dbg_0a[4]), .Y(n516) );
  INVX1 U553 ( .A(dbg_04[0]), .Y(n712) );
  INVX1 U554 ( .A(dbg_07[0]), .Y(n706) );
  INVX1 U555 ( .A(dbg_0a[0]), .Y(n700) );
  INVX1 U556 ( .A(dbg_0c[3]), .Y(n552) );
  INVX1 U557 ( .A(dbg_04[6]), .Y(n445) );
  INVX1 U558 ( .A(dbg_07[6]), .Y(n442) );
  INVX1 U559 ( .A(dbg_0a[6]), .Y(n439) );
  INVX1 U560 ( .A(dbg_04[5]), .Y(n484) );
  INVX1 U561 ( .A(dbg_07[5]), .Y(n481) );
  INVX1 U562 ( .A(dbg_0a[5]), .Y(n478) );
  INVX1 U563 ( .A(dbg_0c[6]), .Y(n436) );
  INVX1 U564 ( .A(dbg_05[3]), .Y(n562) );
  INVX1 U565 ( .A(dbg_08[3]), .Y(n559) );
  INVX1 U566 ( .A(dbg_0b[3]), .Y(n556) );
  INVX1 U567 ( .A(dbg_05[4]), .Y(n523) );
  INVX1 U568 ( .A(dbg_08[4]), .Y(n520) );
  INVX1 U569 ( .A(dbg_0b[4]), .Y(n517) );
  INVX1 U570 ( .A(dbg_05[0]), .Y(n714) );
  INVX1 U571 ( .A(dbg_08[0]), .Y(n708) );
  INVX1 U572 ( .A(dbg_0b[0]), .Y(n702) );
  INVX1 U573 ( .A(dbg_0d[3]), .Y(n553) );
  INVX1 U574 ( .A(dbg_05[6]), .Y(n446) );
  INVX1 U575 ( .A(dbg_08[6]), .Y(n443) );
  INVX1 U576 ( .A(dbg_0b[6]), .Y(n440) );
  INVX1 U577 ( .A(dbg_05[5]), .Y(n485) );
  INVX1 U578 ( .A(dbg_08[5]), .Y(n482) );
  INVX1 U579 ( .A(dbg_0b[5]), .Y(n479) );
  INVX1 U580 ( .A(dbg_0d[6]), .Y(n437) );
  INVX1 U581 ( .A(dbg_03[3]), .Y(n563) );
  INVX1 U582 ( .A(dbg_06[3]), .Y(n560) );
  INVX1 U583 ( .A(dbg_09[3]), .Y(n557) );
  INVX1 U584 ( .A(dbg_03[4]), .Y(n524) );
  INVX1 U585 ( .A(dbg_03[0]), .Y(n716) );
  INVX1 U586 ( .A(dbg_03[6]), .Y(n447) );
  INVX1 U587 ( .A(dbg_06[6]), .Y(n444) );
  INVX1 U588 ( .A(dbg_09[6]), .Y(n441) );
  INVX1 U589 ( .A(dbg_03[5]), .Y(n486) );
  INVX1 U590 ( .A(dbg_06[5]), .Y(n483) );
  INVX1 U591 ( .A(dbg_09[5]), .Y(n480) );
  INVX1 U592 ( .A(wr_buf[0]), .Y(n791) );
  INVX1 U593 ( .A(wr_buf[1]), .Y(n668) );
  INVX1 U594 ( .A(wr_buf[5]), .Y(n499) );
  INVX1 U595 ( .A(wr_buf[3]), .Y(n577) );
  INVX1 U596 ( .A(wr_buf[6]), .Y(n461) );
  INVX1 U597 ( .A(wr_buf[4]), .Y(n538) );
  INVX1 U598 ( .A(dbg_04[2]), .Y(n600) );
  INVX1 U599 ( .A(dbg_07[2]), .Y(n597) );
  INVX1 U600 ( .A(dbg_0a[2]), .Y(n594) );
  INVX1 U601 ( .A(c_buf_21__2_), .Y(n583) );
  INVX1 U602 ( .A(c_buf_18__2_), .Y(n585) );
  INVX1 U603 ( .A(dbg_0c[2]), .Y(n591) );
  INVX1 U604 ( .A(dbg_04[1]), .Y(n640) );
  INVX1 U605 ( .A(dbg_07[1]), .Y(n637) );
  INVX1 U606 ( .A(dbg_0a[1]), .Y(n634) );
  INVX1 U607 ( .A(c_buf_21__1_), .Y(n623) );
  INVX1 U608 ( .A(c_buf_18__1_), .Y(n625) );
  INVX1 U609 ( .A(dbg_0c[1]), .Y(n631) );
  INVX1 U610 ( .A(c_buf_21__3_), .Y(n544) );
  INVX1 U611 ( .A(c_buf_18__3_), .Y(n546) );
  INVX1 U612 ( .A(c_buf_21__4_), .Y(n505) );
  INVX1 U613 ( .A(c_buf_18__4_), .Y(n507) );
  INVX1 U614 ( .A(dbg_0c[4]), .Y(n513) );
  INVX1 U615 ( .A(c_buf_21__0_), .Y(n677) );
  INVX1 U616 ( .A(c_buf_18__0_), .Y(n682) );
  INVX1 U617 ( .A(dbg_0c[0]), .Y(n694) );
  INVX1 U618 ( .A(c_buf_21__6_), .Y(n428) );
  INVX1 U619 ( .A(c_buf_18__6_), .Y(n430) );
  INVX1 U620 ( .A(c_buf_21__5_), .Y(n467) );
  INVX1 U621 ( .A(c_buf_18__5_), .Y(n469) );
  INVX1 U622 ( .A(dbg_0c[5]), .Y(n475) );
  INVX1 U623 ( .A(dbg_05[2]), .Y(n601) );
  INVX1 U624 ( .A(dbg_08[2]), .Y(n598) );
  INVX1 U625 ( .A(dbg_0b[2]), .Y(n595) );
  INVX1 U626 ( .A(c_buf_22__2_), .Y(n584) );
  INVX1 U627 ( .A(c_buf_19__2_), .Y(n586) );
  INVX1 U628 ( .A(dbg_0d[2]), .Y(n592) );
  INVX1 U629 ( .A(dbg_05[1]), .Y(n652) );
  INVX1 U630 ( .A(dbg_08[1]), .Y(n638) );
  INVX1 U631 ( .A(dbg_0b[1]), .Y(n635) );
  INVX1 U632 ( .A(c_buf_22__1_), .Y(n624) );
  INVX1 U633 ( .A(c_buf_19__1_), .Y(n626) );
  INVX1 U634 ( .A(dbg_0d[1]), .Y(n632) );
  INVX1 U635 ( .A(c_buf_22__3_), .Y(n545) );
  INVX1 U636 ( .A(c_buf_19__3_), .Y(n547) );
  INVX1 U637 ( .A(c_buf_22__4_), .Y(n506) );
  INVX1 U638 ( .A(c_buf_19__4_), .Y(n508) );
  INVX1 U639 ( .A(dbg_0d[4]), .Y(n514) );
  INVX1 U640 ( .A(c_buf_22__0_), .Y(n679) );
  INVX1 U641 ( .A(c_buf_19__0_), .Y(n684) );
  INVX1 U642 ( .A(dbg_0d[0]), .Y(n696) );
  INVX1 U643 ( .A(c_buf_22__6_), .Y(n429) );
  INVX1 U644 ( .A(c_buf_19__6_), .Y(n431) );
  INVX1 U645 ( .A(c_buf_22__5_), .Y(n468) );
  INVX1 U646 ( .A(c_buf_19__5_), .Y(n470) );
  INVX1 U647 ( .A(dbg_0d[5]), .Y(n476) );
  INVX1 U648 ( .A(dbg_03[2]), .Y(n602) );
  INVX1 U649 ( .A(dbg_06[2]), .Y(n599) );
  INVX1 U650 ( .A(dbg_09[2]), .Y(n596) );
  INVX1 U651 ( .A(dbg_0e[2]), .Y(n593) );
  INVX1 U652 ( .A(dbg_03[1]), .Y(n653) );
  INVX1 U653 ( .A(dbg_06[1]), .Y(n639) );
  INVX1 U654 ( .A(dbg_09[1]), .Y(n636) );
  INVX1 U655 ( .A(c_buf_20__1_), .Y(n627) );
  INVX1 U656 ( .A(dbg_0e[1]), .Y(n633) );
  INVX1 U657 ( .A(dbg_06[4]), .Y(n521) );
  INVX1 U658 ( .A(dbg_09[4]), .Y(n518) );
  INVX1 U659 ( .A(dbg_06[0]), .Y(n710) );
  INVX1 U660 ( .A(dbg_09[0]), .Y(n704) );
  INVX1 U661 ( .A(c_buf_20__3_), .Y(n548) );
  INVX1 U662 ( .A(dbg_0e[3]), .Y(n554) );
  INVX1 U663 ( .A(c_buf_20__4_), .Y(n509) );
  INVX1 U664 ( .A(dbg_0e[4]), .Y(n515) );
  INVX1 U665 ( .A(c_buf_20__0_), .Y(n686) );
  INVX1 U666 ( .A(dbg_0e[0]), .Y(n698) );
  INVX1 U667 ( .A(c_buf_20__6_), .Y(n432) );
  INVX1 U668 ( .A(dbg_0e[6]), .Y(n438) );
  INVX1 U669 ( .A(c_buf_20__5_), .Y(n471) );
  INVX1 U670 ( .A(dbg_0e[5]), .Y(n477) );
  OR2X1 U671 ( .A(d_psrd), .B(n322), .Y(n308) );
  NAND2X1 U672 ( .A(n3), .B(pre_1_adr[14]), .Y(n809) );
  AO21X1 U673 ( .B(n812), .C(n816), .A(n811), .Y(n646) );
  AND3X1 U674 ( .A(wd_twlb[0]), .B(we_twlb), .C(n813), .Y(n812) );
  MUX2X1 U675 ( .D0(n814), .D1(pmem_twlb[0]), .S(n32), .Y(n811) );
  AO21X1 U676 ( .B(n817), .C(n816), .A(n815), .Y(n645) );
  AND3X1 U677 ( .A(wd_twlb[1]), .B(we_twlb), .C(n813), .Y(n817) );
  MUX2X1 U678 ( .D0(n814), .D1(pmem_twlb[1]), .S(n32), .Y(n815) );
  OAI211X1 U679 ( .C(pre_1_adr[13]), .D(n809), .A(n808), .B(n807), .Y(n814) );
  AOI33X1 U680 ( .A(n806), .B(n805), .C(n804), .D(sfr_psofs[14]), .E(n803), 
        .F(n802), .Y(n807) );
  NAND32X1 U681 ( .B(memaddr_c[13]), .C(n798), .A(n797), .Y(n808) );
  INVX1 U682 ( .A(sfr_psofs[13]), .Y(n802) );
  INVX1 U683 ( .A(wr_buf[2]), .Y(n617) );
  INVX1 U684 ( .A(c_buf_20__2_), .Y(n587) );
  OAI32X1 U685 ( .A(n742), .B(d_psrd), .C(n81), .D(n757), .E(n335), .Y(n797)
         );
  NAND21X1 U686 ( .B(d_psrd), .A(n304), .Y(n756) );
  NAND31X1 U687 ( .C(d_psrd), .A(n55), .B(n289), .Y(n304) );
  NAND3X1 U688 ( .A(n819), .B(n755), .C(n286), .Y(n55) );
  NAND43X1 U689 ( .B(n291), .C(n290), .D(d_psrd), .A(n819), .Y(n335) );
  INVX1 U690 ( .A(n755), .Y(n290) );
  NAND21X1 U691 ( .B(n195), .A(n194), .Y(n306) );
  GEN2XL U692 ( .D(c_adr[14]), .E(n798), .C(n131), .B(n130), .A(n129), .Y(n195) );
  AOI21X1 U693 ( .B(n215), .C(n200), .A(n193), .Y(n194) );
  OAI32X1 U694 ( .A(n92), .B(memaddr_c[12]), .C(n136), .D(memaddr_c[13]), .E(
        n228), .Y(n131) );
  INVX1 U695 ( .A(n770), .Y(n771) );
  NAND21X1 U696 ( .B(c_ptr[2]), .A(n772), .Y(n770) );
  AO2222XL U697 ( .A(memaddr_c[10]), .B(n797), .C(pre_1_adr[10]), .D(n3), .E(
        memaddr[10]), .F(n343), .G(sfr_psofs[10]), .H(n342), .Y(N864) );
  AO2222XL U698 ( .A(memaddr_c[13]), .B(n797), .C(pre_1_adr[13]), .D(n344), 
        .E(memaddr[13]), .F(n343), .G(sfr_psofs[13]), .H(n342), .Y(N867) );
  AO2222XL U699 ( .A(memaddr_c[12]), .B(n797), .C(pre_1_adr[12]), .D(n344), 
        .E(memaddr[12]), .F(n343), .G(sfr_psofs[12]), .H(n342), .Y(N866) );
  AO2222XL U700 ( .A(memaddr_c[11]), .B(n797), .C(pre_1_adr[11]), .D(n3), .E(
        memaddr[11]), .F(n343), .G(sfr_psofs[11]), .H(n342), .Y(N865) );
  AO2222XL U701 ( .A(memaddr_c[9]), .B(n797), .C(pre_1_adr[9]), .D(n3), .E(
        memaddr[9]), .F(n343), .G(sfr_psofs[9]), .H(n342), .Y(N863) );
  AO2222XL U702 ( .A(memaddr_c[8]), .B(n797), .C(pre_1_adr[8]), .D(n344), .E(
        memaddr[8]), .F(n343), .G(sfr_psofs[8]), .H(n342), .Y(N862) );
  AO2222XL U703 ( .A(memaddr_c[7]), .B(n797), .C(pre_1_adr[7]), .D(n344), .E(
        memaddr[7]), .F(n343), .G(sfr_psofs[7]), .H(n342), .Y(N861) );
  AO2222XL U704 ( .A(memaddr_c[5]), .B(n797), .C(pre_1_adr[5]), .D(n3), .E(
        memaddr[5]), .F(n343), .G(sfr_psofs[5]), .H(n342), .Y(N859) );
  AO2222XL U705 ( .A(memaddr_c[2]), .B(n14), .C(pre_1_adr[2]), .D(n344), .E(
        memaddr[2]), .F(n343), .G(sfr_psofs[2]), .H(n342), .Y(N856) );
  AO2222XL U706 ( .A(memaddr_c[1]), .B(n14), .C(pre_1_adr[1]), .D(n3), .E(
        memaddr[1]), .F(n343), .G(sfr_psofs[1]), .H(n342), .Y(N855) );
  OAI21BBX1 U707 ( .A(N445), .B(n749), .C(n56), .Y(N840) );
  AOI21XL U708 ( .B(memaddr_c[14]), .C(n24), .A(n81), .Y(n56) );
  OAI21BBX1 U709 ( .A(N431), .B(n21), .C(n57), .Y(N826) );
  AOI21XL U710 ( .B(memaddr_c[0]), .C(n24), .A(n82), .Y(n57) );
  NAND32X1 U711 ( .B(n753), .C(n749), .A(n748), .Y(N825) );
  NAND31X1 U712 ( .C(n25), .A(n755), .B(n786), .Y(n748) );
  INVX1 U713 ( .A(n769), .Y(n772) );
  NAND43X1 U714 ( .B(c_ptr[3]), .C(n768), .D(n767), .A(n766), .Y(n769) );
  OAI211X1 U715 ( .C(n339), .D(n798), .A(n809), .B(n338), .Y(N868) );
  OA21X1 U716 ( .B(n337), .C(n341), .A(n799), .Y(n338) );
  INVX1 U717 ( .A(n797), .Y(n339) );
  INVX1 U718 ( .A(sfr_psofs[14]), .Y(n337) );
  INVX1 U719 ( .A(c_adr[4]), .Y(n113) );
  AO21XL U720 ( .B(memaddr_c[2]), .C(n360), .A(n101), .Y(n112) );
  OAI211X1 U721 ( .C(n109), .D(n108), .A(n107), .B(n106), .Y(n110) );
  NAND32X1 U722 ( .B(c_ptr[4]), .C(n757), .A(n756), .Y(n764) );
  XOR3X1 U723 ( .A(c_adr[11]), .B(memaddr_c[11]), .C(n265), .Y(n269) );
  NAND21X1 U724 ( .B(n328), .A(n800), .Y(N824) );
  GEN2XL U725 ( .D(n325), .E(n324), .C(n25), .B(n766), .A(n323), .Y(n328) );
  OA21X1 U726 ( .B(n847), .C(n421), .A(n84), .Y(n323) );
  AND3X1 U727 ( .A(n321), .B(cs_ft[0]), .C(n320), .Y(n325) );
  OAI21X1 U728 ( .B(n310), .C(n81), .A(n309), .Y(N822) );
  AND4X1 U729 ( .A(n801), .B(n825), .C(n893), .D(n303), .Y(n310) );
  GEN2XL U730 ( .D(n768), .E(n308), .C(n307), .B(n320), .A(n757), .Y(n309) );
  AOI221XL U731 ( .A(n316), .B(n851), .C(n827), .D(mcu_psw), .E(n786), .Y(n303) );
  NAND6XL U732 ( .A(n277), .B(n276), .C(n275), .D(n274), .E(n273), .F(n272), 
        .Y(n286) );
  OA21X1 U733 ( .B(n234), .C(n264), .A(n233), .Y(n275) );
  XOR3XL U734 ( .A(c_adr[5]), .B(memaddr_c[5]), .C(n51), .Y(n277) );
  GEN2XL U735 ( .D(c_adr[9]), .E(n124), .C(n123), .B(n122), .A(n121), .Y(n125)
         );
  INVX1 U736 ( .A(memaddr_c[9]), .Y(n124) );
  AND3X1 U737 ( .A(c_adr[10]), .B(n120), .C(n119), .Y(n121) );
  OA21X1 U738 ( .B(c_adr[10]), .C(n120), .A(n119), .Y(n122) );
  NAND21X1 U739 ( .B(c_adr[11]), .A(memaddr_c[11]), .Y(n119) );
  AO21X1 U740 ( .B(dbg_01[0]), .C(n79), .A(n675), .Y(N479) );
  AO21X1 U741 ( .B(dbg_02[0]), .C(n79), .A(n28), .Y(N487) );
  AO21X1 U742 ( .B(dbg_03[0]), .C(n79), .A(n29), .Y(N495) );
  AO21X1 U743 ( .B(dbg_04[0]), .C(n79), .A(n675), .Y(N503) );
  AO21X1 U744 ( .B(dbg_05[0]), .C(n79), .A(n28), .Y(N511) );
  AO21X1 U745 ( .B(dbg_06[0]), .C(n79), .A(n29), .Y(N519) );
  AO21X1 U746 ( .B(dbg_07[0]), .C(n78), .A(n675), .Y(N527) );
  AO21X1 U747 ( .B(dbg_01[1]), .C(n77), .A(n622), .Y(N480) );
  AO21X1 U748 ( .B(dbg_02[1]), .C(n77), .A(n22), .Y(N488) );
  AO21X1 U749 ( .B(dbg_03[1]), .C(n77), .A(n23), .Y(N496) );
  AO21X1 U750 ( .B(dbg_04[1]), .C(n76), .A(n622), .Y(N504) );
  AO21X1 U751 ( .B(dbg_05[1]), .C(n76), .A(n22), .Y(N512) );
  AO21X1 U752 ( .B(dbg_06[1]), .C(n76), .A(n23), .Y(N520) );
  AO21X1 U753 ( .B(dbg_07[1]), .C(n76), .A(n622), .Y(N528) );
  AO21X1 U754 ( .B(dbg_01[2]), .C(n74), .A(n582), .Y(N481) );
  AO21X1 U755 ( .B(dbg_02[2]), .C(n74), .A(n18), .Y(N489) );
  AO21X1 U756 ( .B(dbg_03[2]), .C(n74), .A(n19), .Y(N497) );
  AO21X1 U757 ( .B(dbg_04[2]), .C(n74), .A(n582), .Y(N505) );
  AO21X1 U758 ( .B(dbg_05[2]), .C(n74), .A(n18), .Y(N513) );
  AO21X1 U759 ( .B(dbg_06[2]), .C(n74), .A(n19), .Y(N521) );
  AO21X1 U760 ( .B(dbg_07[2]), .C(n74), .A(n582), .Y(N529) );
  AO21X1 U761 ( .B(dbg_01[3]), .C(n72), .A(n543), .Y(N482) );
  AO21X1 U762 ( .B(dbg_02[3]), .C(n72), .A(n15), .Y(N490) );
  AO21X1 U763 ( .B(dbg_03[3]), .C(n72), .A(n16), .Y(N498) );
  AO21X1 U764 ( .B(dbg_04[3]), .C(n72), .A(n543), .Y(N506) );
  AO21X1 U765 ( .B(dbg_05[3]), .C(n72), .A(n15), .Y(N514) );
  AO21X1 U766 ( .B(dbg_06[3]), .C(n72), .A(n16), .Y(N522) );
  AO21X1 U767 ( .B(dbg_07[3]), .C(n72), .A(n543), .Y(N530) );
  AO21X1 U768 ( .B(dbg_01[4]), .C(n70), .A(n504), .Y(N483) );
  AO21X1 U769 ( .B(dbg_02[4]), .C(n70), .A(n12), .Y(N491) );
  AO21X1 U770 ( .B(dbg_03[4]), .C(n70), .A(n13), .Y(N499) );
  AO21X1 U771 ( .B(dbg_04[4]), .C(n70), .A(n504), .Y(N507) );
  AO21X1 U772 ( .B(dbg_05[4]), .C(n69), .A(n12), .Y(N515) );
  AO21X1 U773 ( .B(dbg_06[4]), .C(n69), .A(n13), .Y(N523) );
  AO21X1 U774 ( .B(dbg_07[4]), .C(n69), .A(n504), .Y(N531) );
  AO21X1 U775 ( .B(dbg_01[5]), .C(n68), .A(n466), .Y(N484) );
  AO21X1 U776 ( .B(dbg_02[5]), .C(n67), .A(n10), .Y(N492) );
  AO21X1 U777 ( .B(dbg_03[5]), .C(n67), .A(n11), .Y(N500) );
  AO21X1 U778 ( .B(dbg_04[5]), .C(n67), .A(n466), .Y(N508) );
  AO21X1 U779 ( .B(dbg_05[5]), .C(n67), .A(n10), .Y(N516) );
  AO21X1 U780 ( .B(dbg_06[5]), .C(n67), .A(n11), .Y(N524) );
  AO21X1 U781 ( .B(dbg_07[5]), .C(n67), .A(n466), .Y(N532) );
  AO21X1 U782 ( .B(dbg_01[6]), .C(n65), .A(n427), .Y(N485) );
  AO21X1 U783 ( .B(dbg_02[6]), .C(n65), .A(n7), .Y(N493) );
  AO21X1 U784 ( .B(dbg_03[6]), .C(n65), .A(n8), .Y(N501) );
  AO21X1 U785 ( .B(dbg_04[6]), .C(n65), .A(n427), .Y(N509) );
  AO21X1 U786 ( .B(dbg_05[6]), .C(n65), .A(n7), .Y(N517) );
  AO21X1 U787 ( .B(dbg_06[6]), .C(n65), .A(n8), .Y(N525) );
  AO21X1 U788 ( .B(dbg_07[6]), .C(n65), .A(n427), .Y(N533) );
  AO21X1 U789 ( .B(dbg_01[7]), .C(n79), .A(n358), .Y(N486) );
  AO21X1 U790 ( .B(dbg_02[7]), .C(n79), .A(n4), .Y(N494) );
  AO21X1 U791 ( .B(dbg_03[7]), .C(n79), .A(n5), .Y(N502) );
  AO21X1 U792 ( .B(dbg_04[7]), .C(n79), .A(n358), .Y(N510) );
  AO21X1 U793 ( .B(dbg_05[7]), .C(n676), .A(n4), .Y(N518) );
  AO21X1 U794 ( .B(dbg_06[7]), .C(n63), .A(n5), .Y(N526) );
  AO21X1 U795 ( .B(dbg_07[7]), .C(n63), .A(n358), .Y(N534) );
  AO21X1 U796 ( .B(dbg_08[0]), .C(n78), .A(n28), .Y(N535) );
  AO21X1 U797 ( .B(dbg_08[1]), .C(n76), .A(n22), .Y(N536) );
  AO21X1 U798 ( .B(dbg_08[2]), .C(n74), .A(n18), .Y(N537) );
  AO21X1 U799 ( .B(dbg_08[3]), .C(n71), .A(n15), .Y(N538) );
  AO21X1 U800 ( .B(dbg_08[4]), .C(n69), .A(n12), .Y(N539) );
  AO21X1 U801 ( .B(dbg_08[5]), .C(n67), .A(n10), .Y(N540) );
  AO21X1 U802 ( .B(dbg_08[6]), .C(n65), .A(n7), .Y(N541) );
  AO21X1 U803 ( .B(dbg_08[7]), .C(n63), .A(n4), .Y(N542) );
  AO21X1 U804 ( .B(dbg_09[0]), .C(n78), .A(n29), .Y(N543) );
  AO21X1 U805 ( .B(dbg_09[1]), .C(n76), .A(n23), .Y(N544) );
  AO21X1 U806 ( .B(dbg_09[2]), .C(n74), .A(n19), .Y(N545) );
  AO21X1 U807 ( .B(dbg_09[3]), .C(n71), .A(n16), .Y(N546) );
  AO21X1 U808 ( .B(dbg_09[4]), .C(n69), .A(n13), .Y(N547) );
  AO21X1 U809 ( .B(dbg_09[5]), .C(n67), .A(n11), .Y(N548) );
  AO21X1 U810 ( .B(dbg_09[6]), .C(n64), .A(n8), .Y(N549) );
  AO21X1 U811 ( .B(dbg_09[7]), .C(n63), .A(n5), .Y(N550) );
  AO21X1 U812 ( .B(dbg_0a[0]), .C(n78), .A(n675), .Y(N551) );
  AO21X1 U813 ( .B(dbg_0a[1]), .C(n76), .A(n622), .Y(N552) );
  AO21X1 U814 ( .B(dbg_0a[2]), .C(n74), .A(n582), .Y(N553) );
  AO21X1 U815 ( .B(dbg_0a[3]), .C(n71), .A(n543), .Y(N554) );
  AO21X1 U816 ( .B(dbg_0a[4]), .C(n69), .A(n504), .Y(N555) );
  AO21X1 U817 ( .B(dbg_0a[5]), .C(n67), .A(n466), .Y(N556) );
  AO21X1 U818 ( .B(dbg_0a[6]), .C(n64), .A(n427), .Y(N557) );
  AO21X1 U819 ( .B(dbg_0a[7]), .C(n63), .A(n358), .Y(N558) );
  AO21X1 U820 ( .B(dbg_0b[0]), .C(n78), .A(n28), .Y(N559) );
  AO21X1 U821 ( .B(dbg_0b[1]), .C(n76), .A(n22), .Y(N560) );
  AO21X1 U822 ( .B(dbg_0b[2]), .C(n73), .A(n18), .Y(N561) );
  AO21X1 U823 ( .B(dbg_0b[3]), .C(n71), .A(n15), .Y(N562) );
  AO21X1 U824 ( .B(dbg_0b[4]), .C(n69), .A(n12), .Y(N563) );
  AO21X1 U825 ( .B(dbg_0b[5]), .C(n67), .A(n10), .Y(N564) );
  AO21X1 U826 ( .B(dbg_0b[6]), .C(n64), .A(n7), .Y(N565) );
  AO21X1 U827 ( .B(dbg_0b[7]), .C(n63), .A(n4), .Y(N566) );
  AO21X1 U828 ( .B(dbg_0c[0]), .C(n78), .A(n29), .Y(N567) );
  AO21X1 U829 ( .B(dbg_0c[1]), .C(n76), .A(n23), .Y(N568) );
  AO21X1 U830 ( .B(dbg_0c[2]), .C(n73), .A(n19), .Y(N569) );
  AO21X1 U831 ( .B(dbg_0c[3]), .C(n71), .A(n16), .Y(N570) );
  AO21X1 U832 ( .B(dbg_0c[4]), .C(n69), .A(n13), .Y(N571) );
  AO21X1 U833 ( .B(dbg_0c[5]), .C(n66), .A(n11), .Y(N572) );
  AO21X1 U834 ( .B(dbg_0c[6]), .C(n64), .A(n8), .Y(N573) );
  AO21X1 U835 ( .B(dbg_0c[7]), .C(n63), .A(n5), .Y(N574) );
  AO21X1 U836 ( .B(dbg_0d[0]), .C(n78), .A(n675), .Y(N575) );
  AO21X1 U837 ( .B(dbg_0d[1]), .C(n76), .A(n622), .Y(N576) );
  AO21X1 U838 ( .B(dbg_0d[2]), .C(n73), .A(n582), .Y(N577) );
  AO21X1 U839 ( .B(dbg_0d[3]), .C(n71), .A(n543), .Y(N578) );
  AO21X1 U840 ( .B(dbg_0d[4]), .C(n69), .A(n504), .Y(N579) );
  AO21X1 U841 ( .B(dbg_0d[5]), .C(n66), .A(n466), .Y(N580) );
  AO21X1 U842 ( .B(dbg_0d[6]), .C(n64), .A(n427), .Y(N581) );
  AO21X1 U843 ( .B(dbg_0d[7]), .C(n63), .A(n358), .Y(N582) );
  AO21X1 U844 ( .B(dbg_0e[0]), .C(n78), .A(n28), .Y(N583) );
  AO21X1 U845 ( .B(dbg_0e[1]), .C(n75), .A(n22), .Y(N584) );
  AO21X1 U846 ( .B(dbg_0e[2]), .C(n73), .A(n18), .Y(N585) );
  AO21X1 U847 ( .B(dbg_0e[3]), .C(n71), .A(n15), .Y(N586) );
  AO21X1 U848 ( .B(dbg_0e[4]), .C(n69), .A(n12), .Y(N587) );
  AO21X1 U849 ( .B(dbg_0e[5]), .C(n66), .A(n10), .Y(N588) );
  AO21X1 U850 ( .B(dbg_0e[6]), .C(n64), .A(n7), .Y(N589) );
  AO21X1 U851 ( .B(dbg_0e[7]), .C(n63), .A(n4), .Y(N590) );
  AO21X1 U852 ( .B(dbg_0f[0]), .C(n78), .A(n29), .Y(N591) );
  AO21X1 U853 ( .B(dbg_0f[1]), .C(n75), .A(n23), .Y(N592) );
  AO21X1 U854 ( .B(dbg_0f[2]), .C(n73), .A(n19), .Y(N593) );
  AO21X1 U855 ( .B(dbg_0f[3]), .C(n71), .A(n16), .Y(N594) );
  AO21X1 U856 ( .B(dbg_0f[4]), .C(n68), .A(n13), .Y(N595) );
  AO21X1 U857 ( .B(dbg_0f[5]), .C(n66), .A(n11), .Y(N596) );
  AO21X1 U858 ( .B(dbg_0f[6]), .C(n64), .A(n8), .Y(N597) );
  AO21X1 U859 ( .B(dbg_0f[7]), .C(n63), .A(n5), .Y(N598) );
  AO21X1 U860 ( .B(c_buf_16__0_), .C(n78), .A(n675), .Y(N599) );
  AO21X1 U861 ( .B(c_buf_16__1_), .C(n75), .A(n622), .Y(N600) );
  AO21X1 U862 ( .B(c_buf_16__2_), .C(n73), .A(n582), .Y(N601) );
  AO21X1 U863 ( .B(c_buf_16__3_), .C(n71), .A(n543), .Y(N602) );
  AO21X1 U864 ( .B(c_buf_16__4_), .C(n68), .A(n504), .Y(N603) );
  AO21X1 U865 ( .B(c_buf_16__5_), .C(n66), .A(n466), .Y(N604) );
  AO21X1 U866 ( .B(c_buf_16__6_), .C(n64), .A(n427), .Y(N605) );
  AO21X1 U867 ( .B(c_buf_16__7_), .C(n62), .A(n358), .Y(N606) );
  AO21X1 U868 ( .B(c_buf_17__0_), .C(n77), .A(n28), .Y(N607) );
  AO21X1 U869 ( .B(c_buf_17__1_), .C(n75), .A(n22), .Y(N608) );
  AO21X1 U870 ( .B(c_buf_17__2_), .C(n73), .A(n18), .Y(N609) );
  AO21X1 U871 ( .B(c_buf_17__3_), .C(n71), .A(n15), .Y(N610) );
  AO21X1 U872 ( .B(c_buf_17__4_), .C(n68), .A(n12), .Y(N611) );
  AO21X1 U873 ( .B(c_buf_17__5_), .C(n66), .A(n10), .Y(N612) );
  AO21X1 U874 ( .B(c_buf_17__6_), .C(n64), .A(n7), .Y(N613) );
  AO21X1 U875 ( .B(c_buf_17__7_), .C(n62), .A(n4), .Y(N614) );
  AO21X1 U876 ( .B(c_buf_18__0_), .C(n77), .A(n29), .Y(N615) );
  AO21X1 U877 ( .B(c_buf_18__1_), .C(n75), .A(n23), .Y(N616) );
  AO21X1 U878 ( .B(c_buf_18__2_), .C(n73), .A(n19), .Y(N617) );
  AO21X1 U879 ( .B(c_buf_18__3_), .C(n70), .A(n16), .Y(N618) );
  AO21X1 U880 ( .B(c_buf_18__4_), .C(n68), .A(n13), .Y(N619) );
  AO21X1 U881 ( .B(c_buf_18__5_), .C(n66), .A(n11), .Y(N620) );
  AO21X1 U882 ( .B(c_buf_18__6_), .C(n64), .A(n8), .Y(N621) );
  AO21X1 U883 ( .B(c_buf_18__7_), .C(n62), .A(n5), .Y(N622) );
  AO21X1 U884 ( .B(c_buf_19__0_), .C(n77), .A(n675), .Y(N623) );
  AO21X1 U885 ( .B(c_buf_19__1_), .C(n75), .A(n622), .Y(N624) );
  AO21X1 U886 ( .B(c_buf_19__2_), .C(n73), .A(n582), .Y(N625) );
  AO21X1 U887 ( .B(c_buf_19__3_), .C(n70), .A(n543), .Y(N626) );
  AO21X1 U888 ( .B(c_buf_19__4_), .C(n68), .A(n504), .Y(N627) );
  AO21X1 U889 ( .B(c_buf_19__5_), .C(n66), .A(n466), .Y(N628) );
  AO21X1 U890 ( .B(c_buf_19__6_), .C(n676), .A(n427), .Y(N629) );
  AO21X1 U891 ( .B(c_buf_19__7_), .C(n62), .A(n358), .Y(N630) );
  AO21X1 U892 ( .B(c_buf_20__0_), .C(n77), .A(n28), .Y(N631) );
  AO21X1 U893 ( .B(c_buf_20__1_), .C(n75), .A(n22), .Y(N632) );
  AO21X1 U894 ( .B(c_buf_20__2_), .C(n73), .A(n18), .Y(N633) );
  AO21X1 U895 ( .B(c_buf_20__3_), .C(n70), .A(n15), .Y(N634) );
  AO21X1 U896 ( .B(c_buf_20__4_), .C(n68), .A(n12), .Y(N635) );
  AO21X1 U897 ( .B(c_buf_20__5_), .C(n66), .A(n10), .Y(N636) );
  AO21X1 U898 ( .B(c_buf_20__6_), .C(n676), .A(n7), .Y(N637) );
  AO21X1 U899 ( .B(c_buf_20__7_), .C(n62), .A(n4), .Y(N638) );
  AO21X1 U900 ( .B(c_buf_21__0_), .C(n77), .A(n29), .Y(N639) );
  AO21X1 U901 ( .B(c_buf_21__1_), .C(n75), .A(n23), .Y(N640) );
  AO21X1 U902 ( .B(c_buf_21__2_), .C(n72), .A(n19), .Y(N641) );
  AO21X1 U903 ( .B(c_buf_21__3_), .C(n70), .A(n16), .Y(N642) );
  AO21X1 U904 ( .B(c_buf_21__4_), .C(n68), .A(n13), .Y(N643) );
  AO21X1 U905 ( .B(c_buf_21__5_), .C(n66), .A(n11), .Y(N644) );
  AO21X1 U906 ( .B(c_buf_21__6_), .C(n676), .A(n8), .Y(N645) );
  AO21X1 U907 ( .B(c_buf_21__7_), .C(n62), .A(n5), .Y(N646) );
  AO21X1 U908 ( .B(c_buf_22__0_), .C(n77), .A(n675), .Y(N647) );
  AO21X1 U909 ( .B(c_buf_22__1_), .C(n75), .A(n622), .Y(N648) );
  AO21X1 U910 ( .B(c_buf_22__2_), .C(n72), .A(n582), .Y(N649) );
  AO21X1 U911 ( .B(c_buf_22__3_), .C(n70), .A(n543), .Y(N650) );
  AO21X1 U912 ( .B(c_buf_22__4_), .C(n68), .A(n504), .Y(N651) );
  AO21X1 U913 ( .B(c_buf_22__5_), .C(n65), .A(n466), .Y(N652) );
  AO21X1 U914 ( .B(c_buf_22__6_), .C(n676), .A(n427), .Y(N653) );
  AO21X1 U915 ( .B(c_buf_22__7_), .C(n62), .A(n358), .Y(N654) );
  AO21X1 U916 ( .B(wr_buf[0]), .C(n77), .A(n28), .Y(N655) );
  AO21X1 U917 ( .B(wr_buf[1]), .C(n75), .A(n22), .Y(N656) );
  AO21X1 U918 ( .B(wr_buf[2]), .C(n72), .A(n18), .Y(N657) );
  AO21X1 U919 ( .B(wr_buf[3]), .C(n70), .A(n15), .Y(N658) );
  AO21X1 U920 ( .B(wr_buf[4]), .C(n68), .A(n12), .Y(N659) );
  AO21X1 U921 ( .B(wr_buf[5]), .C(n65), .A(n10), .Y(N660) );
  AO21X1 U922 ( .B(wr_buf[6]), .C(n676), .A(n7), .Y(N661) );
  AO21X1 U923 ( .B(wr_buf[7]), .C(n62), .A(n4), .Y(N662) );
  AO21X1 U924 ( .B(n84), .C(n319), .A(n789), .Y(N823) );
  NAND32X1 U925 ( .B(n847), .C(n741), .A(n317), .Y(n319) );
  AOI32X1 U926 ( .A(n788), .B(mcu_psw), .C(n421), .D(n316), .E(n906), .Y(n317)
         );
  AOI21BX1 U927 ( .C(c_adr[12]), .B(memaddr_c[12]), .A(n58), .Y(n127) );
  AOI21X1 U928 ( .B(c_adr[11]), .C(n126), .A(n125), .Y(n58) );
  AND4X1 U929 ( .A(n271), .B(n270), .C(n269), .D(n268), .Y(n272) );
  XOR3X1 U930 ( .A(memaddr_c[13]), .B(c_adr[13]), .C(n263), .Y(n271) );
  XOR3X1 U931 ( .A(c_adr[14]), .B(memaddr_c[14]), .C(n264), .Y(n270) );
  XOR3X1 U932 ( .A(c_adr[12]), .B(memaddr_c[12]), .C(n267), .Y(n268) );
  OA21X1 U933 ( .B(n905), .C(r_pwdn_en), .A(n322), .Y(n324) );
  OAI32X1 U934 ( .A(n118), .B(memaddr_c[8]), .C(n135), .D(n117), .E(n116), .Y(
        n123) );
  AO21X1 U935 ( .B(memaddr_c[8]), .C(n135), .A(n118), .Y(n116) );
  AOI211X1 U936 ( .C(c_adr[7]), .D(n170), .A(n115), .B(n114), .Y(n117) );
  INVX1 U937 ( .A(n94), .Y(n118) );
  INVX1 U938 ( .A(n758), .Y(n759) );
  NAND32X1 U939 ( .B(c_ptr[3]), .C(n764), .A(n773), .Y(n758) );
  INVX1 U940 ( .A(n95), .Y(n100) );
  NAND21X1 U941 ( .B(c_adr[7]), .A(memaddr_c[7]), .Y(n95) );
  AOI32X1 U942 ( .A(c_adr[4]), .B(n97), .C(n106), .D(c_adr[5]), .E(n96), .Y(
        n98) );
  INVXL U943 ( .A(memaddr_c[5]), .Y(n96) );
  NAND2X1 U944 ( .A(hit_ps_c), .B(mcu_psr_c), .Y(n87) );
  NAND21X1 U945 ( .B(c_adr[13]), .A(memaddr_c[13]), .Y(n128) );
  GEN3XL U946 ( .F(n84), .G(n334), .E(n333), .D(n332), .C(n331), .B(n849), .A(
        n330), .Y(n648) );
  AND2X1 U947 ( .A(n329), .B(n333), .Y(n331) );
  INVXL U948 ( .A(memaddr_c[1]), .Y(n103) );
  AND2XL U949 ( .A(c_adr[0]), .B(n198), .Y(n104) );
  NAND21XL U950 ( .B(c_adr[5]), .A(memaddr_c[5]), .Y(n106) );
  AO21X1 U951 ( .B(n844), .C(n823), .A(n822), .Y(n647) );
  MUX2BXL U952 ( .D0(n821), .D1(n820), .S(n839), .Y(n822) );
  AND2X1 U953 ( .A(pmem_re), .B(n818), .Y(n821) );
  NAND21XL U954 ( .B(n81), .A(n819), .Y(n820) );
  AND2X1 U955 ( .A(n282), .B(n336), .Y(N845) );
  XOR2X1 U956 ( .A(c_ptr[3]), .B(n283), .Y(n282) );
  AND2X1 U957 ( .A(n281), .B(n336), .Y(N844) );
  XOR2X1 U958 ( .A(c_ptr[2]), .B(n781), .Y(n281) );
  NOR5X1 U959 ( .A(c_ptr[3]), .B(n306), .C(n305), .D(n25), .E(n767), .Y(n307)
         );
  OAI22XL U960 ( .A(n81), .B(n801), .C(mcu_psw), .D(n800), .Y(n803) );
  NAND21X1 U961 ( .B(c_adr[9]), .A(memaddr_c[9]), .Y(n94) );
  NAND21X1 U962 ( .B(c_adr[14]), .A(memaddr_c[14]), .Y(n130) );
  MUX2X1 U963 ( .D0(n844), .D1(pmem_pgm), .S(n843), .Y(n644) );
  AND2X1 U964 ( .A(n842), .B(n841), .Y(n843) );
  INVXL U965 ( .A(n840), .Y(n842) );
  NAND21X1 U966 ( .B(n51), .A(c_adr[5]), .Y(n239) );
  NAND21X1 U967 ( .B(n340), .A(memaddr[14]), .Y(n799) );
  XOR3X1 U968 ( .A(c_adr[8]), .B(memaddr_c[8]), .C(n258), .Y(n259) );
  NAND21X1 U969 ( .B(n257), .A(n256), .Y(n258) );
  INVX1 U970 ( .A(c_adr[7]), .Y(n257) );
  MUX2X1 U971 ( .D0(n89), .D1(n25), .S(n818), .Y(n649) );
  AND2X1 U972 ( .A(n844), .B(n87), .Y(n89) );
  AND4X1 U973 ( .A(n262), .B(n261), .C(n260), .D(n259), .Y(n273) );
  XOR3X1 U974 ( .A(c_adr[10]), .B(memaddr_c[10]), .C(n254), .Y(n261) );
  XOR3X1 U975 ( .A(c_adr[9]), .B(memaddr_c[9]), .C(n252), .Y(n262) );
  XOR3X1 U976 ( .A(c_adr[7]), .B(memaddr_c[7]), .C(n255), .Y(n260) );
  INVX1 U977 ( .A(cs_n), .Y(pmem_csb) );
  INVX1 U978 ( .A(n312), .Y(n333) );
  NAND21X1 U979 ( .B(d_psrd), .A(n766), .Y(n312) );
  AO21XL U980 ( .B(n84), .C(n313), .A(n333), .Y(N821) );
  NAND32X1 U981 ( .B(n311), .C(n907), .A(n742), .Y(n313) );
  INVX1 U982 ( .A(n837), .Y(n311) );
  NOR21XL U983 ( .B(n826), .A(n824), .Y(n834) );
  NOR43XL U984 ( .B(n895), .C(r_multi), .D(n896), .A(pmem_re), .Y(n824) );
  MUX2X1 U985 ( .D0(n350), .D1(n349), .S(adr_p[14]), .Y(n666) );
  NAND21X1 U986 ( .B(n351), .A(pmem_a[9]), .Y(n349) );
  NAND32X1 U987 ( .B(cs_ft[0]), .C(cs_ft[1]), .A(n315), .Y(n894) );
  OAI22X1 U988 ( .A(adr_p[14]), .B(adr_p[13]), .C(pmem_a[9]), .D(n351), .Y(
        n829) );
  NAND43X1 U989 ( .B(pmem_a[11]), .C(pmem_a[12]), .D(pmem_a[10]), .A(n348), 
        .Y(n351) );
  AND4X1 U990 ( .A(n350), .B(n347), .C(n346), .D(n345), .Y(n348) );
  INVX1 U991 ( .A(pmem_a[15]), .Y(n347) );
  INVX1 U992 ( .A(pmem_a[14]), .Y(n346) );
  INVX1 U993 ( .A(pmem_a[13]), .Y(n345) );
  INVX1 U994 ( .A(n86), .Y(n315) );
  NAND21X1 U995 ( .B(n298), .A(cs_ft[2]), .Y(n86) );
  INVX1 U996 ( .A(adr_p[13]), .Y(n350) );
  NAND43X1 U997 ( .B(cs_ft[1]), .C(cs_ft[3]), .D(cs_ft[0]), .A(cs_ft[2]), .Y(
        n837) );
  OR2X1 U998 ( .A(cs_ft[3]), .B(n287), .Y(n830) );
  NAND21X1 U999 ( .B(cs_ft[2]), .A(n298), .Y(n294) );
  NAND21X1 U1000 ( .B(n314), .A(cs_ft[0]), .Y(n892) );
  OR2X1 U1001 ( .A(cs_ft[0]), .B(n314), .Y(n836) );
  NAND32X1 U1002 ( .B(cs_ft[1]), .C(n298), .A(n300), .Y(n314) );
  NAND32X1 U1003 ( .B(n297), .C(n296), .A(n295), .Y(n893) );
  INVX1 U1004 ( .A(n294), .Y(n295) );
  INVX1 U1005 ( .A(cs_ft[0]), .Y(n296) );
  NAND21X1 U1006 ( .B(cs_ft[1]), .A(cs_ft[0]), .Y(n299) );
  INVX1 U1007 ( .A(cs_ft[1]), .Y(n297) );
  NAND21XL U1008 ( .B(n148), .A(c_adr[1]), .Y(n149) );
  NAND21XL U1009 ( .B(c_adr[1]), .A(n148), .Y(n217) );
  XOR2X1 U1010 ( .A(n140), .B(c_adr[6]), .Y(n165) );
  NAND21X1 U1011 ( .B(n139), .A(c_adr[5]), .Y(n140) );
  INVX1 U1012 ( .A(c_ptr[0]), .Y(n293) );
  INVX1 U1013 ( .A(c_ptr[1]), .Y(n148) );
  INVX1 U1014 ( .A(n132), .Y(n150) );
  NAND21XL U1015 ( .B(n293), .A(c_adr[0]), .Y(n132) );
  NAND21XL U1016 ( .B(n773), .A(c_adr[2]), .Y(n144) );
  NAND21XL U1017 ( .B(c_adr[2]), .A(n773), .Y(n219) );
  XOR2X1 U1018 ( .A(n159), .B(c_adr[5]), .Y(n164) );
  INVX1 U1019 ( .A(c_ptr[2]), .Y(n773) );
  XOR2X1 U1020 ( .A(n177), .B(c_adr[10]), .Y(n181) );
  NAND21X1 U1021 ( .B(n176), .A(c_adr[9]), .Y(n177) );
  XOR2X1 U1022 ( .A(n767), .B(c_adr[4]), .Y(n242) );
  XOR2XL U1023 ( .A(n148), .B(c_adr[1]), .Y(n237) );
  XOR2XL U1024 ( .A(n773), .B(c_adr[2]), .Y(n231) );
  XOR2XL U1025 ( .A(n293), .B(c_adr[0]), .Y(n196) );
  INVX1 U1026 ( .A(n134), .Y(n222) );
  NAND21X1 U1027 ( .B(n767), .A(c_adr[4]), .Y(n134) );
  NAND21X1 U1028 ( .B(c_adr[4]), .A(n767), .Y(n223) );
  XOR2X1 U1029 ( .A(n172), .B(n135), .Y(n174) );
  NAND21X1 U1030 ( .B(n171), .A(c_adr[7]), .Y(n172) );
  INVX1 U1031 ( .A(c_ptr[3]), .Y(n765) );
  INVX1 U1032 ( .A(c_ptr[4]), .Y(n767) );
  XNOR2XL U1033 ( .A(n176), .B(c_adr[9]), .Y(n59) );
  OAI222XL U1034 ( .A(sfr_wdat[7]), .B(n672), .C(n355), .D(n17), .E(
        memdatao[7]), .F(n671), .Y(N793) );
  INVX1 U1035 ( .A(n356), .Y(n355) );
  OAI221XL U1036 ( .A(sfr_wdat[1]), .B(n672), .C(memdatao[1]), .D(n671), .E(
        n619), .Y(N787) );
  OA22X1 U1037 ( .A(n618), .B(n751), .C(n846), .D(n617), .Y(n619) );
  INVX1 U1038 ( .A(n620), .Y(n618) );
  OAI221X1 U1039 ( .A(sfr_wdat[2]), .B(n672), .C(memdatao[2]), .D(n671), .E(
        n579), .Y(N788) );
  OA22X1 U1040 ( .A(n578), .B(n751), .C(n846), .D(n577), .Y(n579) );
  INVX1 U1041 ( .A(n580), .Y(n578) );
  OAI221XL U1042 ( .A(sfr_wdat[3]), .B(n672), .C(memdatao[3]), .D(n671), .E(
        n540), .Y(N789) );
  OA22X1 U1043 ( .A(n539), .B(n751), .C(n846), .D(n538), .Y(n540) );
  INVX1 U1044 ( .A(n541), .Y(n539) );
  OAI221X1 U1045 ( .A(sfr_wdat[4]), .B(n672), .C(memdatao[4]), .D(n671), .E(
        n501), .Y(N790) );
  OA22X1 U1046 ( .A(n500), .B(n751), .C(n846), .D(n499), .Y(n501) );
  INVX1 U1047 ( .A(n502), .Y(n500) );
  OAI221X1 U1048 ( .A(sfr_wdat[5]), .B(n672), .C(memdatao[5]), .D(n671), .E(
        n463), .Y(N791) );
  OA22X1 U1049 ( .A(n462), .B(n17), .C(n846), .D(n461), .Y(n463) );
  INVX1 U1050 ( .A(n464), .Y(n462) );
  OAI221X1 U1051 ( .A(sfr_wdat[6]), .B(n672), .C(memdatao[6]), .D(n671), .E(
        n424), .Y(N792) );
  OA22X1 U1052 ( .A(n423), .B(n17), .C(n846), .D(n422), .Y(n424) );
  INVX1 U1053 ( .A(n425), .Y(n423) );
  OAI221XL U1054 ( .A(sfr_wdat[0]), .B(n672), .C(memdatao[0]), .D(n671), .E(
        n670), .Y(N786) );
  OA22X1 U1055 ( .A(n669), .B(n751), .C(n846), .D(n668), .Y(n670) );
  INVX1 U1056 ( .A(n673), .Y(n669) );
  XNOR2XL U1057 ( .A(n171), .B(c_adr[7]), .Y(n60) );
  INVX1 U1058 ( .A(n133), .Y(n220) );
  XOR2X1 U1059 ( .A(n186), .B(c_adr[12]), .Y(n188) );
  NAND21X1 U1060 ( .B(n185), .A(c_adr[11]), .Y(n186) );
  XOR2X1 U1061 ( .A(n185), .B(c_adr[11]), .Y(n184) );
  XOR2X1 U1062 ( .A(n138), .B(c_adr[13]), .Y(n191) );
  NAND21X1 U1063 ( .B(n138), .A(c_adr[13]), .Y(n137) );
  NAND21X1 U1064 ( .B(n135), .A(c_adr[7]), .Y(n225) );
  NAND21XL U1065 ( .B(c_adr[0]), .A(n293), .Y(n236) );
  NAND2X1 U1066 ( .A(c_adr[11]), .B(n266), .Y(n267) );
  NAND2X1 U1067 ( .A(c_adr[9]), .B(n253), .Y(n254) );
  AND2X1 U1068 ( .A(c_adr[5]), .B(c_adr[6]), .Y(n61) );
  INVX1 U1069 ( .A(c_adr[8]), .Y(n135) );
  INVX1 U1070 ( .A(c_adr[6]), .Y(n99) );
  NAND2X1 U1071 ( .A(c_adr[10]), .B(c_adr[9]), .Y(n226) );
  NAND5XL U1072 ( .A(o_inst[7]), .B(o_inst[6]), .C(o_inst[5]), .D(n738), .E(
        n737), .Y(n859) );
  AND4X1 U1073 ( .A(n860), .B(r_rdy), .C(n861), .D(n733), .Y(n738) );
  AND4X1 U1074 ( .A(o_inst[0]), .B(n736), .C(n735), .D(n734), .Y(n737) );
  NAND21X1 U1075 ( .B(n136), .A(c_adr[11]), .Y(n227) );
  INVX1 U1076 ( .A(c_adr[12]), .Y(n136) );
  INVX1 U1077 ( .A(c_adr[13]), .Y(n228) );
  NAND21X1 U1078 ( .B(c_ptr[1]), .A(n293), .Y(n278) );
  INVX1 U1079 ( .A(c_adr[14]), .Y(n234) );
  NAND43X1 U1080 ( .B(c_ptr[2]), .C(n278), .D(n767), .A(c_ptr[3]), .Y(n289) );
  NAND32X1 U1081 ( .B(cs_ft[0]), .C(n294), .A(n297), .Y(n739) );
  INVX1 U1082 ( .A(d_psrd), .Y(n848) );
  NAND21X1 U1083 ( .B(n616), .A(n353), .Y(n356) );
  MUX2X1 U1084 ( .D0(pmem_q0[7]), .D1(pmem_q1[7]), .S(n667), .Y(n353) );
  NAND21X1 U1085 ( .B(n616), .A(n615), .Y(n620) );
  MUX2X1 U1086 ( .D0(pmem_q0[1]), .D1(pmem_q1[1]), .S(n667), .Y(n615) );
  NAND21X1 U1087 ( .B(n616), .A(n576), .Y(n580) );
  MUX2X1 U1088 ( .D0(pmem_q0[2]), .D1(pmem_q1[2]), .S(n667), .Y(n576) );
  NAND21X1 U1089 ( .B(n616), .A(n537), .Y(n541) );
  MUX2X1 U1090 ( .D0(pmem_q0[3]), .D1(pmem_q1[3]), .S(n667), .Y(n537) );
  NAND21X1 U1091 ( .B(n616), .A(n460), .Y(n464) );
  MUX2X1 U1092 ( .D0(pmem_q0[5]), .D1(pmem_q1[5]), .S(n667), .Y(n460) );
  NAND21X1 U1093 ( .B(n616), .A(n420), .Y(n425) );
  MUX2X1 U1094 ( .D0(pmem_q0[6]), .D1(pmem_q1[6]), .S(n667), .Y(n420) );
  OAI22X1 U1095 ( .A(pmem_q0[4]), .B(n667), .C(pmem_q1[4]), .D(n666), .Y(n502)
         );
  OAI22X1 U1096 ( .A(pmem_q0[0]), .B(n667), .C(pmem_q1[0]), .D(n666), .Y(n673)
         );
  NAND21X1 U1097 ( .B(mcu_psw), .A(n421), .Y(n908) );
  NAND21X1 U1098 ( .B(mcu_psw), .A(n354), .Y(n672) );
  INVX1 U1099 ( .A(memaddr[10]), .Y(n736) );
  INVXL U1100 ( .A(memaddr[0]), .Y(n733) );
  INVX1 U1101 ( .A(memaddr[13]), .Y(n805) );
  INVX1 U1102 ( .A(memaddr[11]), .Y(n735) );
  INVX1 U1103 ( .A(n280), .Y(n781) );
  NAND21X1 U1104 ( .B(n293), .A(c_ptr[1]), .Y(n280) );
  INVX1 U1105 ( .A(n90), .Y(n778) );
  NAND21X1 U1106 ( .B(c_ptr[0]), .A(c_ptr[1]), .Y(n90) );
  INVX1 U1107 ( .A(n91), .Y(n776) );
  NAND21X1 U1108 ( .B(c_ptr[1]), .A(c_ptr[0]), .Y(n91) );
  AO2222XL U1109 ( .A(memaddr_c[0]), .B(n14), .C(pre_1_adr[0]), .D(n344), .E(
        memaddr[0]), .F(n6), .G(sfr_psofs[0]), .H(n9), .Y(N854) );
  XOR2XL U1110 ( .A(memaddr_c[0]), .B(n224), .Y(n276) );
  OA22XL U1111 ( .A(memaddr_c[0]), .B(n196), .C(memaddr_c[1]), .D(n151), .Y(
        n155) );
  INVXL U1112 ( .A(memaddr_c[0]), .Y(n198) );
  AO2222XL U1113 ( .A(memaddr_c[6]), .B(n14), .C(pre_1_adr[6]), .D(n3), .E(
        memaddr[6]), .F(n6), .G(sfr_psofs[6]), .H(n9), .Y(N860) );
  XOR3XL U1114 ( .A(c_adr[6]), .B(memaddr_c[6]), .C(n239), .Y(n250) );
  OAI32XL U1115 ( .A(n100), .B(memaddr_c[6]), .C(n99), .D(n98), .E(n105), .Y(
        n115) );
  AO21XL U1116 ( .B(memaddr_c[6]), .C(n99), .A(n100), .Y(n105) );
  OAI32XL U1117 ( .A(n168), .B(n167), .C(n166), .D(memaddr_c[6]), .E(n165), 
        .Y(n169) );
  AO2222XL U1118 ( .A(memaddr_c[3]), .B(n14), .C(pre_1_adr[3]), .D(n344), .E(
        memaddr[3]), .F(n6), .G(sfr_psofs[3]), .H(n9), .Y(N857) );
  XOR2XL U1119 ( .A(memaddr_c[3]), .B(n247), .Y(n248) );
  NAND21XL U1120 ( .B(c_adr[3]), .A(memaddr_c[3]), .Y(n102) );
  NAND21XL U1121 ( .B(n143), .A(memaddr_c[3]), .Y(n203) );
  OA22XL U1122 ( .A(memaddr_c[3]), .B(n147), .C(memaddr_c[2]), .D(n146), .Y(
        n158) );
  AO2222XL U1123 ( .A(memaddr_c[4]), .B(n14), .C(pre_1_adr[4]), .D(n3), .E(
        memaddr[4]), .F(n6), .G(sfr_psofs[4]), .H(n9), .Y(N858) );
  XOR2XL U1124 ( .A(memaddr_c[4]), .B(n243), .Y(n249) );
  AOI221XL U1125 ( .A(memaddr_c[4]), .B(n113), .C(n112), .D(n111), .E(n110), 
        .Y(n114) );
  INVXL U1126 ( .A(memaddr_c[4]), .Y(n97) );
  NAND21XL U1127 ( .B(n156), .A(memaddr_c[4]), .Y(n205) );
  MAJ3X1 U1128 ( .A(c_adr[1]), .B(n104), .C(n103), .Y(n108) );
  INVX1 U1129 ( .A(wspp_cnt[0]), .Y(N353) );
  OR2X1 U1130 ( .A(wspp_cnt[1]), .B(wspp_cnt[0]), .Y(n852) );
  OAI21BBX1 U1131 ( .A(wspp_cnt[0]), .B(wspp_cnt[1]), .C(n852), .Y(N354) );
  OR2X1 U1132 ( .A(n852), .B(wspp_cnt[2]), .Y(n853) );
  OAI21BBX1 U1133 ( .A(n852), .B(wspp_cnt[2]), .C(n853), .Y(N355) );
  OR2X1 U1134 ( .A(n853), .B(wspp_cnt[3]), .Y(n854) );
  OAI21BBX1 U1135 ( .A(n853), .B(wspp_cnt[3]), .C(n854), .Y(N356) );
  OR2X1 U1136 ( .A(n854), .B(wspp_cnt[4]), .Y(n855) );
  OAI21BBX1 U1137 ( .A(n854), .B(wspp_cnt[4]), .C(n855), .Y(N357) );
  XNOR2XL U1138 ( .A(n855), .B(wspp_cnt[5]), .Y(N358) );
  OR2X1 U1139 ( .A(wspp_cnt[5]), .B(n855), .Y(n856) );
  XNOR2XL U1140 ( .A(wspp_cnt[6]), .B(n856), .Y(N359) );
  NAND2X1 U1141 ( .A(n858), .B(n859), .Y(o_set_hold) );
  NOR4XL U1142 ( .A(n862), .B(memaddr[4]), .C(memaddr[6]), .D(memaddr[5]), .Y(
        n861) );
  OR3XL U1143 ( .A(memaddr[8]), .B(memaddr[9]), .C(memaddr[7]), .Y(n862) );
  NOR4XL U1144 ( .A(n863), .B(memaddr[12]), .C(memaddr[14]), .D(memaddr[13]), 
        .Y(n860) );
  OR3XL U1145 ( .A(memaddr[2]), .B(memaddr[3]), .C(memaddr[1]), .Y(n863) );
  INVX1 U1146 ( .A(n858), .Y(o_bkp_hold) );
  NAND2X1 U1147 ( .A(n864), .B(n865), .Y(n858) );
  NOR4XL U1148 ( .A(n866), .B(n867), .C(n868), .D(n869), .Y(n865) );
  XOR2X1 U1149 ( .A(bkpt_pc[10]), .B(memaddr[10]), .Y(n869) );
  XOR2X1 U1150 ( .A(bkpt_pc[0]), .B(memaddr[0]), .Y(n868) );
  NAND32X1 U1151 ( .B(un_hold), .C(n845), .A(bkpt_ena), .Y(n867) );
  NAND4X1 U1152 ( .A(n870), .B(n871), .C(n872), .D(n873), .Y(n866) );
  XNOR2XL U1153 ( .A(memaddr[11]), .B(bkpt_pc[11]), .Y(n873) );
  XNOR2XL U1154 ( .A(memaddr[12]), .B(bkpt_pc[12]), .Y(n872) );
  XNOR2XL U1155 ( .A(memaddr[13]), .B(bkpt_pc[13]), .Y(n871) );
  XNOR2XL U1156 ( .A(memaddr[14]), .B(bkpt_pc[14]), .Y(n870) );
  NOR4XL U1157 ( .A(n874), .B(n875), .C(n876), .D(n877), .Y(n864) );
  XOR2X1 U1158 ( .A(bkpt_pc[5]), .B(memaddr[5]), .Y(n877) );
  XOR2X1 U1159 ( .A(bkpt_pc[4]), .B(memaddr[4]), .Y(n876) );
  NAND3X1 U1160 ( .A(n878), .B(n879), .C(n880), .Y(n875) );
  XNOR2XL U1161 ( .A(memaddr[2]), .B(bkpt_pc[2]), .Y(n880) );
  XNOR2XL U1162 ( .A(memaddr[3]), .B(bkpt_pc[3]), .Y(n879) );
  XNOR2XL U1163 ( .A(memaddr[1]), .B(bkpt_pc[1]), .Y(n878) );
  NAND4X1 U1164 ( .A(n881), .B(n882), .C(n883), .D(n884), .Y(n874) );
  XNOR2XL U1165 ( .A(memaddr[6]), .B(bkpt_pc[6]), .Y(n884) );
  XNOR2XL U1166 ( .A(memaddr[7]), .B(bkpt_pc[7]), .Y(n883) );
  XNOR2XL U1167 ( .A(memaddr[8]), .B(bkpt_pc[8]), .Y(n882) );
  XNOR2XL U1168 ( .A(memaddr[9]), .B(bkpt_pc[9]), .Y(n881) );
  MUX2IX1 U1169 ( .D0(n885), .D1(n886), .S(n887), .Y(n651) );
  NAND3X1 U1170 ( .A(n888), .B(n85), .C(dummy[0]), .Y(n885) );
  MUX2IX1 U1171 ( .D0(n889), .D1(n890), .S(n887), .Y(n650) );
  AND4X1 U1172 ( .A(dw_ena), .B(sfr_psw), .C(n888), .D(n85), .Y(n887) );
  NAND2X1 U1173 ( .A(dummy[0]), .B(n891), .Y(n890) );
  NAND3X1 U1174 ( .A(n888), .B(n85), .C(dummy[1]), .Y(n889) );
  INVX1 U1175 ( .A(dw_rst), .Y(n888) );
  NAND21X1 U1176 ( .B(wspp_cnt[4]), .A(n897), .Y(n896) );
  OAI21AX1 U1177 ( .B(wspp_cnt[3]), .C(n898), .A(wspp_cnt[6]), .Y(n897) );
  MUX2IX1 U1178 ( .D0(n899), .D1(n900), .S(wspp_cnt[5]), .Y(n895) );
  AND2X1 U1179 ( .A(n901), .B(wspp_cnt[4]), .Y(n900) );
  OAI21X1 U1180 ( .B(wspp_cnt[6]), .C(n898), .A(n901), .Y(n899) );
  NAND2X1 U1181 ( .A(wspp_cnt[6]), .B(wspp_cnt[3]), .Y(n901) );
  MUX2IX1 U1182 ( .D0(n857), .D1(n845), .S(n850), .Y(mempsack) );
  NAND21X1 U1183 ( .B(rd_buf[7]), .A(d_psrd), .Y(d_inst[7]) );
  NAND21X1 U1184 ( .B(rd_buf[6]), .A(n25), .Y(d_inst[6]) );
  NAND21X1 U1185 ( .B(rd_buf[5]), .A(n25), .Y(d_inst[5]) );
  AND2X1 U1186 ( .A(rd_buf[4]), .B(n25), .Y(d_inst[4]) );
  NAND21X1 U1187 ( .B(rd_buf[3]), .A(n25), .Y(d_inst[3]) );
  NAND21X1 U1188 ( .B(rd_buf[2]), .A(d_psrd), .Y(d_inst[2]) );
  NAND21X1 U1189 ( .B(rd_buf[1]), .A(d_psrd), .Y(d_inst[1]) );
  AND2X1 U1190 ( .A(rd_buf[0]), .B(n25), .Y(d_inst[0]) );
  INVX1 U1191 ( .A(n902), .Y(N974) );
  AOI31X1 U1192 ( .A(un_hold), .B(n85), .C(n845), .D(n923), .Y(n902) );
  NOR2X1 U1193 ( .A(n903), .B(srst), .Y(n923) );
  OAI31XL U1194 ( .A(n908), .B(wr_buf[0]), .C(n851), .D(n894), .Y(n907) );
  NAND2X1 U1195 ( .A(n912), .B(n891), .Y(n886) );
  INVX1 U1196 ( .A(dummy[1]), .Y(n891) );
  INVX1 U1197 ( .A(dummy[0]), .Y(n912) );
  OAI31XL U1198 ( .A(n892), .B(n849), .C(n913), .D(n893), .Y(n909) );
  INVX1 U1199 ( .A(n905), .Y(n913) );
  NAND2X1 U1200 ( .A(n910), .B(n911), .Y(n905) );
  NAND2X1 U1201 ( .A(mcu_psw), .B(hit_ps), .Y(n911) );
  NAND4X1 U1202 ( .A(d_hold[3]), .B(d_hold[2]), .C(n914), .D(d_hold[1]), .Y(
        n910) );
  NOR2X1 U1203 ( .A(n903), .B(n915), .Y(n914) );
  INVX1 U1204 ( .A(r_hold_mcu), .Y(n903) );
  NOR41XL U1205 ( .D(n898), .A(wspp_cnt[0]), .B(wspp_cnt[2]), .C(wspp_cnt[1]), 
        .Y(n904) );
  NOR4XL U1206 ( .A(wspp_cnt[3]), .B(wspp_cnt[4]), .C(wspp_cnt[5]), .D(
        wspp_cnt[6]), .Y(n898) );
  OAI21BBX1 U1207 ( .A(N359), .B(n20), .C(n908), .Y(N801) );
  OAI21BBX1 U1208 ( .A(N358), .B(n847), .C(n908), .Y(N800) );
  OAI21BBX1 U1209 ( .A(N357), .B(n847), .C(n908), .Y(N799) );
  AND2X1 U1210 ( .A(N356), .B(n20), .Y(N798) );
  OAI21BBX1 U1211 ( .A(N355), .B(n847), .C(n908), .Y(N797) );
  OAI21BBX1 U1212 ( .A(N354), .B(n847), .C(n908), .Y(N796) );
  OAI21BBX1 U1213 ( .A(N353), .B(n847), .C(n908), .Y(N795) );
  MUX2IX1 U1214 ( .D0(n916), .D1(n917), .S(pmem_a[8]), .Y(N759) );
  AOI21X1 U1215 ( .B(n918), .C(n919), .A(N757), .Y(n917) );
  MUX2BXL U1216 ( .D0(N757), .D1(n920), .S(n919), .Y(N758) );
  INVX1 U1217 ( .A(pmem_a[7]), .Y(n919) );
  NAND2X1 U1218 ( .A(pmem_a[6]), .B(n918), .Y(n920) );
  NOR21XL U1219 ( .B(n918), .A(pmem_a[6]), .Y(N757) );
  NOR2X1 U1220 ( .A(n851), .B(n846), .Y(n918) );
  NAND2X1 U1221 ( .A(n921), .B(n922), .Y(n906) );
  NOR4XL U1222 ( .A(wr_buf[7]), .B(wr_buf[6]), .C(wr_buf[5]), .D(wr_buf[4]), 
        .Y(n922) );
  NOR4XL U1223 ( .A(wr_buf[3]), .B(wr_buf[2]), .C(wr_buf[1]), .D(wr_buf[0]), 
        .Y(n921) );
  AND2X1 U1224 ( .A(d_hold[2]), .B(n85), .Y(N154) );
  AND2X1 U1225 ( .A(d_hold[1]), .B(n85), .Y(N153) );
  NOR2X1 U1226 ( .A(srst), .B(n915), .Y(N152) );
  INVX1 U1227 ( .A(d_hold[0]), .Y(n915) );
  INVX1 U1228 ( .A(n857), .Y(o_ofs_inc) );
endmodule


module ictlr_a0_DW01_inc_2 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1XL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module ictlr_a0_DW01_inc_1 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  HAD1XL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  XOR2X1 U1 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mcu51_a0 ( bclki2c, pc_ini, slp2wakeup, r_hold_mcu, wdt_slow, wdtov, 
        mdubsy, cs_run, t0_intr, clki2c, clkmdu, clkur0, clktm0, clktm1, 
        clkwdt, i2c_autoack, i2c_con_ens1, clkcpu, clkper, reset, ro, port0i, 
        exint_9, exint, clkcpuen, clkperen, port0o, port0ff, rxd0o, txd0, 
        rxd0i, rxd0oe, scli, sdai, sclo, sdao, waitstaten, mempsack, memack, 
        memdatai, memdatao, memaddr, mempswr, mempsrd, memwr, memrd, 
        memdatao_comb, memaddr_comb, mempswr_comb, mempsrd_comb, memwr_comb, 
        memrd_comb, ramdatai, ramdatao, ramaddr, ramwe, ramoe, dbgpo, sfrack, 
        sfrdatai, sfrdatao, sfraddr, sfrwe, sfroe, esfrm_wrdata, esfrm_addr, 
        esfrm_we, esfrm_oe, esfrm_rddata );
  input [15:0] pc_ini;
  output [1:0] wdtov;
  input [7:0] port0i;
  input [7:0] exint;
  output [7:0] port0o;
  output [7:0] port0ff;
  input [7:0] memdatai;
  output [7:0] memdatao;
  output [15:0] memaddr;
  output [7:0] memdatao_comb;
  output [15:0] memaddr_comb;
  input [7:0] ramdatai;
  output [7:0] ramdatao;
  output [7:0] ramaddr;
  output [31:0] dbgpo;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  output [6:0] sfraddr;
  input [7:0] esfrm_wrdata;
  input [6:0] esfrm_addr;
  output [7:0] esfrm_rddata;
  input bclki2c, slp2wakeup, r_hold_mcu, wdt_slow, clki2c, clkmdu, clkur0,
         clktm0, clktm1, clkwdt, i2c_autoack, clkcpu, clkper, reset, exint_9,
         rxd0i, scli, sdai, mempsack, memack, sfrack, esfrm_we, esfrm_oe;
  output mdubsy, cs_run, t0_intr, i2c_con_ens1, ro, clkcpuen, clkperen, rxd0o,
         txd0, rxd0oe, sclo, sdao, waitstaten, mempswr, mempsrd, memwr, memrd,
         mempswr_comb, mempsrd_comb, memwr_comb, memrd_comb, ramwe, ramoe,
         sfrwe, sfroe;
  wire   n122, n123, n124, n125, n126, n127, n128, n129, N7, N8, N9, N10, N11,
         N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, t0_tf1, t1_tf1, t0_tr1,
         t1_tr1, stop_flag, idle_flag, sfroe_s, sfroe_mcu51_per, sfrwe_s,
         sfrwe_mcu51_per, newinstr, intcall_int, cpu_resume, rmwinstr, pmw,
         p2sel, gf0, c, ac, ov, f0, f1, p, rsttowdt, rsttosrst, rst, int0ff,
         int1ff, rxd0ff, sdaiff, rsttowdtff, rsttosrstff, resetff, smod,
         ip0wdts, wdt_tm, bd, ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6,
         iex7, iex8, iex9, isr_tm, i2c_int, i2ccon_o_7, tf1_gate, riti0_gate,
         iex7_gate, iex2_gate, srstflag, int_vect_8b, int_vect_93, int_vect_9b,
         int_vect_a3, wdts, srst, pmuintreq_rev, pmuintreq, t1ov, t0ack, t1ack,
         isr_irq, int0ack, int1ack, iex7ack, iex2ack, iex3ack, iex4ack,
         iex5ack, iex6ack, iex8ack, iex9ack, n6, n7, n8, n9, n10, n11, n1, n2,
         n3, n5, n12, n14, n15, n16, n18, n19, n21, n22, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n45, n46, n48, n49, n50, n52, n53,
         n54, n55, n56, n58, n59, n60, n61, n62, n63, n65, n67, n69, n72, n73,
         n75, n77, n79, n80, n81, n82, n83, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5;
  wire   [13:0] timer_1ms;
  wire   [5:0] ien2;
  wire   [6:0] ramsfraddr;
  wire   [4:0] intvect_int;
  wire   [7:0] ckcon;
  wire   [7:0] dph;
  wire   [7:0] dpl;
  wire   [3:0] dps;
  wire   [7:0] p2;
  wire   [5:0] dpc;
  wire   [7:0] sp;
  wire   [7:0] acc_s;
  wire   [7:0] b;
  wire   [1:0] rs;
  wire   [7:0] arcon;
  wire   [7:0] md0;
  wire   [7:0] md1;
  wire   [7:0] md2;
  wire   [7:0] md3;
  wire   [7:0] md4;
  wire   [7:0] md5;
  wire   [3:0] t0_tmod;
  wire   [7:0] tl0;
  wire   [7:0] th0;
  wire   [3:0] t1_tmod;
  wire   [7:0] tl1;
  wire   [7:0] th1;
  wire   [7:0] wdtrel;
  wire   [6:5] t2con;
  wire   [7:0] s0con;
  wire   [7:0] s0buf;
  wire   [7:0] s0rell;
  wire   [7:0] s0relh;
  wire   [7:0] ien0;
  wire   [5:0] ien1;
  wire   [5:0] ip0;
  wire   [5:0] ip1;
  wire   [7:0] i2cdat_o;
  wire   [7:0] i2cadr_o;
  wire   [5:0] i2ccon_o;
  wire   [7:0] i2csta_o;
  wire   [3:0] isreg;

  mcu51_cpu_a0 u_cpu ( .clkcpu(clkcpu), .rst(dbgpo[22]), .mempsack(mempsack), 
        .memack(memack), .memdatai(memdatai), .memaddr(memaddr), .mempsrd(
        mempsrd), .mempswr(mempswr), .memrd(memrd), .memwr(memwr), 
        .memaddr_comb(memaddr_comb), .mempsrd_comb(mempsrd_comb), 
        .mempswr_comb(mempswr_comb), .memrd_comb(memrd_comb), .memwr_comb(
        memwr_comb), .cpu_hold(r_hold_mcu), .cpu_resume(cpu_resume), .irq(
        dbgpo[20]), .intvect(intvect_int), .intcall(intcall_int), .retiinstr(
        dbgpo[21]), .newinstr(newinstr), .rmwinstr(rmwinstr), .waitstaten(
        waitstaten), .ramdatai(ramdatai), .sfrdatai({esfrm_rddata[7:2], n128, 
        n129}), .ramsfraddr({SYNOPSYS_UNCONNECTED_1, ramsfraddr}), .ramdatao(
        memdatao), .ramoe(), .ramwe(), .sfroe(sfroe_s), .sfrwe(sfrwe_s), 
        .sfroe_r(), .sfrwe_r(), .sfroe_comb_s(), .sfrwe_comb_s(), .pc_o(
        dbgpo[15:0]), .pc_ini(pc_ini), .cs_run(cs_run), .instr(dbgpo[31:24]), 
        .codefetch_s(), .sfrack(sfrack), .ramsfraddr_comb(ramaddr), 
        .ramdatao_comb(ramdatao), .ramoe_comb(ramoe), .ramwe_comb(ramwe), 
        .ckcon(ckcon), .pmw(pmw), .p2sel(p2sel), .gf0(gf0), .stop(stop_flag), 
        .idle(idle_flag), .acc(acc_s), .b(b), .rs(rs), .c(c), .ac(ac), .ov(ov), 
        .p(p), .f0(f0), .f1(f1), .dph(dph), .dpl(dpl), .dps(dps), .dpc(dpc), 
        .p2(p2), .sp(sp) );
  syncneg_a0 u_syncneg ( .clk(clkper), .reset(n79), .rsttowdt(rsttowdt), 
        .rsttosrst(rsttosrst), .rst(rst), .int0(exint[0]), .int1(exint[1]), 
        .port0i(port0i), .rxd0i(rxd0i), .sdai(sdai), .int0ff(int0ff), .int1ff(
        int1ff), .port0ff(port0ff), .t0ff(), .t1ff(), .rxd0ff(rxd0ff), 
        .sdaiff(sdaiff), .rsttowdtff(rsttowdtff), .rsttosrstff(rsttosrstff), 
        .rstff(n122), .resetff(resetff) );
  sfrmux_a0 u_sfrmux ( .isfrwait(n112), .sfraddr({sfraddr[6], n60, n14, n34, 
        sfraddr[2:1], n49}), .c(c), .ac(ac), .f0(f0), .rs(rs), .ov(ov), .f1(f1), .p(p), .acc(acc_s), .b(b), .dpl(dpl), .dph(dph), .dps(dps), .dpc(dpc), .p2(
        p2), .sp(sp), .smod(smod), .pmw(pmw), .p2sel(p2sel), .gf0(gf0), .stop(
        stop_flag), .idle(idle_flag), .ckcon(ckcon), .port0(port0o), .port0ff(
        port0ff), .rmwinstr(rmwinstr), .arcon(arcon), .md0(md0), .md1(md1), 
        .md2(md2), .md3(md3), .md4(md4), .md5(md5), .t0_tmod(t0_tmod), 
        .t0_tf0(dbgpo[17]), .t0_tf1(t0_tf1), .t0_tr0(dbgpo[16]), .t0_tr1(
        t0_tr1), .tl0(tl0), .th0(th0), .t1_tmod(t1_tmod), .t1_tf1(t1_tf1), 
        .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1), .wdtrel(wdtrel), .ip0wdts(
        ip0wdts), .wdt_tm(wdt_tm), .t2con({1'b0, t2con, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .s0con(s0con), .s0buf(s0buf), .s0rell(s0rell), .s0relh(s0relh), 
        .bd(bd), .ie0(ie0), .it0(it0), .ie1(ie1), .it1(it1), .iex2(iex2), 
        .iex3(iex3), .iex4(iex4), .iex5(iex5), .iex6(iex6), .iex7(iex7), 
        .iex8(iex8), .iex9(iex9), .iex10(1'b0), .iex11(1'b0), .iex12(1'b0), 
        .ien0({ien0[7], 1'b0, ien0[5:0]}), .ien1(ien1), .ien2(ien2), .ip0(ip0), 
        .ip1(ip1), .isr_tm(isr_tm), .i2c_int(i2c_int), .i2cdat_o(i2cdat_o), 
        .i2cadr_o(i2cadr_o), .i2ccon_o({i2ccon_o_7, i2c_con_ens1, i2ccon_o}), 
        .i2csta_o({i2csta_o[7:3], 1'b0, 1'b0, 1'b0}), .sfrdatai(sfrdatai), 
        .tf1_gate(tf1_gate), .riti0_gate(riti0_gate), .iex7_gate(iex7_gate), 
        .iex2_gate(iex2_gate), .srstflag(srstflag), .int_vect_8b(int_vect_8b), 
        .int_vect_93(int_vect_93), .int_vect_9b(int_vect_9b), .int_vect_a3(
        int_vect_a3), .ext_sfr_sel(), .sfrdatao({esfrm_rddata[7:2], n128, n129}) );
  pmurstctrl_a0 u_pmurstctrl ( .resetff(resetff), .wdts(wdts), .srst(srst), 
        .pmuintreq(pmuintreq_rev), .stop(stop_flag), .idle(idle_flag), 
        .clkcpu_en(clkcpuen), .clkper_en(clkperen), .cpu_resume(cpu_resume), 
        .rsttowdt(rsttowdt), .rsttosrst(rsttosrst), .rst(rst) );
  wakeupctrl_a0 u_wakeupctrl ( .irq(dbgpo[20]), .int0ff(exint[0]), .int1ff(
        exint[1]), .it0(it0), .it1(it1), .isreg(isreg), .intprior0({ip0[2], 
        ip0[0]}), .intprior1({ip1[2], ip1[0]}), .eal(ien0[7]), .eint0(ien0[0]), 
        .eint1(ien0[2]), .pmuintreq(pmuintreq) );
  mdu_a0 u_mdu ( .clkper(clkmdu), .rst(n81), .mdubsy(mdubsy), .sfrdatai({
        sfrdatao[7], n75, n73, sfrdatao[4], n69, n67, sfrdatao[1:0]}), 
        .sfraddr({n63, n28, n5, sfraddr[3], n56, n52, n3}), .sfrwe(
        sfrwe_mcu51_per), .sfroe(sfroe_mcu51_per), .arcon(arcon), .md0(md0), 
        .md1(md1), .md2(md2), .md3(md3), .md4(md4), .md5(md5) );
  ports_a0 u_ports ( .clkper(clkper), .rst(dbgpo[22]), .port0(port0o), 
        .sfrdatai({sfrdatao[7], n75, sfrdatao[5:4], n69, n67, sfrdatao[1:0]}), 
        .sfraddr({n29, n28, n12, sfraddr[3], n56, n53, n26}), .sfrwe(n32) );
  serial0_a0 u_serial0 ( .t_shift_clk(), .r_shift_clk(), .clkper(clkur0), 
        .rst(dbgpo[22]), .newinstr(newinstr), .rxd0ff(rxd0ff), .t1ov(t1ov), 
        .rxd0o(rxd0o), .rxd0oe(rxd0oe), .txd0(txd0), .sfrdatai({n77, 
        sfrdatao[6:4], n69, n67, sfrdatao[1], n65}), .sfraddr({n63, n61, n12, 
        n58, n55, n53, n2}), .sfrwe(n32), .s0con(s0con), .s0buf(s0buf), 
        .s0rell(s0rell), .s0relh(s0relh), .smod(smod), .bd(bd) );
  timer0_a0 u_timer0 ( .clkper(clktm0), .rst(dbgpo[22]), .newinstr(newinstr), 
        .t0ff(1'b0), .t0ack(t0ack), .t1ack(t1ack), .int0ff(int0ff), .t0_tf0(
        dbgpo[17]), .t0_tf1(t0_tf1), .sfrdatai({sfrdatao[7], n75, 
        sfrdatao[5:2], n125, n126}), .sfraddr({n29, n28, n5, sfraddr[3], n55, 
        n52, n26}), .sfrwe(n32), .t0_tmod(t0_tmod), .t0_tr0(dbgpo[16]), 
        .t0_tr1(t0_tr1), .tl0(tl0), .th0(th0) );
  timer1_a0 u_timer1 ( .clkper(clktm1), .rst(n82), .newinstr(newinstr), .t1ff(
        1'b0), .t1ack(t1ack), .int1ff(int1ff), .t1_tf1(t1_tf1), .t1ov(t1ov), 
        .sfrdatai({sfrdatao[7], n75, sfrdatao[5], n72, n69, n67, sfrdatao[1], 
        n65}), .sfraddr({n29, n28, n12, sfraddr[3], n55, n52, n26}), .sfrwe(
        n32), .t1_tmod(t1_tmod), .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1) );
  watchdog_a0 u_watchdog ( .wdt_slow(wdt_slow), .clkwdt(clkwdt), .clkper(
        clkper), .resetff(rsttowdtff), .newinstr(newinstr), .wdts_s(wdtov), 
        .wdts(wdts), .ip0wdts(ip0wdts), .wdt_tm(wdt_tm), .sfrdatai({
        sfrdatao[7:4], n69, n67, sfrdatao[1:0]}), .sfraddr({n63, n61, n5, n58, 
        n56, n53, n3}), .sfrwe(n32), .wdtrel(wdtrel) );
  isr_a0 u_isr ( .clkper(clkper), .rst(n83), .intcall(intcall_int), 
        .retiinstr(dbgpo[21]), .int_vect_03(ie0), .int_vect_0b(dbgpo[17]), 
        .t0ff(1'b0), .int_vect_13(ie1), .int_vect_1b(tf1_gate), .t1ff(1'b0), 
        .int_vect_23(riti0_gate), .i2c_int(i2c_int), .rxd0ff(rxd0ff), 
        .int_vect_43(iex7_gate), .sdaiff(sdaiff), .int_vect_4b(iex2_gate), 
        .int_vect_53(iex3), .int_vect_5b(iex4), .int_vect_63(iex5), 
        .int_vect_6b(iex6), .int_vect_8b(int_vect_8b), .int_vect_93(
        int_vect_93), .int_vect_9b(int_vect_9b), .int_vect_a3(int_vect_a3), 
        .int_vect_ab(1'b0), .irq(isr_irq), .intvect(intvect_int), .int_ack_03(
        int0ack), .int_ack_0b(t0ack), .int_ack_13(int1ack), .int_ack_1b(t1ack), 
        .int_ack_43(iex7ack), .int_ack_4b(iex2ack), .int_ack_53(iex3ack), 
        .int_ack_5b(iex4ack), .int_ack_63(iex5ack), .int_ack_6b(iex6ack), 
        .int_ack_8b(iex8ack), .int_ack_93(iex9ack), .int_ack_9b(), 
        .int_ack_a3(), .int_ack_ab(), .is_reg(isreg), .ip0(ip0), .ip1(ip1), 
        .ien0({ien0[7], SYNOPSYS_UNCONNECTED_2, ien0[5:0]}), .ien1(ien1), 
        .ien2(ien2), .isr_tm(isr_tm), .sfraddr({n29, n28, n5, n58, n56, n53, 
        n48}), .sfrdatai({sfrdatao[7:6], n73, n72, sfrdatao[3], n124, n125, 
        n126}), .sfrwe(n32) );
  extint_a0 u_extint ( .clkper(clkper), .rst(dbgpo[22]), .newinstr(newinstr), 
        .int0ff(int0ff), .int0ack(int0ack), .int1ff(int1ff), .int1ack(int1ack), 
        .int2ff(exint[2]), .iex2ack(iex2ack), .int3ff(exint[3]), .iex3ack(
        iex3ack), .int4ff(exint[4]), .iex4ack(iex4ack), .int5ff(exint[5]), 
        .iex5ack(iex5ack), .int6ff(exint[6]), .iex6ack(iex6ack), .int7ff(
        exint[7]), .iex7ack(iex7ack), .int8ff(n11), .iex8ack(iex8ack), 
        .int9ff(exint_9), .iex9ack(iex9ack), .ie0(ie0), .it0(it0), .ie1(ie1), 
        .it1(it1), .i2fr(t2con[5]), .iex2(iex2), .i3fr(t2con[6]), .iex3(iex3), 
        .iex4(iex4), .iex5(iex5), .iex6(iex6), .iex7(iex7), .iex8(iex8), 
        .iex9(iex9), .iex10(), .iex11(), .iex12(), .sfraddr({n63, n28, n12, 
        sfraddr[3], n56, n53, n26}), .sfrdatai({sfrdatao[7], n75, 
        sfrdatao[5:3], n67, sfrdatao[1:0]}), .sfrwe(n32) );
  i2c_a0 u_i2c ( .clk(clki2c), .rst(ro), .bclksel(bclki2c), .scli(scli), 
        .sdai(sdai), .sclo(sclo), .sdao(sdao), .intack(i2c_autoack), .si(
        i2c_int), .sfrwe(sfrwe_mcu51_per), .sfraddr({n63, n28, n5, sfraddr[3], 
        n55, n53, n48}), .sfrdatai({n77, sfrdatao[6], n123, sfrdatao[4], n69, 
        sfrdatao[2], n125, n65}), .i2cdat_o(i2cdat_o), .i2cadr_o(i2cadr_o), 
        .i2ccon_o({i2ccon_o_7, i2c_con_ens1, i2ccon_o}), .i2csta_o({
        i2csta_o[7:3], SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5}) );
  softrstctrl_a0 u_softrstctrl ( .clkcpu(clkcpu), .resetff(rsttosrstff), 
        .newinstr(newinstr), .srstreq(srst), .srstflag(srstflag), .sfrdatai({
        sfrdatao[7:6], n73, n72, sfrdatao[3:2], n125, n65}), .sfraddr({n63, 
        n61, n12, n58, n56, n53, n26}), .sfrwe(n32) );
  mcu51_a0_DW01_inc_0 add_268 ( .A(timer_1ms), .SUM({N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7}) );
  DFFQX1 timer_1ms_reg_13_ ( .D(N34), .C(clkper), .Q(timer_1ms[13]) );
  DFFQX1 timer_1ms_reg_8_ ( .D(N29), .C(clkper), .Q(timer_1ms[8]) );
  DFFQX1 timer_1ms_reg_9_ ( .D(N30), .C(clkper), .Q(timer_1ms[9]) );
  DFFQX1 timer_1ms_reg_10_ ( .D(N31), .C(clkper), .Q(timer_1ms[10]) );
  DFFQX1 timer_1ms_reg_11_ ( .D(N32), .C(clkper), .Q(timer_1ms[11]) );
  DFFQX1 timer_1ms_reg_12_ ( .D(N33), .C(clkper), .Q(timer_1ms[12]) );
  DFFQX1 timer_1ms_reg_5_ ( .D(N26), .C(clkper), .Q(timer_1ms[5]) );
  DFFQX1 timer_1ms_reg_6_ ( .D(N27), .C(clkper), .Q(timer_1ms[6]) );
  DFFQX1 timer_1ms_reg_7_ ( .D(N28), .C(clkper), .Q(timer_1ms[7]) );
  DFFQX1 timer_1ms_reg_4_ ( .D(N25), .C(clkper), .Q(timer_1ms[4]) );
  DFFQX1 timer_1ms_reg_3_ ( .D(N24), .C(clkper), .Q(timer_1ms[3]) );
  DFFQX1 timer_1ms_reg_2_ ( .D(N23), .C(clkper), .Q(timer_1ms[2]) );
  DFFQX1 timer_1ms_reg_1_ ( .D(N22), .C(clkper), .Q(timer_1ms[1]) );
  DFFQX1 timer_1ms_reg_0_ ( .D(N21), .C(clkper), .Q(timer_1ms[0]) );
  INVXL U3 ( .A(sfraddr[2]), .Y(n24) );
  INVX3 U4 ( .A(n54), .Y(sfraddr[1]) );
  INVX3 U5 ( .A(n33), .Y(n54) );
  MUX2X2 U6 ( .D0(esfrm_addr[0]), .D1(ramsfraddr[0]), .S(n92), .Y(n19) );
  INVXL U7 ( .A(n34), .Y(n59) );
  INVX2 U8 ( .A(n19), .Y(n50) );
  INVX1 U9 ( .A(ramsfraddr[4]), .Y(n16) );
  INVX1 U10 ( .A(esfrm_addr[4]), .Y(n15) );
  INVX2 U11 ( .A(n50), .Y(sfraddr[0]) );
  INVX2 U12 ( .A(esfrm_we), .Y(n89) );
  INVX2 U13 ( .A(n62), .Y(n60) );
  INVX2 U14 ( .A(n50), .Y(n49) );
  INVX6 U15 ( .A(n93), .Y(sfraddr[6]) );
  INVXL U16 ( .A(n14), .Y(n18) );
  INVXL U17 ( .A(n48), .Y(n1) );
  INVXL U18 ( .A(n1), .Y(n2) );
  INVXL U19 ( .A(n1), .Y(n3) );
  INVXL U20 ( .A(n18), .Y(sfraddr[4]) );
  INVXL U21 ( .A(n18), .Y(n5) );
  INVXL U22 ( .A(n18), .Y(n12) );
  BUFXL U23 ( .A(n128), .Y(esfrm_rddata[1]) );
  MUX2IX4 U24 ( .D0(n15), .D1(n16), .S(n21), .Y(n14) );
  MUX2X1 U25 ( .D0(esfrm_addr[1]), .D1(ramsfraddr[1]), .S(n92), .Y(n33) );
  MUX2X1 U26 ( .D0(esfrm_addr[3]), .D1(ramsfraddr[3]), .S(n92), .Y(n34) );
  MUX2X2 U27 ( .D0(ramsfraddr[2]), .D1(esfrm_addr[2]), .S(n25), .Y(sfraddr[2])
         );
  BUFX1 U28 ( .A(n92), .Y(n21) );
  INVX3 U29 ( .A(n91), .Y(n127) );
  INVX1 U30 ( .A(n92), .Y(n25) );
  INVX2 U31 ( .A(n127), .Y(n62) );
  BUFXL U32 ( .A(n129), .Y(esfrm_rddata[0]) );
  INVX4 U33 ( .A(n90), .Y(n92) );
  NAND21X2 U34 ( .B(esfrm_oe), .A(n89), .Y(n90) );
  MUX2IX4 U35 ( .D0(esfrm_addr[6]), .D1(ramsfraddr[6]), .S(n92), .Y(n93) );
  BUFXL U36 ( .A(n89), .Y(n22) );
  BUFX8 U37 ( .A(n127), .Y(sfraddr[5]) );
  INVXL U38 ( .A(n50), .Y(n26) );
  MUX2IX2 U39 ( .D0(esfrm_addr[5]), .D1(ramsfraddr[5]), .S(n92), .Y(n91) );
  BUFXL U40 ( .A(esfrm_oe), .Y(n27) );
  INVXL U41 ( .A(n62), .Y(n28) );
  INVXL U42 ( .A(n93), .Y(n29) );
  INVX1 U43 ( .A(n6), .Y(n46) );
  INVX1 U44 ( .A(n46), .Y(n30) );
  INVX1 U45 ( .A(sfrwe_mcu51_per), .Y(n31) );
  INVX1 U46 ( .A(n31), .Y(n32) );
  NAND21XL U47 ( .B(n27), .A(n22), .Y(n112) );
  NAND21XL U48 ( .B(n111), .A(n22), .Y(sfrwe_mcu51_per) );
  INVX1 U49 ( .A(n88), .Y(n111) );
  INVXL U50 ( .A(memdatao[3]), .Y(n100) );
  INVX1 U51 ( .A(n112), .Y(n108) );
  INVX1 U52 ( .A(n80), .Y(n79) );
  INVX1 U53 ( .A(reset), .Y(n80) );
  INVXL U54 ( .A(n50), .Y(n48) );
  BUFX3 U55 ( .A(ramdatao[2]), .Y(memdatao_comb[2]) );
  BUFX3 U56 ( .A(ramdatao[4]), .Y(memdatao_comb[4]) );
  BUFX3 U57 ( .A(ramdatao[5]), .Y(memdatao_comb[5]) );
  BUFX3 U58 ( .A(ramdatao[6]), .Y(memdatao_comb[6]) );
  BUFX3 U59 ( .A(ramdatao[7]), .Y(memdatao_comb[7]) );
  INVXL U60 ( .A(n59), .Y(sfraddr[3]) );
  INVX1 U61 ( .A(n101), .Y(sfrdatao[3]) );
  INVX1 U62 ( .A(n86), .Y(ro) );
  INVX1 U63 ( .A(n103), .Y(sfrdatao[4]) );
  INVX1 U64 ( .A(n95), .Y(sfrdatao[0]) );
  INVX1 U65 ( .A(n86), .Y(dbgpo[22]) );
  INVX1 U66 ( .A(n97), .Y(sfrdatao[1]) );
  INVX1 U67 ( .A(n110), .Y(sfrdatao[7]) );
  INVX1 U68 ( .A(n105), .Y(sfrdatao[5]) );
  INVX1 U69 ( .A(n107), .Y(sfrdatao[6]) );
  INVX1 U70 ( .A(n99), .Y(sfrdatao[2]) );
  INVXL U71 ( .A(n24), .Y(n55) );
  INVXL U72 ( .A(n54), .Y(n53) );
  INVXL U73 ( .A(n54), .Y(n52) );
  INVX1 U74 ( .A(n101), .Y(n69) );
  INVX1 U75 ( .A(n99), .Y(n67) );
  INVXL U76 ( .A(n24), .Y(n56) );
  INVX1 U77 ( .A(n95), .Y(n65) );
  INVX1 U78 ( .A(n105), .Y(n73) );
  INVX1 U79 ( .A(n107), .Y(n75) );
  INVX1 U80 ( .A(n110), .Y(n77) );
  INVXL U81 ( .A(n59), .Y(n58) );
  NOR21XL U82 ( .B(N19), .A(n30), .Y(N33) );
  NOR21XL U83 ( .B(N18), .A(n30), .Y(N32) );
  NOR21XL U84 ( .B(N17), .A(n30), .Y(N31) );
  NOR21XL U85 ( .B(N16), .A(n30), .Y(N30) );
  NOR21XL U86 ( .B(N15), .A(n30), .Y(N29) );
  NOR21XL U87 ( .B(N14), .A(n30), .Y(N28) );
  NOR21XL U88 ( .B(N13), .A(n6), .Y(N27) );
  NOR21XL U89 ( .B(N12), .A(n6), .Y(N26) );
  NOR21XL U90 ( .B(N11), .A(n6), .Y(N25) );
  NOR21XL U91 ( .B(N10), .A(n6), .Y(N24) );
  NOR21XL U92 ( .B(N9), .A(n6), .Y(N23) );
  NOR21XL U93 ( .B(N8), .A(n30), .Y(N22) );
  INVX1 U94 ( .A(n87), .Y(n81) );
  INVX1 U95 ( .A(n86), .Y(n83) );
  INVX1 U96 ( .A(n87), .Y(n82) );
  INVX1 U97 ( .A(n103), .Y(n72) );
  BUFX3 U98 ( .A(ramdatao[0]), .Y(memdatao_comb[0]) );
  BUFX3 U99 ( .A(ramdatao[1]), .Y(memdatao_comb[1]) );
  BUFX3 U100 ( .A(ramdatao[3]), .Y(memdatao_comb[3]) );
  BUFX3 U101 ( .A(rxd0i), .Y(dbgpo[23]) );
  NAND21XL U102 ( .B(n112), .A(sfrwe_s), .Y(n88) );
  OR2X1 U103 ( .A(pmuintreq), .B(slp2wakeup), .Y(pmuintreq_rev) );
  INVX1 U104 ( .A(n122), .Y(n86) );
  INVX1 U105 ( .A(n95), .Y(n126) );
  INVXL U106 ( .A(memdatao[0]), .Y(n94) );
  INVX1 U107 ( .A(memdatao[4]), .Y(n102) );
  NOR21XL U108 ( .B(isr_irq), .A(r_hold_mcu), .Y(dbgpo[20]) );
  OR2X1 U109 ( .A(t0_tf1), .B(t1_tf1), .Y(dbgpo[19]) );
  OR2X1 U110 ( .A(t0_tr1), .B(t1_tr1), .Y(dbgpo[18]) );
  INVX1 U111 ( .A(memdatao[7]), .Y(n109) );
  INVX1 U112 ( .A(n97), .Y(n125) );
  INVX1 U113 ( .A(memdatao[1]), .Y(n96) );
  INVX1 U114 ( .A(n99), .Y(n124) );
  INVX1 U115 ( .A(memdatao[2]), .Y(n98) );
  INVX1 U116 ( .A(memdatao[6]), .Y(n106) );
  INVX1 U117 ( .A(n105), .Y(n123) );
  INVX1 U118 ( .A(memdatao[5]), .Y(n104) );
  INVX1 U119 ( .A(sfroe_s), .Y(n113) );
  NOR21XL U120 ( .B(N20), .A(n30), .Y(N34) );
  NOR21XL U121 ( .B(N7), .A(n6), .Y(N21) );
  NAND32X1 U122 ( .B(n11), .C(n79), .A(ien2[1]), .Y(n6) );
  INVX1 U123 ( .A(n122), .Y(n87) );
  NAND43X1 U124 ( .B(timer_1ms[8]), .C(timer_1ms[5]), .D(timer_1ms[12]), .A(
        timer_1ms[0]), .Y(n9) );
  NOR4XL U125 ( .A(n7), .B(n8), .C(n9), .D(n10), .Y(n11) );
  NAND4X1 U126 ( .A(timer_1ms[4]), .B(timer_1ms[3]), .C(timer_1ms[2]), .D(
        timer_1ms[1]), .Y(n7) );
  NAND3X1 U127 ( .A(timer_1ms[7]), .B(timer_1ms[6]), .C(timer_1ms[9]), .Y(n8)
         );
  NAND3X1 U128 ( .A(timer_1ms[11]), .B(timer_1ms[10]), .C(timer_1ms[13]), .Y(
        n10) );
  AND2X1 U129 ( .A(ien0[0]), .B(dbgpo[17]), .Y(t0_intr) );
  AO21XL U130 ( .B(n111), .C(n80), .A(esfrm_we), .Y(sfrwe) );
  INVX1 U131 ( .A(n29), .Y(n45) );
  INVXL U132 ( .A(n45), .Y(n63) );
  INVXL U133 ( .A(n62), .Y(n61) );
  MUX2AXL U134 ( .D0(esfrm_wrdata[2]), .D1(n98), .S(n108), .Y(n99) );
  MUX2AXL U135 ( .D0(esfrm_wrdata[6]), .D1(n106), .S(n108), .Y(n107) );
  MUX2AXL U136 ( .D0(esfrm_wrdata[5]), .D1(n104), .S(n108), .Y(n105) );
  MUX2AXL U137 ( .D0(esfrm_wrdata[7]), .D1(n109), .S(n108), .Y(n110) );
  MUX2AXL U138 ( .D0(esfrm_wrdata[1]), .D1(n96), .S(n108), .Y(n97) );
  MUX2AXL U139 ( .D0(esfrm_wrdata[4]), .D1(n102), .S(n108), .Y(n103) );
  MUX2AXL U140 ( .D0(esfrm_wrdata[0]), .D1(n94), .S(n108), .Y(n95) );
  MUX2AXL U141 ( .D0(esfrm_wrdata[3]), .D1(n100), .S(n108), .Y(n101) );
  NAND21XL U142 ( .B(n27), .A(n113), .Y(sfroe_mcu51_per) );
  AO21XL U143 ( .B(sfroe_s), .C(n80), .A(n27), .Y(sfroe) );
endmodule


module mcu51_a0_DW01_inc_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;

  wire   [13:2] carry;

  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module softrstctrl_a0 ( clkcpu, resetff, newinstr, srstreq, srstflag, sfrdatai, 
        sfraddr, sfrwe );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkcpu, resetff, newinstr, sfrwe;
  output srstreq, srstflag;
  wire   srst_ff0, srst_ff1, N37, N38, N39, N40, N41, net11981, n10, n11, n12,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n13, n28, n29;
  wire   [3:0] srst_count;

  SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 clk_gate_srst_count_reg ( .CLK(clkcpu), 
        .EN(N37), .ENCLK(net11981), .TE(1'b0) );
  DFFQX1 srst_ff0_reg ( .D(n26), .C(clkcpu), .Q(srst_ff0) );
  DFFQX1 srst_ff1_reg ( .D(n24), .C(clkcpu), .Q(srst_ff1) );
  DFFQX1 srst_count_reg_1_ ( .D(N39), .C(net11981), .Q(srst_count[1]) );
  DFFQX1 srst_count_reg_0_ ( .D(N38), .C(net11981), .Q(srst_count[0]) );
  DFFQX1 srst_count_reg_3_ ( .D(N41), .C(net11981), .Q(srst_count[3]) );
  DFFQX1 srst_count_reg_2_ ( .D(N40), .C(net11981), .Q(srst_count[2]) );
  DFFQX1 srst_r_reg ( .D(n27), .C(clkcpu), .Q(srstreq) );
  DFFQX1 srstflag_reg ( .D(n25), .C(clkcpu), .Q(srstflag) );
  INVX1 U3 ( .A(n14), .Y(n6) );
  NAND21X1 U4 ( .B(n1), .A(n6), .Y(n15) );
  NAND42XL U5 ( .C(sfraddr[3]), .D(n17), .A(sfraddr[0]), .B(n18), .Y(n14) );
  NAND2X1 U6 ( .A(sfraddr[2]), .B(sfraddr[1]), .Y(n17) );
  INVX1 U7 ( .A(sfrdatai[0]), .Y(n1) );
  NAND42X1 U8 ( .C(newinstr), .D(n6), .A(n4), .B(n9), .Y(n11) );
  INVX1 U9 ( .A(n12), .Y(n13) );
  NAND2X1 U10 ( .A(n4), .B(n12), .Y(N37) );
  OAI32X1 U11 ( .A(n28), .B(resetff), .C(n10), .D(n11), .E(n29), .Y(n24) );
  AOI21X1 U12 ( .B(newinstr), .C(n9), .A(n6), .Y(n10) );
  OAI33XL U13 ( .A(n16), .B(resetff), .C(n5), .D(n15), .E(resetff), .F(n29), 
        .Y(n27) );
  OAI21X1 U14 ( .B(n19), .C(n8), .A(srstreq), .Y(n16) );
  INVX1 U15 ( .A(n15), .Y(n5) );
  OAI22X1 U16 ( .A(n28), .B(n11), .C(resetff), .D(n15), .Y(n26) );
  NAND21X1 U17 ( .B(n3), .A(n12), .Y(n25) );
  AOI211X1 U18 ( .C(n6), .D(n1), .A(resetff), .B(n2), .Y(n3) );
  INVX1 U19 ( .A(srstflag), .Y(n2) );
  NAND21X1 U20 ( .B(resetff), .A(srstreq), .Y(n12) );
  AOI21BBXL U21 ( .B(srst_count[1]), .C(n12), .A(N38), .Y(n21) );
  OAI32X1 U22 ( .A(n19), .B(srst_count[3]), .C(n12), .D(n20), .E(n8), .Y(N41)
         );
  AOI21AX1 U23 ( .B(n13), .C(n7), .A(n21), .Y(n20) );
  NOR2X1 U24 ( .A(n12), .B(srst_count[0]), .Y(N38) );
  OAI21X1 U25 ( .B(n21), .C(n7), .A(n22), .Y(N40) );
  NAND4X1 U26 ( .A(srst_count[1]), .B(srst_count[0]), .C(n13), .D(n7), .Y(n22)
         );
  NAND3X1 U27 ( .A(srst_count[1]), .B(srst_count[0]), .C(srst_count[2]), .Y(
        n19) );
  INVX1 U28 ( .A(srst_count[3]), .Y(n8) );
  INVX1 U29 ( .A(resetff), .Y(n4) );
  INVX1 U30 ( .A(srstreq), .Y(n9) );
  INVX1 U31 ( .A(srst_count[2]), .Y(n7) );
  NOR2X1 U32 ( .A(n23), .B(n12), .Y(N39) );
  XNOR2XL U33 ( .A(srst_count[1]), .B(srst_count[0]), .Y(n23) );
  INVX1 U34 ( .A(srst_ff0), .Y(n28) );
  INVX1 U35 ( .A(srst_ff1), .Y(n29) );
  AND4XL U36 ( .A(sfrwe), .B(sfraddr[6]), .C(sfraddr[5]), .D(sfraddr[4]), .Y(
        n18) );
endmodule


module SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2c_a0 ( clk, rst, bclksel, scli, sdai, sclo, sdao, intack, si, sfrwe, 
        sfraddr, sfrdatai, i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  output [7:0] i2cdat_o;
  output [7:0] i2cadr_o;
  output [7:0] i2ccon_o;
  output [7:0] i2csta_o;
  input clk, rst, bclksel, scli, sdai, intack, sfrwe;
  output sclo, sdao, si;
  wire   scli_ff, N180, sdai_ff, N181, sclo_int, wait_for_setup_r, adrcomp,
         adrcompen, nedetect, ack_bit, bsd7, pedetect, N224, N225, N226, N227,
         N232, N233, N234, sclint, ack, sdaint, bsd7_tmp, write_data_r, N296,
         N297, N298, N299, N300, N301, N302, N303, N304, N332, N333, N334,
         N335, N336, N342, N343, N344, N345, N346, N347, N348, N349, N350,
         N406, N407, N408, N409, N410, N412, N413, N414, N431, N432, N433,
         N468, N469, N470, N471, N491, N492, N493, N494, N495, busfree, N510,
         N511, rst_delay, clk_count1_ov, N653, N654, N655, N656, N657,
         clk_count2_ov, N685, N686, N687, N688, N689, N690, clkint, clkint_ff,
         N700, N746, N747, N748, N749, N1022, N1023, N1024, N1025, N1026,
         N1027, N1063, N1064, N1065, sclscl, starto_en, N1124, N1125, N1126,
         net12020, net12026, net12031, net12036, net12041, net12046, net12051,
         net12056, net12061, n141, n142, n143, n144, n147, n154, n155, n157,
         n160, n161, n162, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n181, n182, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n200, n202, n203, n216, n217, n218, n219, n220,
         n222, n223, n224, n226, n227, n228, n229, n232, n234, n235, n236,
         n237, n238, n239, n240, n243, n249, n251, n252, n253, n254, n255,
         n256, n257, n259, n260, n261, n262, n263, n264, n267, n268, n269,
         n270, n271, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n288, n289, n291, n293, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n308, n309, n310, n311, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n328,
         n329, n330, n331, n332, n334, n335, n336, n337, n340, n341, n344,
         n348, n350, n351, n352, n353, n354, n355, n356, n357, n362, n364,
         n365, n366, n367, n368, n369, n372, n374, n377, n379, n381, n382,
         n383, n385, n386, n387, n388, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n454, n455, n456, n457, n458, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n483, n484, n485, n486, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n145, n146, n148,
         n149, n150, n151, n152, n153, n156, n158, n159, n163, n164, n165,
         n166, n167, n168, n169, n170, n180, n183, n195, n196, n197, n198,
         n199, n201, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n221, n225, n230, n231, n233, n241, n242, n244,
         n245, n246, n247, n248, n250, n258, n265, n266, n272, n273, n274,
         n286, n287, n290, n292, n294, n305, n306, n307, n312, n325, n326,
         n327, n333, n338, n339, n342, n343, n345, n346, n347, n349, n358,
         n359, n360, n361, n363, n370, n371, n373, n375, n376, n378, n380,
         n384, n389, n433, n453, n459, n460, n461, n462, n482, n487, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545;
  wire   [2:0] fsmmod;
  wire   [4:0] fsmsta;
  wire   [3:0] framesync;
  wire   [2:0] fsmdet;
  wire   [2:0] setup_counter_r;
  wire   [2:0] scli_ff_reg0;
  wire   [2:0] sdai_ff_reg0;
  wire   [2:0] indelay;
  wire   [2:0] fsmsync;
  wire   [1:0] bclkcnt;
  wire   [3:0] clk_count1;
  wire   [3:0] clk_count2;

  SNPS_CLOCK_GATE_HIGH_i2c_a0_0 clk_gate_i2ccon_reg ( .CLK(clk), .EN(N224), 
        .ENCLK(net12020), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_8 clk_gate_i2cdat_reg ( .CLK(clk), .EN(N296), 
        .ENCLK(net12026), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_7 clk_gate_setup_counter_r_reg ( .CLK(clk), .EN(
        N332), .ENCLK(net12031), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_6 clk_gate_i2cadr_reg ( .CLK(clk), .EN(N342), 
        .ENCLK(net12036), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_5 clk_gate_indelay_reg ( .CLK(clk), .EN(N468), 
        .ENCLK(net12041), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_4 clk_gate_framesync_reg ( .CLK(clk), .EN(N491), 
        .ENCLK(net12046), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_3 clk_gate_clk_count1_reg ( .CLK(clk), .EN(N653), 
        .ENCLK(net12051), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_2 clk_gate_clk_count2_reg ( .CLK(clk), .EN(N689), 
        .ENCLK(net12056), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_1 clk_gate_fsmsta_reg ( .CLK(clk), .EN(N1022), 
        .ENCLK(net12061), .TE(1'b0) );
  DFFQX1 i2ccon_reg_3_ ( .D(n495), .C(clk), .Q(i2ccon_o[3]) );
  DFFQX1 scli_ff_reg ( .D(N180), .C(clk), .Q(scli_ff) );
  DFFQX1 sdai_ff_reg ( .D(N181), .C(clk), .Q(sdai_ff) );
  DFFQX1 clk_count2_ov_reg ( .D(N690), .C(clk), .Q(clk_count2_ov) );
  DFFQX1 sdai_ff_reg_reg_2_ ( .D(N433), .C(clk), .Q(sdai_ff_reg0[2]) );
  DFFQX1 sdai_ff_reg_reg_0_ ( .D(N431), .C(clk), .Q(sdai_ff_reg0[0]) );
  DFFQX1 sdai_ff_reg_reg_1_ ( .D(N432), .C(clk), .Q(sdai_ff_reg0[1]) );
  DFFQX1 setup_counter_r_reg_2_ ( .D(N335), .C(net12031), .Q(
        setup_counter_r[2]) );
  DFFQX1 rst_delay_reg ( .D(n37), .C(clk), .Q(rst_delay) );
  DFFQX1 clk_count1_ov_reg ( .D(n505), .C(clk), .Q(clk_count1_ov) );
  DFFQX1 bsd7_reg ( .D(n491), .C(clk), .Q(bsd7) );
  DFFQX1 ack_bit_reg ( .D(n494), .C(net12020), .Q(ack_bit) );
  DFFQX1 clk_count2_reg_3_ ( .D(N688), .C(net12056), .Q(clk_count2[3]) );
  DFFQX1 setup_counter_r_reg_1_ ( .D(N334), .C(net12031), .Q(
        setup_counter_r[1]) );
  DFFQX1 scli_ff_reg_reg_2_ ( .D(N414), .C(clk), .Q(scli_ff_reg0[2]) );
  DFFQX1 starto_en_reg ( .D(n490), .C(clk), .Q(starto_en) );
  DFFQX1 sclscl_reg ( .D(n482), .C(clk), .Q(sclscl) );
  DFFQX1 indelay_reg_2_ ( .D(N471), .C(net12041), .Q(indelay[2]) );
  DFFQX1 clk_count2_reg_1_ ( .D(N686), .C(net12056), .Q(clk_count2[1]) );
  DFFQX1 scli_ff_reg_reg_1_ ( .D(N413), .C(clk), .Q(scli_ff_reg0[1]) );
  DFFQX1 scli_ff_reg_reg_0_ ( .D(N412), .C(clk), .Q(scli_ff_reg0[0]) );
  DFFQX1 setup_counter_r_reg_0_ ( .D(N333), .C(net12031), .Q(
        setup_counter_r[0]) );
  DFFQX1 clk_count2_reg_0_ ( .D(N685), .C(net12056), .Q(clk_count2[0]) );
  DFFQX1 write_data_r_reg ( .D(n500), .C(clk), .Q(write_data_r) );
  DFFQX1 bsd7_tmp_reg ( .D(n492), .C(clk), .Q(bsd7_tmp) );
  DFFQX1 clk_count2_reg_2_ ( .D(N687), .C(net12056), .Q(clk_count2[2]) );
  DFFQX1 indelay_reg_1_ ( .D(N470), .C(net12041), .Q(indelay[1]) );
  DFFQX1 indelay_reg_0_ ( .D(N469), .C(net12041), .Q(indelay[0]) );
  DFFQX1 clkint_ff_reg ( .D(N700), .C(clk), .Q(clkint_ff) );
  DFFQX1 bclkcnt_reg_1_ ( .D(N511), .C(clk), .Q(bclkcnt[1]) );
  DFFQX1 busfree_reg ( .D(n506), .C(clk), .Q(busfree) );
  DFFQX1 adrcompen_reg ( .D(n496), .C(clk), .Q(adrcompen) );
  DFFQX1 fsmsync_reg_1_ ( .D(N747), .C(clk), .Q(fsmsync[1]) );
  DFFQX1 clkint_reg ( .D(n504), .C(clk), .Q(clkint) );
  DFFQX1 clk_count1_reg_0_ ( .D(N654), .C(net12051), .Q(clk_count1[0]) );
  DFFQX1 pedetect_reg ( .D(n497), .C(clk), .Q(pedetect) );
  DFFQX1 fsmsync_reg_2_ ( .D(N748), .C(clk), .Q(fsmsync[2]) );
  DFFQX1 fsmsync_reg_0_ ( .D(N746), .C(clk), .Q(fsmsync[0]) );
  DFFQX1 adrcomp_reg ( .D(n501), .C(clk), .Q(adrcomp) );
  DFFQX1 sclint_reg ( .D(n499), .C(clk), .Q(sclint) );
  DFFQX1 nedetect_reg ( .D(n498), .C(clk), .Q(nedetect) );
  DFFQX1 bclkcnt_reg_0_ ( .D(N510), .C(clk), .Q(bclkcnt[0]) );
  DFFQX1 clk_count1_reg_2_ ( .D(N656), .C(net12051), .Q(clk_count1[2]) );
  DFFQX1 clk_count1_reg_3_ ( .D(N657), .C(net12051), .Q(clk_count1[3]) );
  DFFQX1 clk_count1_reg_1_ ( .D(N655), .C(net12051), .Q(clk_count1[1]) );
  DFFQX1 fsmmod_reg_1_ ( .D(N1125), .C(clk), .Q(fsmmod[1]) );
  DFFQX1 fsmmod_reg_0_ ( .D(N1124), .C(clk), .Q(fsmmod[0]) );
  DFFQX1 sdaint_reg ( .D(n507), .C(clk), .Q(sdaint) );
  DFFQX1 fsmmod_reg_2_ ( .D(N1126), .C(clk), .Q(fsmmod[2]) );
  DFFQX1 ack_reg ( .D(n493), .C(clk), .Q(ack) );
  DFFQX1 fsmdet_reg_0_ ( .D(N1063), .C(clk), .Q(fsmdet[0]) );
  DFFQX1 framesync_reg_0_ ( .D(N492), .C(net12046), .Q(framesync[0]) );
  DFFQX1 fsmdet_reg_1_ ( .D(N1064), .C(clk), .Q(fsmdet[1]) );
  DFFQX1 fsmdet_reg_2_ ( .D(N1065), .C(clk), .Q(fsmdet[2]) );
  DFFQX1 framesync_reg_3_ ( .D(N495), .C(net12046), .Q(framesync[3]) );
  DFFQX1 fsmsta_reg_0_ ( .D(N1023), .C(net12061), .Q(fsmsta[0]) );
  DFFQX1 fsmsta_reg_2_ ( .D(N1025), .C(net12061), .Q(fsmsta[2]) );
  DFFQX1 framesync_reg_1_ ( .D(N493), .C(net12046), .Q(framesync[1]) );
  DFFQX1 framesync_reg_2_ ( .D(N494), .C(net12046), .Q(framesync[2]) );
  DFFQX1 fsmsta_reg_3_ ( .D(N1026), .C(net12061), .Q(fsmsta[3]) );
  DFFQX1 fsmsta_reg_4_ ( .D(N1027), .C(net12061), .Q(fsmsta[4]) );
  DFFQX1 fsmsta_reg_1_ ( .D(N1024), .C(net12061), .Q(fsmsta[1]) );
  DFFQX1 i2csta_reg_4_ ( .D(N410), .C(clk), .Q(i2csta_o[7]) );
  DFFQX1 i2cadr_reg_6_ ( .D(N349), .C(net12036), .Q(i2cadr_o[6]) );
  DFFQX1 i2csta_reg_3_ ( .D(N409), .C(clk), .Q(i2csta_o[6]) );
  DFFQX1 i2cdat_reg_7_ ( .D(N304), .C(net12026), .Q(i2cdat_o[7]) );
  DFFQX1 i2cadr_reg_7_ ( .D(N350), .C(net12036), .Q(i2cadr_o[7]) );
  DFFQX1 i2cdat_reg_6_ ( .D(N303), .C(net12026), .Q(i2cdat_o[6]) );
  DFFQX1 i2ccon_reg_6_ ( .D(N233), .C(net12020), .Q(i2ccon_o[6]) );
  DFFQX1 i2ccon_reg_7_ ( .D(N234), .C(net12020), .Q(i2ccon_o[7]) );
  DFFQX1 i2csta_reg_2_ ( .D(N408), .C(clk), .Q(i2csta_o[5]) );
  DFFQX1 i2csta_reg_1_ ( .D(N407), .C(clk), .Q(i2csta_o[4]) );
  DFFQX1 i2cadr_reg_4_ ( .D(N347), .C(net12036), .Q(i2cadr_o[4]) );
  DFFQX1 i2cadr_reg_5_ ( .D(N348), .C(net12036), .Q(i2cadr_o[5]) );
  DFFQX1 i2ccon_reg_5_ ( .D(N232), .C(net12020), .Q(i2ccon_o[5]) );
  DFFQX1 i2cdat_reg_4_ ( .D(N301), .C(net12026), .Q(i2cdat_o[4]) );
  DFFQX1 i2cdat_reg_5_ ( .D(N302), .C(net12026), .Q(i2cdat_o[5]) );
  DFFQX1 i2ccon_reg_4_ ( .D(n503), .C(clk), .Q(i2ccon_o[4]) );
  DFFQX1 i2csta_reg_0_ ( .D(N406), .C(clk), .Q(i2csta_o[3]) );
  DFFQX1 i2cdat_reg_3_ ( .D(N300), .C(net12026), .Q(i2cdat_o[3]) );
  DFFQX1 i2cadr_reg_3_ ( .D(N346), .C(net12036), .Q(i2cadr_o[3]) );
  DFFQX1 sclo_int_reg ( .D(N749), .C(clk), .Q(sclo_int) );
  DFFQX1 wait_for_setup_r_reg ( .D(N336), .C(clk), .Q(wait_for_setup_r) );
  DFFQX1 sdao_int_reg ( .D(n502), .C(clk), .Q(sdao) );
  DFFQX1 i2cadr_reg_2_ ( .D(N345), .C(net12036), .Q(i2cadr_o[2]) );
  DFFQX1 i2cadr_reg_0_ ( .D(N343), .C(net12036), .Q(i2cadr_o[0]) );
  DFFQX1 i2ccon_reg_2_ ( .D(N227), .C(net12020), .Q(i2ccon_o[2]) );
  DFFQX1 i2cdat_reg_0_ ( .D(N297), .C(net12026), .Q(i2cdat_o[0]) );
  DFFQX1 i2cdat_reg_2_ ( .D(N299), .C(net12026), .Q(i2cdat_o[2]) );
  DFFQX1 i2ccon_reg_0_ ( .D(N225), .C(net12020), .Q(i2ccon_o[0]) );
  DFFQX1 i2cadr_reg_1_ ( .D(N344), .C(net12036), .Q(i2cadr_o[1]) );
  DFFQX1 i2cdat_reg_1_ ( .D(N298), .C(net12026), .Q(i2cdat_o[1]) );
  DFFQX1 i2ccon_reg_1_ ( .D(N226), .C(net12020), .Q(i2ccon_o[1]) );
  INVX1 U3 ( .A(1'b1), .Y(i2csta_o[0]) );
  INVX1 U5 ( .A(1'b1), .Y(i2csta_o[1]) );
  INVX1 U7 ( .A(1'b1), .Y(i2csta_o[2]) );
  GEN2XL U9 ( .D(n205), .E(n7), .C(n195), .B(n183), .A(n251), .Y(n197) );
  AO21X1 U10 ( .B(n269), .C(n520), .A(n270), .Y(n150) );
  OA21X1 U11 ( .B(n309), .C(n528), .A(n529), .Y(n7) );
  INVX1 U12 ( .A(n373), .Y(n8) );
  INVX1 U13 ( .A(n164), .Y(n9) );
  AOI221XL U14 ( .A(n365), .B(n345), .C(n366), .D(n360), .E(n513), .Y(n364) );
  GEN2XL U15 ( .D(n178), .E(n268), .C(n542), .B(i2ccon_o[4]), .A(n14), .Y(n149) );
  AOI21AX1 U16 ( .B(n286), .C(n292), .A(n139), .Y(n10) );
  INVX1 U17 ( .A(N224), .Y(n43) );
  AO21X1 U18 ( .B(sfrdatai[0]), .C(n90), .A(n38), .Y(N343) );
  AND2X1 U19 ( .A(sfrdatai[2]), .B(n90), .Y(N345) );
  AND2X1 U20 ( .A(n29), .B(n90), .Y(N347) );
  AND2X1 U21 ( .A(sfrdatai[6]), .B(n90), .Y(N349) );
  INVX1 U22 ( .A(n45), .Y(n42) );
  AND2X1 U23 ( .A(sfrdatai[0]), .B(n39), .Y(N225) );
  AND2X1 U24 ( .A(sfrdatai[2]), .B(n40), .Y(N227) );
  AND2X1 U25 ( .A(sfrdatai[6]), .B(n40), .Y(N233) );
  INVX1 U26 ( .A(n36), .Y(n34) );
  INVX1 U27 ( .A(n36), .Y(n35) );
  NAND21X1 U28 ( .B(n89), .A(n305), .Y(n139) );
  NAND32X1 U29 ( .B(n36), .C(n28), .A(n230), .Y(n45) );
  NAND21X1 U30 ( .B(n36), .A(n247), .Y(N224) );
  AO21X1 U31 ( .B(n89), .C(n138), .A(n292), .Y(n88) );
  INVX1 U32 ( .A(n247), .Y(n230) );
  INVX1 U33 ( .A(n157), .Y(n292) );
  INVX1 U34 ( .A(n352), .Y(n81) );
  INVX1 U35 ( .A(n350), .Y(n90) );
  AND2X1 U36 ( .A(n25), .B(n90), .Y(N344) );
  AND2X1 U37 ( .A(sfrdatai[5]), .B(n90), .Y(N348) );
  NAND2X1 U38 ( .A(n34), .B(n350), .Y(N342) );
  INVX1 U39 ( .A(n23), .Y(n22) );
  INVX1 U40 ( .A(sfraddr[0]), .Y(n21) );
  INVX1 U41 ( .A(n30), .Y(n29) );
  AND2X1 U42 ( .A(n25), .B(n40), .Y(N226) );
  AND2X1 U43 ( .A(sfrdatai[5]), .B(n40), .Y(N232) );
  INVX1 U44 ( .A(n40), .Y(n36) );
  INVX1 U45 ( .A(n274), .Y(n225) );
  INVX1 U46 ( .A(n138), .Y(n286) );
  NOR2X1 U47 ( .A(n486), .B(n488), .Y(n398) );
  INVX1 U48 ( .A(n287), .Y(n333) );
  NAND21X1 U49 ( .B(n286), .A(n274), .Y(n287) );
  NOR21XL U50 ( .B(n431), .A(n513), .Y(n458) );
  INVX1 U51 ( .A(n39), .Y(n37) );
  INVX1 U52 ( .A(n488), .Y(n522) );
  OR2X1 U53 ( .A(n407), .B(n412), .Y(n411) );
  INVX1 U54 ( .A(n39), .Y(n38) );
  OR2X1 U55 ( .A(sdai), .B(n37), .Y(N181) );
  NOR42XL U56 ( .C(n22), .D(n352), .A(sfraddr[0]), .B(sfraddr[2]), .Y(n157) );
  NOR42XL U57 ( .C(sfraddr[4]), .D(sfraddr[3]), .A(sfraddr[5]), .B(n369), .Y(
        n352) );
  INVX1 U58 ( .A(n272), .Y(n305) );
  NAND43X1 U59 ( .B(n22), .C(sfraddr[0]), .D(n81), .A(sfraddr[2]), .Y(n247) );
  NAND43X1 U60 ( .B(n21), .C(n23), .D(n81), .A(n351), .Y(n350) );
  NOR2X1 U61 ( .A(sfraddr[2]), .B(n38), .Y(n351) );
  AO21X1 U62 ( .B(sfrdatai[3]), .C(n90), .A(n38), .Y(N346) );
  AO21X1 U63 ( .B(sfrdatai[7]), .C(n90), .A(n37), .Y(N350) );
  INVX1 U64 ( .A(sfraddr[1]), .Y(n23) );
  INVX1 U65 ( .A(sfrdatai[4]), .Y(n30) );
  INVX1 U66 ( .A(sfrdatai[3]), .Y(n28) );
  INVX1 U67 ( .A(sfrdatai[7]), .Y(n33) );
  INVX1 U68 ( .A(n26), .Y(n25) );
  INVX1 U69 ( .A(sfrdatai[2]), .Y(n27) );
  INVX1 U70 ( .A(sfrdatai[0]), .Y(n24) );
  INVX1 U71 ( .A(sfrdatai[6]), .Y(n32) );
  AND2X1 U72 ( .A(sfrdatai[7]), .B(n40), .Y(N234) );
  NAND21X1 U73 ( .B(n364), .A(n87), .Y(n274) );
  NAND21X1 U74 ( .B(n371), .A(n87), .Y(n138) );
  INVX1 U75 ( .A(n181), .Y(n523) );
  INVX1 U76 ( .A(n86), .Y(n89) );
  NAND21X1 U77 ( .B(n225), .A(n307), .Y(n86) );
  INVX1 U78 ( .A(rst), .Y(n40) );
  INVX1 U79 ( .A(n127), .Y(n380) );
  OAI221X1 U80 ( .A(n435), .B(n134), .C(n535), .D(n340), .E(n454), .Y(n127) );
  AOI211X1 U81 ( .C(n433), .D(n455), .A(n515), .B(n456), .Y(n454) );
  INVX1 U82 ( .A(n457), .Y(n515) );
  INVX1 U83 ( .A(n404), .Y(n513) );
  NOR32XL U84 ( .B(n489), .C(n488), .A(n486), .Y(n402) );
  NAND4X1 U85 ( .A(n442), .B(n434), .C(n438), .D(n444), .Y(n465) );
  NAND3X1 U86 ( .A(n172), .B(n35), .C(n173), .Y(n486) );
  NAND2X1 U87 ( .A(n475), .B(n360), .Y(n457) );
  INVX1 U88 ( .A(n307), .Y(n250) );
  OAI211X1 U89 ( .C(n535), .D(n429), .A(n380), .B(n445), .Y(n439) );
  OA222X1 U90 ( .A(n434), .B(n134), .C(n446), .D(n428), .E(n536), .F(n431), 
        .Y(n445) );
  AOI21X1 U91 ( .B(n423), .C(n432), .A(n536), .Y(n456) );
  INVX1 U92 ( .A(n137), .Y(n134) );
  INVX1 U93 ( .A(n203), .Y(n511) );
  INVX1 U94 ( .A(n364), .Y(n371) );
  NOR2X1 U95 ( .A(n79), .B(n334), .Y(n488) );
  NAND2X1 U96 ( .A(n434), .B(n435), .Y(n407) );
  INVX1 U97 ( .A(n249), .Y(n529) );
  NOR2X1 U98 ( .A(n468), .B(n478), .Y(n442) );
  INVX1 U99 ( .A(rst), .Y(n39) );
  NAND2X1 U100 ( .A(n475), .B(n348), .Y(n435) );
  NAND2X1 U101 ( .A(n343), .B(n514), .Y(n431) );
  INVX1 U102 ( .A(n236), .Y(n461) );
  NAND3X1 U103 ( .A(n428), .B(n340), .C(n429), .Y(n409) );
  NAND3X1 U104 ( .A(n203), .B(n443), .C(n444), .Y(n440) );
  NAND4X1 U105 ( .A(n458), .B(n427), .C(n423), .D(n340), .Y(n473) );
  NAND2X1 U106 ( .A(n431), .B(n432), .Y(n412) );
  INVX1 U107 ( .A(n336), .Y(n540) );
  INVX1 U108 ( .A(n62), .Y(n68) );
  NAND21X1 U109 ( .B(n242), .A(n533), .Y(n62) );
  INVX1 U110 ( .A(n320), .Y(n518) );
  INVX1 U111 ( .A(n281), .Y(n145) );
  INVX1 U112 ( .A(n377), .Y(n61) );
  OR2X1 U113 ( .A(scli), .B(n37), .Y(N180) );
  NAND21X1 U114 ( .B(n157), .A(n290), .Y(n272) );
  OAI21X1 U115 ( .B(n154), .C(n376), .A(n155), .Y(n492) );
  GEN2XL U116 ( .D(n272), .E(n33), .C(n307), .B(n39), .A(n266), .Y(n155) );
  INVX1 U117 ( .A(n154), .Y(n266) );
  AO21X1 U118 ( .B(n157), .C(n265), .A(n273), .Y(n154) );
  INVX1 U119 ( .A(n273), .Y(n338) );
  OAI21X1 U120 ( .B(n160), .C(n358), .A(n161), .Y(n493) );
  OAI21BBX1 U121 ( .A(n453), .B(n162), .C(n160), .Y(n161) );
  OAI21X1 U122 ( .B(n10), .C(n521), .A(n162), .Y(n160) );
  INVX1 U123 ( .A(n248), .Y(n162) );
  NAND32X1 U124 ( .B(n307), .C(n292), .A(n290), .Y(n327) );
  NAND21X1 U125 ( .B(n17), .A(n157), .Y(n194) );
  OA21X1 U126 ( .B(n157), .C(n294), .A(n327), .Y(n147) );
  OAI211X1 U127 ( .C(n362), .D(n521), .A(n194), .B(n35), .Y(N296) );
  AND2X1 U128 ( .A(n139), .B(n138), .Y(n362) );
  OAI22X1 U129 ( .A(n17), .B(n30), .C(n10), .D(n102), .Y(N301) );
  OAI22X1 U130 ( .A(n17), .B(n28), .C(n10), .D(n103), .Y(N300) );
  OAI22X1 U131 ( .A(n17), .B(n27), .C(n10), .D(n104), .Y(N299) );
  OAI22X1 U132 ( .A(n17), .B(n26), .C(n10), .D(n105), .Y(N298) );
  OAI22X1 U133 ( .A(n17), .B(n24), .C(n358), .D(n10), .Y(N297) );
  INVX1 U134 ( .A(sfrdatai[1]), .Y(n26) );
  INVX1 U135 ( .A(sfrdatai[5]), .Y(n31) );
  OR3XL U136 ( .A(n359), .B(n85), .C(n181), .Y(n307) );
  NAND2X1 U137 ( .A(n34), .B(n182), .Y(n181) );
  INVX1 U138 ( .A(n331), .Y(n514) );
  INVX1 U139 ( .A(n184), .Y(n536) );
  NAND2X1 U140 ( .A(n483), .B(n360), .Y(n423) );
  NAND2X1 U141 ( .A(n514), .B(n479), .Y(n404) );
  INVX1 U142 ( .A(n84), .Y(n87) );
  NAND32X1 U143 ( .B(n181), .C(n85), .A(n359), .Y(n84) );
  NAND2X1 U144 ( .A(n480), .B(n514), .Y(n427) );
  OAI221X1 U145 ( .A(n536), .B(n390), .C(n184), .D(n427), .E(n423), .Y(n455)
         );
  INVX1 U146 ( .A(n125), .Y(n345) );
  OAI211X1 U147 ( .C(n545), .D(n432), .A(n380), .B(n389), .Y(n451) );
  INVX1 U148 ( .A(n452), .Y(n389) );
  OAI211X1 U149 ( .C(n349), .D(n413), .A(n447), .B(n448), .Y(N1024) );
  AOI31X1 U150 ( .A(n402), .B(n358), .C(n136), .D(n460), .Y(n448) );
  OAI31XL U151 ( .A(n449), .B(n450), .C(n451), .D(n400), .Y(n447) );
  INVX1 U152 ( .A(n414), .Y(n460) );
  NAND31X1 U153 ( .C(n174), .A(n398), .B(n179), .Y(n414) );
  NAND31X1 U154 ( .C(n330), .A(n370), .B(n366), .Y(n432) );
  NAND21X1 U155 ( .B(n36), .A(n294), .Y(n248) );
  AOI22X1 U156 ( .A(n514), .B(n475), .C(n475), .D(n481), .Y(n434) );
  OR2X1 U157 ( .A(n184), .B(n131), .Y(n137) );
  AOI21X1 U158 ( .B(n358), .C(n402), .A(n37), .Y(n417) );
  NAND4X1 U159 ( .A(n413), .B(n173), .C(n417), .D(n469), .Y(N1023) );
  INVX1 U160 ( .A(n264), .Y(n360) );
  INVX1 U161 ( .A(n294), .Y(n265) );
  NAND2X1 U162 ( .A(n348), .B(n483), .Y(n203) );
  OAI21X1 U163 ( .B(n200), .C(n536), .A(n371), .Y(n224) );
  AND2X1 U164 ( .A(n224), .B(n218), .Y(n223) );
  AOI221XL U165 ( .A(n407), .B(n408), .C(n535), .D(n409), .E(n410), .Y(n406)
         );
  INVX1 U166 ( .A(n120), .Y(n343) );
  NAND21X1 U167 ( .B(n347), .A(n366), .Y(n120) );
  NOR2X1 U168 ( .A(n341), .B(n375), .Y(n475) );
  NOR3XL U169 ( .A(n390), .B(n358), .C(n184), .Y(n430) );
  OAI221X1 U170 ( .A(n203), .B(n133), .C(n425), .D(n458), .E(n132), .Y(n450)
         );
  INVX1 U171 ( .A(n426), .Y(n133) );
  AOI32X1 U172 ( .A(n131), .B(n164), .C(n130), .D(n129), .E(n358), .Y(n132) );
  INVX1 U173 ( .A(n434), .Y(n130) );
  OAI22X1 U174 ( .A(n184), .B(n390), .C(n203), .D(n128), .Y(n129) );
  NAND41X1 U175 ( .D(n476), .A(n403), .B(n443), .C(n477), .Y(n452) );
  NAND3X1 U176 ( .A(n184), .B(n408), .C(n478), .Y(n477) );
  OAI22X1 U177 ( .A(n429), .B(n446), .C(n428), .D(n535), .Y(n476) );
  OAI21BX1 U178 ( .C(n400), .B(n436), .A(n437), .Y(N1025) );
  AO21X1 U179 ( .B(n136), .C(n358), .A(n135), .Y(n437) );
  NOR41XL U180 ( .D(n438), .A(n439), .B(n440), .C(n441), .Y(n436) );
  INVX1 U181 ( .A(n402), .Y(n135) );
  NAND2X1 U182 ( .A(n480), .B(n360), .Y(n428) );
  NAND2X1 U183 ( .A(n481), .B(n343), .Y(n429) );
  NAND2X1 U184 ( .A(n536), .B(n545), .Y(n446) );
  NAND2X1 U185 ( .A(n430), .B(n453), .Y(n443) );
  INVX1 U186 ( .A(n425), .Y(n535) );
  NAND21X1 U187 ( .B(n246), .A(n79), .Y(n258) );
  NAND32X1 U188 ( .B(n85), .C(n334), .A(n168), .Y(n198) );
  GEN2XL U189 ( .D(n165), .E(n164), .C(n329), .B(n163), .A(n159), .Y(n321) );
  AOI31X1 U190 ( .A(n330), .B(n331), .C(n332), .D(n537), .Y(n329) );
  OAI211X1 U191 ( .C(n156), .D(n153), .A(n290), .B(n152), .Y(n163) );
  NAND21X1 U192 ( .B(n181), .A(n158), .Y(n159) );
  NAND21X1 U193 ( .B(n264), .A(n343), .Y(n340) );
  NAND42X1 U194 ( .C(n402), .D(n400), .A(n414), .B(n485), .Y(N1022) );
  NOR21XL U195 ( .B(n413), .A(n486), .Y(n485) );
  AOI22BXL U196 ( .B(n427), .A(n408), .D(n137), .C(n407), .Y(n418) );
  NOR2X1 U197 ( .A(n310), .B(rst), .Y(n236) );
  NAND43X1 U198 ( .B(n165), .C(n50), .D(n181), .A(n537), .Y(N491) );
  AO21X1 U199 ( .B(n533), .C(n232), .A(n198), .Y(n56) );
  NOR4XL U200 ( .A(n486), .B(n522), .C(n521), .D(n489), .Y(n400) );
  NOR2X1 U201 ( .A(n524), .B(n395), .Y(n334) );
  AND2X1 U202 ( .A(n368), .B(n360), .Y(n478) );
  NAND3X1 U203 ( .A(n342), .B(n35), .C(n260), .Y(n336) );
  AND2X1 U204 ( .A(n368), .B(n348), .Y(n468) );
  NOR2X1 U205 ( .A(n530), .B(n309), .Y(n249) );
  INVX1 U206 ( .A(n365), .Y(n363) );
  NAND2X1 U207 ( .A(n346), .B(n365), .Y(n263) );
  INVX1 U208 ( .A(n115), .Y(n346) );
  INVX1 U209 ( .A(n124), .Y(n348) );
  NAND3X1 U210 ( .A(n79), .B(n462), .C(n282), .Y(n173) );
  AND2X1 U211 ( .A(n80), .B(n168), .Y(n496) );
  AO21X1 U212 ( .B(n39), .C(n79), .A(n78), .Y(n80) );
  INVX1 U213 ( .A(n182), .Y(n79) );
  AOI211X1 U214 ( .C(n164), .D(nedetect), .A(n181), .B(n106), .Y(n78) );
  INVX1 U215 ( .A(n341), .Y(n361) );
  NOR3XL U216 ( .A(n521), .B(n511), .C(n426), .Y(n489) );
  NOR2X1 U217 ( .A(n527), .B(n509), .Y(n282) );
  OAI221X1 U218 ( .A(n252), .B(n181), .C(n539), .D(n181), .E(n35), .Y(n506) );
  OA21X1 U219 ( .B(n253), .C(n201), .A(n199), .Y(n252) );
  INVX1 U220 ( .A(n232), .Y(n201) );
  INVX1 U221 ( .A(n198), .Y(n199) );
  INVX1 U222 ( .A(n313), .Y(n378) );
  OAI31XL U223 ( .A(n353), .B(n355), .C(n526), .D(n354), .Y(N335) );
  NAND3X1 U224 ( .A(n381), .B(n382), .C(n227), .Y(n202) );
  NOR2X1 U225 ( .A(n229), .B(n282), .Y(n381) );
  NAND2X1 U226 ( .A(n481), .B(n483), .Y(n444) );
  NAND2X1 U227 ( .A(n483), .B(n514), .Y(n438) );
  NAND2X1 U228 ( .A(n360), .B(n479), .Y(n403) );
  NAND2X1 U229 ( .A(n383), .B(n79), .Y(n172) );
  NOR2X1 U230 ( .A(n297), .B(n291), .Y(N687) );
  XNOR2XL U231 ( .A(n293), .B(n532), .Y(n297) );
  INVX1 U232 ( .A(n184), .Y(n164) );
  INVX1 U233 ( .A(n142), .Y(n508) );
  INVX1 U234 ( .A(n408), .Y(n433) );
  NAND2X1 U235 ( .A(n353), .B(n354), .Y(N336) );
  NAND2X1 U236 ( .A(n236), .B(n534), .Y(N700) );
  NAND2X1 U237 ( .A(n236), .B(n531), .Y(N689) );
  NOR2X1 U238 ( .A(n197), .B(n12), .Y(n11) );
  OAI22X1 U239 ( .A(n215), .B(n196), .C(n204), .D(n249), .Y(n12) );
  INVX1 U240 ( .A(n178), .Y(n537) );
  OA21X1 U241 ( .B(n268), .C(n542), .A(n152), .Y(n140) );
  OR2X1 U242 ( .A(n123), .B(n13), .Y(N407) );
  AOI21X1 U243 ( .B(n124), .C(n331), .A(n346), .Y(n13) );
  OA21X1 U244 ( .B(n240), .C(n205), .A(n212), .Y(n195) );
  NOR42XL U245 ( .C(n67), .D(n390), .A(n382), .B(n388), .Y(n70) );
  NAND21X1 U246 ( .B(n382), .A(n67), .Y(n63) );
  INVX1 U247 ( .A(n123), .Y(n119) );
  INVX1 U248 ( .A(n50), .Y(n158) );
  NOR2X1 U249 ( .A(n328), .B(n164), .Y(n320) );
  NAND2X1 U250 ( .A(n289), .B(n339), .Y(n281) );
  OR2X1 U251 ( .A(n228), .B(n38), .Y(n267) );
  AOI21X1 U252 ( .B(n408), .C(n9), .A(n442), .Y(n441) );
  INVX1 U253 ( .A(n76), .Y(n67) );
  NOR2X1 U254 ( .A(n528), .B(n530), .Y(n302) );
  NOR2X1 U255 ( .A(n280), .B(n283), .Y(n268) );
  OAI21X1 U256 ( .B(n323), .C(n518), .A(n523), .Y(N494) );
  XNOR2XL U257 ( .A(n322), .B(n538), .Y(n323) );
  INVX1 U258 ( .A(n328), .Y(n165) );
  INVX1 U259 ( .A(n388), .Y(n533) );
  NAND2X1 U260 ( .A(n34), .B(n313), .Y(n317) );
  AOI211X1 U261 ( .C(n114), .D(n349), .A(n113), .B(n522), .Y(n501) );
  NAND43X1 U262 ( .B(n111), .C(n126), .D(n110), .A(n109), .Y(n114) );
  OAI211X1 U263 ( .C(n112), .D(n290), .A(n168), .B(n35), .Y(n113) );
  INVX1 U264 ( .A(n200), .Y(n111) );
  INVX1 U265 ( .A(n204), .Y(n211) );
  OAI21AX1 U266 ( .B(n520), .C(n190), .A(n186), .Y(n499) );
  NOR2X1 U267 ( .A(n290), .B(n15), .Y(n14) );
  NOR2X1 U268 ( .A(n268), .B(n542), .Y(n15) );
  NAND2X1 U269 ( .A(n34), .B(n187), .Y(n186) );
  NAND2X1 U270 ( .A(n540), .B(n271), .Y(N468) );
  INVX1 U271 ( .A(n218), .Y(n244) );
  INVX1 U272 ( .A(n285), .Y(n542) );
  INVX1 U273 ( .A(n229), .Y(n241) );
  INVX1 U274 ( .A(n228), .Y(n242) );
  INVX1 U275 ( .A(n177), .Y(n74) );
  INVX1 U276 ( .A(n390), .Y(n153) );
  NOR21XL U277 ( .B(n260), .A(n271), .Y(n278) );
  NAND2X1 U278 ( .A(n388), .B(n280), .Y(n377) );
  NOR2X1 U279 ( .A(n524), .B(n525), .Y(n394) );
  NOR2X1 U280 ( .A(n339), .B(n541), .Y(n260) );
  NOR2X1 U281 ( .A(n342), .B(n339), .Y(n270) );
  INVX1 U282 ( .A(n190), .Y(n384) );
  NAND2X1 U283 ( .A(n283), .B(n285), .Y(n284) );
  INVX1 U284 ( .A(n243), .Y(n196) );
  AND2X1 U285 ( .A(sclo_int), .B(n519), .Y(sclo) );
  INVX1 U286 ( .A(wait_for_setup_r), .Y(n519) );
  NAND31X1 U287 ( .C(n36), .A(n16), .B(n258), .Y(n273) );
  NAND4X1 U288 ( .A(n521), .B(nedetect), .C(n305), .D(n250), .Y(n16) );
  AO22AXL U289 ( .A(n143), .B(n144), .C(bsd7), .D(n144), .Y(n491) );
  OAI211X1 U290 ( .C(n327), .D(n33), .A(n326), .B(n325), .Y(n143) );
  NAND3X1 U291 ( .A(n338), .B(n333), .C(n147), .Y(n144) );
  AO21X1 U292 ( .B(n520), .C(n376), .A(n294), .Y(n326) );
  MUX2X1 U293 ( .D0(n59), .D1(i2ccon_o[4]), .S(n58), .Y(n503) );
  AND2X1 U294 ( .A(n230), .B(n39), .Y(n59) );
  NOR21XL U295 ( .B(n35), .A(n57), .Y(n58) );
  MUX2X1 U296 ( .D0(n56), .D1(n29), .S(n230), .Y(n57) );
  MUX2X1 U297 ( .D0(n48), .D1(i2ccon_o[3]), .S(n47), .Y(n495) );
  AO21X1 U298 ( .B(n44), .C(n43), .A(n42), .Y(n48) );
  AOI21X1 U299 ( .B(n46), .C(n45), .A(n44), .Y(n47) );
  NOR21XL U300 ( .B(i2ccon_o[6]), .A(n41), .Y(n44) );
  AND3X1 U301 ( .A(n333), .B(n39), .C(n312), .Y(n325) );
  NAND32X1 U302 ( .B(n307), .C(n306), .A(n305), .Y(n312) );
  INVX1 U303 ( .A(i2cdat_o[7]), .Y(n306) );
  AND3X1 U304 ( .A(n258), .B(n18), .C(n88), .Y(n17) );
  OA22X1 U305 ( .A(i2ccon_o[6]), .B(n37), .C(n89), .D(n290), .Y(n18) );
  OAI22AX1 U306 ( .D(i2cdat_o[6]), .C(n10), .A(n17), .B(n33), .Y(N304) );
  OAI22AX1 U307 ( .D(i2cdat_o[5]), .C(n10), .A(n17), .B(n32), .Y(N303) );
  OAI22AX1 U308 ( .D(i2cdat_o[4]), .C(n10), .A(n17), .B(n31), .Y(N302) );
  OAI21X1 U309 ( .B(n192), .C(n193), .A(n194), .Y(n500) );
  NAND43X1 U310 ( .B(n286), .C(n250), .D(n247), .A(write_data_r), .Y(n193) );
  NAND32X1 U311 ( .B(n305), .C(n246), .A(n258), .Y(n192) );
  NAND21X1 U312 ( .B(intack), .A(n43), .Y(n46) );
  MUX2X1 U313 ( .D0(n233), .D1(ack_bit), .S(n231), .Y(n494) );
  NAND21X1 U314 ( .B(sfrdatai[2]), .A(n34), .Y(n233) );
  AOI31X1 U315 ( .A(n230), .B(i2ccon_o[3]), .C(n225), .D(n37), .Y(n231) );
  NOR21XL U316 ( .B(n366), .A(fsmsta[3]), .Y(n483) );
  NOR21XL U317 ( .B(n345), .A(fsmsta[2]), .Y(n480) );
  NAND21X1 U318 ( .B(fsmsta[3]), .A(fsmsta[4]), .Y(n341) );
  NAND21X1 U319 ( .B(n8), .A(fsmsta[0]), .Y(n331) );
  NAND21X1 U320 ( .B(fsmsta[4]), .A(fsmsta[3]), .Y(n125) );
  NAND2X1 U321 ( .A(framesync[3]), .B(n177), .Y(n184) );
  NOR3XL U322 ( .A(framesync[1]), .B(framesync[2]), .C(framesync[0]), .Y(n177)
         );
  NOR2X1 U323 ( .A(n375), .B(fsmsta[4]), .Y(n366) );
  NOR2X1 U324 ( .A(n341), .B(fsmsta[2]), .Y(n479) );
  NAND21X1 U325 ( .B(n307), .A(i2ccon_o[3]), .Y(n294) );
  NOR21XL U326 ( .B(n83), .A(n82), .Y(n359) );
  INVX1 U327 ( .A(n368), .Y(n83) );
  AND3X1 U328 ( .A(fsmsta[2]), .B(n347), .C(n367), .Y(n82) );
  OAI21X1 U329 ( .B(n517), .C(fsmsta[0]), .A(fsmsta[1]), .Y(n367) );
  OR4X1 U330 ( .A(i2cdat_o[5]), .B(i2cdat_o[4]), .C(i2cdat_o[6]), .D(n19), .Y(
        n136) );
  NAND4X1 U331 ( .A(n105), .B(n104), .C(n103), .D(n102), .Y(n19) );
  NAND21X1 U332 ( .B(n370), .A(fsmsta[1]), .Y(n264) );
  NAND21X1 U333 ( .B(fsmsta[0]), .A(n375), .Y(n365) );
  GEN2XL U334 ( .D(framesync[3]), .E(n222), .C(bsd7), .B(n223), .A(n38), .Y(
        n220) );
  NOR3XL U335 ( .A(fsmsta[3]), .B(fsmsta[4]), .C(fsmsta[2]), .Y(n368) );
  NAND21X1 U336 ( .B(n136), .A(i2cadr_o[0]), .Y(n128) );
  NAND3X1 U337 ( .A(fsmdet[0]), .B(n524), .C(fsmdet[1]), .Y(n182) );
  NAND32X1 U338 ( .B(n398), .C(n36), .A(n399), .Y(N1027) );
  AOI22X1 U339 ( .A(n400), .B(n401), .C(n402), .D(ack), .Y(n399) );
  NAND4X1 U340 ( .A(n403), .B(n404), .C(n405), .D(n406), .Y(n401) );
  AOI22X1 U341 ( .A(n363), .B(fsmsta[4]), .C(n536), .D(n411), .Y(n405) );
  INVX1 U342 ( .A(fsmsta[2]), .Y(n375) );
  NAND2X1 U343 ( .A(n368), .B(n373), .Y(n390) );
  INVX1 U344 ( .A(fsmsta[1]), .Y(n373) );
  NAND2X1 U345 ( .A(sdao), .B(n536), .Y(n425) );
  INVX1 U346 ( .A(fsmsta[4]), .Y(n517) );
  INVX1 U347 ( .A(fsmsta[0]), .Y(n370) );
  OAI22AX1 U348 ( .D(n216), .C(n217), .A(n216), .B(n545), .Y(n502) );
  NAND32X1 U349 ( .B(n244), .C(n245), .A(n226), .Y(n216) );
  AOI211X1 U350 ( .C(n219), .D(n218), .A(n220), .B(n245), .Y(n217) );
  OAI211X1 U351 ( .C(adrcomp), .D(n242), .A(i2ccon_o[6]), .B(n241), .Y(n245)
         );
  INVX1 U352 ( .A(fsmdet[2]), .Y(n524) );
  ENOX1 U353 ( .A(ack_bit), .B(n224), .C(n224), .D(n359), .Y(n219) );
  OAI211X1 U354 ( .C(ack), .D(n390), .A(n435), .B(n512), .Y(n484) );
  INVX1 U355 ( .A(n465), .Y(n512) );
  OAI211X1 U356 ( .C(n425), .D(n427), .A(n463), .B(n464), .Y(n449) );
  AOI32X1 U357 ( .A(n363), .B(fsmsta[1]), .C(n346), .D(n468), .E(n184), .Y(
        n463) );
  AOI31X1 U358 ( .A(n465), .B(n9), .C(n433), .D(n466), .Y(n464) );
  OAI21X1 U359 ( .B(n545), .C(n423), .A(n467), .Y(n466) );
  NAND2X1 U360 ( .A(n400), .B(n470), .Y(n469) );
  OAI211X1 U361 ( .C(n446), .D(n432), .A(n471), .B(n472), .Y(n470) );
  AOI33X1 U362 ( .A(n9), .B(n408), .C(n514), .D(sdaint), .E(n484), .F(n536), 
        .Y(n471) );
  AOI211X1 U363 ( .C(n473), .D(n425), .A(n452), .B(n410), .Y(n472) );
  OAI211X1 U364 ( .C(adrcomp), .D(n413), .A(n414), .B(n415), .Y(N1026) );
  AOI21AX1 U365 ( .B(n400), .C(n416), .A(n417), .Y(n415) );
  NAND4X1 U366 ( .A(n418), .B(n419), .C(n420), .D(n421), .Y(n416) );
  AOI22X1 U367 ( .A(n430), .B(sdaint), .C(n412), .D(n9), .Y(n419) );
  NAND2X1 U368 ( .A(fsmsta[3]), .B(fsmsta[1]), .Y(n330) );
  INVX1 U369 ( .A(i2cdat_o[3]), .Y(n102) );
  INVX1 U370 ( .A(i2cdat_o[2]), .Y(n103) );
  OAI211X1 U371 ( .C(n426), .D(n474), .A(n457), .B(n263), .Y(n410) );
  NAND2X1 U372 ( .A(n511), .B(ack), .Y(n474) );
  NOR21XL U373 ( .B(framesync[3]), .A(n222), .Y(n178) );
  INVX1 U374 ( .A(i2ccon_o[3]), .Y(n290) );
  NAND21X1 U375 ( .B(n202), .A(i2ccon_o[4]), .Y(n168) );
  AO21X1 U376 ( .B(n77), .C(n76), .A(n75), .Y(n413) );
  NAND32X1 U377 ( .B(i2ccon_o[3]), .C(n74), .A(n73), .Y(n77) );
  INVX1 U378 ( .A(n398), .Y(n75) );
  INVX1 U379 ( .A(framesync[3]), .Y(n73) );
  NAND21X1 U380 ( .B(rst), .A(i2ccon_o[6]), .Y(n246) );
  NAND31X1 U381 ( .C(framesync[1]), .A(n538), .B(framesync[0]), .Y(n222) );
  NAND32X1 U382 ( .B(n334), .C(n169), .A(n314), .Y(n310) );
  AOI22AXL U383 ( .A(n315), .B(n520), .D(n289), .C(n339), .Y(n314) );
  INVX1 U384 ( .A(n168), .Y(n169) );
  ENOX1 U385 ( .A(n508), .B(n539), .C(sclo_int), .D(n232), .Y(n315) );
  NAND21X1 U386 ( .B(sdaint), .A(n126), .Y(n131) );
  NAND21X1 U387 ( .B(fsmsta[0]), .A(fsmsta[1]), .Y(n124) );
  NAND21X1 U388 ( .B(n347), .A(fsmsta[4]), .Y(n115) );
  AO22AXL U389 ( .A(n355), .B(n526), .C(n188), .D(n357), .Y(n353) );
  NOR2X1 U390 ( .A(write_data_r), .B(n36), .Y(n357) );
  AOI21AX1 U391 ( .B(adrcomp), .C(adrcompen), .A(n227), .Y(n218) );
  GEN2XL U392 ( .D(n540), .E(n544), .C(N469), .B(indelay[2]), .A(n335), .Y(
        N471) );
  NOR4XL U393 ( .A(indelay[2]), .B(n544), .C(n336), .D(n543), .Y(n335) );
  INVX1 U394 ( .A(indelay[1]), .Y(n544) );
  INVX1 U395 ( .A(indelay[0]), .Y(n543) );
  GEN2XL U396 ( .D(framesync[3]), .E(n319), .C(n200), .B(n320), .A(n321), .Y(
        N495) );
  OR2X1 U397 ( .A(n322), .B(n538), .Y(n319) );
  NAND2X1 U398 ( .A(sdao), .B(n453), .Y(n408) );
  MUX2X1 U399 ( .D0(n209), .D1(n208), .S(i2ccon_o[7]), .Y(n210) );
  AND4X1 U400 ( .A(clk_count1[0]), .B(n212), .C(n205), .D(n249), .Y(n209) );
  AND3X1 U401 ( .A(n378), .B(n207), .C(n206), .Y(n208) );
  INVX1 U402 ( .A(n251), .Y(n206) );
  NAND21X1 U403 ( .B(scli_ff_reg0[1]), .A(n34), .Y(N414) );
  NOR3XL U404 ( .A(n462), .B(fsmmod[2]), .C(n527), .Y(n229) );
  NAND21X1 U405 ( .B(scli_ff_reg0[0]), .A(n34), .Y(N413) );
  NOR3XL U406 ( .A(n322), .B(framesync[3]), .C(n538), .Y(n200) );
  NOR3XL U407 ( .A(fsmmod[0]), .B(fsmmod[1]), .C(n509), .Y(n232) );
  AND3X1 U408 ( .A(n173), .B(n172), .C(n171), .Y(n41) );
  OA22X1 U409 ( .A(n174), .B(n175), .C(n349), .D(n176), .Y(n171) );
  OAI21X1 U410 ( .B(n177), .C(n178), .A(n522), .Y(n176) );
  AOI22X1 U411 ( .A(n536), .B(pedetect), .C(n179), .D(n522), .Y(n175) );
  NAND2X1 U412 ( .A(clk_count1_ov), .B(n236), .Y(n291) );
  OAI21X1 U413 ( .B(framesync[3]), .C(n177), .A(n184), .Y(n179) );
  AOI211X1 U414 ( .C(n200), .D(nedetect), .A(n36), .B(n223), .Y(n226) );
  INVX1 U415 ( .A(sdaint), .Y(n453) );
  NOR3XL U416 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(n462), .Y(n383) );
  NAND2X1 U417 ( .A(bclkcnt[1]), .B(n318), .Y(n313) );
  XOR2X1 U418 ( .A(bclksel), .B(bclkcnt[0]), .Y(n318) );
  NAND3X1 U419 ( .A(n462), .B(n509), .C(fsmmod[1]), .Y(n382) );
  NAND3X1 U420 ( .A(n536), .B(adrcomp), .C(adrcompen), .Y(n426) );
  INVX1 U421 ( .A(fsmsta[3]), .Y(n347) );
  AOI221XL U422 ( .A(n363), .B(fsmsta[3]), .C(n422), .D(n516), .E(n510), .Y(
        n421) );
  INVX1 U423 ( .A(n263), .Y(n510) );
  NOR2X1 U424 ( .A(n433), .B(n184), .Y(n422) );
  INVX1 U425 ( .A(n423), .Y(n516) );
  AND2X1 U426 ( .A(n55), .B(n54), .Y(N690) );
  AO22X1 U427 ( .A(i2ccon_o[7]), .B(n53), .C(n52), .D(n51), .Y(n55) );
  INVX1 U428 ( .A(n291), .Y(n54) );
  INVX1 U429 ( .A(n293), .Y(n51) );
  NAND3X1 U430 ( .A(fsmmod[0]), .B(n527), .C(fsmmod[2]), .Y(n142) );
  OAI32X1 U431 ( .A(n461), .B(n11), .C(n303), .D(n36), .E(n285), .Y(N656) );
  XNOR2XL U432 ( .A(n302), .B(clk_count1[2]), .Y(n303) );
  OAI32X1 U433 ( .A(n521), .B(n185), .C(n186), .D(sclint), .E(n187), .Y(n497)
         );
  INVX1 U434 ( .A(ack), .Y(n358) );
  EORX1 U435 ( .A(n424), .B(n425), .C(n426), .D(ack), .Y(n420) );
  NAND21X1 U436 ( .B(n409), .A(n427), .Y(n424) );
  INVX1 U437 ( .A(sdao), .Y(n545) );
  AOI21X1 U438 ( .B(n462), .C(fsmmod[2]), .A(n383), .Y(n227) );
  NOR2X1 U439 ( .A(fsmsta[1]), .B(fsmsta[0]), .Y(n481) );
  NAND2X1 U440 ( .A(sclint), .B(n34), .Y(n188) );
  AOI31X1 U441 ( .A(scli_ff_reg0[2]), .B(N414), .C(N413), .D(n190), .Y(n185)
         );
  INVX1 U442 ( .A(fsmmod[0]), .Y(n462) );
  OAI22X1 U443 ( .A(i2ccon_o[7]), .B(n221), .C(n243), .D(n215), .Y(n239) );
  MUX2X1 U444 ( .D0(n214), .D1(n213), .S(i2ccon_o[1]), .Y(n221) );
  NAND21X1 U445 ( .B(n240), .A(n212), .Y(n213) );
  NAND21X1 U446 ( .B(n7), .A(i2ccon_o[0]), .Y(n214) );
  OAI21X1 U447 ( .B(n534), .C(n234), .A(n235), .Y(n504) );
  OAI21X1 U448 ( .B(n461), .C(n534), .A(n234), .Y(n235) );
  NAND21X1 U449 ( .B(clk_count2_ov), .A(n236), .Y(n234) );
  INVX1 U450 ( .A(fsmmod[2]), .Y(n509) );
  INVX1 U451 ( .A(clk_count1[1]), .Y(n530) );
  OAI21X1 U452 ( .B(clk_count2[0]), .C(n461), .A(n299), .Y(N685) );
  NAND4X1 U453 ( .A(fsmsync[2]), .B(n541), .C(n339), .D(n34), .Y(n299) );
  OAI21X1 U454 ( .B(n384), .C(n188), .A(n189), .Y(n498) );
  NAND42X1 U455 ( .C(n185), .D(n190), .A(nedetect), .B(n34), .Y(n189) );
  INVX1 U456 ( .A(framesync[2]), .Y(n538) );
  OAI21X1 U457 ( .B(rst_delay), .C(n311), .A(n35), .Y(N653) );
  AND4X1 U458 ( .A(n215), .B(n180), .C(n207), .D(n313), .Y(n311) );
  INVX1 U459 ( .A(n310), .Y(n180) );
  INVX1 U460 ( .A(fsmmod[1]), .Y(n527) );
  INVX1 U461 ( .A(i2ccon_o[6]), .Y(n85) );
  INVX1 U462 ( .A(fsmdet[1]), .Y(n525) );
  NAND2X1 U463 ( .A(fsmdet[0]), .B(n525), .Y(n395) );
  OAI2B11X1 U464 ( .D(write_data_r), .C(sclint), .A(n353), .B(n35), .Y(N332)
         );
  NAND2X1 U465 ( .A(clk_count1[3]), .B(clk_count1[2]), .Y(n309) );
  NOR3XL U466 ( .A(n461), .B(n11), .C(n300), .Y(N657) );
  XNOR2XL U467 ( .A(clk_count1[3]), .B(n301), .Y(n300) );
  AND2X1 U468 ( .A(clk_count1[2]), .B(n302), .Y(n301) );
  NOR3XL U469 ( .A(n461), .B(n11), .C(n304), .Y(N655) );
  XNOR2XL U470 ( .A(clk_count1[1]), .B(clk_count1[0]), .Y(n304) );
  NOR3XL U471 ( .A(n461), .B(clk_count1[0]), .C(n11), .Y(N654) );
  OAI31XL U472 ( .A(n459), .B(n37), .C(n531), .D(n237), .Y(n505) );
  OAI211X1 U473 ( .C(n238), .D(n239), .A(n459), .B(n236), .Y(n237) );
  INVX1 U474 ( .A(rst_delay), .Y(n459) );
  AO21X1 U475 ( .B(n249), .C(n211), .A(n210), .Y(n238) );
  OAI211X1 U476 ( .C(n345), .D(n361), .A(fsmsta[1]), .B(n363), .Y(n467) );
  NAND2X1 U477 ( .A(framesync[1]), .B(framesync[0]), .Y(n322) );
  NOR2X1 U478 ( .A(n202), .B(adrcomp), .Y(n174) );
  NOR2X1 U479 ( .A(n336), .B(indelay[0]), .Y(N469) );
  OAI21AX1 U480 ( .B(framesync[0]), .C(n518), .A(n321), .Y(N492) );
  INVX1 U481 ( .A(i2cdat_o[1]), .Y(n104) );
  NOR2X1 U482 ( .A(n356), .B(n353), .Y(N334) );
  AOI21X1 U483 ( .B(setup_counter_r[1]), .C(setup_counter_r[0]), .A(n355), .Y(
        n356) );
  NOR2X1 U484 ( .A(setup_counter_r[0]), .B(n353), .Y(N333) );
  NOR2X1 U485 ( .A(n295), .B(n291), .Y(N688) );
  XNOR2XL U486 ( .A(clk_count2[3]), .B(n296), .Y(n295) );
  NOR2X1 U487 ( .A(n532), .B(n293), .Y(n296) );
  NOR2X1 U488 ( .A(n298), .B(n291), .Y(N686) );
  XNOR2XL U489 ( .A(clk_count2[1]), .B(clk_count2[0]), .Y(n298) );
  INVX1 U490 ( .A(i2cdat_o[0]), .Y(n105) );
  INVX1 U491 ( .A(n254), .Y(n482) );
  AOI32X1 U492 ( .A(n508), .B(n39), .C(n255), .D(n487), .E(sclscl), .Y(n254)
         );
  INVX1 U493 ( .A(n255), .Y(n487) );
  NAND3X1 U494 ( .A(n521), .B(n35), .C(n508), .Y(n255) );
  NAND21X1 U495 ( .B(n37), .A(i2ccon_o[3]), .Y(n123) );
  NAND21X1 U496 ( .B(i2ccon_o[3]), .A(n178), .Y(n76) );
  NAND31X1 U497 ( .C(clk_count1[2]), .A(n530), .B(n528), .Y(n308) );
  AO21X1 U498 ( .B(n520), .C(i2ccon_o[3]), .A(n334), .Y(n50) );
  NAND21X1 U499 ( .B(clkint_ff), .A(clkint), .Y(n280) );
  NAND32X1 U500 ( .B(n49), .C(n178), .A(n158), .Y(n328) );
  INVX1 U501 ( .A(nedetect), .Y(n49) );
  NAND21X1 U502 ( .B(n207), .A(i2ccon_o[7]), .Y(n204) );
  NAND42X1 U503 ( .C(n361), .D(n123), .A(n122), .B(n340), .Y(N410) );
  NAND21X1 U504 ( .B(n121), .A(fsmsta[4]), .Y(n122) );
  AOI21BBXL U505 ( .B(n150), .C(n149), .A(n267), .Y(N748) );
  NAND32X1 U506 ( .B(n334), .C(n246), .A(n387), .Y(n71) );
  NAND3X1 U507 ( .A(n164), .B(pedetect), .C(n511), .Y(n387) );
  AND4X1 U508 ( .A(n97), .B(n96), .C(n95), .D(n94), .Y(n98) );
  XOR2X1 U509 ( .A(n91), .B(i2cdat_o[4]), .Y(n97) );
  XOR2X1 U510 ( .A(n92), .B(i2cdat_o[0]), .Y(n96) );
  XOR2X1 U511 ( .A(n93), .B(i2cdat_o[6]), .Y(n95) );
  NAND2X1 U512 ( .A(clkint_ff), .B(n534), .Y(n388) );
  XOR2X1 U513 ( .A(n104), .B(i2cadr_o[2]), .Y(n94) );
  XOR2X1 U514 ( .A(i2cadr_o[3]), .B(i2cdat_o[2]), .Y(n99) );
  AO21X1 U515 ( .B(n107), .C(n128), .A(n106), .Y(n110) );
  NAND43X1 U516 ( .B(n101), .C(n100), .D(n99), .A(n98), .Y(n107) );
  XOR2X1 U517 ( .A(i2cadr_o[6]), .B(i2cdat_o[5]), .Y(n101) );
  XOR2X1 U518 ( .A(i2cadr_o[4]), .B(i2cdat_o[3]), .Y(n100) );
  AO21X1 U519 ( .B(n116), .C(n115), .A(n123), .Y(N408) );
  XOR2X1 U520 ( .A(fsmsta[2]), .B(n360), .Y(n116) );
  NOR3XL U521 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(fsmmod[0]), .Y(n228) );
  INVX1 U522 ( .A(sclint), .Y(n520) );
  AOI221XL U523 ( .A(n108), .B(ack), .C(n203), .D(n202), .E(n49), .Y(n109) );
  INVX1 U524 ( .A(n136), .Y(n108) );
  INVX1 U525 ( .A(fsmsync[1]), .Y(n339) );
  NOR2X1 U526 ( .A(n308), .B(clk_count1[3]), .Y(n251) );
  NAND5XL U527 ( .A(starto_en), .B(i2ccon_o[5]), .C(n290), .D(n453), .E(n68), 
        .Y(n64) );
  NAND3X1 U528 ( .A(fsmsync[0]), .B(n339), .C(fsmsync[2]), .Y(n285) );
  AND3X1 U529 ( .A(starto_en), .B(n290), .C(n68), .Y(n69) );
  INVX1 U530 ( .A(n170), .Y(n207) );
  NAND21X1 U531 ( .B(n212), .A(i2ccon_o[1]), .Y(n170) );
  INVX1 U532 ( .A(pedetect), .Y(n521) );
  NOR2X1 U533 ( .A(fsmsync[2]), .B(fsmsync[0]), .Y(n289) );
  INVX1 U534 ( .A(i2ccon_o[0]), .Y(n212) );
  AOI21AX1 U535 ( .B(clk_count1[3]), .C(n302), .A(n309), .Y(n240) );
  INVX1 U536 ( .A(clkint), .Y(n534) );
  AOI221XL U537 ( .A(n361), .B(n360), .C(fsmsta[4]), .D(n363), .E(n511), .Y(
        n112) );
  INVX1 U538 ( .A(clk_count1[0]), .Y(n528) );
  NAND2X1 U539 ( .A(n289), .B(fsmsync[1]), .Y(n283) );
  OAI21X1 U540 ( .B(n259), .C(n167), .A(n166), .Y(N749) );
  AOI21X1 U541 ( .B(n541), .C(n339), .A(n260), .Y(n259) );
  INVX1 U542 ( .A(n246), .Y(n166) );
  AOI211X1 U543 ( .C(n346), .D(fsmsta[1]), .A(n261), .B(n290), .Y(n167) );
  OAI21X1 U544 ( .B(n256), .C(n453), .A(n257), .Y(n507) );
  NOR3XL U545 ( .A(sdai_ff_reg0[0]), .B(sdai_ff_reg0[2]), .C(sdai_ff_reg0[1]), 
        .Y(n256) );
  AOI31X1 U546 ( .A(sdai_ff_reg0[1]), .B(sdai_ff_reg0[0]), .C(sdai_ff_reg0[2]), 
        .D(n37), .Y(n257) );
  OAI21X1 U547 ( .B(n324), .C(n518), .A(n523), .Y(N493) );
  XNOR2XL U548 ( .A(framesync[1]), .B(framesync[0]), .Y(n324) );
  NOR4XL U549 ( .A(n279), .B(n520), .C(n280), .D(n281), .Y(n277) );
  AOI221XL U550 ( .A(fsmmod[0]), .B(n527), .C(n462), .D(n509), .E(n282), .Y(
        n279) );
  NAND4X1 U551 ( .A(scli_ff_reg0[1]), .B(scli_ff_reg0[0]), .C(n191), .D(n384), 
        .Y(n187) );
  NOR21XL U552 ( .B(scli_ff_reg0[2]), .A(n38), .Y(n191) );
  AOI21X1 U553 ( .B(fsmsta[2]), .C(n370), .A(n517), .Y(n332) );
  INVX1 U554 ( .A(i2ccon_o[1]), .Y(n205) );
  AOI31X1 U555 ( .A(n275), .B(n276), .C(n151), .D(n267), .Y(N747) );
  NAND21X1 U556 ( .B(n283), .A(n280), .Y(n275) );
  AOI32X1 U557 ( .A(fsmsync[0]), .B(n339), .C(n342), .D(n284), .E(n290), .Y(
        n151) );
  NOR3XL U558 ( .A(n277), .B(n278), .C(n270), .Y(n276) );
  NOR3XL U559 ( .A(n141), .B(n539), .C(n520), .Y(n490) );
  OAI211X1 U560 ( .C(n533), .D(starto_en), .A(n142), .B(n35), .Y(n141) );
  AOI21X1 U561 ( .B(n148), .C(n146), .A(n267), .Y(N746) );
  AOI211X1 U562 ( .C(n268), .D(n537), .A(n278), .B(n288), .Y(n146) );
  AOI211X1 U563 ( .C(n520), .D(n145), .A(n14), .B(n140), .Y(n148) );
  AOI21AX1 U564 ( .B(sdaint), .C(n541), .A(n270), .Y(n288) );
  NAND3X1 U565 ( .A(n39), .B(n520), .C(write_data_r), .Y(n354) );
  OAI211X1 U566 ( .C(fsmsta[4]), .D(n262), .A(n263), .B(n520), .Y(n261) );
  AOI21X1 U567 ( .B(n264), .C(n375), .A(n347), .Y(n262) );
  INVX1 U568 ( .A(i2ccon_o[2]), .Y(n126) );
  OAI211X1 U569 ( .C(n344), .D(n125), .A(n119), .B(n118), .Y(N409) );
  MUX2X1 U570 ( .D0(n117), .D1(n121), .S(fsmsta[3]), .Y(n118) );
  INVX1 U571 ( .A(n344), .Y(n117) );
  NOR2X1 U572 ( .A(n264), .B(n375), .Y(n344) );
  OAI211X1 U573 ( .C(fsmsta[0]), .D(n346), .A(n119), .B(n121), .Y(N406) );
  AOI21BX1 U574 ( .C(n396), .B(n397), .A(n188), .Y(N1063) );
  NAND2X1 U575 ( .A(n394), .B(n453), .Y(n397) );
  OAI32X1 U576 ( .A(n394), .B(fsmdet[0]), .C(n453), .D(n395), .E(fsmdet[2]), 
        .Y(n396) );
  AOI31X1 U577 ( .A(n372), .B(n66), .C(n65), .D(n71), .Y(N1126) );
  NAND32X1 U578 ( .B(n61), .C(n241), .A(sclint), .Y(n66) );
  AOI222XL U579 ( .A(n508), .B(n374), .C(n282), .D(n49), .E(n232), .F(n253), 
        .Y(n372) );
  MUX2X1 U580 ( .D0(n64), .D1(n63), .S(i2ccon_o[4]), .Y(n65) );
  AOI31X1 U581 ( .A(n381), .B(n379), .C(n60), .D(n71), .Y(N1125) );
  NAND2X1 U582 ( .A(n383), .B(nedetect), .Y(n379) );
  AO21X1 U583 ( .B(n67), .C(i2ccon_o[4]), .A(n382), .Y(n60) );
  AOI31X1 U584 ( .A(n385), .B(n386), .C(n72), .D(n71), .Y(N1124) );
  OAI21BBX1 U585 ( .A(n377), .B(sclint), .C(n229), .Y(n385) );
  AOI22X1 U586 ( .A(n383), .B(n49), .C(n508), .D(n374), .Y(n386) );
  OAI211X1 U587 ( .C(n70), .D(n69), .A(i2ccon_o[5]), .B(n152), .Y(n72) );
  NOR2X1 U588 ( .A(n337), .B(n336), .Y(N470) );
  XNOR2XL U589 ( .A(indelay[1]), .B(indelay[0]), .Y(n337) );
  NOR2X1 U590 ( .A(n316), .B(n317), .Y(N511) );
  XNOR2XL U591 ( .A(bclkcnt[1]), .B(bclkcnt[0]), .Y(n316) );
  NOR2X1 U592 ( .A(bclkcnt[0]), .B(n317), .Y(N510) );
  NOR2X1 U593 ( .A(n392), .B(n188), .Y(N1064) );
  AOI221XL U594 ( .A(fsmdet[2]), .B(fsmdet[0]), .C(n393), .D(n453), .E(n394), 
        .Y(n392) );
  OAI21X1 U595 ( .B(fsmdet[2]), .C(fsmdet[0]), .A(n395), .Y(n393) );
  NOR2X1 U596 ( .A(n391), .B(n188), .Y(N1065) );
  AOI221XL U597 ( .A(sdaint), .B(fsmdet[1]), .C(fsmdet[2]), .D(n525), .E(n79), 
        .Y(n391) );
  INVX1 U598 ( .A(busfree), .Y(n539) );
  INVX1 U599 ( .A(i2cadr_o[7]), .Y(n93) );
  INVX1 U600 ( .A(i2cadr_o[1]), .Y(n92) );
  INVX1 U601 ( .A(i2cadr_o[5]), .Y(n91) );
  NOR32XL U602 ( .B(indelay[1]), .C(indelay[2]), .A(indelay[0]), .Y(n271) );
  OAI31XL U603 ( .A(scli_ff_reg0[0]), .B(scli_ff_reg0[2]), .C(scli_ff_reg0[1]), 
        .D(n519), .Y(n190) );
  NAND21X1 U604 ( .B(fsmsta[1]), .A(n363), .Y(n121) );
  NAND21X1 U605 ( .B(i2ccon_o[7]), .A(n207), .Y(n215) );
  AO21X1 U606 ( .B(clk_count2[0]), .C(i2ccon_o[0]), .A(i2ccon_o[1]), .Y(n53)
         );
  AO21X1 U607 ( .B(clk_count2[3]), .C(clk_count2[2]), .A(n183), .Y(n52) );
  NAND2X1 U608 ( .A(clk_count2[1]), .B(clk_count2[0]), .Y(n293) );
  NAND2X1 U609 ( .A(clk_count1[3]), .B(n308), .Y(n243) );
  INVX1 U610 ( .A(fsmsync[0]), .Y(n541) );
  INVX1 U611 ( .A(fsmsync[2]), .Y(n342) );
  INVX1 U612 ( .A(i2ccon_o[4]), .Y(n152) );
  INVX1 U613 ( .A(i2ccon_o[7]), .Y(n183) );
  NOR2X1 U614 ( .A(setup_counter_r[1]), .B(setup_counter_r[0]), .Y(n355) );
  INVX1 U615 ( .A(adrcomp), .Y(n349) );
  ENOX1 U616 ( .A(fsmsync[0]), .B(n342), .C(n271), .D(n260), .Y(n269) );
  INVX1 U617 ( .A(clk_count2[2]), .Y(n532) );
  NAND2X1 U618 ( .A(n533), .B(sclint), .Y(n253) );
  NAND2X1 U619 ( .A(sclscl), .B(pedetect), .Y(n374) );
  INVX1 U620 ( .A(adrcompen), .Y(n106) );
  INVX1 U621 ( .A(i2ccon_o[5]), .Y(n156) );
  INVX1 U622 ( .A(bsd7_tmp), .Y(n376) );
  OR2X1 U623 ( .A(sdai_ff_reg0[1]), .B(n38), .Y(N433) );
  OR2X1 U624 ( .A(sdai_ff_reg0[0]), .B(n38), .Y(N432) );
  OR2X1 U625 ( .A(sdai_ff), .B(n38), .Y(N431) );
  OR2X1 U626 ( .A(scli_ff), .B(n38), .Y(N412) );
  INVX1 U627 ( .A(clk_count1_ov), .Y(n531) );
  INVX1 U628 ( .A(setup_counter_r[2]), .Y(n526) );
  BUFX3 U629 ( .A(i2ccon_o[3]), .Y(si) );
  NAND2X1 U630 ( .A(sfrwe), .B(sfraddr[6]), .Y(n369) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module extint_a0 ( clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, 
        int2ff, iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, 
        int6ff, iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, 
        ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7, 
        iex8, iex9, iex10, iex11, iex12, sfraddr, sfrdatai, sfrwe );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, int2ff,
         iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, int6ff,
         iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, sfrwe;
  output ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12;
  wire   int0_ff1, int0_fall, int0_clr, N23, int1_ff1, int1_fall, int1_clr,
         N51, int2_ff1, iex2_set, N71, int3_ff1, iex3_set, N90, iex4_set,
         int4_ff1, iex5_set, int5_ff1, iex6_set, int6_ff1, iex7_set, int7_ff1,
         iex8_set, int8_ff1, iex9_set, int9_ff1, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n56, n57, n58, n61, n64, n67, n74, n84, n91, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n54, n55, n59,
         n60, n62, n63, n65, n66, n68, n69, n70, n71, n72, n73, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n92, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133;

  DFFQX1 int4_ff1_reg ( .D(n86), .C(clkper), .Q(int4_ff1) );
  DFFQX1 int5_ff1_reg ( .D(n80), .C(clkper), .Q(int5_ff1) );
  DFFQX1 int6_ff1_reg ( .D(n83), .C(clkper), .Q(int6_ff1) );
  DFFQX1 int7_ff1_reg ( .D(n85), .C(clkper), .Q(int7_ff1) );
  DFFQX1 int8_ff1_reg ( .D(n131), .C(clkper), .Q(int8_ff1) );
  DFFQX1 int9_ff1_reg ( .D(n79), .C(clkper), .Q(int9_ff1) );
  DFFQX1 iex2_set_reg ( .D(n110), .C(clkper), .Q(iex2_set) );
  DFFQX1 iex3_set_reg ( .D(n107), .C(clkper), .Q(iex3_set) );
  DFFQX1 iex6_set_reg ( .D(n101), .C(clkper), .Q(iex6_set) );
  DFFQX1 iex7_set_reg ( .D(n99), .C(clkper), .Q(iex7_set) );
  DFFQX1 iex8_set_reg ( .D(n97), .C(clkper), .Q(iex8_set) );
  DFFQX1 iex9_set_reg ( .D(n95), .C(clkper), .Q(iex9_set) );
  DFFQX1 int2_ff1_reg ( .D(N71), .C(clkper), .Q(int2_ff1) );
  DFFQX1 int3_ff1_reg ( .D(N90), .C(clkper), .Q(int3_ff1) );
  DFFQX1 iex4_set_reg ( .D(n105), .C(clkper), .Q(iex4_set) );
  DFFQX1 iex5_set_reg ( .D(n103), .C(clkper), .Q(iex5_set) );
  DFFQX1 int0_fall_reg ( .D(n116), .C(clkper), .Q(int0_fall) );
  DFFQX1 int1_fall_reg ( .D(n112), .C(clkper), .Q(int1_fall) );
  DFFQX1 int0_clr_reg ( .D(n118), .C(clkper), .Q(int0_clr) );
  DFFQX1 int1_clr_reg ( .D(n114), .C(clkper), .Q(int1_clr) );
  DFFQX1 int0_ff1_reg ( .D(N23), .C(clkper), .Q(int0_ff1) );
  DFFQX1 int1_ff1_reg ( .D(N51), .C(clkper), .Q(int1_ff1) );
  DFFQX1 i3fr_s_reg ( .D(n108), .C(clkper), .Q(i3fr) );
  DFFQX1 i2fr_s_reg ( .D(n81), .C(clkper), .Q(i2fr) );
  DFFQX1 iex5_s_reg ( .D(n102), .C(clkper), .Q(iex5) );
  DFFQX1 iex6_s_reg ( .D(n100), .C(clkper), .Q(iex6) );
  DFFQX1 iex8_s_reg ( .D(n96), .C(clkper), .Q(iex8) );
  DFFQX1 iex9_s_reg ( .D(n94), .C(clkper), .Q(iex9) );
  DFFQX1 iex4_s_reg ( .D(n104), .C(clkper), .Q(iex4) );
  DFFQX1 ie1_s_reg ( .D(n111), .C(clkper), .Q(ie1) );
  DFFQX1 iex7_s_reg ( .D(n98), .C(clkper), .Q(iex7) );
  DFFQX1 it1_s_reg ( .D(n113), .C(clkper), .Q(it1) );
  DFFQX1 it0_s_reg ( .D(n117), .C(clkper), .Q(it0) );
  DFFQX1 iex3_s_reg ( .D(n106), .C(clkper), .Q(iex3) );
  DFFQX1 ie0_s_reg ( .D(n115), .C(clkper), .Q(ie0) );
  DFFQX1 iex2_s_reg ( .D(n109), .C(clkper), .Q(iex2) );
  INVX1 U3 ( .A(1'b1), .Y(iex12) );
  INVX1 U5 ( .A(1'b1), .Y(iex11) );
  INVX1 U7 ( .A(1'b1), .Y(iex10) );
  NOR2X1 U9 ( .A(newinstr), .B(n19), .Y(n47) );
  INVX1 U10 ( .A(n47), .Y(n7) );
  INVX1 U11 ( .A(n47), .Y(n8) );
  NAND32XL U12 ( .B(sfraddr[3]), .C(n12), .A(n74), .Y(n57) );
  AND2XL U13 ( .A(n74), .B(sfraddr[3]), .Y(n10) );
  AND4XL U14 ( .A(sfraddr[3]), .B(sfraddr[4]), .C(sfraddr[5]), .D(sfrwe), .Y(
        n51) );
  INVX1 U15 ( .A(n62), .Y(n24) );
  INVX1 U16 ( .A(n56), .Y(n59) );
  INVX1 U17 ( .A(n12), .Y(n11) );
  INVX1 U18 ( .A(rst), .Y(n16) );
  INVX1 U19 ( .A(n19), .Y(n17) );
  NAND21X1 U20 ( .B(n18), .A(n57), .Y(n62) );
  AOI21X1 U21 ( .B(n10), .C(n11), .A(n18), .Y(n9) );
  NOR2X1 U22 ( .A(rst), .B(n78), .Y(n56) );
  INVX1 U23 ( .A(n57), .Y(n78) );
  INVX1 U24 ( .A(n66), .Y(n75) );
  NAND21X1 U25 ( .B(n11), .A(n10), .Y(n66) );
  INVX1 U26 ( .A(n46), .Y(n82) );
  NAND21X1 U27 ( .B(n57), .A(n16), .Y(n63) );
  INVX1 U28 ( .A(n20), .Y(n18) );
  INVX1 U29 ( .A(n20), .Y(n19) );
  NOR42XL U30 ( .C(sfrwe), .D(n93), .A(sfraddr[0]), .B(sfraddr[1]), .Y(n74) );
  NOR3XL U31 ( .A(sfraddr[2]), .B(sfraddr[5]), .C(sfraddr[4]), .Y(n93) );
  NAND2X1 U32 ( .A(n51), .B(n52), .Y(n46) );
  NOR43XL U33 ( .B(sfraddr[2]), .C(sfraddr[0]), .D(sfraddr[1]), .A(n11), .Y(
        n52) );
  INVX1 U34 ( .A(sfrdatai[3]), .Y(n15) );
  INVX1 U35 ( .A(sfrdatai[1]), .Y(n13) );
  INVX1 U36 ( .A(n58), .Y(n85) );
  NAND2X1 U37 ( .A(n16), .B(n41), .Y(N71) );
  INVX1 U38 ( .A(int0ack), .Y(n127) );
  INVX1 U39 ( .A(int1ack), .Y(n128) );
  INVX1 U40 ( .A(rst), .Y(n20) );
  NAND2X1 U41 ( .A(n17), .B(n87), .Y(N90) );
  INVX1 U42 ( .A(n53), .Y(n131) );
  INVX1 U43 ( .A(n64), .Y(n80) );
  INVX1 U44 ( .A(n48), .Y(n79) );
  INVX1 U45 ( .A(n67), .Y(n86) );
  OAI32X1 U46 ( .A(n89), .B(int0ack), .C(n7), .D(n18), .E(n91), .Y(n116) );
  OAI32X1 U47 ( .A(n92), .B(int1ack), .C(n7), .D(n18), .E(n84), .Y(n112) );
  OAI22X1 U48 ( .A(n19), .B(n128), .C(n8), .D(n90), .Y(n114) );
  OAI22X1 U49 ( .A(n19), .B(n127), .C(n8), .D(n88), .Y(n118) );
  NAND2X1 U50 ( .A(int7ff), .B(n16), .Y(n58) );
  INVX1 U51 ( .A(int2ff), .Y(n41) );
  INVX1 U52 ( .A(int3ff), .Y(n87) );
  INVX1 U53 ( .A(n61), .Y(n83) );
  NAND2X1 U54 ( .A(n84), .B(n92), .Y(n69) );
  NAND2X1 U55 ( .A(n91), .B(n89), .Y(n73) );
  NAND2X1 U56 ( .A(int8ff), .B(n16), .Y(n53) );
  NOR2X1 U57 ( .A(rst), .B(n133), .Y(N51) );
  NOR2X1 U58 ( .A(n19), .B(n132), .Y(N23) );
  NAND2X1 U59 ( .A(int5ff), .B(n16), .Y(n64) );
  OAI32X1 U60 ( .A(n122), .B(iex5ack), .C(n7), .D(int5_ff1), .E(n64), .Y(n103)
         );
  INVX1 U61 ( .A(iex5_set), .Y(n122) );
  NAND2X1 U62 ( .A(int9ff), .B(n16), .Y(n48) );
  NAND2X1 U63 ( .A(int4ff), .B(n16), .Y(n67) );
  OAI32X1 U64 ( .A(n8), .B(iex9ack), .C(n126), .D(int9_ff1), .E(n48), .Y(n95)
         );
  INVX1 U65 ( .A(iex9_set), .Y(n126) );
  OAI32X1 U66 ( .A(n121), .B(iex4ack), .C(n7), .D(int4_ff1), .E(n67), .Y(n105)
         );
  INVX1 U67 ( .A(iex4_set), .Y(n121) );
  NOR21XL U68 ( .B(n17), .A(n71), .Y(n111) );
  MUX3X1 U69 ( .D0(int1ff), .D1(n70), .D2(n15), .S0(it1), .S1(n75), .Y(n71) );
  AOI33X1 U70 ( .A(n90), .B(n128), .C(n69), .D(ie1), .E(n90), .F(n128), .Y(n70) );
  NOR21XL U71 ( .B(n17), .A(n77), .Y(n115) );
  MUX3X1 U72 ( .D0(int0ff), .D1(n76), .D2(n13), .S0(it0), .S1(n75), .Y(n77) );
  AOI33X1 U73 ( .A(n88), .B(n127), .C(n73), .D(ie0), .E(n88), .F(n127), .Y(n76) );
  NAND21X1 U74 ( .B(n27), .A(n26), .Y(n100) );
  NOR21XL U75 ( .B(sfrdatai[5]), .A(n63), .Y(n27) );
  NAND21X1 U76 ( .B(iex6ack), .A(n25), .Y(n26) );
  AO22X1 U77 ( .A(n24), .B(iex6_set), .C(n56), .D(iex6), .Y(n25) );
  AND2X1 U78 ( .A(n68), .B(n17), .Y(n113) );
  MUX2X1 U79 ( .D0(it1), .D1(sfrdatai[2]), .S(n75), .Y(n68) );
  AND2X1 U80 ( .A(n72), .B(n17), .Y(n117) );
  MUX2X1 U81 ( .D0(it0), .D1(sfrdatai[0]), .S(n75), .Y(n72) );
  MUX2X1 U82 ( .D0(n33), .D1(i3fr), .S(n9), .Y(n108) );
  AND2X1 U83 ( .A(sfrdatai[6]), .B(n17), .Y(n33) );
  MUX2X1 U84 ( .D0(n40), .D1(i2fr), .S(n9), .Y(n81) );
  AND2X1 U85 ( .A(sfrdatai[5]), .B(n17), .Y(n40) );
  NAND21X1 U86 ( .B(n23), .A(n22), .Y(n98) );
  NOR21XL U87 ( .B(sfrdatai[0]), .A(n63), .Y(n23) );
  NAND21X1 U88 ( .B(iex7ack), .A(n21), .Y(n22) );
  AO22X1 U89 ( .A(n24), .B(iex7_set), .C(n56), .D(iex7), .Y(n21) );
  NAND21X1 U90 ( .B(n30), .A(n29), .Y(n102) );
  NOR21XL U91 ( .B(sfrdatai[4]), .A(n63), .Y(n30) );
  NAND21X1 U92 ( .B(iex5ack), .A(n28), .Y(n29) );
  ENOX1 U93 ( .A(n62), .B(n122), .C(iex5), .D(n56), .Y(n28) );
  OAI22X1 U94 ( .A(iex3ack), .B(n39), .C(n63), .D(n14), .Y(n106) );
  INVX1 U95 ( .A(sfrdatai[2]), .Y(n14) );
  OA22X1 U96 ( .A(n62), .B(n38), .C(n59), .D(n37), .Y(n39) );
  INVX1 U97 ( .A(iex3), .Y(n37) );
  OAI22X1 U98 ( .A(iex4ack), .B(n32), .C(n15), .D(n63), .Y(n104) );
  OA22X1 U99 ( .A(n62), .B(n121), .C(n59), .D(n31), .Y(n32) );
  INVX1 U100 ( .A(iex4), .Y(n31) );
  OAI22X1 U101 ( .A(iex2ack), .B(n65), .C(n13), .D(n63), .Y(n109) );
  OA22X1 U102 ( .A(n62), .B(n60), .C(n59), .D(n55), .Y(n65) );
  INVX1 U103 ( .A(iex2), .Y(n55) );
  OAI21X1 U104 ( .B(n19), .C(n44), .A(n45), .Y(n94) );
  NAND4X1 U105 ( .A(iex9), .B(n46), .C(n129), .D(n16), .Y(n45) );
  AOI32X1 U106 ( .A(n46), .B(n129), .C(iex9_set), .D(sfrdatai[1]), .E(n82), 
        .Y(n44) );
  INVX1 U107 ( .A(iex9ack), .Y(n129) );
  OAI21X1 U108 ( .B(n19), .C(n49), .A(n50), .Y(n96) );
  NAND4X1 U109 ( .A(iex8), .B(n46), .C(n130), .D(n16), .Y(n50) );
  AOI32X1 U110 ( .A(n46), .B(n130), .C(iex8_set), .D(sfrdatai[0]), .E(n82), 
        .Y(n49) );
  INVX1 U111 ( .A(iex8ack), .Y(n130) );
  OAI32X1 U112 ( .A(iex3ack), .B(n8), .C(n38), .D(n19), .E(n36), .Y(n107) );
  MUX2X1 U113 ( .D0(n35), .D1(n34), .S(i3fr), .Y(n36) );
  NAND21X1 U114 ( .B(n87), .A(n120), .Y(n34) );
  NAND21X1 U115 ( .B(int3ff), .A(int3_ff1), .Y(n35) );
  OAI32X1 U116 ( .A(n125), .B(iex8ack), .C(n7), .D(int8_ff1), .E(n53), .Y(n97)
         );
  INVX1 U117 ( .A(iex8_set), .Y(n125) );
  OAI32X1 U118 ( .A(n124), .B(iex7ack), .C(n7), .D(int7_ff1), .E(n58), .Y(n99)
         );
  INVX1 U119 ( .A(iex7_set), .Y(n124) );
  OAI32X1 U120 ( .A(n123), .B(iex6ack), .C(n8), .D(int6_ff1), .E(n61), .Y(n101) );
  INVX1 U121 ( .A(iex6_set), .Y(n123) );
  OAI32X1 U122 ( .A(n8), .B(iex2ack), .C(n60), .D(n18), .E(n54), .Y(n110) );
  MUX2X1 U123 ( .D0(n43), .D1(n42), .S(i2fr), .Y(n54) );
  NAND21X1 U124 ( .B(int2ff), .A(int2_ff1), .Y(n43) );
  NAND21X1 U125 ( .B(n41), .A(n119), .Y(n42) );
  NAND2X1 U126 ( .A(int6ff), .B(n16), .Y(n61) );
  NAND2X1 U127 ( .A(int1_ff1), .B(n133), .Y(n84) );
  NAND2X1 U128 ( .A(int0_ff1), .B(n132), .Y(n91) );
  INVX1 U129 ( .A(int0ff), .Y(n132) );
  INVX1 U130 ( .A(int1ff), .Y(n133) );
  INVX1 U131 ( .A(int1_clr), .Y(n90) );
  INVX1 U132 ( .A(int0_clr), .Y(n88) );
  INVX1 U133 ( .A(int1_fall), .Y(n92) );
  INVX1 U134 ( .A(int0_fall), .Y(n89) );
  INVX1 U135 ( .A(int3_ff1), .Y(n120) );
  INVX1 U136 ( .A(int2_ff1), .Y(n119) );
  INVX1 U137 ( .A(iex3_set), .Y(n38) );
  INVX1 U138 ( .A(iex2_set), .Y(n60) );
  INVX1 U139 ( .A(sfraddr[6]), .Y(n12) );
endmodule


module isr_a0 ( clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, 
        t0ff, int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff, 
        int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b, 
        int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, int_vect_ab, irq, intvect, int_ack_03, int_ack_0b, 
        int_ack_13, int_ack_1b, int_ack_43, int_ack_4b, int_ack_53, int_ack_5b, 
        int_ack_63, int_ack_6b, int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, 
        int_ack_ab, is_reg, ip0, ip1, ien0, ien1, ien2, isr_tm, sfraddr, 
        sfrdatai, sfrwe );
  output [4:0] intvect;
  output [3:0] is_reg;
  output [5:0] ip0;
  output [5:0] ip1;
  output [7:0] ien0;
  output [5:0] ien1;
  output [5:0] ien2;
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, t0ff,
         int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff,
         int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b,
         int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b,
         int_vect_a3, int_vect_ab, sfrwe;
  output irq, int_ack_03, int_ack_0b, int_ack_13, int_ack_1b, int_ack_43,
         int_ack_4b, int_ack_53, int_ack_5b, int_ack_63, int_ack_6b,
         int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, int_ack_ab, isr_tm;
  wire   N38, N39, N40, N41, N42, N43, N44, N45, N49, N50, N51, N52, N53, N54,
         N55, N58, N59, N60, N61, N62, N63, N64, N67, N68, N69, N70, N71, N72,
         N73, N76, N77, N78, N79, N80, N81, N82, irq_r, N200, N207, N208, N209,
         N210, N211, N212, net12078, net12084, net12089, net12094, net12099,
         net12104, n42, n43, n47, n48, n49, n50, n53, n56, n57, n60, n61, n62,
         n63, n64, n65, n66, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n125, n126, n128, n129,
         n130, n196, n197, n198, n199, n200, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n44, n45, n46, n51, n52, n54, n55, n58, n59, n68, n78,
         n95, n124, n127, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248;

  SNPS_CLOCK_GATE_HIGH_isr_a0_0 clk_gate_ien0_reg_reg ( .CLK(clkper), .EN(N38), 
        .ENCLK(net12078), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_5 clk_gate_ien1_reg_reg ( .CLK(clkper), .EN(N49), 
        .ENCLK(net12084), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_4 clk_gate_ien2_reg_reg ( .CLK(clkper), .EN(N58), 
        .ENCLK(net12089), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_3 clk_gate_ip0_reg_reg ( .CLK(clkper), .EN(N67), 
        .ENCLK(net12094), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_2 clk_gate_ip1_reg_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12099), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_1 clk_gate_intvect_reg_reg ( .CLK(clkper), .EN(
        N207), .ENCLK(net12104), .TE(1'b0) );
  DFFQX1 intvect_reg_reg_2_ ( .D(N210), .C(net12104), .Q(intvect[2]) );
  DFFQX1 intvect_reg_reg_1_ ( .D(N209), .C(net12104), .Q(intvect[1]) );
  DFFQX1 intvect_reg_reg_0_ ( .D(N208), .C(net12104), .Q(intvect[0]) );
  DFFQX1 intvect_reg_reg_4_ ( .D(N212), .C(net12104), .Q(intvect[4]) );
  DFFQX1 intvect_reg_reg_3_ ( .D(N211), .C(net12104), .Q(intvect[3]) );
  DFFQX1 is_reg_s_reg_0_ ( .D(n199), .C(clkper), .Q(is_reg[0]) );
  DFFQX1 is_reg_s_reg_1_ ( .D(n196), .C(clkper), .Q(is_reg[1]) );
  DFFQX1 ien2_reg_reg_5_ ( .D(N64), .C(net12089), .Q(ien2[5]) );
  DFFQX1 is_reg_s_reg_2_ ( .D(n197), .C(clkper), .Q(is_reg[2]) );
  DFFQX1 ip1_reg_reg_5_ ( .D(N82), .C(net12099), .Q(ip1[5]) );
  DFFQX1 ip0_reg_reg_5_ ( .D(N73), .C(net12094), .Q(ip0[5]) );
  DFFQX1 ien0_reg_reg_4_ ( .D(N43), .C(net12078), .Q(ien0[4]) );
  DFFQX1 ien0_reg_reg_5_ ( .D(N44), .C(net12078), .Q(ien0[5]) );
  DFFQX1 ien2_reg_reg_4_ ( .D(N63), .C(net12089), .Q(ien2[4]) );
  DFFQX1 ien1_reg_reg_5_ ( .D(N55), .C(net12084), .Q(ien1[5]) );
  DFFQX1 ien1_reg_reg_4_ ( .D(N54), .C(net12084), .Q(ien1[4]) );
  DFFQX1 ip1_reg_reg_4_ ( .D(N81), .C(net12099), .Q(ip1[4]) );
  DFFQX1 ip0_reg_reg_4_ ( .D(N72), .C(net12094), .Q(ip0[4]) );
  DFFQX1 is_reg_s_reg_3_ ( .D(n198), .C(clkper), .Q(is_reg[3]) );
  DFFQX1 isr_tm_reg_reg ( .D(n200), .C(clkper), .Q(isr_tm) );
  DFFQX1 ien2_reg_reg_3_ ( .D(N62), .C(net12089), .Q(ien2[3]) );
  DFFQX1 ien0_reg_reg_3_ ( .D(N42), .C(net12078), .Q(ien0[3]) );
  DFFQX1 ip1_reg_reg_3_ ( .D(N80), .C(net12099), .Q(ip1[3]) );
  DFFQX1 ien1_reg_reg_3_ ( .D(N53), .C(net12084), .Q(ien1[3]) );
  DFFQX1 ip0_reg_reg_3_ ( .D(N71), .C(net12094), .Q(ip0[3]) );
  DFFQX1 irq_r_reg ( .D(N200), .C(clkper), .Q(irq_r) );
  DFFQX1 ien0_reg_reg_6_ ( .D(N45), .C(net12078), .Q(ien0[7]) );
  DFFQX1 ien2_reg_reg_0_ ( .D(N59), .C(net12089), .Q(ien2[0]) );
  DFFQX1 ien2_reg_reg_2_ ( .D(N61), .C(net12089), .Q(ien2[2]) );
  DFFQX1 ien0_reg_reg_1_ ( .D(N40), .C(net12078), .Q(ien0[1]) );
  DFFQX1 ien1_reg_reg_0_ ( .D(N50), .C(net12084), .Q(ien1[0]) );
  DFFQX1 ien0_reg_reg_2_ ( .D(N41), .C(net12078), .Q(ien0[2]) );
  DFFQX1 ien2_reg_reg_1_ ( .D(N60), .C(net12089), .Q(ien2[1]) );
  DFFQX1 ien0_reg_reg_0_ ( .D(N39), .C(net12078), .Q(ien0[0]) );
  DFFQX1 ip1_reg_reg_2_ ( .D(N79), .C(net12099), .Q(ip1[2]) );
  DFFQX1 ip1_reg_reg_0_ ( .D(N77), .C(net12099), .Q(ip1[0]) );
  DFFQX1 ip0_reg_reg_0_ ( .D(N68), .C(net12094), .Q(ip0[0]) );
  DFFQX1 ien1_reg_reg_2_ ( .D(N52), .C(net12084), .Q(ien1[2]) );
  DFFQX1 ien1_reg_reg_1_ ( .D(N51), .C(net12084), .Q(ien1[1]) );
  DFFQX1 ip0_reg_reg_1_ ( .D(N69), .C(net12094), .Q(ip0[1]) );
  DFFQX1 ip1_reg_reg_1_ ( .D(N78), .C(net12099), .Q(ip1[1]) );
  DFFQX1 ip0_reg_reg_2_ ( .D(N70), .C(net12094), .Q(ip0[2]) );
  INVX1 U3 ( .A(1'b1), .Y(ien0[6]) );
  MUX2X1 U5 ( .D0(int_vect_43), .D1(sdaiff), .S(isr_tm), .Y(n136) );
  AO21X1 U6 ( .B(ip0[5]), .C(n154), .A(n16), .Y(n155) );
  OA222X1 U7 ( .A(n216), .B(n215), .C(n214), .D(n213), .E(n212), .F(n211), .Y(
        n3) );
  NAND31XL U8 ( .C(sfraddr[6]), .A(n26), .B(sfrwe), .Y(n70) );
  NAND3X1 U9 ( .A(sfraddr[5]), .B(n23), .C(n84), .Y(n4) );
  INVX1 U10 ( .A(n77), .Y(n34) );
  NAND21X1 U11 ( .B(n20), .A(n33), .Y(n77) );
  INVX1 U12 ( .A(n83), .Y(n32) );
  INVX1 U13 ( .A(n79), .Y(n35) );
  INVX1 U14 ( .A(n82), .Y(n31) );
  NAND21X1 U15 ( .B(sfraddr[0]), .A(n33), .Y(n82) );
  NAND32X1 U16 ( .B(n20), .C(n4), .A(n25), .Y(n79) );
  NAND32X1 U17 ( .B(sfraddr[4]), .C(n4), .A(n20), .Y(n83) );
  INVX1 U18 ( .A(n30), .Y(n33) );
  NAND21X1 U19 ( .B(n4), .A(sfraddr[4]), .Y(n30) );
  NAND2X1 U20 ( .A(n26), .B(n79), .Y(N67) );
  NAND2X1 U21 ( .A(n26), .B(n83), .Y(N38) );
  NAND2X1 U22 ( .A(n26), .B(n82), .Y(N49) );
  NAND2X1 U23 ( .A(n26), .B(n77), .Y(N76) );
  INVX1 U24 ( .A(n80), .Y(n29) );
  NAND2X1 U25 ( .A(n26), .B(n80), .Y(N58) );
  INVX1 U26 ( .A(n22), .Y(n21) );
  NOR32XL U27 ( .B(n106), .C(n107), .A(n108), .Y(n92) );
  AND4X1 U28 ( .A(n107), .B(n88), .C(n114), .D(n109), .Y(n85) );
  NOR21XL U29 ( .B(n97), .A(n105), .Y(n114) );
  NAND21X1 U30 ( .B(n201), .A(n157), .Y(n214) );
  INVX1 U31 ( .A(sfraddr[4]), .Y(n25) );
  INVX1 U32 ( .A(n24), .Y(n23) );
  INVX1 U33 ( .A(n201), .Y(n202) );
  INVX1 U34 ( .A(sfraddr[0]), .Y(n20) );
  INVX1 U35 ( .A(n95), .Y(n59) );
  INVX1 U36 ( .A(n48), .Y(n247) );
  NAND2X1 U37 ( .A(n248), .B(n26), .Y(n43) );
  NAND2X1 U38 ( .A(n115), .B(n239), .Y(n109) );
  INVX1 U39 ( .A(n121), .Y(n239) );
  AND2X1 U40 ( .A(sfrdatai[0]), .B(n34), .Y(N77) );
  AND2X1 U41 ( .A(sfrdatai[1]), .B(n34), .Y(N78) );
  AND2X1 U42 ( .A(sfrdatai[2]), .B(n34), .Y(N79) );
  AND2X1 U43 ( .A(sfrdatai[3]), .B(n34), .Y(N80) );
  AND2X1 U44 ( .A(sfrdatai[4]), .B(n34), .Y(N81) );
  AND2X1 U45 ( .A(sfrdatai[5]), .B(n34), .Y(N82) );
  AND2X1 U46 ( .A(sfrdatai[0]), .B(n35), .Y(N68) );
  AND2X1 U47 ( .A(sfrdatai[1]), .B(n35), .Y(N69) );
  AND2X1 U48 ( .A(sfrdatai[2]), .B(n35), .Y(N70) );
  AND2X1 U49 ( .A(sfrdatai[3]), .B(n35), .Y(N71) );
  AND2X1 U50 ( .A(sfrdatai[4]), .B(n35), .Y(N72) );
  AND2X1 U51 ( .A(sfrdatai[5]), .B(n35), .Y(N73) );
  AND2X1 U52 ( .A(sfrdatai[0]), .B(n31), .Y(N50) );
  AND2X1 U53 ( .A(sfrdatai[1]), .B(n31), .Y(N51) );
  AND2X1 U54 ( .A(sfrdatai[2]), .B(n31), .Y(N52) );
  AND2X1 U55 ( .A(sfrdatai[3]), .B(n31), .Y(N53) );
  AND2X1 U56 ( .A(sfrdatai[4]), .B(n31), .Y(N54) );
  AND2X1 U57 ( .A(sfrdatai[5]), .B(n31), .Y(N55) );
  AND2X1 U58 ( .A(sfrdatai[0]), .B(n32), .Y(N39) );
  AND2X1 U59 ( .A(sfrdatai[1]), .B(n32), .Y(N40) );
  AND2X1 U60 ( .A(sfrdatai[2]), .B(n32), .Y(N41) );
  AND2X1 U61 ( .A(sfrdatai[3]), .B(n32), .Y(N42) );
  AND2X1 U62 ( .A(sfrdatai[4]), .B(n32), .Y(N43) );
  AND2X1 U63 ( .A(sfrdatai[5]), .B(n32), .Y(N44) );
  AND2X1 U64 ( .A(sfrdatai[7]), .B(n32), .Y(N45) );
  NOR3XL U65 ( .A(n70), .B(sfraddr[2]), .C(n21), .Y(n84) );
  NAND43X1 U66 ( .B(n22), .C(n24), .D(n25), .A(n81), .Y(n80) );
  NOR4XL U67 ( .A(sfraddr[5]), .B(sfraddr[2]), .C(sfraddr[0]), .D(n70), .Y(n81) );
  AND2X1 U68 ( .A(sfrdatai[0]), .B(n29), .Y(N59) );
  AND2X1 U69 ( .A(sfrdatai[1]), .B(n29), .Y(N60) );
  AND2X1 U70 ( .A(sfrdatai[2]), .B(n29), .Y(N61) );
  AND2X1 U71 ( .A(sfrdatai[3]), .B(n29), .Y(N62) );
  AND2X1 U72 ( .A(sfrdatai[4]), .B(n29), .Y(N63) );
  AND2X1 U73 ( .A(sfrdatai[5]), .B(n29), .Y(N64) );
  INVX1 U74 ( .A(sfraddr[1]), .Y(n22) );
  NOR32XL U75 ( .B(n113), .C(n112), .A(n7), .Y(n125) );
  NOR32XL U76 ( .B(n91), .C(n93), .A(n90), .Y(n117) );
  NOR32XL U77 ( .B(n126), .C(n117), .A(n116), .Y(n119) );
  NAND31X1 U78 ( .C(n8), .A(n129), .B(n125), .Y(n90) );
  NOR32XL U79 ( .B(n94), .C(n96), .A(n6), .Y(n112) );
  NAND32X1 U80 ( .B(n190), .C(n156), .A(n172), .Y(n201) );
  OAI211X1 U81 ( .C(n90), .D(n93), .A(n109), .B(n110), .Y(n101) );
  NAND21X1 U82 ( .B(n126), .A(n117), .Y(n106) );
  NAND21X1 U83 ( .B(n118), .A(n119), .Y(n97) );
  AND2X1 U84 ( .A(n8), .B(n125), .Y(n104) );
  AND2X1 U85 ( .A(n116), .B(n117), .Y(n105) );
  NAND2X1 U86 ( .A(n119), .B(n118), .Y(n121) );
  INVX1 U87 ( .A(n189), .Y(n172) );
  INVX1 U88 ( .A(sfraddr[3]), .Y(n24) );
  NOR43XL U89 ( .B(n98), .C(n123), .D(n106), .A(n104), .Y(n86) );
  AOI21X1 U90 ( .B(n7), .C(n112), .A(n128), .Y(n123) );
  AOI21X1 U91 ( .B(n93), .C(n91), .A(n90), .Y(n128) );
  NOR3XL U92 ( .A(n130), .B(rst), .C(intcall), .Y(N200) );
  NOR4XL U93 ( .A(n115), .B(n120), .C(n122), .D(n121), .Y(n130) );
  AOI31X1 U94 ( .A(n87), .B(n88), .C(n237), .D(rst), .Y(N210) );
  NAND32X1 U95 ( .B(n94), .C(n6), .A(n96), .Y(n87) );
  INVX1 U96 ( .A(n89), .Y(n237) );
  OAI31XL U97 ( .A(n90), .B(n241), .C(n91), .D(n92), .Y(n89) );
  AOI31X1 U98 ( .A(n238), .B(n92), .C(n102), .D(rst), .Y(N208) );
  INVX1 U99 ( .A(n101), .Y(n238) );
  NOR3XL U100 ( .A(n103), .B(n104), .C(n105), .Y(n102) );
  INVX1 U101 ( .A(n232), .Y(n103) );
  AOI31X1 U102 ( .A(n97), .B(n98), .C(n99), .D(rst), .Y(N209) );
  NOR2X1 U103 ( .A(n100), .B(n101), .Y(n99) );
  INVX1 U104 ( .A(n233), .Y(n100) );
  NOR2X1 U105 ( .A(rst), .B(n86), .Y(N211) );
  NOR2X1 U106 ( .A(rst), .B(n85), .Y(N212) );
  NAND4X1 U107 ( .A(n86), .B(n96), .C(n85), .D(n111), .Y(N207) );
  NOR43XL U108 ( .B(n94), .C(n110), .D(n26), .A(n108), .Y(n111) );
  INVX1 U109 ( .A(n184), .Y(n175) );
  NOR21XL U110 ( .B(n112), .A(n113), .Y(n108) );
  NAND21X1 U111 ( .B(n129), .A(n125), .Y(n98) );
  INVX1 U112 ( .A(n153), .Y(n157) );
  INVX1 U113 ( .A(n156), .Y(n144) );
  NAND2X1 U114 ( .A(n6), .B(n96), .Y(n110) );
  INVX1 U115 ( .A(n93), .Y(n241) );
  INVX1 U116 ( .A(n171), .Y(n173) );
  NAND21X1 U117 ( .B(n55), .A(n48), .Y(n95) );
  INVX1 U118 ( .A(intcall), .Y(n248) );
  NOR2X1 U119 ( .A(n248), .B(rst), .Y(n48) );
  INVX1 U120 ( .A(rst), .Y(n26) );
  NAND42X1 U121 ( .C(n120), .D(n121), .A(n122), .B(n240), .Y(n107) );
  INVX1 U122 ( .A(n240), .Y(n115) );
  INVX1 U123 ( .A(n231), .Y(n122) );
  NAND21X1 U124 ( .B(n3), .A(n230), .Y(n231) );
  NAND3X1 U125 ( .A(n239), .B(n240), .C(n120), .Y(n88) );
  NAND21X1 U126 ( .B(n224), .A(n178), .Y(n232) );
  OR2X1 U127 ( .A(n226), .B(n192), .Y(n233) );
  NAND21X1 U128 ( .B(n165), .A(n5), .Y(n189) );
  NAND2X1 U129 ( .A(n142), .B(n205), .Y(n149) );
  NAND21X1 U130 ( .B(n152), .A(n151), .Y(n171) );
  INVX1 U131 ( .A(n148), .Y(n152) );
  INVX1 U132 ( .A(n166), .Y(n151) );
  OA22X1 U133 ( .A(n16), .B(n210), .C(n212), .D(n209), .Y(n216) );
  OAI211X1 U134 ( .C(n5), .D(n168), .A(n163), .B(n11), .Y(n184) );
  NAND21X1 U135 ( .B(n3), .A(n13), .Y(n113) );
  NAND21X1 U136 ( .B(n228), .A(n162), .Y(n94) );
  INVX1 U137 ( .A(n194), .Y(n96) );
  OAI211X1 U138 ( .C(n218), .D(n193), .A(n232), .B(n233), .Y(n194) );
  AND2X1 U139 ( .A(n193), .B(n217), .Y(n5) );
  NOR2X1 U140 ( .A(n227), .B(n208), .Y(n6) );
  INVX1 U141 ( .A(n145), .Y(n205) );
  OAI211X1 U142 ( .C(n144), .D(n181), .A(n175), .B(n180), .Y(n145) );
  INVX1 U143 ( .A(n191), .Y(n226) );
  OAI221X1 U144 ( .A(n190), .B(n189), .C(n188), .D(n187), .E(n186), .Y(n191)
         );
  GEN2XL U145 ( .D(n185), .E(n184), .C(n183), .B(n182), .A(n181), .Y(n186) );
  INVX1 U146 ( .A(n180), .Y(n183) );
  NAND32X1 U147 ( .B(n178), .C(n14), .A(n219), .Y(n190) );
  NAND21X1 U148 ( .B(n227), .A(n222), .Y(n93) );
  NAND32X1 U149 ( .B(n162), .C(n19), .A(n221), .Y(n213) );
  NAND32X1 U150 ( .B(n12), .C(n220), .A(n192), .Y(n156) );
  NAND32X1 U151 ( .B(n15), .C(n13), .A(n223), .Y(n154) );
  NAND32X1 U152 ( .B(n18), .C(n222), .A(n208), .Y(n153) );
  NAND21X1 U153 ( .B(n226), .A(n220), .Y(n129) );
  OR3XL U154 ( .A(n19), .B(n228), .C(n221), .Y(n91) );
  NAND32X1 U155 ( .B(n230), .C(n3), .A(n15), .Y(n126) );
  INVX1 U156 ( .A(n225), .Y(n116) );
  NAND21X1 U157 ( .B(n224), .A(n14), .Y(n225) );
  NOR2X1 U158 ( .A(n218), .B(n217), .Y(n7) );
  NOR2X1 U159 ( .A(n224), .B(n219), .Y(n8) );
  NAND21X1 U160 ( .B(n226), .A(n12), .Y(n118) );
  ENOX1 U161 ( .A(n244), .B(n75), .C(n76), .D(intcall), .Y(int_ack_03) );
  OAI21X1 U162 ( .B(n246), .C(n245), .A(n60), .Y(n76) );
  AOI211X1 U163 ( .C(n66), .D(n67), .A(int_ack_03), .B(int_ack_43), .Y(n50) );
  OAI22AX1 U164 ( .D(n124), .C(n95), .A(n47), .B(n164), .Y(n198) );
  OAI21X1 U165 ( .B(n43), .C(n131), .A(n127), .Y(n197) );
  AO21X1 U166 ( .B(n47), .C(n164), .A(n234), .Y(n131) );
  AO21X1 U167 ( .B(n124), .C(n234), .A(n95), .Y(n127) );
  NOR2X1 U168 ( .A(n73), .B(n244), .Y(int_ack_43) );
  INVX1 U169 ( .A(n54), .Y(n55) );
  NAND31X1 U170 ( .C(retiinstr), .A(n247), .B(n26), .Y(n47) );
  NOR2X1 U171 ( .A(n65), .B(n75), .Y(int_ack_13) );
  NOR2X1 U172 ( .A(n63), .B(n75), .Y(int_ack_1b) );
  NAND3X1 U173 ( .A(n60), .B(n61), .C(n243), .Y(n9) );
  AND2X1 U174 ( .A(n60), .B(n245), .Y(n62) );
  NOR2X1 U175 ( .A(n64), .B(n75), .Y(int_ack_0b) );
  NOR2X1 U176 ( .A(n65), .B(n242), .Y(int_ack_93) );
  NOR2X1 U177 ( .A(n64), .B(n242), .Y(int_ack_8b) );
  INVX1 U178 ( .A(n53), .Y(n44) );
  NOR21XL U179 ( .B(n62), .A(n63), .Y(n53) );
  INVX1 U180 ( .A(n57), .Y(n40) );
  NOR21XL U181 ( .B(n62), .A(n64), .Y(n57) );
  NOR2X1 U182 ( .A(n243), .B(n72), .Y(int_ack_6b) );
  NOR2X1 U183 ( .A(n65), .B(n73), .Y(int_ack_53) );
  NOR2X1 U184 ( .A(n63), .B(n73), .Y(int_ack_5b) );
  NOR2X1 U185 ( .A(n64), .B(n73), .Y(int_ack_4b) );
  INVX1 U186 ( .A(n67), .Y(n242) );
  INVX1 U187 ( .A(n66), .Y(n244) );
  INVX1 U188 ( .A(n56), .Y(n52) );
  NOR21XL U189 ( .B(n62), .A(n65), .Y(n56) );
  NAND21X1 U190 ( .B(n227), .A(n18), .Y(n240) );
  INVX1 U191 ( .A(n223), .Y(n230) );
  INVX1 U192 ( .A(n229), .Y(n120) );
  NAND21X1 U193 ( .B(n228), .A(n19), .Y(n229) );
  NOR3XL U194 ( .A(n71), .B(n245), .C(n244), .Y(int_ack_a3) );
  NOR3XL U195 ( .A(n71), .B(n245), .C(n64), .Y(int_ack_ab) );
  NOR2X1 U196 ( .A(n63), .B(n242), .Y(int_ack_9b) );
  AND2X1 U197 ( .A(irq_r), .B(ien0[7]), .Y(irq) );
  MUX2X1 U198 ( .D0(n28), .D1(sfrdatai[5]), .S(n27), .Y(n200) );
  AND2X1 U199 ( .A(isr_tm), .B(n26), .Y(n28) );
  AND4XL U200 ( .A(sfraddr[2]), .B(n69), .C(n21), .D(sfraddr[0]), .Y(n27) );
  NOR4XL U201 ( .A(sfraddr[5]), .B(sfraddr[4]), .C(n23), .D(n70), .Y(n69) );
  INVX1 U202 ( .A(n177), .Y(n224) );
  GEN2XL U203 ( .D(n176), .E(ip0[1]), .C(n175), .B(ip1[1]), .A(n174), .Y(n177)
         );
  INVX1 U204 ( .A(n179), .Y(n176) );
  AO21X1 U205 ( .B(n173), .C(ip0[1]), .A(n172), .Y(n174) );
  INVX1 U206 ( .A(n207), .Y(n227) );
  GEN2XL U207 ( .D(n206), .E(ip0[3]), .C(n205), .B(ip1[3]), .A(n204), .Y(n207)
         );
  AO21X1 U208 ( .B(n203), .C(ip0[3]), .A(n202), .Y(n204) );
  INVX1 U209 ( .A(n195), .Y(n203) );
  NAND2X1 U210 ( .A(ien1[0]), .B(n136), .Y(n217) );
  AO21X1 U211 ( .B(ip0[3]), .C(n153), .A(n195), .Y(n210) );
  AO21X1 U212 ( .B(ip0[2]), .C(n156), .A(n187), .Y(n195) );
  NAND21X1 U213 ( .B(n5), .A(ip0[0]), .Y(n148) );
  NAND2X1 U214 ( .A(ien0[0]), .B(int_vect_03), .Y(n193) );
  NAND32X1 U215 ( .B(is_reg[1]), .C(n211), .A(n150), .Y(n166) );
  NAND3X1 U216 ( .A(n147), .B(n10), .C(n206), .Y(n209) );
  NAND3X1 U217 ( .A(ip1[4]), .B(ip0[4]), .C(n213), .Y(n10) );
  OAI211X1 U218 ( .C(n148), .D(n168), .A(ien0[7]), .B(n164), .Y(n179) );
  INVX1 U219 ( .A(n161), .Y(n228) );
  OAI221X1 U220 ( .A(n160), .B(n159), .C(n158), .D(n210), .E(n214), .Y(n161)
         );
  AOI31X1 U221 ( .A(ip0[4]), .B(n206), .C(n147), .D(n146), .Y(n160) );
  INVX1 U222 ( .A(n149), .Y(n146) );
  AO21X1 U223 ( .B(ip1[4]), .C(n213), .A(n149), .Y(n211) );
  AO21X1 U224 ( .B(ip0[1]), .C(n190), .A(n171), .Y(n187) );
  OR3XL U225 ( .A(is_reg[0]), .B(n155), .C(n210), .Y(n165) );
  INVX1 U226 ( .A(n138), .Y(n206) );
  OAI31XL U227 ( .A(n144), .B(n188), .C(n181), .D(n137), .Y(n138) );
  AOI31X1 U228 ( .A(ip1[1]), .B(ip0[1]), .C(n190), .D(n179), .Y(n137) );
  NOR2X1 U229 ( .A(is_reg[2]), .B(n209), .Y(n11) );
  NOR21XL U230 ( .B(ien0[4]), .A(n143), .Y(n162) );
  MUX2IX1 U231 ( .D0(int_vect_23), .D1(rxd0ff), .S(isr_tm), .Y(n143) );
  NAND42X1 U232 ( .C(isr_tm), .D(n14), .A(ien1[1]), .B(int_vect_4b), .Y(n219)
         );
  NAND32X1 U233 ( .B(n141), .C(isr_tm), .A(int_vect_1b), .Y(n208) );
  INVX1 U234 ( .A(ien0[3]), .Y(n141) );
  NAND21X1 U235 ( .B(n142), .A(ip0[3]), .Y(n147) );
  NAND21X1 U236 ( .B(n157), .A(ip1[3]), .Y(n142) );
  NAND2X1 U237 ( .A(n154), .B(ip1[5]), .Y(n150) );
  NAND21X1 U238 ( .B(n150), .A(ip0[5]), .Y(n163) );
  INVX1 U239 ( .A(ip1[0]), .Y(n168) );
  INVX1 U240 ( .A(n133), .Y(n220) );
  NAND32X1 U241 ( .B(n132), .C(n12), .A(int_vect_53), .Y(n133) );
  INVX1 U242 ( .A(ien1[2]), .Y(n132) );
  INVX1 U243 ( .A(n140), .Y(n222) );
  NAND32X1 U244 ( .B(n139), .C(n18), .A(int_vect_5b), .Y(n140) );
  INVX1 U245 ( .A(ien1[3]), .Y(n139) );
  INVX1 U246 ( .A(n135), .Y(n178) );
  NAND32X1 U247 ( .B(n134), .C(isr_tm), .A(int_vect_0b), .Y(n135) );
  INVX1 U248 ( .A(ien0[1]), .Y(n134) );
  AND2X1 U249 ( .A(ien2[2]), .B(int_vect_93), .Y(n12) );
  AND2X1 U250 ( .A(ien0[5]), .B(i2c_int), .Y(n13) );
  INVX1 U251 ( .A(is_reg[3]), .Y(n164) );
  AND2X1 U252 ( .A(ien2[1]), .B(int_vect_8b), .Y(n14) );
  INVX1 U253 ( .A(n170), .Y(n218) );
  OAI221X1 U254 ( .A(n169), .B(n168), .C(n167), .D(n166), .E(n165), .Y(n170)
         );
  AOI32X1 U255 ( .A(ien0[7]), .B(ip0[0]), .C(n164), .D(n11), .E(n163), .Y(n169) );
  NAND2X1 U256 ( .A(ien1[4]), .B(int_vect_63), .Y(n221) );
  NAND2X1 U257 ( .A(n190), .B(ip1[1]), .Y(n180) );
  INVX1 U258 ( .A(ip0[2]), .Y(n188) );
  INVX1 U259 ( .A(ip1[2]), .Y(n181) );
  AND2X1 U260 ( .A(ien1[5]), .B(int_vect_6b), .Y(n15) );
  NAND2X1 U261 ( .A(ien0[2]), .B(int_vect_13), .Y(n192) );
  AND2X1 U262 ( .A(n213), .B(ip0[4]), .Y(n16) );
  NAND21X1 U263 ( .B(n179), .A(ip0[2]), .Y(n185) );
  OR2X1 U264 ( .A(ip0[1]), .B(n185), .Y(n182) );
  NAND21X1 U265 ( .B(intvect[3]), .A(n74), .Y(n75) );
  OAI211X1 U266 ( .C(n181), .D(n52), .A(n39), .B(n38), .Y(n54) );
  OA222X1 U267 ( .A(n212), .B(n17), .C(n37), .D(n44), .E(n159), .F(n9), .Y(n38) );
  OA22X1 U268 ( .A(n50), .B(n168), .C(n36), .D(n40), .Y(n39) );
  INVX1 U269 ( .A(ip1[3]), .Y(n37) );
  GEN2XL U270 ( .D(n78), .E(n68), .C(n59), .B(is_reg[1]), .A(n58), .Y(n196) );
  INVX1 U271 ( .A(n43), .Y(n78) );
  INVX1 U272 ( .A(n42), .Y(n68) );
  AND3X1 U273 ( .A(n55), .B(n124), .C(n48), .Y(n58) );
  NOR3XL U274 ( .A(intvect[2]), .B(intvect[4]), .C(n248), .Y(n74) );
  INVX1 U275 ( .A(ip0[0]), .Y(n167) );
  NAND2X1 U276 ( .A(n74), .B(intvect[3]), .Y(n73) );
  NOR32XL U277 ( .B(n234), .C(n47), .A(is_reg[3]), .Y(n42) );
  NAND31X1 U278 ( .C(intvect[3]), .A(intcall), .B(intvect[4]), .Y(n71) );
  OAI211X1 U279 ( .C(n188), .D(n52), .A(n51), .B(n46), .Y(n124) );
  OA222X1 U280 ( .A(n215), .B(n17), .C(n45), .D(n44), .E(n158), .F(n9), .Y(n46) );
  OA22X1 U281 ( .A(n50), .B(n167), .C(n41), .D(n40), .Y(n51) );
  INVX1 U282 ( .A(ip0[3]), .Y(n45) );
  NOR2X1 U283 ( .A(n71), .B(intvect[2]), .Y(n67) );
  NOR3XL U284 ( .A(n248), .B(intvect[1]), .C(n245), .Y(n61) );
  OAI31XL U285 ( .A(n247), .B(n54), .C(n124), .D(n49), .Y(n199) );
  GEN2XL U286 ( .D(n42), .E(n235), .C(n43), .B(n247), .A(n236), .Y(n49) );
  INVX1 U287 ( .A(is_reg[0]), .Y(n236) );
  INVX1 U288 ( .A(is_reg[1]), .Y(n235) );
  NAND2X1 U289 ( .A(intvect[4]), .B(intvect[3]), .Y(n60) );
  INVX1 U290 ( .A(ip0[4]), .Y(n158) );
  INVX1 U291 ( .A(ip1[5]), .Y(n212) );
  INVX1 U292 ( .A(ip0[5]), .Y(n215) );
  INVX1 U293 ( .A(ip1[4]), .Y(n159) );
  NAND3X1 U294 ( .A(n61), .B(n60), .C(intvect[0]), .Y(n17) );
  NAND31X1 U295 ( .C(intvect[4]), .A(intvect[3]), .B(n61), .Y(n72) );
  NOR2X1 U296 ( .A(intvect[0]), .B(intvect[1]), .Y(n66) );
  INVX1 U297 ( .A(intvect[0]), .Y(n243) );
  NAND2X1 U298 ( .A(intvect[1]), .B(intvect[0]), .Y(n63) );
  INVX1 U299 ( .A(intvect[1]), .Y(n246) );
  INVX1 U300 ( .A(intvect[2]), .Y(n245) );
  NOR2X1 U301 ( .A(intvect[0]), .B(n72), .Y(int_ack_63) );
  NAND2X1 U302 ( .A(intvect[0]), .B(n246), .Y(n64) );
  NAND2X1 U303 ( .A(intvect[1]), .B(n243), .Y(n65) );
  INVX1 U304 ( .A(ip1[1]), .Y(n36) );
  INVX1 U305 ( .A(is_reg[2]), .Y(n234) );
  INVX1 U306 ( .A(ip0[1]), .Y(n41) );
  NAND2X1 U307 ( .A(ien2[5]), .B(int_vect_ab), .Y(n223) );
  AND2X1 U308 ( .A(ien2[3]), .B(int_vect_9b), .Y(n18) );
  AND2X1 U309 ( .A(ien2[4]), .B(int_vect_a3), .Y(n19) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module watchdog_a0 ( wdt_slow, clkwdt, clkper, resetff, newinstr, wdts_s, wdts, 
        ip0wdts, wdt_tm, sfrdatai, sfraddr, sfrwe, wdtrel );
  output [1:0] wdts_s;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] wdtrel;
  input wdt_slow, clkwdt, clkper, resetff, newinstr, sfrwe;
  output wdts, ip0wdts, wdt_tm;
  wire   wdt_tm_sync, wdt_act_sync, wdt_act, wdtrefresh_sync, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N67, N68, N69, N70, N71, pres_2, N112,
         N113, N114, N115, N116, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, wdt_normal, wdt_normal_ff, N212, net12127, net12133,
         net12138, net12143, net12148, n21, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n59, n60, n61, n62, n63, n64,
         n65, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n107, n108, n109, n110,
         n111, n112, n113, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n58,
         n66, n78, n79, n92, n93, n106, n114, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145;
  wire   [1:0] pres_8;
  wire   [3:0] cycles_reg;
  wire   [3:0] pres_16;
  wire   [6:0] wdth;
  wire   [7:0] wdtl;

  SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 clk_gate_wdtrel_s_reg ( .CLK(clkper), 
        .EN(N26), .ENCLK(net12127), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 clk_gate_cycles_reg_reg ( .CLK(clkwdt), 
        .EN(N67), .ENCLK(net12133), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 clk_gate_pres_16_reg ( .CLK(clkwdt), .EN(
        N112), .ENCLK(net12138), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 clk_gate_wdth_reg ( .CLK(clkwdt), .EN(
        N165), .ENCLK(net12143), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 clk_gate_wdtl_reg ( .CLK(clkwdt), .EN(n21), .ENCLK(net12148), .TE(1'b0) );
  watchdog_a0_DW01_inc_0 add_278 ( .A(wdtl), .SUM({N144, N143, N142, N141, 
        N140, N139, N138, N137}) );
  watchdog_a0_DW01_inc_1 add_272 ( .A(wdth), .SUM({N136, N135, N134, N133, 
        N132, N131, N130}) );
  DFFQX1 wdts_s_reg_1_ ( .D(n126), .C(net12148), .Q(wdts_s[1]) );
  DFFQX1 wdt_act_reg ( .D(n130), .C(clkper), .Q(wdt_act) );
  DFFQX1 wdts_reg ( .D(wdts_s[0]), .C(clkper), .Q(wdts) );
  DFFQX1 wdt_normal_ff_reg ( .D(n78), .C(clkper), .Q(wdt_normal_ff) );
  DFFQX1 wdt_normal_reg ( .D(n133), .C(clkper), .Q(wdt_normal) );
  DFFQX1 wdts_s_reg_0_ ( .D(n132), .C(net12148), .Q(wdts_s[0]) );
  DFFQX1 wdt_act_sync_reg ( .D(wdt_act), .C(clkwdt), .Q(wdt_act_sync) );
  DFFQX1 pres_16_reg_3_ ( .D(N116), .C(net12138), .Q(pres_16[3]) );
  DFFQX1 wdth_reg_6_ ( .D(N172), .C(net12143), .Q(wdth[6]) );
  DFFQX1 pres_16_reg_1_ ( .D(N114), .C(net12138), .Q(pres_16[1]) );
  DFFQX1 pres_16_reg_0_ ( .D(N113), .C(net12138), .Q(pres_16[0]) );
  DFFQX1 pres_16_reg_2_ ( .D(N115), .C(net12138), .Q(pres_16[2]) );
  DFFQX1 pres_8_reg_0_ ( .D(n129), .C(net12133), .Q(pres_8[0]) );
  DFFQX1 pres_8_reg_1_ ( .D(n128), .C(net12133), .Q(pres_8[1]) );
  DFFQX1 wdt_tm_sync_reg ( .D(wdt_tm), .C(clkwdt), .Q(wdt_tm_sync) );
  DFFQX1 pres_2_reg ( .D(n127), .C(net12133), .Q(pres_2) );
  DFFQX1 wdtl_reg_2_ ( .D(N175), .C(net12148), .Q(wdtl[2]) );
  DFFQX1 wdtrefresh_reg ( .D(N212), .C(clkper), .Q(wdtrefresh_sync) );
  DFFQX1 cycles_reg_reg_2_ ( .D(N70), .C(net12133), .Q(cycles_reg[2]) );
  DFFQX1 cycles_reg_reg_1_ ( .D(N69), .C(net12133), .Q(cycles_reg[1]) );
  DFFQX1 wdtl_reg_1_ ( .D(N174), .C(net12148), .Q(wdtl[1]) );
  DFFQX1 wdtl_reg_0_ ( .D(N173), .C(net12148), .Q(wdtl[0]) );
  DFFQX1 cycles_reg_reg_0_ ( .D(N68), .C(net12133), .Q(cycles_reg[0]) );
  DFFQX1 wdtl_reg_3_ ( .D(N176), .C(net12148), .Q(wdtl[3]) );
  DFFQX1 cycles_reg_reg_3_ ( .D(N71), .C(net12133), .Q(cycles_reg[3]) );
  DFFQX1 wdtl_reg_4_ ( .D(N177), .C(net12148), .Q(wdtl[4]) );
  DFFQX1 wdth_reg_1_ ( .D(N167), .C(net12143), .Q(wdth[1]) );
  DFFQX1 wdtl_reg_7_ ( .D(N180), .C(net12148), .Q(wdtl[7]) );
  DFFQX1 wdth_reg_3_ ( .D(N169), .C(net12143), .Q(wdth[3]) );
  DFFQX1 wdth_reg_0_ ( .D(N166), .C(net12143), .Q(wdth[0]) );
  DFFQX1 wdth_reg_4_ ( .D(N170), .C(net12143), .Q(wdth[4]) );
  DFFQX1 wdth_reg_5_ ( .D(N171), .C(net12143), .Q(wdth[5]) );
  DFFQX1 wdth_reg_2_ ( .D(N168), .C(net12143), .Q(wdth[2]) );
  DFFQX1 wdtl_reg_5_ ( .D(N178), .C(net12148), .Q(wdtl[5]) );
  DFFQX1 wdtl_reg_6_ ( .D(N179), .C(net12148), .Q(wdtl[6]) );
  DFFQX1 ip0wdts_reg ( .D(n131), .C(clkper), .Q(ip0wdts) );
  DFFQX1 wdtrel_s_reg_7_ ( .D(N34), .C(net12127), .Q(wdtrel[7]) );
  DFFQX1 wdt_tm_s_reg ( .D(n134), .C(clkper), .Q(wdt_tm) );
  DFFQX1 wdtrel_s_reg_6_ ( .D(N33), .C(net12127), .Q(wdtrel[6]) );
  DFFQX1 wdtrel_s_reg_4_ ( .D(N31), .C(net12127), .Q(wdtrel[4]) );
  DFFQX1 wdtrel_s_reg_5_ ( .D(N32), .C(net12127), .Q(wdtrel[5]) );
  DFFQX1 wdtrel_s_reg_3_ ( .D(N30), .C(net12127), .Q(wdtrel[3]) );
  DFFQX1 wdtrel_s_reg_2_ ( .D(N29), .C(net12127), .Q(wdtrel[2]) );
  DFFQX1 wdtrel_s_reg_0_ ( .D(N27), .C(net12127), .Q(wdtrel[0]) );
  DFFQX1 wdtrel_s_reg_1_ ( .D(N28), .C(net12127), .Q(wdtrel[1]) );
  NAND4XL U3 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(n41), .D(n91), .Y(n90) );
  NOR31XL U4 ( .C(sfraddr[3]), .A(n5), .B(n3), .Y(n81) );
  INVX1 U5 ( .A(n95), .Y(n41) );
  INVX1 U6 ( .A(n4), .Y(n3) );
  INVX1 U7 ( .A(n6), .Y(n5) );
  NOR43XL U8 ( .B(n107), .C(n108), .D(sfraddr[3]), .A(sfraddr[0]), .Y(n77) );
  NOR3XL U9 ( .A(n3), .B(sfraddr[6]), .C(n5), .Y(n107) );
  AND4X1 U10 ( .A(sfraddr[4]), .B(sfraddr[5]), .C(sfrwe), .D(sfrdatai[6]), .Y(
        n108) );
  INVX1 U11 ( .A(n89), .Y(n79) );
  AND2X1 U12 ( .A(sfrdatai[0]), .B(n11), .Y(N27) );
  AND2X1 U13 ( .A(sfrdatai[7]), .B(n11), .Y(N34) );
  AND2X1 U14 ( .A(sfrdatai[1]), .B(n11), .Y(N28) );
  AND2X1 U15 ( .A(sfrdatai[2]), .B(n11), .Y(N29) );
  AND2X1 U16 ( .A(sfrdatai[3]), .B(n11), .Y(N30) );
  AND2X1 U17 ( .A(sfrdatai[4]), .B(n11), .Y(N31) );
  AND2X1 U18 ( .A(sfrdatai[5]), .B(n11), .Y(N32) );
  AND2X1 U19 ( .A(n11), .B(sfrdatai[6]), .Y(N33) );
  NOR3XL U20 ( .A(sfraddr[0]), .B(n5), .C(n3), .Y(n91) );
  INVX1 U21 ( .A(sfrdatai[6]), .Y(n7) );
  INVX1 U22 ( .A(sfraddr[1]), .Y(n4) );
  INVX1 U23 ( .A(sfraddr[2]), .Y(n6) );
  NAND2X1 U24 ( .A(n69), .B(n137), .Y(n121) );
  NOR32XL U25 ( .B(n42), .C(n90), .A(newinstr), .Y(n89) );
  INVX1 U26 ( .A(n105), .Y(n11) );
  NAND2X1 U27 ( .A(n42), .B(n105), .Y(N26) );
  INVX1 U28 ( .A(n28), .Y(n24) );
  INVX1 U29 ( .A(n32), .Y(n27) );
  INVX1 U30 ( .A(n23), .Y(n31) );
  NAND4X1 U31 ( .A(n59), .B(n60), .C(n61), .D(n62), .Y(n54) );
  XOR2X1 U32 ( .A(n26), .B(n25), .Y(n60) );
  XOR2X1 U33 ( .A(n30), .B(n29), .Y(n61) );
  XOR2X1 U34 ( .A(n34), .B(n33), .Y(n62) );
  OR2X1 U35 ( .A(n69), .B(n19), .Y(n68) );
  NAND2X1 U36 ( .A(n110), .B(n50), .Y(n43) );
  NAND21X1 U37 ( .B(n19), .A(n17), .Y(n70) );
  AND2X1 U38 ( .A(n73), .B(n115), .Y(n69) );
  INVX1 U39 ( .A(n73), .Y(n17) );
  OAI21X1 U40 ( .B(n123), .C(n121), .A(n103), .Y(N115) );
  XNOR2XL U41 ( .A(n122), .B(n135), .Y(n123) );
  OAI211X1 U42 ( .C(n50), .D(n113), .A(n106), .B(n42), .Y(N165) );
  INVX1 U43 ( .A(n112), .Y(n106) );
  NAND2X1 U44 ( .A(n111), .B(n110), .Y(n113) );
  NAND21X1 U45 ( .B(n18), .A(n137), .Y(n103) );
  NOR21XL U46 ( .B(N143), .A(n43), .Y(N179) );
  NOR21XL U47 ( .B(N142), .A(n43), .Y(N178) );
  NOR21XL U48 ( .B(N141), .A(n43), .Y(N177) );
  NOR21XL U49 ( .B(N140), .A(n43), .Y(N176) );
  NOR21XL U50 ( .B(N139), .A(n43), .Y(N175) );
  NOR21XL U51 ( .B(N138), .A(n43), .Y(N174) );
  NOR2X1 U52 ( .A(n135), .B(n122), .Y(n116) );
  NAND2X1 U53 ( .A(n99), .B(n137), .Y(n96) );
  INVX1 U54 ( .A(n72), .Y(n137) );
  NOR2X1 U55 ( .A(n140), .B(n58), .Y(n115) );
  INVX1 U56 ( .A(n101), .Y(n138) );
  NAND2X1 U57 ( .A(n42), .B(n72), .Y(N67) );
  OR4X1 U58 ( .A(n95), .B(n4), .C(n6), .D(n1), .Y(n105) );
  OR4XL U59 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(sfraddr[0]), .D(resetff), .Y(
        n1) );
  MUX2X1 U60 ( .D0(n9), .D1(sfrdatai[6]), .S(n8), .Y(n134) );
  AND2X1 U61 ( .A(wdt_tm), .B(n42), .Y(n9) );
  AND4X1 U62 ( .A(n94), .B(n5), .C(sfraddr[0]), .D(n3), .Y(n8) );
  NOR4XL U63 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(resetff), .D(n95), .Y(n94)
         );
  OAI32X1 U64 ( .A(n90), .B(resetff), .C(n7), .D(n93), .E(n79), .Y(n133) );
  INVX1 U65 ( .A(wdt_normal), .Y(n93) );
  ENOX1 U66 ( .A(resetff), .B(n76), .C(wdt_act), .D(n76), .Y(n130) );
  OAI21X1 U67 ( .B(n77), .C(resetff), .A(n136), .Y(n76) );
  AND2X1 U68 ( .A(n13), .B(n42), .Y(n131) );
  MUX2X1 U69 ( .D0(sfrdatai[6]), .D1(n12), .S(n80), .Y(n13) );
  NAND21X1 U70 ( .B(ip0wdts), .A(n136), .Y(n12) );
  NAND4X1 U71 ( .A(n41), .B(sfraddr[5]), .C(sfraddr[0]), .D(n81), .Y(n80) );
  INVX1 U72 ( .A(n88), .Y(n78) );
  AOI32X1 U73 ( .A(wdt_normal), .B(n42), .C(n79), .D(n89), .E(wdt_normal_ff), 
        .Y(n88) );
  AND3X1 U74 ( .A(n77), .B(wdt_normal_ff), .C(n42), .Y(N212) );
  OR2X1 U75 ( .A(wdtrel[0]), .B(wdtrel[1]), .Y(n28) );
  NAND21X1 U76 ( .B(wdtrel[2]), .A(n24), .Y(n32) );
  NAND21X1 U77 ( .B(wdtrel[3]), .A(n27), .Y(n23) );
  INVX1 U78 ( .A(n22), .Y(n40) );
  NAND21X1 U79 ( .B(wdtrel[4]), .A(n31), .Y(n22) );
  XOR2X1 U80 ( .A(wdth[3]), .B(n2), .Y(n59) );
  AOI21X1 U81 ( .B(wdtrel[4]), .C(n23), .A(n40), .Y(n2) );
  AO21X1 U82 ( .B(wdtrel[3]), .C(n32), .A(n31), .Y(n33) );
  AO21X1 U83 ( .B(wdtrel[2]), .C(n28), .A(n27), .Y(n29) );
  NAND21X1 U84 ( .B(wdtrel[5]), .A(n40), .Y(n38) );
  OAI21X1 U85 ( .B(n43), .C(n44), .A(n45), .Y(n126) );
  NAND41X1 U86 ( .D(n46), .A(wdts_s[1]), .B(n47), .C(n44), .Y(n45) );
  OAI31XL U87 ( .A(n141), .B(n48), .C(n49), .D(n50), .Y(n46) );
  NAND3X1 U88 ( .A(n51), .B(n52), .C(n53), .Y(n44) );
  NOR4XL U89 ( .A(n54), .B(n55), .C(n56), .D(n57), .Y(n53) );
  XOR2X1 U90 ( .A(n37), .B(n36), .Y(n55) );
  XOR3X1 U91 ( .A(wdth[4]), .B(wdtrel[5]), .C(n40), .Y(n57) );
  XOR3X1 U92 ( .A(n39), .B(wdth[5]), .C(n38), .Y(n56) );
  AO21X1 U93 ( .B(wdtrel[0]), .C(wdtrel[1]), .A(n24), .Y(n25) );
  OAI22AX1 U94 ( .D(n82), .C(n43), .A(n136), .B(n82), .Y(n132) );
  OAI211X1 U95 ( .C(n83), .D(n84), .A(n50), .B(n47), .Y(n82) );
  NAND4X1 U96 ( .A(n86), .B(n141), .C(wdth[2]), .D(n87), .Y(n83) );
  NAND3X1 U97 ( .A(n48), .B(wdth[6]), .C(n85), .Y(n84) );
  NOR3XL U98 ( .A(n49), .B(n144), .C(n143), .Y(n85) );
  INVX1 U99 ( .A(wdth[4]), .Y(n143) );
  INVX1 U100 ( .A(wdth[5]), .Y(n144) );
  NAND4X1 U101 ( .A(n117), .B(n118), .C(wdtl[3]), .D(n119), .Y(n49) );
  AND2X1 U102 ( .A(wdtl[0]), .B(wdtl[1]), .Y(n119) );
  XNOR2XL U103 ( .A(n145), .B(wdtl[5]), .Y(n117) );
  XNOR2XL U104 ( .A(n145), .B(wdtl[6]), .Y(n118) );
  NOR21XL U105 ( .B(n104), .A(wdtrefresh_sync), .Y(n73) );
  NAND42X1 U106 ( .C(n49), .D(n141), .A(wdtl[4]), .B(n86), .Y(n50) );
  NOR43XL U107 ( .B(n115), .C(n104), .D(pres_2), .A(n16), .Y(n111) );
  NOR21XL U108 ( .B(wdtrel[7]), .A(n15), .Y(n16) );
  NOR21XL U109 ( .B(pres_16[3]), .A(n14), .Y(n15) );
  INVX1 U110 ( .A(n116), .Y(n14) );
  NOR21XL U111 ( .B(N144), .A(n43), .Y(N180) );
  XNOR2XL U112 ( .A(wdtl[4]), .B(wdt_slow), .Y(n48) );
  AO22X1 U113 ( .A(wdtrel[6]), .B(n112), .C(N136), .D(n110), .Y(N172) );
  AO22X1 U114 ( .A(wdtrel[5]), .B(n112), .C(N135), .D(n110), .Y(N171) );
  OAI22X1 U115 ( .A(n58), .B(n70), .C(n75), .D(n72), .Y(n129) );
  OA21X1 U116 ( .B(pres_8[0]), .C(n17), .A(n18), .Y(n75) );
  NAND2X1 U117 ( .A(cycles_reg[1]), .B(cycles_reg[0]), .Y(n101) );
  NOR3XL U118 ( .A(n101), .B(cycles_reg[2]), .C(n139), .Y(n104) );
  OAI32X1 U119 ( .A(n67), .B(resetff), .C(n92), .D(n68), .E(n66), .Y(n127) );
  INVX1 U120 ( .A(pres_2), .Y(n66) );
  OA21X1 U121 ( .B(pres_2), .C(wdtrefresh_sync), .A(n18), .Y(n67) );
  INVX1 U122 ( .A(n68), .Y(n92) );
  NOR42XL U123 ( .C(wdtl[2]), .D(wdtl[0]), .A(n64), .B(n65), .Y(n51) );
  XOR2X1 U124 ( .A(n20), .B(wdtl[4]), .Y(n64) );
  XNOR2XL U125 ( .A(n145), .B(wdtl[3]), .Y(n65) );
  NAND21X1 U126 ( .B(n35), .A(wdt_slow), .Y(n20) );
  INVX1 U127 ( .A(wdtrel[0]), .Y(n35) );
  AOI211X1 U128 ( .C(n145), .D(n142), .A(n63), .B(wdtl[1]), .Y(n52) );
  ENOX1 U129 ( .A(wdtl[5]), .B(n142), .C(wdt_slow), .D(wdtl[5]), .Y(n63) );
  INVX1 U130 ( .A(wdtl[6]), .Y(n142) );
  OAI22X1 U131 ( .A(n140), .B(n70), .C(n71), .D(n72), .Y(n128) );
  AOI21X1 U132 ( .B(n74), .C(n73), .A(wdt_tm_sync), .Y(n71) );
  XNOR2XL U133 ( .A(n58), .B(pres_8[1]), .Y(n74) );
  OAI21X1 U134 ( .B(n120), .C(n121), .A(n103), .Y(N116) );
  XNOR2XL U135 ( .A(pres_16[3]), .B(n116), .Y(n120) );
  OAI21X1 U136 ( .B(n124), .C(n121), .A(n103), .Y(N114) );
  XNOR2XL U137 ( .A(pres_16[1]), .B(pres_16[0]), .Y(n124) );
  OAI21X1 U138 ( .B(pres_16[0]), .C(n121), .A(n103), .Y(N113) );
  OAI31XL U139 ( .A(n96), .B(n138), .C(n139), .D(n97), .Y(N71) );
  OAI21X1 U140 ( .B(n98), .C(wdt_tm_sync), .A(n137), .Y(n97) );
  AND4X1 U141 ( .A(n139), .B(cycles_reg[2]), .C(n99), .D(n138), .Y(n98) );
  NAND21X1 U142 ( .B(wdt_slow), .A(n35), .Y(n36) );
  NOR2X1 U143 ( .A(n104), .B(wdtrefresh_sync), .Y(n99) );
  OAI211X1 U144 ( .C(n125), .D(n72), .A(n103), .B(n42), .Y(N112) );
  AOI21X1 U145 ( .B(n69), .C(pres_2), .A(wdtrefresh_sync), .Y(n125) );
  INVX1 U146 ( .A(wdth[2]), .Y(n34) );
  INVX1 U147 ( .A(wdth[0]), .Y(n26) );
  INVX1 U148 ( .A(cycles_reg[3]), .Y(n139) );
  INVX1 U149 ( .A(wdtl[7]), .Y(n37) );
  INVX1 U150 ( .A(wdth[1]), .Y(n30) );
  INVX1 U151 ( .A(wdtrel[6]), .Y(n39) );
  INVX1 U152 ( .A(n109), .Y(n21) );
  AOI211X1 U153 ( .C(n110), .D(n111), .A(n112), .B(resetff), .Y(n109) );
  NAND21X1 U154 ( .B(wdt_tm_sync), .A(n47), .Y(n19) );
  NOR32XL U155 ( .B(n18), .C(n10), .A(n100), .Y(N70) );
  XNOR2XL U156 ( .A(n138), .B(cycles_reg[2]), .Y(n100) );
  INVX1 U157 ( .A(n96), .Y(n10) );
  XNOR2XL U158 ( .A(wdtl[7]), .B(n145), .Y(n86) );
  NOR21XL U159 ( .B(N137), .A(n43), .Y(N173) );
  INVX1 U160 ( .A(resetff), .Y(n42) );
  NOR2X1 U161 ( .A(n114), .B(resetff), .Y(n112) );
  NAND2X1 U162 ( .A(wdt_act_sync), .B(n42), .Y(n72) );
  AO22X1 U163 ( .A(n112), .B(wdtrel[4]), .C(N134), .D(n110), .Y(N170) );
  AO22X1 U164 ( .A(n112), .B(wdtrel[3]), .C(N133), .D(n110), .Y(N169) );
  AO22X1 U165 ( .A(n112), .B(wdtrel[2]), .C(N132), .D(n110), .Y(N168) );
  AO22X1 U166 ( .A(n112), .B(wdtrel[1]), .C(N131), .D(n110), .Y(N167) );
  AO22X1 U167 ( .A(n112), .B(wdtrel[0]), .C(N130), .D(n110), .Y(N166) );
  NOR2X1 U168 ( .A(n72), .B(wdtrefresh_sync), .Y(n110) );
  AND3X1 U169 ( .A(wdth[3]), .B(wdth[1]), .C(wdth[0]), .Y(n87) );
  NOR2X1 U170 ( .A(wdtrefresh_sync), .B(resetff), .Y(n47) );
  OAI21X1 U171 ( .B(n102), .C(n96), .A(n103), .Y(N69) );
  XNOR2XL U172 ( .A(cycles_reg[1]), .B(cycles_reg[0]), .Y(n102) );
  OAI21X1 U173 ( .B(cycles_reg[0]), .C(n96), .A(n103), .Y(N68) );
  INVX1 U174 ( .A(wdtl[2]), .Y(n141) );
  NAND2X1 U175 ( .A(pres_16[1]), .B(pres_16[0]), .Y(n122) );
  INVX1 U176 ( .A(pres_8[0]), .Y(n58) );
  INVX1 U177 ( .A(pres_16[2]), .Y(n135) );
  INVX1 U178 ( .A(pres_8[1]), .Y(n140) );
  INVX1 U179 ( .A(wdtrefresh_sync), .Y(n114) );
  INVX1 U180 ( .A(wdts_s[0]), .Y(n136) );
  INVX1 U181 ( .A(wdt_tm_sync), .Y(n18) );
  INVX1 U182 ( .A(wdt_slow), .Y(n145) );
  NAND32XL U183 ( .B(sfraddr[4]), .C(sfraddr[6]), .A(sfrwe), .Y(n95) );
endmodule


module watchdog_a0_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module watchdog_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer1_a0 ( clkper, rst, newinstr, t1ff, t1ack, int1ff, t1_tf1, t1ov, 
        sfrdatai, sfraddr, sfrwe, t1_tmod, t1_tr1, tl1, th1 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t1_tmod;
  output [7:0] tl1;
  output [7:0] th1;
  input clkper, rst, newinstr, t1ff, t1ack, int1ff, sfrwe;
  output t1_tf1, t1ov, t1_tr1;
  wire   t1clr, th1_ov_ff, tl1_ov_ff, N31, N32, N33, N34, N35, N36, N37, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N95, N96, N97, N98, clk_ov12, N100, net12165,
         net12171, net12176, n20, n21, n23, n24, n27, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n46, n52, n53, n54, n55, n56, n57, n58, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n22, n25, n26, n28, n29, n30, n31, n32, n43, n44, n45,
         n47, n48, n49, n50, n51, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70;
  wire   [1:0] t0_mode;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer1_a0_0 clk_gate_t1_mode_reg ( .CLK(clkper), .EN(
        N31), .ENCLK(net12165), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_2 clk_gate_tl1_s_reg ( .CLK(clkper), .EN(N50), 
        .ENCLK(net12171), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_1 clk_gate_th1_s_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12176), .TE(1'b0) );
  timer1_a0_DW01_inc_0 add_278 ( .A(th1), .SUM({N75, N74, N73, N72, N71, N70, 
        N69, N68}) );
  timer1_a0_DW01_inc_1 add_244 ( .A(tl1), .SUM({N49, N48, N47, N46, N45, N44, 
        N43, N42}) );
  DFFQX1 clk_count_reg_1_ ( .D(N96), .C(clkper), .Q(clk_count[1]) );
  DFFQX1 th1_ov_ff_reg ( .D(n55), .C(clkper), .Q(th1_ov_ff) );
  DFFQX1 clk_count_reg_2_ ( .D(N97), .C(clkper), .Q(clk_count[2]) );
  DFFQX1 clk_count_reg_0_ ( .D(N95), .C(clkper), .Q(clk_count[0]) );
  DFFQX1 clk_count_reg_3_ ( .D(N98), .C(clkper), .Q(clk_count[3]) );
  DFFQX1 tl1_ov_ff_reg ( .D(n56), .C(clkper), .Q(tl1_ov_ff) );
  DFFQX1 t1clr_reg ( .D(n57), .C(clkper), .Q(t1clr) );
  DFFQX1 clk_ov12_reg ( .D(N100), .C(clkper), .Q(clk_ov12) );
  DFFQX1 t0_mode_reg_1_ ( .D(N37), .C(net12165), .Q(t0_mode[1]) );
  DFFQX1 t0_mode_reg_0_ ( .D(N36), .C(net12165), .Q(t0_mode[0]) );
  DFFQX1 tl1_s_reg_7_ ( .D(N58), .C(net12171), .Q(tl1[7]) );
  DFFQX1 tl1_s_reg_6_ ( .D(N57), .C(net12171), .Q(tl1[6]) );
  DFFQX1 t1_gate_reg ( .D(N32), .C(net12165), .Q(t1_tmod[3]) );
  DFFQX1 t1_ct_reg ( .D(N33), .C(net12165), .Q(t1_tmod[2]) );
  DFFQX1 tl1_s_reg_5_ ( .D(N56), .C(net12171), .Q(tl1[5]) );
  DFFQX1 th1_s_reg_7_ ( .D(N84), .C(net12176), .Q(th1[7]) );
  DFFQX1 th1_s_reg_6_ ( .D(N83), .C(net12176), .Q(th1[6]) );
  DFFQX1 th1_s_reg_5_ ( .D(N82), .C(net12176), .Q(th1[5]) );
  DFFQX1 th1_s_reg_4_ ( .D(N81), .C(net12176), .Q(th1[4]) );
  DFFQX1 t1_mode_reg_0_ ( .D(N34), .C(net12165), .Q(t1_tmod[0]) );
  DFFQX1 tl1_s_reg_4_ ( .D(N55), .C(net12171), .Q(tl1[4]) );
  DFFQX1 t1_mode_reg_1_ ( .D(N35), .C(net12165), .Q(t1_tmod[1]) );
  DFFQX1 tl1_s_reg_3_ ( .D(N54), .C(net12171), .Q(tl1[3]) );
  DFFQX1 th1_s_reg_3_ ( .D(N80), .C(net12176), .Q(th1[3]) );
  DFFQX1 t1_tr1_s_reg ( .D(n58), .C(clkper), .Q(t1_tr1) );
  DFFQX1 t1_tf1_s_reg ( .D(n54), .C(clkper), .Q(t1_tf1) );
  DFFQX1 tl1_s_reg_2_ ( .D(N53), .C(net12171), .Q(tl1[2]) );
  DFFQX1 tl1_s_reg_0_ ( .D(N51), .C(net12171), .Q(tl1[0]) );
  DFFQX1 th1_s_reg_2_ ( .D(N79), .C(net12176), .Q(th1[2]) );
  DFFQX1 th1_s_reg_0_ ( .D(N77), .C(net12176), .Q(th1[0]) );
  DFFQX1 tl1_s_reg_1_ ( .D(N52), .C(net12171), .Q(tl1[1]) );
  DFFQX1 th1_s_reg_1_ ( .D(N78), .C(net12176), .Q(th1[1]) );
  AND2X1 U3 ( .A(n5), .B(n9), .Y(N32) );
  INVX1 U4 ( .A(n39), .Y(n45) );
  NAND31X1 U5 ( .C(sfraddr[0]), .A(n1), .B(n33), .Y(n20) );
  INVX1 U6 ( .A(n52), .Y(n9) );
  INVX1 U7 ( .A(n31), .Y(n66) );
  NAND21X1 U8 ( .B(n46), .A(n7), .Y(n31) );
  NOR2X1 U9 ( .A(n2), .B(n52), .Y(N36) );
  NOR2X1 U10 ( .A(n4), .B(n52), .Y(N37) );
  NAND2X1 U11 ( .A(n7), .B(n52), .Y(N31) );
  NAND21X1 U12 ( .B(n41), .A(n7), .Y(n39) );
  INVX1 U13 ( .A(n6), .Y(n5) );
  INVX1 U14 ( .A(n4), .Y(n3) );
  NOR21XL U15 ( .B(n42), .A(sfraddr[2]), .Y(n33) );
  AND3XL U16 ( .A(sfrwe), .B(sfraddr[3]), .C(n53), .Y(n42) );
  NOR3XL U17 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n53) );
  INVX1 U18 ( .A(n22), .Y(n28) );
  NAND21X1 U19 ( .B(rst), .A(n46), .Y(n22) );
  NAND3X1 U20 ( .A(sfraddr[0]), .B(n33), .C(sfraddr[1]), .Y(n46) );
  NAND42X1 U21 ( .C(sfraddr[1]), .D(rst), .A(n33), .B(sfraddr[0]), .Y(n52) );
  OR4X1 U22 ( .A(n68), .B(n67), .C(n66), .D(rst), .Y(N50) );
  NAND4X1 U23 ( .A(sfraddr[2]), .B(sfraddr[0]), .C(n42), .D(n1), .Y(n41) );
  INVX1 U24 ( .A(n40), .Y(n44) );
  INVX1 U25 ( .A(n25), .Y(n67) );
  NAND21X1 U26 ( .B(n26), .A(n28), .Y(n25) );
  AND2X1 U27 ( .A(sfrdatai[6]), .B(n9), .Y(N33) );
  AND2X1 U28 ( .A(sfrdatai[4]), .B(n9), .Y(N34) );
  AND2X1 U29 ( .A(sfrdatai[5]), .B(n9), .Y(N35) );
  NAND3X1 U30 ( .A(n39), .B(n7), .C(n40), .Y(N76) );
  INVX1 U31 ( .A(sfrdatai[1]), .Y(n4) );
  INVX1 U32 ( .A(sfrdatai[7]), .Y(n6) );
  INVX1 U33 ( .A(sfraddr[1]), .Y(n1) );
  INVX1 U34 ( .A(sfrdatai[0]), .Y(n2) );
  INVX1 U35 ( .A(t1ov), .Y(n61) );
  INVX1 U36 ( .A(n26), .Y(n49) );
  INVX1 U37 ( .A(rst), .Y(n7) );
  INVX1 U38 ( .A(n30), .Y(n68) );
  NAND32X1 U39 ( .B(n49), .C(n29), .A(n28), .Y(n30) );
  AO22X1 U40 ( .A(sfrdatai[6]), .B(n45), .C(N74), .D(n44), .Y(N83) );
  AO22X1 U41 ( .A(sfrdatai[5]), .B(n45), .C(N73), .D(n44), .Y(N82) );
  AO22X1 U42 ( .A(sfrdatai[4]), .B(n45), .C(N72), .D(n44), .Y(N81) );
  AO22X1 U43 ( .A(sfrdatai[3]), .B(n45), .C(N71), .D(n44), .Y(N80) );
  AO22X1 U44 ( .A(sfrdatai[2]), .B(n45), .C(N70), .D(n44), .Y(N79) );
  AO22X1 U45 ( .A(n45), .B(n3), .C(N69), .D(n44), .Y(N78) );
  NAND3X1 U46 ( .A(n24), .B(n20), .C(n23), .Y(n21) );
  NAND31X1 U47 ( .C(rst), .A(n41), .B(n47), .Y(n40) );
  NAND21X1 U48 ( .B(newinstr), .A(n7), .Y(n27) );
  OAI22X1 U49 ( .A(rst), .B(n50), .C(n27), .D(n60), .Y(n55) );
  NAND21X1 U50 ( .B(n49), .A(n50), .Y(t1ov) );
  INVX1 U51 ( .A(n51), .Y(n32) );
  INVX1 U52 ( .A(n24), .Y(n12) );
  NAND21X1 U53 ( .B(n19), .A(n32), .Y(n26) );
  NAND2X1 U54 ( .A(n38), .B(n7), .Y(n36) );
  NOR2X1 U55 ( .A(rst), .B(n38), .Y(N100) );
  AO222X1 U56 ( .A(n67), .B(th1[0]), .C(N42), .D(n68), .E(n66), .F(sfrdatai[0]), .Y(N51) );
  AO222X1 U57 ( .A(n67), .B(th1[7]), .C(N49), .D(n68), .E(n66), .F(n5), .Y(N58) );
  AO222X1 U58 ( .A(n67), .B(th1[6]), .C(N48), .D(n68), .E(sfrdatai[6]), .F(n66), .Y(N57) );
  AO222X1 U59 ( .A(n67), .B(th1[5]), .C(N47), .D(n68), .E(sfrdatai[5]), .F(n66), .Y(N56) );
  AO222X1 U60 ( .A(n67), .B(th1[4]), .C(N46), .D(n68), .E(sfrdatai[4]), .F(n66), .Y(N55) );
  AO222X1 U61 ( .A(n67), .B(th1[3]), .C(N45), .D(n68), .E(sfrdatai[3]), .F(n66), .Y(N54) );
  AO222X1 U62 ( .A(n67), .B(th1[2]), .C(N44), .D(n68), .E(sfrdatai[2]), .F(n66), .Y(N53) );
  AO222X1 U63 ( .A(n67), .B(th1[1]), .C(N43), .D(n68), .E(n66), .F(n3), .Y(N52) );
  MUX2X1 U64 ( .D0(n65), .D1(t1_tf1), .S(n64), .Y(n54) );
  OAI31XL U65 ( .A(n20), .B(rst), .C(n6), .D(n21), .Y(n65) );
  AND3X1 U66 ( .A(n23), .B(n20), .C(n63), .Y(n64) );
  AO21X1 U67 ( .B(n62), .C(n61), .A(n21), .Y(n63) );
  AO22X1 U68 ( .A(n5), .B(n45), .C(N75), .D(n44), .Y(N84) );
  AO22X1 U69 ( .A(n45), .B(sfrdatai[0]), .C(N68), .D(n44), .Y(N77) );
  AND2X1 U70 ( .A(n8), .B(n7), .Y(n58) );
  MUX2X1 U71 ( .D0(sfrdatai[6]), .D1(t1_tr1), .S(n20), .Y(n8) );
  AO22AXL U72 ( .A(t1ack), .B(n7), .C(t1clr), .D(n27), .Y(n57) );
  OAI22AX1 U73 ( .D(tl1_ov_ff), .C(n27), .A(rst), .B(n51), .Y(n56) );
  NAND43X1 U74 ( .B(n29), .C(n18), .D(n17), .A(n16), .Y(n51) );
  AND4X1 U75 ( .A(tl1[1]), .B(tl1[0]), .C(tl1[3]), .D(tl1[2]), .Y(n16) );
  INVX1 U76 ( .A(tl1[4]), .Y(n18) );
  AOI32X1 U77 ( .A(tl1[6]), .B(tl1[5]), .C(tl1[7]), .D(n19), .E(n15), .Y(n17)
         );
  NAND6XL U78 ( .A(th1[0]), .B(th1[1]), .C(th1[2]), .D(th1[3]), .E(th1[4]), 
        .F(n48), .Y(n50) );
  AND4X1 U79 ( .A(th1[5]), .B(th1[6]), .C(th1[7]), .D(n47), .Y(n48) );
  NAND2X1 U80 ( .A(t0_mode[1]), .B(t0_mode[0]), .Y(n24) );
  OAI211X1 U81 ( .C(n19), .D(n15), .A(n14), .B(n13), .Y(n29) );
  OA21X1 U82 ( .B(int1ff), .C(n10), .A(clk_ov12), .Y(n14) );
  OA21X1 U83 ( .B(t1_tr1), .C(n12), .A(n11), .Y(n13) );
  INVX1 U84 ( .A(t1_tmod[3]), .Y(n10) );
  INVX1 U85 ( .A(n43), .Y(n47) );
  NAND21X1 U86 ( .B(t1_tmod[1]), .A(n32), .Y(n43) );
  NOR3XL U87 ( .A(rst), .B(t1clr), .C(t1ack), .Y(n23) );
  INVX1 U88 ( .A(t1_tmod[1]), .Y(n19) );
  INVX1 U89 ( .A(t1_tmod[0]), .Y(n15) );
  INVX1 U90 ( .A(t1_tmod[2]), .Y(n11) );
  NAND31X1 U91 ( .C(n36), .A(clk_count[1]), .B(clk_count[0]), .Y(n34) );
  AOI21BBXL U92 ( .B(clk_count[1]), .C(n36), .A(N95), .Y(n35) );
  OAI32X1 U93 ( .A(n69), .B(clk_count[3]), .C(n34), .D(n35), .E(n70), .Y(N98)
         );
  INVX1 U94 ( .A(clk_count[3]), .Y(n70) );
  NOR2X1 U95 ( .A(n36), .B(clk_count[0]), .Y(N95) );
  OAI22X1 U96 ( .A(n35), .B(n69), .C(clk_count[2]), .D(n34), .Y(N97) );
  MUX2X1 U97 ( .D0(n60), .D1(n59), .S(t1_tmod[1]), .Y(n62) );
  NAND21X1 U98 ( .B(t1_tmod[0]), .A(tl1_ov_ff), .Y(n59) );
  NAND4X1 U99 ( .A(clk_count[3]), .B(clk_count[1]), .C(clk_count[0]), .D(n69), 
        .Y(n38) );
  INVX1 U100 ( .A(clk_count[2]), .Y(n69) );
  NOR2X1 U101 ( .A(n37), .B(n36), .Y(N96) );
  XNOR2XL U102 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n37) );
  INVX1 U103 ( .A(th1_ov_ff), .Y(n60) );
endmodule


module timer1_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module timer1_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer0_a0 ( clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, t0_tf0, 
        t0_tf1, sfrdatai, sfraddr, sfrwe, t0_tmod, t0_tr0, t0_tr1, tl0, th0 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t0_tmod;
  output [7:0] tl0;
  output [7:0] th0;
  input clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, sfrwe;
  output t0_tf0, t0_tf1, t0_tr0, t0_tr1;
  wire   t0clr, th0_ov_ff, tl0_ov_ff, t1clr, N39, N40, N41, N42, N43, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N101, N102, N103, N104, clk_ov12, N106, net12193,
         net12199, net12204, n26, n27, n30, n39, n45, n47, n48, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n28, n29, n31, n32, n33,
         n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n46, n49, n50, n51,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer0_a0_0 clk_gate_t0_ct_reg ( .CLK(clkper), .EN(N39), 
        .ENCLK(net12193), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_2 clk_gate_th0_s_reg ( .CLK(clkper), .EN(N55), 
        .ENCLK(net12199), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_1 clk_gate_tl0_s_reg ( .CLK(clkper), .EN(N79), 
        .ENCLK(net12204), .TE(1'b0) );
  timer0_a0_DW01_inc_0 add_347 ( .A(tl0), .SUM({N78, N77, N76, N75, N74, N73, 
        N72, N71}) );
  timer0_a0_DW01_inc_1 add_309 ( .A(th0), .SUM({N54, N53, N52, N51, N50, N49, 
        N48, N47}) );
  DFFQX1 t1clr_reg ( .D(n63), .C(clkper), .Q(t1clr) );
  DFFQX1 clk_count_reg_1_ ( .D(N102), .C(clkper), .Q(clk_count[1]) );
  DFFQX1 clk_count_reg_2_ ( .D(N103), .C(clkper), .Q(clk_count[2]) );
  DFFQX1 clk_count_reg_0_ ( .D(N101), .C(clkper), .Q(clk_count[0]) );
  DFFQX1 t0clr_reg ( .D(n65), .C(clkper), .Q(t0clr) );
  DFFQX1 tl0_ov_ff_reg ( .D(n64), .C(clkper), .Q(tl0_ov_ff) );
  DFFQX1 th0_ov_ff_reg ( .D(n61), .C(clkper), .Q(th0_ov_ff) );
  DFFQX1 clk_count_reg_3_ ( .D(N104), .C(clkper), .Q(clk_count[3]) );
  DFFQX1 clk_ov12_reg ( .D(N106), .C(clkper), .Q(clk_ov12) );
  DFFQX1 tl0_s_reg_7_ ( .D(N87), .C(net12204), .Q(tl0[7]) );
  DFFQX1 tl0_s_reg_6_ ( .D(N86), .C(net12204), .Q(tl0[6]) );
  DFFQX1 th0_s_reg_7_ ( .D(N63), .C(net12199), .Q(th0[7]) );
  DFFQX1 tl0_s_reg_5_ ( .D(N85), .C(net12204), .Q(tl0[5]) );
  DFFQX1 th0_s_reg_5_ ( .D(N61), .C(net12199), .Q(th0[5]) );
  DFFQX1 th0_s_reg_6_ ( .D(N62), .C(net12199), .Q(th0[6]) );
  DFFQX1 th0_s_reg_4_ ( .D(N60), .C(net12199), .Q(th0[4]) );
  DFFQX1 tl0_s_reg_4_ ( .D(N84), .C(net12204), .Q(tl0[4]) );
  DFFQX1 t0_gate_reg ( .D(N40), .C(net12193), .Q(t0_tmod[3]) );
  DFFQX1 th0_s_reg_3_ ( .D(N59), .C(net12199), .Q(th0[3]) );
  DFFQX1 tl0_s_reg_3_ ( .D(N83), .C(net12204), .Q(tl0[3]) );
  DFFQX1 t0_tf0_s_reg ( .D(n60), .C(clkper), .Q(t0_tf0) );
  DFFQX1 t0_tr0_s_reg ( .D(n67), .C(clkper), .Q(t0_tr0) );
  DFFQX1 t0_tr1_s_reg ( .D(n66), .C(clkper), .Q(t0_tr1) );
  DFFQX1 t0_tf1_s_reg ( .D(n62), .C(clkper), .Q(t0_tf1) );
  DFFQX1 t0_ct_reg ( .D(N41), .C(net12193), .Q(t0_tmod[2]) );
  DFFQX1 tl0_s_reg_2_ ( .D(N82), .C(net12204), .Q(tl0[2]) );
  DFFQX1 th0_s_reg_2_ ( .D(N58), .C(net12199), .Q(th0[2]) );
  DFFQX1 th0_s_reg_1_ ( .D(N57), .C(net12199), .Q(th0[1]) );
  DFFQX1 th0_s_reg_0_ ( .D(N56), .C(net12199), .Q(th0[0]) );
  DFFQX1 tl0_s_reg_0_ ( .D(N80), .C(net12204), .Q(tl0[0]) );
  DFFQX1 t0_mode_reg_0_ ( .D(N42), .C(net12193), .Q(t0_tmod[0]) );
  DFFQX1 t0_mode_reg_1_ ( .D(N43), .C(net12193), .Q(t0_tmod[1]) );
  DFFQX1 tl0_s_reg_1_ ( .D(N81), .C(net12204), .Q(tl0[1]) );
  OR2X1 U3 ( .A(t1clr), .B(t1ack), .Y(n1) );
  NAND21X1 U4 ( .B(n14), .A(n74), .Y(n69) );
  NAND21X1 U5 ( .B(n26), .A(n13), .Y(n74) );
  INVX1 U6 ( .A(n26), .Y(n40) );
  INVX1 U7 ( .A(n47), .Y(n38) );
  INVX1 U8 ( .A(n14), .Y(n13) );
  NAND21X1 U9 ( .B(n14), .A(n45), .Y(n31) );
  NAND3X1 U10 ( .A(n3), .B(n4), .C(n39), .Y(n26) );
  INVX1 U11 ( .A(n53), .Y(n17) );
  INVX1 U12 ( .A(n29), .Y(n77) );
  NAND21X1 U13 ( .B(n45), .A(n13), .Y(n29) );
  NAND2X1 U14 ( .A(n13), .B(n53), .Y(N39) );
  NAND21X1 U15 ( .B(n48), .A(n13), .Y(n47) );
  INVX1 U16 ( .A(sfraddr[0]), .Y(n3) );
  INVX1 U17 ( .A(n12), .Y(n11) );
  INVX1 U18 ( .A(n10), .Y(n9) );
  INVX1 U19 ( .A(n8), .Y(n7) );
  INVX1 U20 ( .A(n6), .Y(n5) );
  INVX1 U21 ( .A(n16), .Y(n14) );
  INVX1 U22 ( .A(n16), .Y(n15) );
  NOR21XL U23 ( .B(n52), .A(sfraddr[2]), .Y(n39) );
  AND3XL U24 ( .A(sfrwe), .B(sfraddr[3]), .C(n54), .Y(n52) );
  NOR3XL U25 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n54) );
  NAND3X1 U26 ( .A(n39), .B(n3), .C(sfraddr[1]), .Y(n45) );
  NAND42X1 U27 ( .C(sfraddr[1]), .D(n14), .A(n39), .B(sfraddr[0]), .Y(n53) );
  INVX1 U28 ( .A(n28), .Y(n76) );
  NAND21X1 U29 ( .B(n31), .A(n33), .Y(n28) );
  OR4X1 U30 ( .A(n77), .B(n76), .C(n2), .D(n15), .Y(N79) );
  AND2X1 U31 ( .A(sfrdatai[3]), .B(n17), .Y(N40) );
  AND2X1 U32 ( .A(sfrdatai[0]), .B(n17), .Y(N42) );
  AND2X1 U33 ( .A(sfrdatai[1]), .B(n17), .Y(N43) );
  AND2X1 U34 ( .A(sfrdatai[2]), .B(n17), .Y(N41) );
  NAND32X1 U35 ( .B(n75), .C(n15), .A(n47), .Y(N55) );
  NAND4X1 U36 ( .A(sfraddr[2]), .B(n52), .C(n3), .D(n4), .Y(n48) );
  INVX1 U37 ( .A(sfraddr[1]), .Y(n4) );
  INVX1 U38 ( .A(sfrdatai[6]), .Y(n10) );
  INVX1 U39 ( .A(sfrdatai[4]), .Y(n6) );
  INVX1 U40 ( .A(sfrdatai[7]), .Y(n12) );
  INVX1 U41 ( .A(sfrdatai[5]), .Y(n8) );
  INVX1 U42 ( .A(rst), .Y(n16) );
  INVX1 U43 ( .A(t0ack), .Y(n78) );
  NOR3XL U44 ( .A(n33), .B(n32), .C(n31), .Y(n2) );
  OAI22X1 U45 ( .A(n19), .B(n69), .C(n74), .D(n6), .Y(n67) );
  AO22X1 U46 ( .A(N53), .B(n75), .C(n9), .D(n38), .Y(N62) );
  AO22X1 U47 ( .A(N52), .B(n75), .C(n7), .D(n38), .Y(N61) );
  AO22X1 U48 ( .A(N51), .B(n75), .C(n5), .D(n38), .Y(N60) );
  AO22X1 U49 ( .A(N50), .B(n75), .C(sfrdatai[3]), .D(n38), .Y(N59) );
  AO22X1 U50 ( .A(N49), .B(n75), .C(sfrdatai[2]), .D(n38), .Y(N58) );
  AO22X1 U51 ( .A(N48), .B(n75), .C(sfrdatai[1]), .D(n38), .Y(N57) );
  INVX1 U52 ( .A(n37), .Y(n75) );
  NAND32X1 U53 ( .B(n15), .C(n36), .A(n41), .Y(n37) );
  INVX1 U54 ( .A(n48), .Y(n36) );
  NAND21X1 U55 ( .B(newinstr), .A(n13), .Y(n30) );
  OAI22X1 U56 ( .A(n15), .B(n78), .C(n30), .D(n79), .Y(n65) );
  INVX1 U57 ( .A(n49), .Y(n43) );
  INVX1 U58 ( .A(n25), .Y(n33) );
  NAND32X1 U59 ( .B(n50), .C(n24), .A(n23), .Y(n25) );
  NAND2X1 U60 ( .A(n55), .B(n13), .Y(n58) );
  NOR2X1 U61 ( .A(n15), .B(n55), .Y(N106) );
  AO222X1 U62 ( .A(n76), .B(th0[7]), .C(n77), .D(n11), .E(N78), .F(n2), .Y(N87) );
  AO222X1 U63 ( .A(n76), .B(th0[6]), .C(n77), .D(n9), .E(N77), .F(n2), .Y(N86)
         );
  AO222X1 U64 ( .A(n76), .B(th0[5]), .C(n77), .D(n7), .E(N76), .F(n2), .Y(N85)
         );
  AO222X1 U65 ( .A(n76), .B(th0[4]), .C(n5), .D(n77), .E(N75), .F(n2), .Y(N84)
         );
  AO222X1 U66 ( .A(n76), .B(th0[3]), .C(sfrdatai[3]), .D(n77), .E(N74), .F(n2), 
        .Y(N83) );
  AO222X1 U67 ( .A(n76), .B(th0[2]), .C(sfrdatai[2]), .D(n77), .E(N73), .F(n2), 
        .Y(N82) );
  AO222X1 U68 ( .A(n76), .B(th0[1]), .C(sfrdatai[1]), .D(n77), .E(N72), .F(n2), 
        .Y(N81) );
  AO222X1 U69 ( .A(n76), .B(th0[0]), .C(n77), .D(sfrdatai[0]), .E(N71), .F(n2), 
        .Y(N80) );
  OAI21X1 U70 ( .B(n74), .C(n8), .A(n73), .Y(n60) );
  AOI31X1 U71 ( .A(n27), .B(n26), .C(n72), .D(n71), .Y(n73) );
  NOR3XL U72 ( .A(n15), .B(t0clr), .C(t0ack), .Y(n27) );
  MUX2X1 U73 ( .D0(n68), .D1(n51), .S(t0_tmod[1]), .Y(n72) );
  AND4X1 U74 ( .A(t0_tf0), .B(n79), .C(n70), .D(n78), .Y(n71) );
  INVX1 U75 ( .A(n69), .Y(n70) );
  MUX2X1 U76 ( .D0(n46), .D1(t0_tf1), .S(n44), .Y(n62) );
  OAI32X1 U77 ( .A(n15), .B(n40), .C(n1), .D(n74), .E(n12), .Y(n46) );
  AOI211X1 U78 ( .C(n43), .D(t0_tmod[1]), .A(n69), .B(n1), .Y(n44) );
  OAI22AX1 U79 ( .D(t0_tr1), .C(n69), .A(n74), .B(n10), .Y(n66) );
  AO22X1 U80 ( .A(N54), .B(n75), .C(n11), .D(n38), .Y(N63) );
  AO22X1 U81 ( .A(N47), .B(n75), .C(sfrdatai[0]), .D(n38), .Y(N56) );
  AO22AXL U82 ( .A(t1ack), .B(n13), .C(t1clr), .D(n30), .Y(n63) );
  OAI22AX1 U83 ( .D(th0_ov_ff), .C(n30), .A(n15), .B(n49), .Y(n61) );
  OAI22AX1 U84 ( .D(tl0_ov_ff), .C(n30), .A(n15), .B(n50), .Y(n64) );
  NAND43X1 U85 ( .B(n32), .C(n22), .D(n21), .A(n20), .Y(n50) );
  AND4X1 U86 ( .A(tl0[1]), .B(tl0[0]), .C(tl0[3]), .D(tl0[2]), .Y(n20) );
  INVX1 U87 ( .A(tl0[4]), .Y(n22) );
  AOI32X1 U88 ( .A(tl0[6]), .B(tl0[5]), .C(tl0[7]), .D(n24), .E(n23), .Y(n21)
         );
  NAND42X1 U89 ( .C(t0_tmod[2]), .D(n19), .A(clk_ov12), .B(n18), .Y(n32) );
  NAND21X1 U90 ( .B(int0ff), .A(t0_tmod[3]), .Y(n18) );
  NAND6XL U91 ( .A(th0[1]), .B(th0[0]), .C(th0[2]), .D(th0[3]), .E(th0[4]), 
        .F(n42), .Y(n49) );
  AND4X1 U92 ( .A(th0[5]), .B(th0[6]), .C(th0[7]), .D(n41), .Y(n42) );
  NAND21X1 U93 ( .B(th0_ov_ff), .A(n49), .Y(n68) );
  INVX1 U94 ( .A(n35), .Y(n41) );
  MUX2BXL U95 ( .D0(n50), .D1(n34), .S(t0_tmod[1]), .Y(n35) );
  AND3X1 U96 ( .A(t0_tr1), .B(t0_tmod[0]), .C(clk_ov12), .Y(n34) );
  INVX1 U97 ( .A(t0_tmod[0]), .Y(n23) );
  INVX1 U98 ( .A(t0_tmod[1]), .Y(n24) );
  INVX1 U99 ( .A(t0_tr0), .Y(n19) );
  NAND31X1 U100 ( .C(n58), .A(clk_count[1]), .B(clk_count[0]), .Y(n56) );
  AOI21BBXL U101 ( .B(clk_count[1]), .C(n58), .A(N101), .Y(n57) );
  OAI32X1 U102 ( .A(n80), .B(clk_count[3]), .C(n56), .D(n57), .E(n81), .Y(N104) );
  INVX1 U103 ( .A(clk_count[3]), .Y(n81) );
  NOR2X1 U104 ( .A(n58), .B(clk_count[0]), .Y(N101) );
  OAI22X1 U105 ( .A(n57), .B(n80), .C(clk_count[2]), .D(n56), .Y(N103) );
  NAND21X1 U106 ( .B(tl0_ov_ff), .A(n50), .Y(n51) );
  NOR2X1 U107 ( .A(n59), .B(n58), .Y(N102) );
  XNOR2XL U108 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n59) );
  NAND4X1 U109 ( .A(clk_count[3]), .B(clk_count[1]), .C(clk_count[0]), .D(n80), 
        .Y(n55) );
  INVX1 U110 ( .A(clk_count[2]), .Y(n80) );
  INVX1 U111 ( .A(t0clr), .Y(n79) );
endmodule


module timer0_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module timer0_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module serial0_a0 ( t_shift_clk, r_shift_clk, clkper, rst, newinstr, rxd0ff, 
        t1ov, rxd0o, rxd0oe, txd0, sfrdatai, sfraddr, sfrwe, s0con, s0buf, 
        s0rell, s0relh, smod, bd );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] s0con;
  output [7:0] s0buf;
  output [7:0] s0rell;
  output [7:0] s0relh;
  input clkper, rst, newinstr, rxd0ff, t1ov, sfrwe;
  output t_shift_clk, r_shift_clk, rxd0o, rxd0oe, txd0, smod, bd;
  wire   r_clk_ov2, t1ov_ff, N59, ri_tmp, rxd0_val, s0con2_val, s0con2_tmp,
         ti_tmp, N108, N109, N110, N111, N112, N113, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, baud_rate_ov, N142, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N166, N169, N170, N185, N186, N187,
         N188, N190, clk_ov12, N191, r_start, baud_r_count, baud_r2_clk, N207,
         t_baud_ov, t_start, N223, N224, N225, N226, N227, N230, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N281,
         N282, N283, N284, N303, rxd0_fall, rxd0_ff, rxd0_fall_fl,
         receive_11_bits, N306, N307, N324, N325, N326, N327, N333, ri0_fall,
         ri0_ff, N348, N360, N361, N362, N363, N364, N375, N376, N377, N378,
         N379, N380, N381, N382, N424, N425, N426, N427, N428, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, net12232, net12238,
         net12243, net12248, net12253, net12258, net12263, net12268, net12273,
         net12278, net12283, n13, n92, n98, n102, n103, n104, n105, n108, n114,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n130, n131, n134, n135, n136, n137, n138, n140, n141, n142, n146,
         n149, n151, n152, n153, n155, n156, n157, n158, n159, n164, n165,
         n166, n167, n168, n169, n172, n173, n174, n175, n176, n177, n178,
         n179, n181, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n199, n200, n202, n203, n207,
         n208, n209, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97, n99,
         n100, n101, n106, n107, n109, n110, n111, n112, n113, n115, n127,
         n128, n129, n132, n133, n139, n143, n144, n145, n147, n148, n150,
         n154, n160, n161, n162, n163, n170, n171, n180, n182, n198, n201,
         n204, n205, n206, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294;
  wire   [3:0] r_baud_count;
  wire   [3:0] r_shift_count;
  wire   [3:0] t_shift_count;
  wire   [9:0] tim_baud;
  wire   [3:0] clk_count;
  wire   [3:0] t_baud_count;
  wire   [10:0] t_shift_reg;
  wire   [1:0] fluctuation_conter;
  wire   [2:0] rxd0_vec;
  wire   [7:0] r_shift_reg;

  MAJ3X1 U336 ( .A(rxd0_vec[1]), .B(rxd0_vec[0]), .C(rxd0_vec[2]), .Y(n172) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_0 clk_gate_s0con_s_reg ( .CLK(clkper), .EN(
        N108), .ENCLK(net12232), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_10 clk_gate_s0rell_s_reg ( .CLK(clkper), 
        .EN(N117), .ENCLK(net12238), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_9 clk_gate_s0relh_s_reg ( .CLK(clkper), .EN(
        N128), .ENCLK(net12243), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_8 clk_gate_tim_baud_reg ( .CLK(clkper), .EN(
        N166), .ENCLK(net12248), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_7 clk_gate_t_baud_count_reg ( .CLK(clkper), 
        .EN(N223), .ENCLK(net12253), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_6 clk_gate_t_shift_reg_reg ( .CLK(clkper), 
        .EN(N257), .ENCLK(net12258), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_5 clk_gate_rxd0_vec_reg ( .CLK(clkper), .EN(
        N324), .ENCLK(net12263), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_4 clk_gate_r_baud_count_reg ( .CLK(clkper), 
        .EN(N360), .ENCLK(net12268), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_3 clk_gate_r_shift_reg_reg ( .CLK(clkper), 
        .EN(n13), .ENCLK(net12273), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_2 clk_gate_r_shift_count_reg ( .CLK(clkper), 
        .EN(N428), .ENCLK(net12278), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_1 clk_gate_s0buf_r_reg ( .CLK(clkper), .EN(
        N471), .ENCLK(net12283), .TE(1'b0) );
  serial0_a0_DW01_inc_0 add_584 ( .A(tim_baud), .SUM({N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145}) );
  DFFQX1 t_shift_reg_reg_9_ ( .D(N267), .C(net12258), .Q(t_shift_reg[9]) );
  DFFQX1 t_shift_reg_reg_8_ ( .D(N266), .C(net12258), .Q(t_shift_reg[8]) );
  DFFQX1 t_shift_reg_reg_7_ ( .D(N265), .C(net12258), .Q(t_shift_reg[7]) );
  DFFQX1 t_shift_reg_reg_6_ ( .D(N264), .C(net12258), .Q(t_shift_reg[6]) );
  DFFQX1 t_shift_reg_reg_5_ ( .D(N263), .C(net12258), .Q(t_shift_reg[5]) );
  DFFQX1 t_shift_reg_reg_4_ ( .D(N262), .C(net12258), .Q(t_shift_reg[4]) );
  DFFQX1 t_shift_reg_reg_3_ ( .D(N261), .C(net12258), .Q(t_shift_reg[3]) );
  DFFQX1 t_shift_reg_reg_10_ ( .D(N268), .C(net12258), .Q(t_shift_reg[10]) );
  DFFQX1 r_shift_reg_reg_0_ ( .D(N375), .C(net12273), .Q(r_shift_reg[0]) );
  DFFQX1 t_shift_reg_reg_1_ ( .D(N259), .C(net12258), .Q(t_shift_reg[1]) );
  DFFQX1 rxd0_vec_reg_2_ ( .D(N327), .C(net12263), .Q(rxd0_vec[2]) );
  DFFQX1 rxd0_vec_reg_1_ ( .D(N326), .C(net12263), .Q(rxd0_vec[1]) );
  DFFQX1 rxd0_ff_reg ( .D(N307), .C(clkper), .Q(rxd0_ff) );
  DFFQX1 t_shift_reg_reg_2_ ( .D(N260), .C(net12258), .Q(t_shift_reg[2]) );
  DFFQX1 rxd0_vec_reg_0_ ( .D(N325), .C(net12263), .Q(rxd0_vec[0]) );
  DFFQX1 s0con2_tmp_reg ( .D(n232), .C(clkper), .Q(s0con2_tmp) );
  DFFQX1 ri_tmp_reg ( .D(n238), .C(clkper), .Q(ri_tmp) );
  DFFQX1 baud_r_count_reg ( .D(n245), .C(clkper), .Q(baud_r_count) );
  DFFQX1 t_shift_reg_reg_0_ ( .D(N258), .C(net12258), .Q(t_shift_reg[0]) );
  DFFQX1 r_shift_reg_reg_7_ ( .D(N382), .C(net12273), .Q(r_shift_reg[7]) );
  DFFQX1 r_shift_reg_reg_6_ ( .D(N381), .C(net12273), .Q(r_shift_reg[6]) );
  DFFQX1 r_shift_reg_reg_5_ ( .D(N380), .C(net12273), .Q(r_shift_reg[5]) );
  DFFQX1 r_shift_reg_reg_4_ ( .D(N379), .C(net12273), .Q(r_shift_reg[4]) );
  DFFQX1 r_shift_reg_reg_3_ ( .D(N378), .C(net12273), .Q(r_shift_reg[3]) );
  DFFQX1 r_shift_reg_reg_2_ ( .D(N377), .C(net12273), .Q(r_shift_reg[2]) );
  DFFQX1 r_shift_reg_reg_1_ ( .D(N376), .C(net12273), .Q(r_shift_reg[1]) );
  DFFQX1 fluctuation_conter_reg_0_ ( .D(n234), .C(clkper), .Q(
        fluctuation_conter[0]) );
  DFFQX1 ti_tmp_reg ( .D(n242), .C(clkper), .Q(ti_tmp) );
  DFFQX1 ri0_ff_reg ( .D(N348), .C(clkper), .Q(ri0_ff) );
  DFFQX1 receive_11_bits_reg ( .D(n229), .C(clkper), .Q(receive_11_bits) );
  DFFQX1 fluctuation_conter_reg_1_ ( .D(n233), .C(clkper), .Q(
        fluctuation_conter[1]) );
  DFFQX1 s0con2_val_reg ( .D(n231), .C(net12263), .Q(s0con2_val) );
  DFFQX1 rxd0_fall_fl_reg ( .D(n235), .C(clkper), .Q(rxd0_fall_fl) );
  DFFQX1 t_shift_count_reg_3_ ( .D(N284), .C(net12258), .Q(t_shift_count[3])
         );
  DFFQX1 clk_count_reg_1_ ( .D(N186), .C(clkper), .Q(clk_count[1]) );
  DFFQX1 clk_count_reg_0_ ( .D(N185), .C(clkper), .Q(clk_count[0]) );
  DFFQX1 rxd0_val_reg ( .D(N333), .C(clkper), .Q(rxd0_val) );
  DFFQX1 clk_count_reg_3_ ( .D(N188), .C(clkper), .Q(clk_count[3]) );
  DFFQX1 clk_count_reg_2_ ( .D(N187), .C(clkper), .Q(clk_count[2]) );
  DFFQX1 t_shift_count_reg_1_ ( .D(N282), .C(net12258), .Q(t_shift_count[1])
         );
  DFFQX1 t_shift_count_reg_2_ ( .D(N283), .C(net12258), .Q(t_shift_count[2])
         );
  DFFQX1 t_shift_count_reg_0_ ( .D(N281), .C(net12258), .Q(t_shift_count[0])
         );
  DFFQX1 rxd0_fall_reg ( .D(N306), .C(clkper), .Q(rxd0_fall) );
  DFFQX1 baud_r2_clk_reg ( .D(N207), .C(clkper), .Q(baud_r2_clk) );
  DFFQX1 clk_ov12_reg ( .D(N191), .C(clkper), .Q(clk_ov12) );
  DFFQX1 t_baud_ov_reg ( .D(N230), .C(clkper), .Q(t_baud_ov) );
  DFFQX1 tim_baud_reg_3_ ( .D(N170), .C(net12248), .Q(tim_baud[3]) );
  DFFQX1 tim_baud_reg_4_ ( .D(n277), .C(net12248), .Q(tim_baud[4]) );
  DFFQX1 t_baud_count_reg_3_ ( .D(N227), .C(net12253), .Q(t_baud_count[3]) );
  DFFQX1 r_shift_count_reg_1_ ( .D(N425), .C(net12278), .Q(r_shift_count[1])
         );
  DFFQX1 r_shift_count_reg_3_ ( .D(N427), .C(net12278), .Q(r_shift_count[3])
         );
  DFFQX1 r_shift_count_reg_2_ ( .D(N426), .C(net12278), .Q(r_shift_count[2])
         );
  DFFQX1 ri0_fall_reg ( .D(n236), .C(clkper), .Q(ri0_fall) );
  DFFQX1 r_baud_count_reg_2_ ( .D(N363), .C(net12268), .Q(r_baud_count[2]) );
  DFFQX1 r_baud_count_reg_3_ ( .D(N364), .C(net12268), .Q(r_baud_count[3]) );
  DFFQX1 t_baud_count_reg_1_ ( .D(N225), .C(net12253), .Q(t_baud_count[1]) );
  DFFQX1 t_baud_count_reg_0_ ( .D(N224), .C(net12253), .Q(t_baud_count[0]) );
  DFFQX1 r_start_reg ( .D(n240), .C(clkper), .Q(r_start) );
  DFFQX1 t_baud_count_reg_2_ ( .D(N226), .C(net12253), .Q(t_baud_count[2]) );
  DFFQX1 t1ov_ff_reg ( .D(N59), .C(clkper), .Q(t1ov_ff) );
  DFFQX1 tim_baud_reg_2_ ( .D(N169), .C(net12248), .Q(tim_baud[2]) );
  DFFQX1 tim_baud_reg_7_ ( .D(n274), .C(net12248), .Q(tim_baud[7]) );
  DFFQX1 tim_baud_reg_5_ ( .D(n276), .C(net12248), .Q(tim_baud[5]) );
  DFFQX1 tim_baud_reg_1_ ( .D(n278), .C(net12248), .Q(tim_baud[1]) );
  DFFQX1 tim_baud_reg_6_ ( .D(n275), .C(net12248), .Q(tim_baud[6]) );
  DFFQX1 tim_baud_reg_0_ ( .D(n279), .C(net12248), .Q(tim_baud[0]) );
  DFFQX1 r_baud_count_reg_1_ ( .D(N362), .C(net12268), .Q(r_baud_count[1]) );
  DFFQX1 r_shift_count_reg_0_ ( .D(N424), .C(net12278), .Q(r_shift_count[0])
         );
  DFFQX1 tim_baud_reg_9_ ( .D(n281), .C(net12248), .Q(tim_baud[9]) );
  DFFQX1 tim_baud_reg_8_ ( .D(n280), .C(net12248), .Q(tim_baud[8]) );
  DFFQX1 r_baud_count_reg_0_ ( .D(N361), .C(net12268), .Q(r_baud_count[0]) );
  DFFQX1 r_clk_ov2_reg ( .D(N190), .C(clkper), .Q(r_clk_ov2) );
  DFFQX1 baud_rate_ov_reg ( .D(N142), .C(clkper), .Q(baud_rate_ov) );
  DFFQX1 s0rell_s_reg_7_ ( .D(N125), .C(net12238), .Q(s0rell[7]) );
  DFFQX1 s0relh_s_reg_6_ ( .D(N135), .C(net12243), .Q(s0relh[6]) );
  DFFQX1 s0buf_r_reg_7_ ( .D(N479), .C(net12283), .Q(s0buf[7]) );
  DFFQX1 s0buf_r_reg_6_ ( .D(N478), .C(net12283), .Q(s0buf[6]) );
  DFFQX1 s0relh_s_reg_5_ ( .D(N134), .C(net12243), .Q(s0relh[5]) );
  DFFQX1 smod_s_reg ( .D(n244), .C(clkper), .Q(smod) );
  DFFQX1 bd_s_reg ( .D(n271), .C(clkper), .Q(bd) );
  DFFQX1 s0relh_s_reg_7_ ( .D(N136), .C(net12243), .Q(s0relh[7]) );
  DFFQX1 s0buf_r_reg_5_ ( .D(N477), .C(net12283), .Q(s0buf[5]) );
  DFFQX1 s0relh_s_reg_4_ ( .D(N133), .C(net12243), .Q(s0relh[4]) );
  DFFQX1 s0rell_s_reg_6_ ( .D(N124), .C(net12238), .Q(s0rell[6]) );
  DFFQX1 s0rell_s_reg_5_ ( .D(N123), .C(net12238), .Q(s0rell[5]) );
  DFFQX1 s0con_s_reg_5_ ( .D(N111), .C(net12232), .Q(s0con[5]) );
  DFFQX1 s0buf_r_reg_4_ ( .D(N476), .C(net12283), .Q(s0buf[4]) );
  DFFQX1 s0rell_s_reg_4_ ( .D(N122), .C(net12238), .Q(s0rell[4]) );
  DFFQX1 s0con_s_reg_4_ ( .D(N110), .C(net12232), .Q(s0con[4]) );
  DFFQX1 s0rell_s_reg_3_ ( .D(N121), .C(net12238), .Q(s0rell[3]) );
  DFFQX1 s0relh_s_reg_3_ ( .D(N132), .C(net12243), .Q(s0relh[3]) );
  DFFQX1 s0buf_r_reg_3_ ( .D(N475), .C(net12283), .Q(s0buf[3]) );
  DFFQX1 s0con_s_reg_3_ ( .D(N109), .C(net12232), .Q(s0con[3]) );
  DFFQX1 rxd0o_reg ( .D(N303), .C(clkper), .Q(rxd0o) );
  DFFQX1 t_start_reg ( .D(n243), .C(clkper), .Q(t_start) );
  DFFQX1 txd0_reg ( .D(n239), .C(clkper), .Q(txd0) );
  DFFQX1 s0con_s_reg_6_ ( .D(N112), .C(net12232), .Q(s0con[6]) );
  DFFQX1 s0con_s_reg_7_ ( .D(N113), .C(net12232), .Q(s0con[7]) );
  DFFQX1 s0relh_s_reg_2_ ( .D(N131), .C(net12243), .Q(s0relh[2]) );
  DFFQX1 s0buf_r_reg_2_ ( .D(N474), .C(net12283), .Q(s0buf[2]) );
  DFFQX1 s0rell_s_reg_0_ ( .D(N118), .C(net12238), .Q(s0rell[0]) );
  DFFQX1 s0rell_s_reg_1_ ( .D(N119), .C(net12238), .Q(s0rell[1]) );
  DFFQX1 s0rell_s_reg_2_ ( .D(N120), .C(net12238), .Q(s0rell[2]) );
  DFFQX1 s0buf_r_reg_0_ ( .D(N472), .C(net12283), .Q(s0buf[0]) );
  DFFQX1 s0relh_s_reg_0_ ( .D(N129), .C(net12243), .Q(s0relh[0]) );
  DFFQX1 s0con_s_reg_0_ ( .D(n237), .C(clkper), .Q(s0con[0]) );
  DFFQX1 s0buf_r_reg_1_ ( .D(N473), .C(net12283), .Q(s0buf[1]) );
  DFFQX1 s0relh_s_reg_1_ ( .D(N130), .C(net12243), .Q(s0relh[1]) );
  DFFQX1 s0con_s_reg_2_ ( .D(n230), .C(clkper), .Q(s0con[2]) );
  DFFQX1 s0con_s_reg_1_ ( .D(n241), .C(clkper), .Q(s0con[1]) );
  NOR32XL U3 ( .B(tim_baud[4]), .C(tim_baud[3]), .A(n225), .Y(n224) );
  NAND21XL U4 ( .B(n60), .A(sfraddr[4]), .Y(n226) );
  OR2XL U5 ( .A(sfraddr[4]), .B(n60), .Y(n228) );
  BUFX3 U6 ( .A(n8), .Y(n1) );
  INVX1 U7 ( .A(n258), .Y(n2) );
  NOR41XL U8 ( .D(r_shift_count[0]), .A(r_shift_count[1]), .B(r_shift_count[2]), .C(r_shift_count[3]), .Y(n98) );
  INVX1 U9 ( .A(N108), .Y(n148) );
  NAND21X1 U10 ( .B(n37), .A(n115), .Y(N108) );
  INVX1 U11 ( .A(n115), .Y(n162) );
  INVX1 U12 ( .A(n49), .Y(n36) );
  INVX1 U13 ( .A(n48), .Y(n37) );
  INVX1 U14 ( .A(n49), .Y(n38) );
  INVX1 U15 ( .A(n48), .Y(n39) );
  INVX1 U16 ( .A(n49), .Y(n40) );
  NAND21X1 U17 ( .B(n134), .A(n42), .Y(n115) );
  NAND21X1 U18 ( .B(n37), .A(n134), .Y(n150) );
  AO21X1 U19 ( .B(n96), .C(n22), .A(n39), .Y(N129) );
  AO21X1 U20 ( .B(n96), .C(n24), .A(n40), .Y(N130) );
  AO21X1 U21 ( .B(n162), .C(n34), .A(n55), .Y(N112) );
  INVX1 U22 ( .A(n226), .Y(n96) );
  AND2X1 U23 ( .A(n162), .B(n28), .Y(N109) );
  AND2X1 U24 ( .A(n162), .B(n30), .Y(N110) );
  AND2X1 U25 ( .A(n162), .B(n32), .Y(N111) );
  AO21X1 U26 ( .B(n93), .C(n22), .A(n39), .Y(N118) );
  AO21X1 U27 ( .B(n93), .C(n28), .A(n39), .Y(N121) );
  AO21X1 U28 ( .B(n93), .C(n30), .A(n40), .Y(N122) );
  AO21X1 U29 ( .B(n93), .C(n34), .A(n40), .Y(N124) );
  INVX1 U30 ( .A(n228), .Y(n93) );
  AND2X1 U31 ( .A(n96), .B(n26), .Y(N131) );
  AND2X1 U32 ( .A(n96), .B(n28), .Y(N132) );
  AND2X1 U33 ( .A(n96), .B(n30), .Y(N133) );
  AND2X1 U34 ( .A(n96), .B(n32), .Y(N134) );
  AND2X1 U35 ( .A(n96), .B(n34), .Y(N135) );
  AND2X1 U36 ( .A(n93), .B(n24), .Y(N119) );
  AND2X1 U37 ( .A(n93), .B(n26), .Y(N120) );
  AND2X1 U38 ( .A(n93), .B(n32), .Y(N123) );
  INVX1 U39 ( .A(n181), .Y(n267) );
  NAND2X1 U40 ( .A(n44), .B(n226), .Y(N128) );
  NAND2X1 U41 ( .A(n45), .B(n228), .Y(N117) );
  INVX1 U42 ( .A(n54), .Y(n48) );
  INVX1 U43 ( .A(n54), .Y(n49) );
  INVX1 U44 ( .A(n57), .Y(n41) );
  INVX1 U45 ( .A(n53), .Y(n50) );
  INVX1 U46 ( .A(n56), .Y(n43) );
  INVX1 U47 ( .A(n56), .Y(n42) );
  INVX1 U48 ( .A(n53), .Y(n51) );
  INVX1 U49 ( .A(n55), .Y(n45) );
  INVX1 U50 ( .A(n55), .Y(n44) );
  INVX1 U51 ( .A(n55), .Y(n46) );
  INVX1 U52 ( .A(n54), .Y(n47) );
  INVX1 U53 ( .A(n53), .Y(n52) );
  NOR32XL U54 ( .B(n227), .C(sfraddr[4]), .A(sfraddr[5]), .Y(n146) );
  NAND3X1 U55 ( .A(n140), .B(n227), .C(sfraddr[5]), .Y(n60) );
  NOR2X1 U56 ( .A(n193), .B(n36), .Y(n181) );
  INVX1 U57 ( .A(n176), .Y(n270) );
  NAND3X1 U58 ( .A(n267), .B(n50), .C(n176), .Y(N257) );
  INVX1 U59 ( .A(n176), .Y(n211) );
  INVX1 U60 ( .A(n27), .Y(n26) );
  INVX1 U61 ( .A(n25), .Y(n24) );
  NOR3XL U62 ( .A(n38), .B(sfraddr[6]), .C(n20), .Y(n140) );
  INVX1 U63 ( .A(n33), .Y(n32) );
  INVX1 U64 ( .A(n29), .Y(n28) );
  INVX1 U65 ( .A(n31), .Y(n30) );
  INVX1 U66 ( .A(n35), .Y(n34) );
  INVX1 U67 ( .A(n23), .Y(n22) );
  INVX1 U68 ( .A(n59), .Y(n54) );
  INVX1 U69 ( .A(n58), .Y(n56) );
  INVX1 U70 ( .A(n59), .Y(n53) );
  INVX1 U71 ( .A(n58), .Y(n57) );
  INVX1 U72 ( .A(n58), .Y(n55) );
  INVX1 U73 ( .A(sfrwe), .Y(n272) );
  NOR4XL U74 ( .A(n272), .B(n21), .C(sfraddr[0]), .D(sfraddr[2]), .Y(n227) );
  NAND21X1 U75 ( .B(n262), .A(n181), .Y(n179) );
  NAND3X1 U76 ( .A(n193), .B(n50), .C(t_shift_clk), .Y(n176) );
  AND2X1 U77 ( .A(sfrdatai[7]), .B(n162), .Y(N113) );
  INVX1 U78 ( .A(n183), .Y(n268) );
  NAND4XL U79 ( .A(sfraddr[0]), .B(sfraddr[4]), .C(n194), .D(n195), .Y(n193)
         );
  NOR4XL U80 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[2]), .D(sfraddr[1]), 
        .Y(n195) );
  NOR2X1 U81 ( .A(n21), .B(n272), .Y(n194) );
  AO21X1 U82 ( .B(sfrdatai[7]), .C(n93), .A(n40), .Y(N125) );
  AND2X1 U83 ( .A(sfrdatai[7]), .B(n96), .Y(N136) );
  INVXL U84 ( .A(sfraddr[3]), .Y(n21) );
  INVX1 U85 ( .A(sfraddr[1]), .Y(n20) );
  INVX1 U86 ( .A(sfrdatai[1]), .Y(n25) );
  INVX1 U87 ( .A(sfrdatai[2]), .Y(n27) );
  INVX1 U88 ( .A(sfrdatai[0]), .Y(n23) );
  INVX1 U89 ( .A(sfrdatai[6]), .Y(n35) );
  INVX1 U90 ( .A(sfrdatai[3]), .Y(n29) );
  INVX1 U91 ( .A(sfrdatai[4]), .Y(n31) );
  INVX1 U92 ( .A(sfrdatai[5]), .Y(n33) );
  INVX1 U93 ( .A(rst), .Y(n59) );
  INVX1 U94 ( .A(n249), .Y(n157) );
  OAI31XL U95 ( .A(n255), .B(n262), .C(n3), .D(n248), .Y(n249) );
  NAND21X1 U96 ( .B(n82), .A(n149), .Y(n111) );
  NAND21X1 U97 ( .B(n36), .A(n127), .Y(n133) );
  NOR21XL U98 ( .B(t1ov), .A(n36), .Y(N59) );
  INVX1 U99 ( .A(n204), .Y(n265) );
  INVX1 U100 ( .A(rst), .Y(n58) );
  INVX1 U101 ( .A(n254), .Y(n114) );
  NAND2X1 U102 ( .A(n264), .B(n151), .Y(N428) );
  INVX1 U103 ( .A(n13), .Y(n151) );
  INVX1 U104 ( .A(n258), .Y(n262) );
  NOR21XL U105 ( .B(n262), .A(n286), .Y(rxd0oe) );
  NAND21X1 U106 ( .B(n258), .A(n181), .Y(n183) );
  NAND21X1 U107 ( .B(n36), .A(n7), .Y(n204) );
  NAND21X1 U108 ( .B(n37), .A(n128), .Y(N382) );
  OA21X1 U109 ( .B(n38), .C(n130), .A(N382), .Y(n3) );
  NOR21XL U110 ( .B(n98), .A(n36), .Y(n149) );
  NAND21X1 U111 ( .B(n131), .A(n262), .Y(n82) );
  NAND32X1 U112 ( .B(n221), .C(n251), .A(n7), .Y(n77) );
  NAND21X1 U113 ( .B(n82), .A(n98), .Y(n254) );
  OAI221X1 U114 ( .A(n82), .B(n251), .C(n2), .D(n77), .E(n52), .Y(n13) );
  AOI21X1 U115 ( .B(n286), .C(n251), .A(n39), .Y(n116) );
  NAND21X1 U116 ( .B(n7), .A(n41), .Y(N324) );
  OAI21X1 U117 ( .B(n284), .C(n121), .A(n51), .Y(n207) );
  NAND32X1 U118 ( .B(n38), .C(n258), .A(n252), .Y(n248) );
  INVX1 U119 ( .A(n78), .Y(n94) );
  INVX1 U120 ( .A(n143), .Y(n127) );
  INVX1 U121 ( .A(n256), .Y(n221) );
  AND2X1 U122 ( .A(n180), .B(n182), .Y(N224) );
  INVX1 U123 ( .A(n201), .Y(n180) );
  OAI32X1 U124 ( .A(n283), .B(n121), .C(n207), .D(n208), .E(n284), .Y(N188) );
  OAI22X1 U125 ( .A(n111), .B(n99), .C(n110), .D(n97), .Y(N473) );
  OAI22X1 U126 ( .A(n111), .B(n100), .C(n110), .D(n99), .Y(N474) );
  OAI22X1 U127 ( .A(n111), .B(n101), .C(n110), .D(n100), .Y(N475) );
  OAI22X1 U128 ( .A(n111), .B(n106), .C(n110), .D(n101), .Y(N476) );
  OAI22X1 U129 ( .A(n111), .B(n107), .C(n110), .D(n106), .Y(N477) );
  OAI22X1 U130 ( .A(n111), .B(n109), .C(n110), .D(n107), .Y(N478) );
  OAI22X1 U131 ( .A(n128), .B(n111), .C(n110), .D(n109), .Y(N479) );
  INVX1 U132 ( .A(n98), .Y(n220) );
  NOR2X1 U133 ( .A(n286), .B(n131), .Y(t_shift_clk) );
  OAI21X1 U134 ( .B(n251), .C(n123), .A(n124), .Y(n240) );
  OAI211X1 U135 ( .C(n108), .D(n125), .A(n123), .B(n52), .Y(n124) );
  NAND42X1 U136 ( .C(n125), .D(n114), .A(n126), .B(n52), .Y(n123) );
  INVX1 U137 ( .A(n253), .Y(n125) );
  OAI211X1 U138 ( .C(n139), .D(n110), .A(n111), .B(n52), .Y(N471) );
  NOR2X1 U139 ( .A(n168), .B(n166), .Y(N363) );
  XNOR2XL U140 ( .A(n92), .B(n290), .Y(n168) );
  NAND3X1 U141 ( .A(n45), .B(n291), .C(n166), .Y(N360) );
  NAND2X1 U142 ( .A(n44), .B(n203), .Y(N223) );
  NAND31X1 U143 ( .C(n258), .A(n116), .B(n263), .Y(N303) );
  NAND32X1 U144 ( .B(n258), .C(n252), .A(n251), .Y(n253) );
  MUX2X1 U145 ( .D0(n250), .D1(n252), .S(n262), .Y(n264) );
  AO21X1 U146 ( .B(n7), .C(rxd0ff), .A(n39), .Y(N325) );
  NAND32X1 U147 ( .B(n38), .C(n8), .A(n78), .Y(N166) );
  NAND21X1 U148 ( .B(n37), .A(n99), .Y(N376) );
  NAND21X1 U149 ( .B(n37), .A(n100), .Y(N377) );
  NAND21X1 U150 ( .B(n37), .A(n101), .Y(N378) );
  NAND21X1 U151 ( .B(n37), .A(n106), .Y(N379) );
  NAND21X1 U152 ( .B(n37), .A(n107), .Y(N380) );
  NAND21X1 U153 ( .B(n37), .A(n109), .Y(N381) );
  NAND21X1 U154 ( .B(n36), .A(n97), .Y(N375) );
  AND3X1 U155 ( .A(n63), .B(n47), .C(n68), .Y(N142) );
  INVX1 U156 ( .A(n61), .Y(n63) );
  INVX1 U157 ( .A(n250), .Y(n255) );
  NOR3XL U158 ( .A(n285), .B(n38), .C(n266), .Y(N207) );
  NOR2X1 U159 ( .A(n36), .B(n142), .Y(n245) );
  XNOR2XL U160 ( .A(n266), .B(n285), .Y(n142) );
  NOR2X1 U161 ( .A(n36), .B(n213), .Y(N307) );
  NAND21X1 U162 ( .B(r_baud_count[2]), .A(n289), .Y(n218) );
  INVX1 U163 ( .A(n92), .Y(n289) );
  NAND21X1 U164 ( .B(s0con[6]), .A(n214), .Y(n258) );
  INVX1 U165 ( .A(s0con[7]), .Y(n214) );
  INVX1 U166 ( .A(t_start), .Y(n286) );
  OAI21BX1 U167 ( .C(ri_tmp), .B(n150), .A(n4), .Y(n237) );
  MUX2IX1 U168 ( .D0(N348), .D1(n22), .S(n162), .Y(n4) );
  AO21X1 U169 ( .B(n162), .C(n26), .A(n161), .Y(n230) );
  MUX2BXL U170 ( .D0(n160), .D1(n154), .S(s0con2_tmp), .Y(n161) );
  NAND21X1 U171 ( .B(n150), .A(s0con2_val), .Y(n154) );
  AND2X1 U172 ( .A(s0con[2]), .B(n148), .Y(n160) );
  OAI222XL U173 ( .A(n25), .B(n115), .C(n150), .D(n113), .E(N108), .F(n112), 
        .Y(n241) );
  INVX1 U174 ( .A(ti_tmp), .Y(n113) );
  INVX1 U175 ( .A(s0con[1]), .Y(n112) );
  GEN2XL U176 ( .D(t_shift_count[1]), .E(t_shift_count[0]), .C(n178), .B(n270), 
        .A(n269), .Y(N282) );
  INVX1 U177 ( .A(n179), .Y(n269) );
  AO21X1 U178 ( .B(n211), .C(n210), .A(n206), .Y(N281) );
  INVX1 U179 ( .A(t_shift_count[0]), .Y(n210) );
  OA21X1 U180 ( .B(s0con[7]), .C(n205), .A(n181), .Y(n206) );
  INVX1 U181 ( .A(s0con[6]), .Y(n205) );
  OAI211X1 U182 ( .C(n23), .D(n179), .A(n51), .B(n191), .Y(N260) );
  AOI22X1 U183 ( .A(n268), .B(n24), .C(t_shift_reg[3]), .D(n270), .Y(n191) );
  OAI211X1 U184 ( .C(n25), .D(n179), .A(n47), .B(n190), .Y(N261) );
  AOI22X1 U185 ( .A(n268), .B(n26), .C(t_shift_reg[4]), .D(n270), .Y(n190) );
  OAI211X1 U186 ( .C(n179), .D(n33), .A(n51), .B(n186), .Y(N265) );
  AOI22X1 U187 ( .A(n268), .B(n34), .C(t_shift_reg[8]), .D(n270), .Y(n186) );
  OAI211X1 U188 ( .C(n179), .D(n35), .A(n43), .B(n185), .Y(N266) );
  AOI22X1 U189 ( .A(n268), .B(sfrdatai[7]), .C(t_shift_reg[9]), .D(n270), .Y(
        n185) );
  OAI2B11X1 U190 ( .D(t_shift_reg[1]), .C(n176), .A(n267), .B(n44), .Y(N258)
         );
  OAI211X1 U191 ( .C(n27), .D(n179), .A(n46), .B(n189), .Y(N262) );
  AOI22X1 U192 ( .A(n28), .B(n268), .C(t_shift_reg[5]), .D(n270), .Y(n189) );
  OAI211X1 U193 ( .C(n179), .D(n29), .A(n48), .B(n188), .Y(N263) );
  AOI22X1 U194 ( .A(n30), .B(n268), .C(t_shift_reg[6]), .D(n270), .Y(n188) );
  OAI211X1 U195 ( .C(n179), .D(n31), .A(n42), .B(n187), .Y(N264) );
  AOI22X1 U196 ( .A(n32), .B(n268), .C(t_shift_reg[7]), .D(n270), .Y(n187) );
  NAND3X1 U197 ( .A(n183), .B(n50), .C(n184), .Y(N267) );
  AOI22X1 U198 ( .A(t_shift_reg[10]), .B(n270), .C(sfrdatai[7]), .D(n181), .Y(
        n184) );
  OAI211X1 U199 ( .C(n23), .D(n183), .A(n49), .B(n192), .Y(N259) );
  NAND2X1 U200 ( .A(t_shift_reg[2]), .B(n270), .Y(n192) );
  MUX2BXL U201 ( .D0(sfrdatai[7]), .D1(n5), .S(n6), .Y(n271) );
  NAND2X1 U202 ( .A(bd), .B(n43), .Y(n5) );
  NAND4X1 U203 ( .A(sfraddr[6]), .B(n146), .C(n41), .D(n20), .Y(n6) );
  MUX2X1 U204 ( .D0(n65), .D1(sfrdatai[7]), .S(n64), .Y(n244) );
  AND2X1 U205 ( .A(smod), .B(n52), .Y(n65) );
  AND4X1 U206 ( .A(n141), .B(n140), .C(sfraddr[0]), .D(sfraddr[2]), .Y(n64) );
  NOR4XL U207 ( .A(sfraddr[5]), .B(sfraddr[4]), .C(sfraddr[3]), .D(n272), .Y(
        n141) );
  NAND32X1 U208 ( .B(n211), .C(n38), .A(n90), .Y(N268) );
  NAND21X1 U209 ( .B(n267), .A(n89), .Y(n90) );
  NAND21X1 U210 ( .B(s0con[3]), .A(s0con[7]), .Y(n89) );
  OAI21X1 U211 ( .B(n175), .C(n176), .A(n267), .Y(N284) );
  XOR2X1 U212 ( .A(n138), .B(t_shift_count[3]), .Y(n175) );
  AOI21X1 U213 ( .B(n138), .C(n177), .A(n176), .Y(N283) );
  NAND21X1 U214 ( .B(n178), .A(t_shift_count[2]), .Y(n177) );
  NAND2X1 U215 ( .A(n137), .B(n267), .Y(n243) );
  OAI211X1 U216 ( .C(t_shift_count[3]), .D(n138), .A(n51), .B(t_start), .Y(
        n137) );
  AOI21X1 U217 ( .B(n74), .C(n254), .A(n39), .Y(n238) );
  MUX2X1 U218 ( .D0(n73), .D1(n139), .S(n127), .Y(n74) );
  NAND21X1 U219 ( .B(newinstr), .A(ri_tmp), .Y(n73) );
  MUX2X1 U220 ( .D0(s0con2_tmp), .D1(n147), .S(n145), .Y(n232) );
  AOI32X1 U221 ( .A(n48), .B(n144), .C(n143), .D(n147), .E(n139), .Y(n145) );
  INVX1 U222 ( .A(n133), .Y(n147) );
  INVX1 U223 ( .A(newinstr), .Y(n144) );
  NOR2X1 U224 ( .A(n36), .B(n135), .Y(n242) );
  AOI32X1 U225 ( .A(t_shift_clk), .B(t_shift_count[0]), .C(n136), .D(ti_tmp), 
        .E(n144), .Y(n135) );
  NOR3XL U226 ( .A(t_shift_count[1]), .B(t_shift_count[3]), .C(
        t_shift_count[2]), .Y(n136) );
  AO21X1 U227 ( .B(s0relh[6]), .C(n163), .A(n203), .Y(n201) );
  AO21X1 U228 ( .B(t_baud_count[1]), .C(t_baud_count[0]), .A(n201), .Y(n199)
         );
  MUX2X1 U229 ( .D0(n68), .D1(baud_rate_ov), .S(s0con[6]), .Y(n69) );
  MUX2BXL U230 ( .D0(n72), .D1(t1ov_ff), .S(n71), .Y(n266) );
  AND2X1 U231 ( .A(s0con[6]), .B(n70), .Y(n71) );
  NAND21X1 U232 ( .B(n262), .A(n69), .Y(n72) );
  INVX1 U233 ( .A(bd), .Y(n70) );
  NAND21X1 U234 ( .B(n204), .A(t_start), .Y(n203) );
  NAND21X1 U235 ( .B(r_clk_ov2), .A(n62), .Y(n68) );
  AO22X1 U236 ( .A(n180), .B(n171), .C(t_baud_count[3]), .D(n170), .Y(N227) );
  AO21X1 U237 ( .B(t_baud_count[3]), .C(n287), .A(n163), .Y(n171) );
  INVX1 U238 ( .A(n199), .Y(n170) );
  MUX2BXL U239 ( .D0(baud_r2_clk), .D1(n266), .S(smod), .Y(n7) );
  OAI22X1 U240 ( .A(n2), .B(n88), .C(n159), .D(n248), .Y(N425) );
  OA22X1 U241 ( .A(n38), .B(n250), .C(n159), .D(n3), .Y(n88) );
  AOI21X1 U242 ( .B(r_shift_count[1]), .C(r_shift_count[0]), .A(n158), .Y(n159) );
  OAI21X1 U243 ( .B(n199), .C(n287), .A(n200), .Y(N226) );
  NAND43X1 U244 ( .B(n201), .C(n198), .D(n182), .A(n287), .Y(n200) );
  INVX1 U245 ( .A(t_baud_count[2]), .Y(n287) );
  INVX1 U246 ( .A(t_baud_count[1]), .Y(n198) );
  AOI21X1 U247 ( .B(n155), .C(n156), .A(n157), .Y(N426) );
  NAND21X1 U248 ( .B(n158), .A(r_shift_count[2]), .Y(n156) );
  INVX1 U249 ( .A(s0relh[7]), .Y(n62) );
  NOR2X1 U250 ( .A(r_shift_count[0]), .B(n157), .Y(N424) );
  MUX2IX1 U251 ( .D0(t_baud_ov), .D1(clk_ov12), .S(n262), .Y(n131) );
  NOR21XL U252 ( .B(rxd0_fall_fl), .A(N324), .Y(n102) );
  NAND43X1 U253 ( .B(s0con[0]), .C(n76), .D(n77), .A(n149), .Y(n110) );
  INVX1 U254 ( .A(n82), .Y(n76) );
  AO21X1 U255 ( .B(r_clk_ov2), .C(n62), .A(n8), .Y(n78) );
  MUX2X1 U256 ( .D0(n67), .D1(n18), .S(s0relh[6]), .Y(n256) );
  AND3X1 U257 ( .A(n290), .B(n164), .C(r_baud_count[3]), .Y(n67) );
  OR4X1 U258 ( .A(s0con[0]), .B(n262), .C(n220), .D(n77), .Y(n143) );
  INVX1 U259 ( .A(n77), .Y(r_shift_clk) );
  NAND41X1 U260 ( .D(n223), .A(tim_baud[9]), .B(tim_baud[8]), .C(n224), .Y(n61) );
  AOI21BBXL U261 ( .B(clk_count[1]), .C(n207), .A(N185), .Y(n208) );
  NOR21XL U262 ( .B(n180), .A(n202), .Y(N225) );
  XNOR2XL U263 ( .A(t_baud_count[1]), .B(t_baud_count[0]), .Y(n202) );
  GEN2XL U264 ( .D(n292), .E(n293), .C(n102), .B(fluctuation_conter[1]), .A(
        n103), .Y(n233) );
  INVX1 U265 ( .A(n104), .Y(n292) );
  NOR4XL U266 ( .A(fluctuation_conter[1]), .B(n102), .C(n104), .D(n293), .Y(
        n103) );
  NAND21X1 U267 ( .B(n259), .A(n258), .Y(n126) );
  AOI32X1 U268 ( .A(n257), .B(n256), .C(n7), .D(n108), .E(n255), .Y(n259) );
  AO21X1 U269 ( .B(n130), .C(rxd0_val), .A(n98), .Y(n257) );
  AND2X1 U270 ( .A(n91), .B(n45), .Y(N170) );
  AO22X1 U271 ( .A(s0rell[3]), .B(n8), .C(N148), .D(n94), .Y(n91) );
  AND2X1 U272 ( .A(n95), .B(n46), .Y(N169) );
  AO22X1 U273 ( .A(s0rell[2]), .B(n8), .C(N147), .D(n94), .Y(n95) );
  MUX2BXL U274 ( .D0(baud_rate_ov), .D1(n61), .S(s0relh[7]), .Y(n8) );
  OAI21BBX1 U275 ( .A(s0relh[1]), .B(n1), .C(n9), .Y(n281) );
  AOI21X1 U276 ( .B(N154), .C(n94), .A(n40), .Y(n9) );
  OAI21BBX1 U277 ( .A(s0relh[0]), .B(n1), .C(n10), .Y(n280) );
  AOI21X1 U278 ( .B(N153), .C(n94), .A(n39), .Y(n10) );
  OAI21BBX1 U279 ( .A(s0rell[7]), .B(n8), .C(n11), .Y(n274) );
  AOI21X1 U280 ( .B(N152), .C(n94), .A(n40), .Y(n11) );
  OAI21BBX1 U281 ( .A(s0rell[6]), .B(n8), .C(n12), .Y(n275) );
  AOI21X1 U282 ( .B(N151), .C(n94), .A(n40), .Y(n12) );
  OAI21BBX1 U283 ( .A(s0rell[5]), .B(n8), .C(n14), .Y(n276) );
  AOI21X1 U284 ( .B(N150), .C(n94), .A(n40), .Y(n14) );
  OAI21BBX1 U285 ( .A(s0rell[4]), .B(n1), .C(n15), .Y(n277) );
  AOI21X1 U286 ( .B(N149), .C(n94), .A(n39), .Y(n15) );
  OAI21BBX1 U287 ( .A(s0rell[1]), .B(n8), .C(n16), .Y(n278) );
  AOI21X1 U288 ( .B(N146), .C(n94), .A(n40), .Y(n16) );
  OAI21BBX1 U289 ( .A(s0rell[0]), .B(n8), .C(n17), .Y(n279) );
  AOI21X1 U290 ( .B(N145), .C(n94), .A(n40), .Y(n17) );
  NAND2X1 U291 ( .A(rxd0_fall_fl), .B(n43), .Y(n104) );
  OAI22BX1 U292 ( .B(r_shift_reg[1]), .A(n111), .D(r_shift_reg[0]), .C(n110), 
        .Y(N472) );
  AND2X1 U293 ( .A(s0con[7]), .B(n247), .Y(n229) );
  OAI33XL U294 ( .A(n246), .B(n38), .C(n222), .D(n221), .E(n38), .F(n220), .Y(
        n247) );
  INVX1 U295 ( .A(receive_11_bits), .Y(n222) );
  MUX2BXL U296 ( .D0(n219), .D1(n218), .S(s0relh[6]), .Y(n246) );
  OAI32X1 U297 ( .A(n207), .B(clk_count[2]), .C(n121), .D(n208), .E(n283), .Y(
        N187) );
  OAI32X1 U298 ( .A(n104), .B(fluctuation_conter[0]), .C(n102), .D(n293), .E(
        n273), .Y(n234) );
  INVX1 U299 ( .A(n102), .Y(n273) );
  OAI32X1 U300 ( .A(n132), .B(n38), .C(n129), .D(n128), .E(n133), .Y(n231) );
  INVX1 U301 ( .A(s0con2_val), .Y(n129) );
  NOR6XL U302 ( .A(n251), .B(s0con[0]), .C(n139), .D(n262), .E(n221), .F(n220), 
        .Y(n132) );
  OAI32X1 U303 ( .A(n291), .B(n104), .C(n294), .D(n169), .E(n166), .Y(N362) );
  INVX1 U304 ( .A(fluctuation_conter[1]), .Y(n294) );
  AOI21X1 U305 ( .B(r_baud_count[1]), .C(n288), .A(n164), .Y(n169) );
  OAI32X1 U306 ( .A(n291), .B(n104), .C(n293), .D(r_baud_count[0]), .E(n166), 
        .Y(N361) );
  NAND3X1 U307 ( .A(r_start), .B(n291), .C(n265), .Y(n166) );
  NOR2X1 U308 ( .A(n207), .B(clk_count[0]), .Y(N185) );
  NOR2X1 U309 ( .A(n288), .B(r_baud_count[1]), .Y(n164) );
  NOR4XL U310 ( .A(n196), .B(t_baud_count[1]), .C(t_baud_count[3]), .D(
        t_baud_count[2]), .Y(N230) );
  NAND2X1 U311 ( .A(t_baud_count[0]), .B(n265), .Y(n196) );
  INVX1 U312 ( .A(n75), .Y(N348) );
  NAND21X1 U313 ( .B(n37), .A(s0con[0]), .Y(n75) );
  INVX1 U314 ( .A(r_baud_count[0]), .Y(n288) );
  NOR2X1 U315 ( .A(n165), .B(n166), .Y(N364) );
  XNOR2XL U316 ( .A(r_baud_count[3]), .B(n167), .Y(n165) );
  NOR2X1 U317 ( .A(n290), .B(n92), .Y(n167) );
  NAND3X1 U318 ( .A(tim_baud[6]), .B(tim_baud[5]), .C(tim_baud[7]), .Y(n223)
         );
  NAND3X1 U319 ( .A(n116), .B(n117), .C(n118), .Y(n239) );
  NAND4X1 U320 ( .A(t_shift_count[3]), .B(t_shift_count[0]), .C(txd0), .D(n122), .Y(n117) );
  MUX2BXL U321 ( .D0(n263), .D1(n119), .S(n262), .Y(n118) );
  AND3X1 U322 ( .A(n2), .B(n261), .C(n260), .Y(n122) );
  AND2X1 U323 ( .A(r_baud_count[2]), .B(n164), .Y(n18) );
  NAND21X1 U324 ( .B(n87), .A(rxd0_fall), .Y(n250) );
  NOR32XL U325 ( .B(n216), .C(n46), .A(n215), .Y(n235) );
  MUX2X1 U326 ( .D0(r_baud_count[3]), .D1(r_baud_count[2]), .S(s0relh[6]), .Y(
        n216) );
  AOI32X1 U327 ( .A(n214), .B(n213), .C(n212), .D(rxd0_fall_fl), .E(n105), .Y(
        n215) );
  INVX1 U328 ( .A(rxd0ff), .Y(n213) );
  NAND32X1 U329 ( .B(n87), .C(n86), .A(n85), .Y(n252) );
  INVX1 U330 ( .A(ri0_fall), .Y(n86) );
  INVX1 U331 ( .A(n131), .Y(n85) );
  INVX1 U332 ( .A(n197), .Y(n163) );
  NAND41X1 U333 ( .D(t_baud_count[3]), .A(t_baud_count[2]), .B(t_baud_count[1]), .C(t_baud_count[0]), .Y(n197) );
  NAND21X1 U334 ( .B(r_shift_count[2]), .A(n158), .Y(n155) );
  MUX2X1 U335 ( .D0(n84), .D1(ri0_fall), .S(n83), .Y(n236) );
  AND3X1 U337 ( .A(ri0_ff), .B(n47), .C(n79), .Y(n84) );
  AND3X1 U338 ( .A(n82), .B(n47), .C(n81), .Y(n83) );
  NAND32X1 U339 ( .B(n258), .C(n80), .A(n79), .Y(n81) );
  AO21X1 U340 ( .B(rxd0_vec[1]), .C(n7), .A(n39), .Y(N327) );
  AO21X1 U341 ( .B(rxd0_vec[0]), .C(n7), .A(n39), .Y(N326) );
  INVX1 U342 ( .A(r_baud_count[2]), .Y(n290) );
  AND2X1 U343 ( .A(clk_count[0]), .B(n46), .Y(N190) );
  NOR42XL U344 ( .C(r_shift_count[3]), .D(r_shift_count[1]), .A(
        r_shift_count[0]), .B(r_shift_count[2]), .Y(n130) );
  INVX1 U345 ( .A(r_start), .Y(n251) );
  AND2X1 U346 ( .A(n217), .B(n18), .Y(n219) );
  INVX1 U347 ( .A(r_baud_count[3]), .Y(n217) );
  NOR2X1 U348 ( .A(r_shift_count[1]), .B(r_shift_count[0]), .Y(n158) );
  NOR2X1 U349 ( .A(n155), .B(r_shift_count[3]), .Y(n108) );
  OAI21X1 U350 ( .B(N382), .C(n152), .A(n153), .Y(N427) );
  GEN2XL U351 ( .D(n130), .E(n258), .C(n152), .B(n264), .A(n55), .Y(n153) );
  AOI21X1 U352 ( .B(n155), .C(r_shift_count[3]), .A(n108), .Y(n152) );
  NOR42XL U353 ( .C(n283), .D(N190), .A(n284), .B(clk_count[1]), .Y(N191) );
  NOR4XL U354 ( .A(n173), .B(receive_11_bits), .C(rxd0_fall), .D(n36), .Y(N306) );
  OAI21X1 U355 ( .B(n174), .C(rxd0_fall_fl), .A(n251), .Y(n173) );
  NOR21XL U356 ( .B(rxd0_ff), .A(rxd0ff), .Y(n174) );
  NAND3X1 U357 ( .A(tim_baud[1]), .B(tim_baud[0]), .C(tim_baud[2]), .Y(n225)
         );
  NOR2X1 U358 ( .A(n209), .B(n207), .Y(N186) );
  XNOR2XL U359 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n209) );
  INVX1 U360 ( .A(s0con[4]), .Y(n87) );
  NAND21X1 U361 ( .B(t_shift_count[2]), .A(n178), .Y(n138) );
  NAND2X1 U362 ( .A(n19), .B(n45), .Y(N333) );
  MUX2IX1 U363 ( .D0(n172), .D1(rxd0ff), .S(n2), .Y(n19) );
  NAND2X1 U364 ( .A(r_baud_count[1]), .B(r_baud_count[0]), .Y(n92) );
  NAND2X1 U365 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n121) );
  AND3X1 U366 ( .A(n98), .B(s0con[6]), .C(rxd0_ff), .Y(n212) );
  NOR2X1 U367 ( .A(t_shift_count[1]), .B(t_shift_count[0]), .Y(n178) );
  OAI31XL U368 ( .A(n282), .B(clk_count[3]), .C(clk_count[2]), .D(n120), .Y(
        n119) );
  INVX1 U369 ( .A(n121), .Y(n282) );
  OAI31XL U370 ( .A(clk_count[0]), .B(clk_count[2]), .C(clk_count[1]), .D(
        clk_count[3]), .Y(n120) );
  INVX1 U371 ( .A(rxd0_val), .Y(n128) );
  INVX1 U372 ( .A(n66), .Y(n139) );
  NAND21X1 U373 ( .B(rxd0_val), .A(s0con[5]), .Y(n66) );
  INVX1 U374 ( .A(clk_count[3]), .Y(n284) );
  INVX1 U375 ( .A(t_shift_count[2]), .Y(n260) );
  INVX1 U376 ( .A(t_shift_count[1]), .Y(n261) );
  NAND2X1 U377 ( .A(rxd0_fall), .B(n108), .Y(n105) );
  INVX1 U378 ( .A(s0con[0]), .Y(n79) );
  INVX1 U379 ( .A(rxd0_fall), .Y(n291) );
  INVX1 U380 ( .A(r_shift_reg[2]), .Y(n99) );
  INVX1 U381 ( .A(r_shift_reg[3]), .Y(n100) );
  INVX1 U382 ( .A(r_shift_reg[4]), .Y(n101) );
  INVX1 U383 ( .A(r_shift_reg[5]), .Y(n106) );
  INVX1 U384 ( .A(r_shift_reg[6]), .Y(n107) );
  INVX1 U385 ( .A(r_shift_reg[7]), .Y(n109) );
  INVX1 U386 ( .A(fluctuation_conter[0]), .Y(n293) );
  INVX1 U387 ( .A(t_baud_count[0]), .Y(n182) );
  INVX1 U388 ( .A(r_shift_reg[1]), .Y(n97) );
  INVX1 U389 ( .A(clk_count[2]), .Y(n283) );
  INVX1 U390 ( .A(t_shift_reg[0]), .Y(n263) );
  INVX1 U391 ( .A(baud_r_count), .Y(n285) );
  INVX1 U392 ( .A(ri0_ff), .Y(n80) );
  NAND31X1 U393 ( .C(sfraddr[6]), .A(n20), .B(n146), .Y(n134) );
endmodule


module serial0_a0_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ports_a0 ( clkper, rst, port0, sfrdatai, sfraddr, sfrwe );
  output [7:0] port0;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkper, rst, sfrwe;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, net12300, n2, n3, n4, n1, n5;

  SNPS_CLOCK_GATE_HIGH_ports_a0 clk_gate_p0_reg ( .CLK(clkper), .EN(N2), 
        .ENCLK(net12300), .TE(1'b0) );
  DFFQX1 p0_reg_7_ ( .D(N10), .C(net12300), .Q(port0[7]) );
  DFFQX1 p0_reg_6_ ( .D(N9), .C(net12300), .Q(port0[6]) );
  DFFQX1 p0_reg_4_ ( .D(N7), .C(net12300), .Q(port0[4]) );
  DFFQX1 p0_reg_5_ ( .D(N8), .C(net12300), .Q(port0[5]) );
  DFFQX1 p0_reg_3_ ( .D(N6), .C(net12300), .Q(port0[3]) );
  DFFQX1 p0_reg_0_ ( .D(N3), .C(net12300), .Q(port0[0]) );
  DFFQX1 p0_reg_2_ ( .D(N5), .C(net12300), .Q(port0[2]) );
  DFFQX1 p0_reg_1_ ( .D(N4), .C(net12300), .Q(port0[1]) );
  INVX1 U2 ( .A(n2), .Y(n5) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(N2) );
  NAND42X1 U4 ( .C(sfraddr[3]), .D(sfraddr[2]), .A(n3), .B(n4), .Y(n2) );
  NOR3XL U5 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n3) );
  NOR42XL U6 ( .C(sfrwe), .D(n1), .A(sfraddr[1]), .B(sfraddr[0]), .Y(n4) );
  AND2X1 U7 ( .A(sfrdatai[0]), .B(n5), .Y(N3) );
  AND2X1 U8 ( .A(sfrdatai[1]), .B(n5), .Y(N4) );
  AND2X1 U9 ( .A(sfrdatai[2]), .B(n5), .Y(N5) );
  AND2X1 U10 ( .A(sfrdatai[3]), .B(n5), .Y(N6) );
  AND2X1 U11 ( .A(sfrdatai[4]), .B(n5), .Y(N7) );
  AND2X1 U12 ( .A(sfrdatai[5]), .B(n5), .Y(N8) );
  AND2X1 U13 ( .A(sfrdatai[6]), .B(n5), .Y(N9) );
  AND2X1 U14 ( .A(sfrdatai[7]), .B(n5), .Y(N10) );
  INVX1 U15 ( .A(rst), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ports_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mdu_a0 ( clkper, rst, mdubsy, sfrdatai, sfraddr, sfrwe, sfroe, arcon, 
        md0, md1, md2, md3, md4, md5 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] arcon;
  output [7:0] md0;
  output [7:0] md1;
  output [7:0] md2;
  output [7:0] md3;
  output [7:0] md4;
  output [7:0] md5;
  input clkper, rst, sfrwe, sfroe;
  output mdubsy;
  wire   N104, N105, N106, N107, N108, N109, setmdef, N190, N191, N192, N193,
         N194, N195, N196, N197, N198, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N332, N333, N334, N335, N336, N337, N338, N339,
         N340, N405, N406, N407, N408, N409, N410, N411, N412, N413, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N566, N567, N568, N569, N570,
         N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581,
         N610, N612, N613, N614, N674, N675, N676, N677, N678, set_div16,
         set_div32, N802, N892, N893, N894, N895, net12318, net12324, net12329,
         net12334, net12339, net12344, net12349, n166, n167, n171, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n195, n197,
         n198, n200, n201, n202, n204, n206, n208, n209, n210, n211, n212,
         n213, n214, n217, n218, n220, n221, n222, n223, n225, n227, n228,
         n229, n231, n232, n233, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n248, n253, n254, n255, n256, n257,
         n258, n260, n263, n264, n265, n267, n277, n278, n291, n294, n296,
         n297, n299, n302, n306, n317, n318, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n364, n365, n366, n367, n384, n386,
         n387, n388, n389, n390, n391, n394, n396, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n168, n169, n170, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n193, n194, n196, n199, n203, n205, n207, n215, n216,
         n219, n224, n226, n230, n234, n247, n249, n250, n251, n252, n259,
         n261, n262, n266, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n292, n293, n295, n298, n300, n301, n303, n304, n305,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n385, n392, n393, n395, n397,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2;
  wire   [3:0] oper_reg;
  wire   [4:1] counter_st;
  wire   [17:1] sum1;
  wire   [17:1] sum;
  wire   [15:0] norm_reg;
  wire   [1:0] mdu_op;
  wire   [17:0] arg_a;
  wire   [16:1] arg_b;
  wire   [17:0] arg_c;
  wire   [16:1] arg_d;
  wire   [4:3] r384_carry;

  SNPS_CLOCK_GATE_HIGH_mdu_a0_0 clk_gate_arcon_s_reg ( .CLK(clkper), .EN(N104), 
        .ENCLK(net12318), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_6 clk_gate_md0_s_reg ( .CLK(clkper), .EN(N190), 
        .ENCLK(net12324), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_5 clk_gate_md1_s_reg ( .CLK(clkper), .EN(N258), 
        .ENCLK(net12329), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_4 clk_gate_md2_s_reg ( .CLK(clkper), .EN(N332), 
        .ENCLK(net12334), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_3 clk_gate_md3_s_reg ( .CLK(clkper), .EN(N405), 
        .ENCLK(net12339), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_2 clk_gate_md4_s_reg ( .CLK(clkper), .EN(N453), 
        .ENCLK(net12344), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_1 clk_gate_md5_s_reg ( .CLK(clkper), .EN(N483), 
        .ENCLK(net12349), .TE(1'b0) );
  mdu_a0_DW01_add_0 add_1040 ( .A(arg_c), .B({1'b0, arg_d, n87}), .CI(1'b0), 
        .SUM({sum, SYNOPSYS_UNCONNECTED_1}), .CO() );
  mdu_a0_DW01_add_1 add_961 ( .A({arg_a[17:1], n31}), .B({1'b0, arg_b, n87}), 
        .CI(1'b0), .SUM({sum1, SYNOPSYS_UNCONNECTED_2}), .CO() );
  DFFQX1 setmdef_reg ( .D(N802), .C(clkper), .Q(setmdef) );
  DFFQX1 set_div16_reg ( .D(n414), .C(clkper), .Q(set_div16) );
  DFFQX1 set_div32_reg ( .D(n413), .C(clkper), .Q(set_div32) );
  DFFQX1 counter_st_reg_0_ ( .D(N674), .C(clkper), .Q(N610) );
  DFFQX1 counter_st_reg_4_ ( .D(N678), .C(clkper), .Q(counter_st[4]) );
  DFFQX1 counter_st_reg_2_ ( .D(N676), .C(clkper), .Q(counter_st[2]) );
  DFFQX1 counter_st_reg_3_ ( .D(N677), .C(clkper), .Q(counter_st[3]) );
  DFFQX1 counter_st_reg_1_ ( .D(N675), .C(clkper), .Q(counter_st[1]) );
  DFFQX1 oper_reg_reg_1_ ( .D(N893), .C(clkper), .Q(oper_reg[1]) );
  DFFQX1 oper_reg_reg_0_ ( .D(N892), .C(clkper), .Q(oper_reg[0]) );
  DFFQX1 oper_reg_reg_2_ ( .D(N894), .C(clkper), .Q(oper_reg[2]) );
  DFFQX1 oper_reg_reg_3_ ( .D(N895), .C(clkper), .Q(oper_reg[3]) );
  DFFQX1 arcon_s_reg_6_ ( .D(n408), .C(clkper), .Q(arcon[6]) );
  DFFQX1 arcon_s_reg_7_ ( .D(n410), .C(clkper), .Q(arcon[7]) );
  DFFQX1 md0_s_reg_6_ ( .D(N197), .C(net12324), .Q(md0[6]) );
  DFFQX1 md0_s_reg_7_ ( .D(N198), .C(net12324), .Q(md0[7]) );
  DFFQX1 md1_s_reg_5_ ( .D(N264), .C(net12329), .Q(md1[5]) );
  DFFQX1 arcon_s_reg_5_ ( .D(n409), .C(net12318), .Q(arcon[5]) );
  DFFQX1 md0_s_reg_5_ ( .D(N196), .C(net12324), .Q(md0[5]) );
  DFFQX1 md1_s_reg_4_ ( .D(N263), .C(net12329), .Q(md1[4]) );
  DFFQX1 arcon_s_reg_4_ ( .D(N109), .C(net12318), .Q(arcon[4]) );
  DFFQX1 md0_s_reg_4_ ( .D(N195), .C(net12324), .Q(md0[4]) );
  DFFQX1 norm_reg_reg_15_ ( .D(N581), .C(clkper), .Q(norm_reg[15]) );
  DFFQX1 md1_s_reg_6_ ( .D(N265), .C(net12329), .Q(md1[6]) );
  DFFQX1 norm_reg_reg_14_ ( .D(N580), .C(clkper), .Q(norm_reg[14]) );
  DFFQX1 arcon_s_reg_3_ ( .D(N108), .C(net12318), .Q(arcon[3]) );
  DFFQX1 md5_s_reg_6_ ( .D(N490), .C(net12349), .Q(md5[6]) );
  DFFQX1 norm_reg_reg_13_ ( .D(N579), .C(clkper), .Q(norm_reg[13]) );
  DFFQX1 md1_s_reg_3_ ( .D(N262), .C(net12329), .Q(md1[3]) );
  DFFQX1 md0_s_reg_3_ ( .D(N194), .C(net12324), .Q(md0[3]) );
  DFFQX1 md5_s_reg_7_ ( .D(N491), .C(net12349), .Q(md5[7]) );
  DFFQX1 md3_s_reg_6_ ( .D(N412), .C(net12339), .Q(md3[6]) );
  DFFQX1 norm_reg_reg_12_ ( .D(N578), .C(clkper), .Q(norm_reg[12]) );
  DFFQX1 md3_s_reg_5_ ( .D(N411), .C(net12339), .Q(md3[5]) );
  DFFQX1 md5_s_reg_5_ ( .D(N489), .C(net12349), .Q(md5[5]) );
  DFFQX1 md5_s_reg_3_ ( .D(N487), .C(net12349), .Q(md5[3]) );
  DFFQX1 md5_s_reg_4_ ( .D(N488), .C(net12349), .Q(md5[4]) );
  DFFQX1 norm_reg_reg_10_ ( .D(N576), .C(clkper), .Q(norm_reg[10]) );
  DFFQX1 norm_reg_reg_11_ ( .D(N577), .C(clkper), .Q(norm_reg[11]) );
  DFFQX1 md3_s_reg_3_ ( .D(N409), .C(net12339), .Q(md3[3]) );
  DFFQX1 md3_s_reg_4_ ( .D(N410), .C(net12339), .Q(md3[4]) );
  DFFQX1 norm_reg_reg_9_ ( .D(N575), .C(clkper), .Q(norm_reg[9]) );
  DFFQX1 norm_reg_reg_8_ ( .D(N574), .C(clkper), .Q(norm_reg[8]) );
  DFFQX1 norm_reg_reg_7_ ( .D(N573), .C(clkper), .Q(norm_reg[7]) );
  DFFQX1 md4_s_reg_7_ ( .D(N461), .C(net12344), .Q(md4[7]) );
  DFFQX1 norm_reg_reg_6_ ( .D(N572), .C(clkper), .Q(norm_reg[6]) );
  DFFQX1 md2_s_reg_7_ ( .D(N340), .C(net12334), .Q(md2[7]) );
  DFFQX1 md4_s_reg_6_ ( .D(N460), .C(net12344), .Q(md4[6]) );
  DFFQX1 norm_reg_reg_4_ ( .D(N570), .C(clkper), .Q(norm_reg[4]) );
  DFFQX1 norm_reg_reg_5_ ( .D(N571), .C(clkper), .Q(norm_reg[5]) );
  DFFQX1 md2_s_reg_5_ ( .D(N338), .C(net12334), .Q(md2[5]) );
  DFFQX1 md2_s_reg_6_ ( .D(N339), .C(net12334), .Q(md2[6]) );
  DFFQX1 md4_s_reg_5_ ( .D(N459), .C(net12344), .Q(md4[5]) );
  DFFQX1 md4_s_reg_4_ ( .D(N458), .C(net12344), .Q(md4[4]) );
  DFFQX1 norm_reg_reg_3_ ( .D(N569), .C(clkper), .Q(norm_reg[3]) );
  DFFQX1 md2_s_reg_4_ ( .D(N337), .C(net12334), .Q(md2[4]) );
  DFFQX1 md4_s_reg_3_ ( .D(N457), .C(net12344), .Q(md4[3]) );
  DFFQX1 norm_reg_reg_2_ ( .D(N568), .C(clkper), .Q(norm_reg[2]) );
  DFFQX1 norm_reg_reg_1_ ( .D(N567), .C(clkper), .Q(norm_reg[1]) );
  DFFQX1 md2_s_reg_3_ ( .D(N336), .C(net12334), .Q(md2[3]) );
  DFFQX1 norm_reg_reg_0_ ( .D(N566), .C(clkper), .Q(norm_reg[0]) );
  DFFQX1 md1_s_reg_7_ ( .D(N266), .C(net12329), .Q(md1[7]) );
  DFFQX1 md3_s_reg_7_ ( .D(N413), .C(net12339), .Q(md3[7]) );
  DFFQX1 mdu_op_reg_0_ ( .D(n411), .C(clkper), .Q(mdu_op[0]) );
  DFFQX1 mdu_op_reg_1_ ( .D(n412), .C(clkper), .Q(mdu_op[1]) );
  DFFQX1 md4_s_reg_0_ ( .D(N454), .C(net12344), .Q(md4[0]) );
  DFFQX1 md4_s_reg_2_ ( .D(N456), .C(net12344), .Q(md4[2]) );
  DFFQX1 md1_s_reg_0_ ( .D(N259), .C(net12329), .Q(md1[0]) );
  DFFQX1 arcon_s_reg_1_ ( .D(N106), .C(net12318), .Q(arcon[1]) );
  DFFQX1 arcon_s_reg_0_ ( .D(N105), .C(net12318), .Q(arcon[0]) );
  DFFQX1 arcon_s_reg_2_ ( .D(N107), .C(net12318), .Q(arcon[2]) );
  DFFQX1 md3_s_reg_0_ ( .D(N406), .C(net12339), .Q(md3[0]) );
  DFFQX1 md2_s_reg_2_ ( .D(N335), .C(net12334), .Q(md2[2]) );
  DFFQX1 md2_s_reg_1_ ( .D(N334), .C(net12334), .Q(md2[1]) );
  DFFQX1 md4_s_reg_1_ ( .D(N455), .C(net12344), .Q(md4[1]) );
  DFFQX1 md5_s_reg_0_ ( .D(N484), .C(net12349), .Q(md5[0]) );
  DFFQX1 md0_s_reg_0_ ( .D(N191), .C(net12324), .Q(md0[0]) );
  DFFQX1 md2_s_reg_0_ ( .D(N333), .C(net12334), .Q(md2[0]) );
  DFFQX1 md5_s_reg_2_ ( .D(N486), .C(net12349), .Q(md5[2]) );
  DFFQX1 md1_s_reg_2_ ( .D(N261), .C(net12329), .Q(md1[2]) );
  DFFQX1 md0_s_reg_2_ ( .D(N193), .C(net12324), .Q(md0[2]) );
  DFFQX1 md1_s_reg_1_ ( .D(N260), .C(net12329), .Q(md1[1]) );
  DFFQX1 md3_s_reg_1_ ( .D(N407), .C(net12339), .Q(md3[1]) );
  DFFQX1 md3_s_reg_2_ ( .D(N408), .C(net12339), .Q(md3[2]) );
  DFFQX1 md5_s_reg_1_ ( .D(N485), .C(net12349), .Q(md5[1]) );
  DFFQX1 md0_s_reg_1_ ( .D(N192), .C(net12324), .Q(md0[1]) );
  OR2X1 U3 ( .A(n342), .B(n387), .Y(n3) );
  BUFX3 U4 ( .A(n185), .Y(n4) );
  INVX1 U5 ( .A(n94), .Y(n5) );
  INVX1 U6 ( .A(n136), .Y(n6) );
  NAND2X1 U7 ( .A(n357), .B(n435), .Y(n7) );
  NAND2X1 U8 ( .A(arg_c[0]), .B(n356), .Y(n8) );
  INVX1 U9 ( .A(n138), .Y(n9) );
  INVX1 U10 ( .A(n358), .Y(n10) );
  BUFX3 U11 ( .A(n393), .Y(n11) );
  INVX1 U12 ( .A(n92), .Y(n12) );
  INVX1 U13 ( .A(n85), .Y(n13) );
  INVX1 U14 ( .A(n357), .Y(n14) );
  NAND2X1 U15 ( .A(n435), .B(sum[17]), .Y(n15) );
  NAND2X1 U16 ( .A(n341), .B(n223), .Y(n16) );
  BUFX3 U17 ( .A(n83), .Y(n17) );
  INVX1 U18 ( .A(n334), .Y(n18) );
  INVX1 U19 ( .A(n56), .Y(n19) );
  INVX1 U20 ( .A(sum[17]), .Y(n20) );
  INVX1 U21 ( .A(n219), .Y(n21) );
  OAI222XL U22 ( .A(counter_st[1]), .B(n269), .C(n268), .D(n266), .E(n262), 
        .F(n283), .Y(n272) );
  NOR4XL U23 ( .A(counter_st[1]), .B(counter_st[2]), .C(counter_st[3]), .D(
        counter_st[4]), .Y(n336) );
  NOR3XL U24 ( .A(n360), .B(n361), .C(n362), .Y(n245) );
  INVX1 U25 ( .A(n190), .Y(n131) );
  INVX1 U28 ( .A(n205), .Y(n181) );
  INVX1 U29 ( .A(n187), .Y(n159) );
  INVX1 U30 ( .A(n186), .Y(n179) );
  INVX1 U31 ( .A(n345), .Y(n130) );
  NOR2X1 U32 ( .A(n363), .B(n359), .Y(n242) );
  INVX1 U33 ( .A(n317), .Y(n360) );
  INVX1 U34 ( .A(n364), .Y(n362) );
  INVX1 U35 ( .A(n339), .Y(n361) );
  INVX1 U36 ( .A(n386), .Y(n363) );
  INVX1 U37 ( .A(n299), .Y(n29) );
  INVX1 U38 ( .A(n337), .Y(n433) );
  AOI21X1 U39 ( .B(n436), .C(n267), .A(n291), .Y(n338) );
  INVX1 U40 ( .A(n384), .Y(n431) );
  INVX1 U41 ( .A(n299), .Y(n30) );
  NOR32XL U42 ( .B(n338), .C(n340), .A(n341), .Y(n318) );
  INVX1 U43 ( .A(n341), .Y(n128) );
  AND3X1 U44 ( .A(n388), .B(n296), .C(n337), .Y(n340) );
  INVX1 U45 ( .A(n264), .Y(n435) );
  INVX1 U46 ( .A(n291), .Y(n430) );
  NAND2X1 U47 ( .A(n358), .B(n435), .Y(n256) );
  NOR2X1 U48 ( .A(n358), .B(n357), .Y(n265) );
  NAND2X1 U49 ( .A(n357), .B(n435), .Y(n257) );
  INVX1 U50 ( .A(n192), .Y(n27) );
  INVX1 U51 ( .A(n192), .Y(n28) );
  AO21X1 U52 ( .B(n134), .C(n362), .A(n133), .Y(n190) );
  NAND21X1 U53 ( .B(n243), .A(n47), .Y(n393) );
  NAND21X1 U54 ( .B(n231), .A(n277), .Y(n185) );
  NAND21X1 U55 ( .B(n364), .A(n277), .Y(n345) );
  NAND21X1 U56 ( .B(n317), .A(n277), .Y(n186) );
  AO21X1 U57 ( .B(n134), .C(n360), .A(n133), .Y(n205) );
  NAND21X1 U58 ( .B(n339), .A(n277), .Y(n187) );
  NAND21X1 U59 ( .B(n386), .A(n277), .Y(n367) );
  AO21X1 U60 ( .B(n134), .C(n359), .A(n133), .Y(n63) );
  AO21X1 U61 ( .B(n134), .C(n363), .A(n133), .Y(n106) );
  NAND21X1 U62 ( .B(n241), .A(n47), .Y(n77) );
  AOI31X1 U63 ( .A(n231), .B(n48), .C(n232), .D(n233), .Y(n201) );
  NAND32X1 U64 ( .B(n438), .C(n215), .A(n47), .Y(n391) );
  AOI21X1 U65 ( .B(n134), .C(n361), .A(n133), .Y(n22) );
  OAI21X1 U66 ( .B(n242), .C(n392), .A(n243), .Y(n189) );
  NOR2X1 U67 ( .A(n246), .B(n392), .Y(n241) );
  NAND4X1 U68 ( .A(n391), .B(n390), .C(n11), .D(n47), .Y(N104) );
  NAND2X1 U69 ( .A(n185), .B(n47), .Y(n183) );
  NAND3X1 U70 ( .A(n187), .B(n48), .C(n318), .Y(N332) );
  NAND3X1 U71 ( .A(n186), .B(n48), .C(n318), .Y(N405) );
  NAND3X1 U72 ( .A(n191), .B(n48), .C(n430), .Y(N453) );
  NAND3X1 U73 ( .A(n4), .B(n47), .C(n430), .Y(N483) );
  NAND3X1 U74 ( .A(n367), .B(n48), .C(n365), .Y(N190) );
  NAND3X1 U75 ( .A(n345), .B(n48), .C(n365), .Y(N258) );
  INVX1 U76 ( .A(n233), .Y(n134) );
  INVX1 U77 ( .A(n243), .Y(n215) );
  NAND2X1 U78 ( .A(n344), .B(sfraddr[0]), .Y(n339) );
  NAND2X1 U79 ( .A(n344), .B(n36), .Y(n364) );
  NAND3X1 U80 ( .A(n36), .B(n37), .C(n278), .Y(n317) );
  INVX1 U81 ( .A(n232), .Y(n395) );
  INVX1 U82 ( .A(n231), .Y(n359) );
  NAND4X1 U83 ( .A(sfraddr[0]), .B(n366), .C(n37), .D(n38), .Y(n386) );
  INVX1 U84 ( .A(sfraddr[0]), .Y(n36) );
  NAND3X1 U85 ( .A(n278), .B(n37), .C(sfraddr[0]), .Y(n246) );
  NAND2X1 U86 ( .A(n387), .B(n342), .Y(n388) );
  NOR2X1 U87 ( .A(n263), .B(n434), .Y(n387) );
  INVX1 U88 ( .A(n299), .Y(n432) );
  NAND3X1 U89 ( .A(n434), .B(n342), .C(n436), .Y(n337) );
  NOR3XL U90 ( .A(n434), .B(n436), .C(n342), .Y(n291) );
  INVX1 U91 ( .A(n343), .Y(n434) );
  INVX1 U92 ( .A(n255), .Y(n438) );
  NOR2X1 U93 ( .A(n342), .B(n343), .Y(n267) );
  NAND3X1 U94 ( .A(n342), .B(n263), .C(n343), .Y(n296) );
  NAND2X1 U95 ( .A(n342), .B(n263), .Y(n396) );
  INVX1 U96 ( .A(n263), .Y(n436) );
  NOR21XL U97 ( .B(n387), .A(n342), .Y(n341) );
  NAND21X1 U98 ( .B(n341), .A(n306), .Y(n384) );
  INVX1 U99 ( .A(n394), .Y(n262) );
  INVX1 U100 ( .A(n299), .Y(n203) );
  NAND2X1 U101 ( .A(n267), .B(n47), .Y(n264) );
  NAND21X1 U102 ( .B(n356), .A(arg_c[0]), .Y(n83) );
  INVX1 U103 ( .A(n332), .Y(n357) );
  INVX1 U104 ( .A(n331), .Y(n358) );
  INVX1 U105 ( .A(n192), .Y(n26) );
  NAND2X1 U106 ( .A(arg_c[0]), .B(n356), .Y(n195) );
  INVX1 U107 ( .A(n34), .Y(n31) );
  INVX1 U108 ( .A(n34), .Y(n32) );
  INVX1 U109 ( .A(n34), .Y(n33) );
  NOR2X1 U110 ( .A(rst), .B(sfrwe), .Y(n233) );
  INVX1 U111 ( .A(n49), .Y(n133) );
  NAND21X1 U112 ( .B(n233), .A(rst), .Y(n49) );
  NAND21X1 U113 ( .B(rst), .A(n241), .Y(n191) );
  OR3XL U114 ( .A(rst), .B(n215), .C(n406), .Y(n390) );
  NOR2X1 U115 ( .A(n392), .B(rst), .Y(n277) );
  INVX1 U116 ( .A(sfrwe), .Y(n392) );
  NAND2X1 U117 ( .A(sfrwe), .B(n395), .Y(n243) );
  AOI211X1 U118 ( .C(n238), .D(n239), .A(n240), .B(rst), .Y(N802) );
  EORX1 U119 ( .A(sfroe), .B(n244), .C(n245), .D(n392), .Y(n238) );
  NOR2X1 U120 ( .A(n241), .B(n189), .Y(n239) );
  NAND3X1 U121 ( .A(n245), .B(n246), .C(n242), .Y(n244) );
  AND3X1 U122 ( .A(n366), .B(n38), .C(sfraddr[1]), .Y(n344) );
  AND2X1 U123 ( .A(n366), .B(sfraddr[2]), .Y(n278) );
  NAND3X1 U124 ( .A(n278), .B(n36), .C(sfraddr[1]), .Y(n231) );
  NAND3X1 U125 ( .A(sfraddr[0]), .B(n278), .C(sfraddr[1]), .Y(n232) );
  INVX1 U126 ( .A(sfraddr[1]), .Y(n37) );
  INVX1 U127 ( .A(sfraddr[2]), .Y(n38) );
  INVX1 U128 ( .A(sfrdatai[1]), .Y(n40) );
  INVX1 U129 ( .A(sfrdatai[0]), .Y(n39) );
  INVX1 U130 ( .A(sfrdatai[4]), .Y(n43) );
  INVX1 U131 ( .A(sfrdatai[3]), .Y(n42) );
  INVX1 U132 ( .A(sfrdatai[2]), .Y(n41) );
  INVX1 U133 ( .A(sfrdatai[7]), .Y(n46) );
  INVX1 U134 ( .A(sfrdatai[6]), .Y(n45) );
  INVX1 U135 ( .A(sfrdatai[5]), .Y(n44) );
  NOR2X1 U136 ( .A(n368), .B(n388), .Y(n299) );
  NAND2X1 U137 ( .A(n398), .B(n206), .Y(n263) );
  NOR42XL U138 ( .C(n401), .D(n212), .A(n437), .B(n166), .Y(n398) );
  INVX1 U139 ( .A(n266), .Y(n273) );
  NOR32XL U140 ( .B(n401), .C(n227), .A(n254), .Y(n343) );
  NAND21X1 U141 ( .B(n388), .A(n368), .Y(n306) );
  NAND4X1 U142 ( .A(n401), .B(n438), .C(n206), .D(n167), .Y(n342) );
  NAND2X1 U143 ( .A(n235), .B(n227), .Y(n255) );
  INVX1 U144 ( .A(n138), .Y(n194) );
  NAND21X1 U145 ( .B(n294), .A(n137), .Y(n138) );
  NAND3X1 U146 ( .A(n212), .B(n206), .C(n210), .Y(n254) );
  INVX1 U147 ( .A(n167), .Y(n437) );
  AND4X1 U148 ( .A(n398), .B(n438), .C(n210), .D(n214), .Y(n394) );
  AND3X1 U149 ( .A(n302), .B(n340), .C(n3), .Y(n365) );
  INVX1 U150 ( .A(rst), .Y(n47) );
  INVX1 U151 ( .A(n206), .Y(n439) );
  INVX1 U152 ( .A(rst), .Y(n48) );
  OAI22X1 U153 ( .A(n209), .B(n210), .C(n218), .D(n227), .Y(n225) );
  INVX1 U154 ( .A(n248), .Y(n279) );
  OAI31XL U155 ( .A(n253), .B(n254), .C(n255), .D(n48), .Y(n248) );
  NAND2X1 U156 ( .A(n214), .B(n167), .Y(n253) );
  INVX1 U157 ( .A(n214), .Y(n441) );
  NAND21X1 U158 ( .B(sum1[17]), .A(n89), .Y(n332) );
  NAND21X1 U159 ( .B(sum[17]), .A(sum1[17]), .Y(n331) );
  INVX1 U160 ( .A(sum[17]), .Y(n89) );
  INVX1 U161 ( .A(sum1[17]), .Y(n356) );
  OAI21BX1 U162 ( .C(sum[2]), .B(n15), .A(n260), .Y(N567) );
  AOI32X1 U163 ( .A(n435), .B(n357), .C(n335), .D(sum1[1]), .E(n334), .Y(n260)
         );
  OAI22X1 U164 ( .A(n436), .B(n333), .C(n263), .D(n350), .Y(n335) );
  INVX1 U165 ( .A(n256), .Y(n334) );
  INVX1 U166 ( .A(n192), .Y(n87) );
  NAND2X1 U167 ( .A(n435), .B(sum[17]), .Y(n258) );
  OAI22X1 U168 ( .A(n197), .B(n333), .C(n350), .D(n74), .Y(n81) );
  OAI222XL U169 ( .A(n415), .B(n256), .C(n461), .D(n257), .E(n258), .F(n371), 
        .Y(N581) );
  OAI222XL U170 ( .A(n417), .B(n256), .C(n460), .D(n7), .E(n15), .F(n373), .Y(
        N579) );
  OAI222XL U171 ( .A(n419), .B(n256), .C(n459), .D(n257), .E(n258), .F(n375), 
        .Y(N577) );
  OAI222XL U172 ( .A(n421), .B(n256), .C(n458), .D(n7), .E(n15), .F(n377), .Y(
        N575) );
  OAI222XL U173 ( .A(n423), .B(n256), .C(n457), .D(n257), .E(n258), .F(n379), 
        .Y(N573) );
  OAI222XL U174 ( .A(n425), .B(n256), .C(n456), .D(n7), .E(n15), .F(n381), .Y(
        N571) );
  OAI222XL U175 ( .A(n427), .B(n256), .C(n455), .D(n257), .E(n258), .F(n383), 
        .Y(N569) );
  OAI222XL U176 ( .A(n416), .B(n256), .C(n451), .D(n7), .E(n15), .F(n372), .Y(
        N580) );
  OAI222XL U177 ( .A(n418), .B(n256), .C(n450), .D(n257), .E(n258), .F(n374), 
        .Y(N578) );
  OAI222XL U178 ( .A(n420), .B(n18), .C(n449), .D(n7), .E(n15), .F(n376), .Y(
        N576) );
  OAI222XL U179 ( .A(n422), .B(n18), .C(n448), .D(n257), .E(n258), .F(n378), 
        .Y(N574) );
  OAI222XL U180 ( .A(n424), .B(n18), .C(n447), .D(n7), .E(n15), .F(n380), .Y(
        N572) );
  OAI222XL U181 ( .A(n426), .B(n18), .C(n446), .D(n257), .E(n258), .F(n382), 
        .Y(N570) );
  OAI222XL U182 ( .A(n428), .B(n18), .C(n443), .D(n7), .E(n15), .F(n385), .Y(
        N568) );
  OAI22X1 U183 ( .A(n62), .B(n63), .C(n185), .D(n40), .Y(N485) );
  OA222X1 U184 ( .A(n377), .B(n89), .C(n421), .D(n331), .E(n458), .F(n332), 
        .Y(n62) );
  OAI22X1 U185 ( .A(n60), .B(n63), .C(n185), .D(n42), .Y(N487) );
  OA222X1 U186 ( .A(n375), .B(n89), .C(n419), .D(n331), .E(n459), .F(n332), 
        .Y(n60) );
  OAI22X1 U187 ( .A(n58), .B(n63), .C(n185), .D(n44), .Y(N489) );
  OA222X1 U188 ( .A(n373), .B(n20), .C(n417), .D(n10), .E(n460), .F(n332), .Y(
        n58) );
  OAI22X1 U189 ( .A(n55), .B(n63), .C(n185), .D(n46), .Y(N491) );
  OA222X1 U190 ( .A(n371), .B(n20), .C(n415), .D(n10), .E(n461), .F(n14), .Y(
        n55) );
  OAI22X1 U191 ( .A(n64), .B(n63), .C(n4), .D(n39), .Y(N484) );
  OA222X1 U192 ( .A(n378), .B(n20), .C(n422), .D(n10), .E(n448), .F(n14), .Y(
        n64) );
  OAI22X1 U193 ( .A(n61), .B(n63), .C(n4), .D(n41), .Y(N486) );
  OA222X1 U194 ( .A(n376), .B(n20), .C(n420), .D(n10), .E(n449), .F(n14), .Y(
        n61) );
  OAI22X1 U195 ( .A(n59), .B(n63), .C(n4), .D(n43), .Y(N488) );
  OA222X1 U196 ( .A(n374), .B(n20), .C(n418), .D(n10), .E(n450), .F(n14), .Y(
        n59) );
  OAI22X1 U197 ( .A(n57), .B(n63), .C(n4), .D(n45), .Y(N490) );
  OA222X1 U198 ( .A(n372), .B(n20), .C(n416), .D(n10), .E(n451), .F(n14), .Y(
        n57) );
  OAI22X1 U199 ( .A(n72), .B(n77), .C(n191), .D(n40), .Y(N455) );
  OA222X1 U200 ( .A(n141), .B(n89), .C(n71), .D(n14), .E(n122), .F(n331), .Y(
        n72) );
  OA22X1 U201 ( .A(n74), .B(n350), .C(n200), .D(n333), .Y(n71) );
  OAI22X1 U202 ( .A(n69), .B(n77), .C(n191), .D(n42), .Y(N457) );
  OA222X1 U203 ( .A(n383), .B(n89), .C(n427), .D(n331), .E(n455), .F(n332), 
        .Y(n69) );
  OAI22X1 U204 ( .A(n67), .B(n77), .C(n191), .D(n44), .Y(N459) );
  OA222X1 U205 ( .A(n381), .B(n89), .C(n425), .D(n331), .E(n456), .F(n332), 
        .Y(n67) );
  OAI22X1 U206 ( .A(n65), .B(n77), .C(n191), .D(n46), .Y(N461) );
  OA222X1 U207 ( .A(n379), .B(n89), .C(n423), .D(n331), .E(n457), .F(n332), 
        .Y(n65) );
  OAI22X1 U208 ( .A(n68), .B(n77), .C(n191), .D(n43), .Y(N458) );
  OA222X1 U209 ( .A(n382), .B(n89), .C(n426), .D(n331), .E(n446), .F(n332), 
        .Y(n68) );
  OAI22X1 U210 ( .A(n66), .B(n77), .C(n191), .D(n45), .Y(N460) );
  OA222X1 U211 ( .A(n380), .B(n89), .C(n424), .D(n331), .E(n447), .F(n332), 
        .Y(n66) );
  OAI22X1 U212 ( .A(n51), .B(n205), .C(n186), .D(n46), .Y(N413) );
  OA2222XL U213 ( .A(n16), .B(n20), .C(n296), .D(n281), .E(n297), .F(n226), 
        .G(n196), .H(n50), .Y(n51) );
  INVX1 U214 ( .A(n294), .Y(n50) );
  OAI22X1 U215 ( .A(n70), .B(n77), .C(n191), .D(n41), .Y(N456) );
  OA222X1 U216 ( .A(n385), .B(n89), .C(n428), .D(n331), .E(n443), .F(n332), 
        .Y(n70) );
  OAI22X1 U217 ( .A(n90), .B(n106), .C(n367), .D(n39), .Y(N191) );
  OA222X1 U218 ( .A(n3), .B(n20), .C(n99), .D(n431), .E(n203), .F(n97), .Y(n90) );
  INVX1 U219 ( .A(n384), .Y(n88) );
  INVX1 U220 ( .A(arg_a[0]), .Y(n34) );
  INVX1 U221 ( .A(n200), .Y(n74) );
  INVX1 U222 ( .A(sum[15]), .Y(n372) );
  INVX1 U223 ( .A(sum[16]), .Y(n371) );
  AO22X1 U224 ( .A(n181), .B(n180), .C(sfrdatai[5]), .D(n179), .Y(N411) );
  OAI221X1 U225 ( .A(n30), .B(n226), .C(n302), .D(n372), .E(n178), .Y(n180) );
  OA222X1 U226 ( .A(n306), .B(n350), .C(n199), .D(n193), .E(n194), .F(n307), 
        .Y(n178) );
  OAI22X1 U227 ( .A(n207), .B(n205), .C(n186), .D(n45), .Y(N412) );
  OA2222XL U228 ( .A(n350), .B(n203), .C(n302), .D(n371), .E(n6), .F(n196), 
        .G(n9), .H(n193), .Y(n207) );
  INVX1 U229 ( .A(arg_a[0]), .Y(n35) );
  INVX1 U230 ( .A(sum[14]), .Y(n373) );
  AO22X1 U231 ( .A(n181), .B(n177), .C(sfrdatai[4]), .D(n179), .Y(N410) );
  OAI221X1 U232 ( .A(n30), .B(n196), .C(n16), .D(n373), .E(n176), .Y(n177) );
  OA222X1 U233 ( .A(n306), .B(n226), .C(n6), .D(n307), .E(n9), .F(n175), .Y(
        n176) );
  INVX1 U234 ( .A(sum[12]), .Y(n375) );
  INVX1 U235 ( .A(sum[13]), .Y(n374) );
  AO22X1 U236 ( .A(n181), .B(n174), .C(sfrdatai[3]), .D(n179), .Y(N409) );
  OAI221X1 U237 ( .A(n21), .B(n196), .C(n302), .D(n374), .E(n173), .Y(n174) );
  OA222X1 U238 ( .A(n29), .B(n193), .C(n6), .D(n175), .E(n9), .F(n304), .Y(
        n173) );
  AO22X1 U239 ( .A(n181), .B(n172), .C(sfrdatai[2]), .D(n179), .Y(N408) );
  OAI221X1 U240 ( .A(n30), .B(n307), .C(n16), .D(n375), .E(n170), .Y(n172) );
  OA222X1 U241 ( .A(n306), .B(n193), .C(n6), .D(n304), .E(n9), .F(n169), .Y(
        n170) );
  INVX1 U242 ( .A(sum[11]), .Y(n376) );
  AO22X1 U243 ( .A(n181), .B(n168), .C(sfrdatai[1]), .D(n179), .Y(N407) );
  OAI221X1 U244 ( .A(n21), .B(n307), .C(n16), .D(n376), .E(n165), .Y(n168) );
  OA222X1 U245 ( .A(n29), .B(n175), .C(n199), .D(n169), .E(n194), .F(n164), 
        .Y(n165) );
  INVX1 U246 ( .A(sum[10]), .Y(n377) );
  INVX1 U247 ( .A(sum[9]), .Y(n378) );
  AO22X1 U248 ( .A(n181), .B(n163), .C(sfrdatai[0]), .D(n179), .Y(N406) );
  OAI221X1 U249 ( .A(n30), .B(n304), .C(n302), .D(n377), .E(n162), .Y(n163) );
  OA222X1 U250 ( .A(n306), .B(n175), .C(n6), .D(n164), .E(n9), .F(n161), .Y(
        n162) );
  AO22X1 U251 ( .A(n22), .B(n160), .C(sfrdatai[7]), .D(n159), .Y(N340) );
  OAI221X1 U252 ( .A(n21), .B(n304), .C(n16), .D(n378), .E(n158), .Y(n160) );
  OA222X1 U253 ( .A(n29), .B(n169), .C(n199), .D(n161), .E(n194), .F(n301), 
        .Y(n158) );
  INVX1 U254 ( .A(sum[8]), .Y(n379) );
  AO22X1 U255 ( .A(n22), .B(n157), .C(sfrdatai[6]), .D(n159), .Y(N339) );
  OAI221X1 U256 ( .A(n30), .B(n164), .C(n16), .D(n379), .E(n156), .Y(n157) );
  OA222X1 U257 ( .A(n306), .B(n169), .C(n199), .D(n301), .E(n194), .F(n155), 
        .Y(n156) );
  INVX1 U258 ( .A(sum[6]), .Y(n381) );
  INVX1 U259 ( .A(sum[7]), .Y(n380) );
  AO22X1 U260 ( .A(n22), .B(n152), .C(sfrdatai[4]), .D(n159), .Y(N337) );
  OAI221X1 U261 ( .A(n30), .B(n301), .C(n16), .D(n381), .E(n151), .Y(n152) );
  OA222X1 U262 ( .A(n306), .B(n161), .C(n199), .D(n303), .E(n194), .F(n150), 
        .Y(n151) );
  AO22X1 U263 ( .A(n22), .B(n154), .C(sfrdatai[5]), .D(n159), .Y(N338) );
  OAI221X1 U264 ( .A(n21), .B(n164), .C(n302), .D(n380), .E(n153), .Y(n154) );
  OA222X1 U265 ( .A(n29), .B(n161), .C(n199), .D(n155), .E(n194), .F(n303), 
        .Y(n153) );
  INVX1 U266 ( .A(sum[5]), .Y(n382) );
  AO22X1 U267 ( .A(n22), .B(n149), .C(sfrdatai[3]), .D(n159), .Y(N336) );
  OAI221X1 U268 ( .A(n21), .B(n301), .C(n302), .D(n382), .E(n148), .Y(n149) );
  OA222X1 U269 ( .A(n29), .B(n155), .C(n199), .D(n150), .E(n194), .F(n147), 
        .Y(n148) );
  INVX1 U270 ( .A(sum1[3]), .Y(n427) );
  INVX1 U271 ( .A(sum1[4]), .Y(n426) );
  INVX1 U272 ( .A(sum1[5]), .Y(n425) );
  INVX1 U273 ( .A(sum1[6]), .Y(n424) );
  INVX1 U274 ( .A(sum1[7]), .Y(n423) );
  INVX1 U275 ( .A(sum1[8]), .Y(n422) );
  INVX1 U276 ( .A(sum1[9]), .Y(n421) );
  INVX1 U277 ( .A(sum1[10]), .Y(n420) );
  INVX1 U278 ( .A(sum1[11]), .Y(n419) );
  INVX1 U279 ( .A(sum1[12]), .Y(n418) );
  INVX1 U280 ( .A(sum1[13]), .Y(n417) );
  INVX1 U281 ( .A(sum1[14]), .Y(n416) );
  INVX1 U282 ( .A(sum1[15]), .Y(n415) );
  INVX1 U283 ( .A(sum1[2]), .Y(n428) );
  INVX1 U284 ( .A(sum[4]), .Y(n383) );
  INVX1 U285 ( .A(sum[3]), .Y(n385) );
  AO22X1 U286 ( .A(n22), .B(n146), .C(sfrdatai[2]), .D(n159), .Y(N335) );
  OAI221X1 U287 ( .A(n30), .B(n303), .C(n16), .D(n383), .E(n145), .Y(n146) );
  OA222X1 U288 ( .A(n306), .B(n155), .C(n199), .D(n147), .E(n194), .F(n305), 
        .Y(n145) );
  AO22X1 U289 ( .A(n22), .B(n144), .C(sfrdatai[1]), .D(n159), .Y(N334) );
  OAI221X1 U290 ( .A(n21), .B(n303), .C(n302), .D(n385), .E(n143), .Y(n144) );
  OA222X1 U291 ( .A(n29), .B(n150), .C(n199), .D(n305), .E(n194), .F(n333), 
        .Y(n143) );
  INVX1 U292 ( .A(sum1[1]), .Y(n122) );
  INVX1 U293 ( .A(sum[2]), .Y(n141) );
  AO22X1 U294 ( .A(n123), .B(n131), .C(sfrdatai[6]), .D(n130), .Y(N265) );
  OAI221X1 U295 ( .A(n30), .B(n333), .C(n122), .D(n128), .E(n121), .Y(n123) );
  OA222X1 U296 ( .A(n21), .B(n305), .C(n126), .D(n124), .E(n125), .F(n120), 
        .Y(n121) );
  AO22X1 U297 ( .A(n132), .B(n131), .C(sfrdatai[7]), .D(n130), .Y(N266) );
  OAI221X1 U298 ( .A(n21), .B(n147), .C(n129), .D(n128), .E(n127), .Y(n132) );
  OA222X1 U299 ( .A(n29), .B(n305), .C(n126), .D(n139), .E(n125), .F(n124), 
        .Y(n127) );
  INVX1 U300 ( .A(sum[1]), .Y(n129) );
  AO22X1 U301 ( .A(n22), .B(n142), .C(sfrdatai[0]), .D(n159), .Y(N333) );
  OAI221X1 U302 ( .A(n30), .B(n147), .C(n302), .D(n141), .E(n140), .Y(n142) );
  OA222X1 U303 ( .A(n306), .B(n150), .C(n199), .D(n333), .E(n194), .F(n139), 
        .Y(n140) );
  OAI22X1 U304 ( .A(n190), .B(n119), .C(n345), .D(n44), .Y(N264) );
  OA2222XL U305 ( .A(n29), .B(n139), .C(n88), .D(n333), .E(n126), .F(n120), 
        .G(n125), .H(n118), .Y(n119) );
  OAI22X1 U306 ( .A(n190), .B(n117), .C(n345), .D(n43), .Y(N263) );
  OA2222XL U307 ( .A(n88), .B(n139), .C(n29), .D(n124), .E(n126), .F(n118), 
        .G(n125), .H(n116), .Y(n117) );
  OAI22X1 U308 ( .A(n190), .B(n115), .C(n345), .D(n42), .Y(N262) );
  OA2222XL U309 ( .A(n431), .B(n124), .C(n203), .D(n120), .E(n126), .F(n116), 
        .G(n125), .H(n114), .Y(n115) );
  OAI22X1 U310 ( .A(n190), .B(n113), .C(n345), .D(n41), .Y(N261) );
  OA2222XL U311 ( .A(n88), .B(n120), .C(n203), .D(n118), .E(n126), .F(n114), 
        .G(n125), .H(n112), .Y(n113) );
  OAI22X1 U312 ( .A(n190), .B(n111), .C(n345), .D(n40), .Y(N260) );
  OA2222XL U313 ( .A(n431), .B(n118), .C(n203), .D(n116), .E(n126), .F(n112), 
        .G(n125), .H(n110), .Y(n111) );
  OAI22X1 U314 ( .A(n190), .B(n109), .C(n345), .D(n39), .Y(N259) );
  OA2222XL U315 ( .A(n88), .B(n116), .C(n203), .D(n114), .E(n126), .F(n110), 
        .G(n125), .H(n108), .Y(n109) );
  OAI222XL U316 ( .A(n390), .B(n276), .C(n391), .D(n275), .E(n393), .F(n41), 
        .Y(N107) );
  INVX1 U317 ( .A(n280), .Y(n275) );
  OAI222XL U318 ( .A(n390), .B(n247), .C(n391), .D(n234), .E(n393), .F(n43), 
        .Y(N109) );
  INVX1 U319 ( .A(n249), .Y(n234) );
  OAI222XL U320 ( .A(n390), .B(n251), .C(n391), .D(n250), .E(n393), .F(n42), 
        .Y(N108) );
  INVX1 U321 ( .A(n252), .Y(n250) );
  OAI222XL U322 ( .A(n393), .B(n40), .C(n391), .D(n271), .E(n390), .F(n270), 
        .Y(N106) );
  INVX1 U323 ( .A(n272), .Y(n271) );
  OAI222XL U324 ( .A(n393), .B(n39), .C(n391), .D(n259), .E(n355), .F(n390), 
        .Y(N105) );
  INVX1 U325 ( .A(n261), .Y(n259) );
  OAI221X1 U326 ( .A(n185), .B(n397), .C(n183), .D(n429), .E(n393), .Y(n412)
         );
  OAI22X1 U327 ( .A(n107), .B(n106), .C(n367), .D(n46), .Y(N198) );
  OA2222XL U328 ( .A(n431), .B(n114), .C(n203), .D(n112), .E(n126), .F(n108), 
        .G(n125), .H(n105), .Y(n107) );
  OAI22X1 U329 ( .A(n104), .B(n106), .C(n367), .D(n45), .Y(N197) );
  OA2222XL U330 ( .A(n88), .B(n112), .C(n203), .D(n110), .E(n126), .F(n105), 
        .G(n125), .H(n103), .Y(n104) );
  OAI22X1 U331 ( .A(n102), .B(n106), .C(n367), .D(n44), .Y(N196) );
  OA2222XL U332 ( .A(n431), .B(n110), .C(n203), .D(n108), .E(n12), .F(n103), 
        .G(n5), .H(n101), .Y(n102) );
  OAI22X1 U333 ( .A(n100), .B(n106), .C(n367), .D(n43), .Y(N195) );
  OA2222XL U334 ( .A(n88), .B(n108), .C(n30), .D(n105), .E(n12), .F(n101), .G(
        n5), .H(n99), .Y(n100) );
  OAI22X1 U335 ( .A(n98), .B(n106), .C(n367), .D(n42), .Y(N194) );
  OA2222XL U336 ( .A(n431), .B(n105), .C(n432), .D(n103), .E(n12), .F(n99), 
        .G(n5), .H(n97), .Y(n98) );
  OAI22X1 U337 ( .A(n96), .B(n106), .C(n367), .D(n41), .Y(N193) );
  OA2222XL U338 ( .A(n88), .B(n103), .C(n432), .D(n101), .E(n12), .F(n97), .G(
        n5), .H(n95), .Y(n96) );
  OAI22X1 U339 ( .A(n93), .B(n106), .C(n367), .D(n40), .Y(N192) );
  OA2222XL U340 ( .A(n203), .B(n99), .C(n356), .D(n3), .E(n12), .F(n95), .G(
        n431), .H(n101), .Y(n93) );
  OAI211X1 U341 ( .C(n201), .D(n202), .A(n185), .B(n393), .Y(N895) );
  AOI211X1 U342 ( .C(n437), .D(n353), .A(n352), .B(n204), .Y(n202) );
  OAI32X1 U343 ( .A(n206), .B(n351), .C(n350), .D(n87), .E(n208), .Y(n352) );
  OAI222XL U344 ( .A(n209), .B(n210), .C(n211), .D(n212), .E(n213), .F(n214), 
        .Y(n204) );
  OAI211X1 U345 ( .C(n201), .D(n289), .A(n185), .B(n11), .Y(N894) );
  AOI211X1 U346 ( .C(n255), .D(n288), .A(n287), .B(n217), .Y(n289) );
  INVX1 U347 ( .A(n218), .Y(n288) );
  OA21X1 U348 ( .B(n300), .C(n298), .A(n295), .Y(N892) );
  OAI22X1 U349 ( .A(n212), .B(n290), .C(n208), .D(n200), .Y(n300) );
  OAI211X1 U350 ( .C(n348), .D(n293), .A(n229), .B(n292), .Y(n298) );
  INVX1 U351 ( .A(n201), .Y(n295) );
  NAND2X1 U352 ( .A(n197), .B(n74), .Y(arg_c[0]) );
  NOR43XL U353 ( .B(n208), .C(n406), .D(n407), .A(n240), .Y(n401) );
  NOR21XL U354 ( .B(n171), .A(n354), .Y(n407) );
  INVX1 U355 ( .A(n330), .Y(n354) );
  NAND21X1 U356 ( .B(n394), .A(n230), .Y(n266) );
  OAI211X1 U357 ( .C(n396), .D(n226), .A(n29), .B(n297), .Y(n230) );
  NAND2X1 U358 ( .A(n402), .B(n405), .Y(n171) );
  NAND2X1 U359 ( .A(n402), .B(n389), .Y(n330) );
  INVX1 U360 ( .A(n92), .Y(n126) );
  AO21X1 U361 ( .B(n336), .C(n433), .A(n135), .Y(n92) );
  OAI21X1 U362 ( .B(n336), .C(n337), .A(n338), .Y(n294) );
  NAND21X1 U363 ( .B(n296), .A(n226), .Y(n137) );
  INVX1 U364 ( .A(n94), .Y(n125) );
  OAI211X1 U365 ( .C(n336), .D(n337), .A(n3), .B(n137), .Y(n94) );
  NAND2X1 U366 ( .A(n403), .B(n404), .Y(n167) );
  NAND2X1 U367 ( .A(n399), .B(n389), .Y(n206) );
  OAI31XL U368 ( .A(n444), .B(n445), .C(n442), .D(mdubsy), .Y(n240) );
  NAND2X1 U369 ( .A(n399), .B(n405), .Y(mdubsy) );
  AND2X1 U370 ( .A(n400), .B(n402), .Y(n166) );
  INVX1 U371 ( .A(n136), .Y(n199) );
  NAND21X1 U372 ( .B(n135), .A(n297), .Y(n136) );
  NAND2X1 U373 ( .A(n404), .B(n402), .Y(n406) );
  NOR2X1 U374 ( .A(n440), .B(n442), .Y(n404) );
  AND2X1 U375 ( .A(n252), .B(n279), .Y(N677) );
  AND2X1 U376 ( .A(n249), .B(n279), .Y(N678) );
  AND2X1 U377 ( .A(n280), .B(n279), .Y(N676) );
  AND2X1 U378 ( .A(n261), .B(n279), .Y(N674) );
  AND2X1 U379 ( .A(n272), .B(n279), .Y(N675) );
  NAND2X1 U380 ( .A(n433), .B(n336), .Y(n297) );
  NAND2X1 U381 ( .A(n399), .B(n404), .Y(n212) );
  NAND2X1 U382 ( .A(n403), .B(n405), .Y(n210) );
  NAND2X1 U383 ( .A(n403), .B(n400), .Y(n227) );
  NAND2X1 U384 ( .A(n403), .B(n389), .Y(n235) );
  INVX1 U385 ( .A(n269), .Y(n274) );
  NAND2X1 U386 ( .A(n341), .B(n223), .Y(n302) );
  INVX1 U387 ( .A(n336), .Y(n368) );
  XOR2X1 U388 ( .A(n454), .B(n370), .Y(n251) );
  NAND2X1 U389 ( .A(n399), .B(n400), .Y(n214) );
  NAND2X1 U390 ( .A(n351), .B(n439), .Y(n348) );
  OA22X1 U391 ( .A(n235), .B(n218), .C(n214), .D(n213), .Y(n229) );
  NAND2X1 U392 ( .A(n368), .B(n237), .Y(n218) );
  NAND4X1 U393 ( .A(n355), .B(n452), .C(n454), .D(n453), .Y(n237) );
  INVX1 U394 ( .A(n84), .Y(n73) );
  INVX1 U395 ( .A(n308), .Y(n281) );
  NAND2X1 U396 ( .A(n228), .B(n453), .Y(n209) );
  INVX1 U397 ( .A(n347), .Y(n292) );
  NOR21XL U398 ( .B(n48), .A(n327), .Y(n408) );
  NOR32XL U399 ( .B(n171), .C(n326), .A(n325), .Y(n327) );
  NAND21X1 U400 ( .B(n330), .A(n312), .Y(n326) );
  MUX2IX1 U401 ( .D0(n324), .D1(n323), .S(n166), .Y(n325) );
  INVX1 U402 ( .A(n211), .Y(n290) );
  AND2X1 U403 ( .A(norm_reg[15]), .B(n31), .Y(arg_a[17]) );
  OAI22X1 U404 ( .A(n35), .B(n443), .C(n32), .D(n147), .Y(arg_a[2]) );
  MUX2X1 U405 ( .D0(n28), .D1(n79), .S(md4[1]), .Y(arg_b[2]) );
  OAI22X1 U406 ( .A(n34), .B(n455), .C(n32), .D(n150), .Y(arg_a[3]) );
  MUX2X1 U407 ( .D0(n28), .D1(n79), .S(md4[2]), .Y(arg_b[3]) );
  MUX2X1 U408 ( .D0(n26), .D1(n86), .S(md4[1]), .Y(arg_d[2]) );
  OAI222XL U409 ( .A(n122), .B(n83), .C(sum1[17]), .D(n82), .E(n31), .F(n427), 
        .Y(arg_c[2]) );
  INVX1 U410 ( .A(n81), .Y(n82) );
  OAI22X1 U411 ( .A(n34), .B(n446), .C(n33), .D(n303), .Y(arg_a[4]) );
  MUX2X1 U412 ( .D0(n28), .D1(n79), .S(md4[3]), .Y(arg_b[4]) );
  MUX2X1 U413 ( .D0(n27), .D1(n86), .S(md4[2]), .Y(arg_d[3]) );
  OAI222XL U414 ( .A(n195), .B(n443), .C(n428), .D(n83), .E(n31), .F(n426), 
        .Y(arg_c[3]) );
  OAI22X1 U415 ( .A(n35), .B(n456), .C(n33), .D(n155), .Y(arg_a[5]) );
  MUX2X1 U416 ( .D0(n28), .D1(n79), .S(md4[4]), .Y(arg_b[5]) );
  MUX2X1 U417 ( .D0(n26), .D1(n86), .S(md4[3]), .Y(arg_d[4]) );
  OAI222XL U418 ( .A(n8), .B(n455), .C(n427), .D(n83), .E(n31), .F(n425), .Y(
        arg_c[4]) );
  OAI22X1 U419 ( .A(n35), .B(n447), .C(n33), .D(n301), .Y(arg_a[6]) );
  MUX2X1 U420 ( .D0(n28), .D1(n79), .S(md4[5]), .Y(arg_b[6]) );
  MUX2X1 U421 ( .D0(n26), .D1(n86), .S(md4[4]), .Y(arg_d[5]) );
  OAI222XL U422 ( .A(n195), .B(n446), .C(n426), .D(n83), .E(n31), .F(n424), 
        .Y(arg_c[5]) );
  OAI22X1 U423 ( .A(n35), .B(n457), .C(n33), .D(n161), .Y(arg_a[7]) );
  MUX2X1 U424 ( .D0(n28), .D1(n79), .S(md4[6]), .Y(arg_b[7]) );
  MUX2X1 U425 ( .D0(n26), .D1(n86), .S(md4[5]), .Y(arg_d[6]) );
  OAI222XL U426 ( .A(n8), .B(n456), .C(n425), .D(n83), .E(n31), .F(n423), .Y(
        arg_c[6]) );
  OAI22X1 U427 ( .A(n35), .B(n448), .C(n33), .D(n164), .Y(arg_a[8]) );
  MUX2X1 U428 ( .D0(n28), .D1(n79), .S(md4[7]), .Y(arg_b[8]) );
  MUX2X1 U429 ( .D0(n26), .D1(n86), .S(md4[6]), .Y(arg_d[7]) );
  OAI222XL U430 ( .A(n195), .B(n447), .C(n424), .D(n83), .E(n31), .F(n422), 
        .Y(arg_c[7]) );
  OAI22X1 U431 ( .A(n35), .B(n458), .C(n33), .D(n169), .Y(arg_a[9]) );
  MUX2X1 U432 ( .D0(n28), .D1(n79), .S(md5[0]), .Y(arg_b[9]) );
  MUX2X1 U433 ( .D0(n26), .D1(n86), .S(md4[7]), .Y(arg_d[8]) );
  OAI222XL U434 ( .A(n8), .B(n457), .C(n423), .D(n83), .E(n31), .F(n421), .Y(
        arg_c[8]) );
  OAI22X1 U435 ( .A(n35), .B(n449), .C(n33), .D(n304), .Y(arg_a[10]) );
  MUX2X1 U436 ( .D0(n28), .D1(n79), .S(md5[1]), .Y(arg_b[10]) );
  MUX2X1 U437 ( .D0(n26), .D1(n86), .S(md5[0]), .Y(arg_d[9]) );
  OAI222XL U438 ( .A(n195), .B(n448), .C(n422), .D(n83), .E(n32), .F(n420), 
        .Y(arg_c[9]) );
  OAI22X1 U439 ( .A(n35), .B(n459), .C(n33), .D(n175), .Y(arg_a[11]) );
  MUX2X1 U440 ( .D0(n28), .D1(n19), .S(md5[2]), .Y(arg_b[11]) );
  MUX2X1 U441 ( .D0(n27), .D1(n86), .S(md5[1]), .Y(arg_d[10]) );
  OAI222XL U442 ( .A(n8), .B(n458), .C(n421), .D(n83), .E(n32), .F(n419), .Y(
        arg_c[10]) );
  OAI22X1 U443 ( .A(n35), .B(n450), .C(n33), .D(n307), .Y(arg_a[12]) );
  MUX2X1 U444 ( .D0(n87), .D1(n19), .S(md5[3]), .Y(arg_b[12]) );
  MUX2X1 U445 ( .D0(n27), .D1(n13), .S(md5[2]), .Y(arg_d[11]) );
  OAI222XL U446 ( .A(n195), .B(n449), .C(n420), .D(n17), .E(n32), .F(n418), 
        .Y(arg_c[11]) );
  OAI22X1 U447 ( .A(n35), .B(n460), .C(n33), .D(n193), .Y(arg_a[13]) );
  MUX2X1 U448 ( .D0(n87), .D1(n19), .S(md5[4]), .Y(arg_b[13]) );
  MUX2X1 U449 ( .D0(n27), .D1(n13), .S(md5[3]), .Y(arg_d[12]) );
  OAI222XL U450 ( .A(n8), .B(n459), .C(n419), .D(n17), .E(n32), .F(n417), .Y(
        arg_c[12]) );
  OAI22X1 U451 ( .A(n34), .B(n451), .C(arg_a[0]), .D(n196), .Y(arg_a[14]) );
  MUX2X1 U452 ( .D0(n87), .D1(n19), .S(md5[5]), .Y(arg_b[14]) );
  MUX2X1 U453 ( .D0(n27), .D1(n13), .S(md5[4]), .Y(arg_d[13]) );
  OAI222XL U454 ( .A(n195), .B(n450), .C(n418), .D(n17), .E(n32), .F(n416), 
        .Y(arg_c[13]) );
  OAI22X1 U455 ( .A(n34), .B(n461), .C(arg_a[0]), .D(n226), .Y(arg_a[15]) );
  MUX2X1 U456 ( .D0(n87), .D1(n19), .S(md5[6]), .Y(arg_b[15]) );
  MUX2X1 U457 ( .D0(n27), .D1(n13), .S(md5[5]), .Y(arg_d[14]) );
  OAI222XL U458 ( .A(n8), .B(n460), .C(n417), .D(n17), .E(n32), .F(n415), .Y(
        arg_c[14]) );
  MUX2X1 U459 ( .D0(n27), .D1(n13), .S(md5[6]), .Y(arg_d[15]) );
  OAI222XL U460 ( .A(n195), .B(n451), .C(n416), .D(n17), .E(n32), .F(n80), .Y(
        arg_c[15]) );
  INVX1 U461 ( .A(sum1[16]), .Y(n80) );
  MUX2X1 U462 ( .D0(md3[7]), .D1(norm_reg[14]), .S(n31), .Y(arg_a[16]) );
  MUX2X1 U463 ( .D0(n26), .D1(n19), .S(md5[7]), .Y(arg_b[16]) );
  MUX2X1 U464 ( .D0(n27), .D1(n13), .S(md5[7]), .Y(arg_d[16]) );
  OAI222XL U465 ( .A(n8), .B(n461), .C(n415), .D(n17), .E(n32), .F(n356), .Y(
        arg_c[16]) );
  NOR21XL U466 ( .B(arg_c[0]), .A(n198), .Y(arg_c[17]) );
  AOI22X1 U467 ( .A(norm_reg[14]), .B(n356), .C(sum1[16]), .D(sum1[17]), .Y(
        n198) );
  NOR2X1 U468 ( .A(mdu_op[0]), .B(mdu_op[1]), .Y(n192) );
  AO21X1 U469 ( .B(md2[0]), .C(n34), .A(n81), .Y(arg_a[1]) );
  MUX2X1 U470 ( .D0(n27), .D1(n79), .S(md4[0]), .Y(arg_b[1]) );
  INVX1 U471 ( .A(n56), .Y(n79) );
  NAND21X1 U472 ( .B(n26), .A(md0[0]), .Y(n56) );
  OAI22X1 U473 ( .A(n78), .B(n77), .C(n191), .D(n39), .Y(N454) );
  AOI22X1 U474 ( .A(n76), .B(n75), .C(sum[17]), .D(sum[1]), .Y(n78) );
  AO21X1 U475 ( .B(md1[6]), .C(n74), .A(n73), .Y(n76) );
  INVX1 U476 ( .A(n265), .Y(n75) );
  NOR2X1 U477 ( .A(n429), .B(mdu_op[0]), .Y(n200) );
  AOI21X1 U478 ( .B(mdu_op[0]), .C(mdu_op[1]), .A(n192), .Y(arg_a[0]) );
  NAND21X1 U479 ( .B(n54), .A(n53), .Y(N566) );
  NOR21XL U480 ( .B(sum[1]), .A(n258), .Y(n54) );
  NAND32X1 U481 ( .B(n264), .C(n265), .A(n52), .Y(n53) );
  AO22X1 U482 ( .A(md1[6]), .B(n263), .C(md3[6]), .D(n436), .Y(n52) );
  NAND2X1 U483 ( .A(mdu_op[0]), .B(n429), .Y(n197) );
  INVX1 U484 ( .A(mdu_op[1]), .Y(n429) );
  INVX1 U485 ( .A(md3[7]), .Y(n350) );
  INVX1 U486 ( .A(md1[7]), .Y(n333) );
  INVX1 U487 ( .A(md2[1]), .Y(n147) );
  INVX1 U488 ( .A(norm_reg[0]), .Y(n443) );
  INVX1 U489 ( .A(md2[3]), .Y(n303) );
  INVX1 U490 ( .A(md2[2]), .Y(n150) );
  INVX1 U491 ( .A(norm_reg[1]), .Y(n455) );
  INVX1 U492 ( .A(norm_reg[2]), .Y(n446) );
  INVX1 U493 ( .A(md2[4]), .Y(n155) );
  INVX1 U494 ( .A(norm_reg[3]), .Y(n456) );
  INVX1 U495 ( .A(md2[5]), .Y(n301) );
  INVX1 U496 ( .A(md2[6]), .Y(n161) );
  INVX1 U497 ( .A(norm_reg[4]), .Y(n447) );
  INVX1 U498 ( .A(norm_reg[5]), .Y(n457) );
  INVX1 U499 ( .A(md2[7]), .Y(n164) );
  INVX1 U500 ( .A(norm_reg[6]), .Y(n448) );
  INVX1 U501 ( .A(md3[1]), .Y(n304) );
  INVX1 U502 ( .A(md3[0]), .Y(n169) );
  INVX1 U503 ( .A(norm_reg[7]), .Y(n458) );
  INVX1 U504 ( .A(norm_reg[8]), .Y(n449) );
  INVX1 U505 ( .A(md3[2]), .Y(n175) );
  INVX1 U506 ( .A(norm_reg[9]), .Y(n459) );
  MUX2X1 U507 ( .D0(n27), .D1(n86), .S(md4[0]), .Y(arg_d[1]) );
  OAI221X1 U508 ( .A(n197), .B(n139), .C(arg_a[0]), .D(n428), .E(n84), .Y(
        arg_c[1]) );
  INVX1 U509 ( .A(md3[3]), .Y(n307) );
  INVX1 U510 ( .A(md3[4]), .Y(n193) );
  INVX1 U511 ( .A(norm_reg[10]), .Y(n450) );
  INVX1 U512 ( .A(norm_reg[11]), .Y(n460) );
  OAI21BX1 U513 ( .C(set_div16), .B(n190), .A(n191), .Y(n414) );
  INVX1 U514 ( .A(md3[5]), .Y(n196) );
  INVX1 U515 ( .A(norm_reg[12]), .Y(n451) );
  NAND3X1 U516 ( .A(n186), .B(n187), .C(n188), .Y(n413) );
  NAND31X1 U517 ( .C(n189), .A(n47), .B(set_div32), .Y(n188) );
  INVX1 U518 ( .A(md3[6]), .Y(n226) );
  MUX2BXL U519 ( .D0(sfrdatai[5]), .D1(n23), .S(n393), .Y(n409) );
  NAND2X1 U520 ( .A(arcon[5]), .B(n47), .Y(n23) );
  OAI2B11X1 U521 ( .D(mdu_op[0]), .C(n183), .A(n184), .B(n393), .Y(n411) );
  NAND31X1 U522 ( .C(n185), .A(n397), .B(set_div16), .Y(n184) );
  AOI21X1 U523 ( .B(n221), .C(n222), .A(n201), .Y(N893) );
  AND3X1 U524 ( .A(n223), .B(n212), .C(n349), .Y(n222) );
  AOI211X1 U525 ( .C(n441), .D(n213), .A(n225), .B(n347), .Y(n221) );
  OA22X1 U526 ( .A(arcon[5]), .B(n348), .C(n208), .D(n197), .Y(n349) );
  INVX1 U527 ( .A(norm_reg[13]), .Y(n461) );
  INVX1 U528 ( .A(n85), .Y(n86) );
  NAND21X1 U529 ( .B(n26), .A(md0[1]), .Y(n85) );
  AND3X1 U530 ( .A(n182), .B(n47), .C(n329), .Y(n410) );
  NAND21X1 U531 ( .B(setmdef), .A(n328), .Y(n329) );
  NAND2X1 U532 ( .A(sfroe), .B(n395), .Y(n182) );
  INVX1 U533 ( .A(arcon[7]), .Y(n328) );
  NAND21X1 U534 ( .B(n74), .A(md3[6]), .Y(n84) );
  INVX1 U535 ( .A(md1[6]), .Y(n139) );
  AO222X1 U536 ( .A(N612), .B(n274), .C(n273), .D(n276), .E(arcon[2]), .F(n394), .Y(n280) );
  AO222X1 U537 ( .A(N614), .B(n274), .C(n273), .D(n247), .E(arcon[4]), .F(n394), .Y(n249) );
  AO222X1 U538 ( .A(N613), .B(n274), .C(n273), .D(n251), .E(arcon[3]), .F(n394), .Y(n252) );
  OAI21BBX1 U539 ( .A(arcon[0]), .B(n394), .C(n24), .Y(n261) );
  MUX2IX1 U540 ( .D0(n273), .D1(n274), .S(N610), .Y(n24) );
  NOR2X1 U541 ( .A(n445), .B(oper_reg[2]), .Y(n402) );
  INVX1 U542 ( .A(oper_reg[3]), .Y(n445) );
  INVX1 U543 ( .A(n270), .Y(n268) );
  NOR2X1 U544 ( .A(n440), .B(oper_reg[1]), .Y(n389) );
  NOR2X1 U545 ( .A(n444), .B(oper_reg[3]), .Y(n403) );
  NOR2X1 U546 ( .A(oper_reg[3]), .B(oper_reg[2]), .Y(n399) );
  NOR2X1 U547 ( .A(oper_reg[1]), .B(oper_reg[0]), .Y(n405) );
  NOR2X1 U548 ( .A(n442), .B(oper_reg[0]), .Y(n400) );
  OAI31XL U549 ( .A(n224), .B(n219), .C(n216), .D(n262), .Y(n269) );
  INVX1 U550 ( .A(n342), .Y(n216) );
  INVX1 U551 ( .A(n306), .Y(n219) );
  OAI22X1 U552 ( .A(n336), .B(n337), .C(n396), .D(md3[6]), .Y(n224) );
  NAND3X1 U553 ( .A(n405), .B(oper_reg[3]), .C(oper_reg[2]), .Y(n208) );
  INVX1 U554 ( .A(oper_reg[1]), .Y(n442) );
  INVX1 U555 ( .A(oper_reg[2]), .Y(n444) );
  INVX1 U556 ( .A(n91), .Y(n135) );
  NAND21X1 U557 ( .B(n296), .A(md3[6]), .Y(n91) );
  INVX1 U558 ( .A(oper_reg[0]), .Y(n440) );
  NAND21X1 U559 ( .B(counter_st[1]), .A(n355), .Y(n369) );
  XNOR2XL U560 ( .A(n453), .B(n25), .Y(n247) );
  NOR2X1 U561 ( .A(counter_st[3]), .B(n370), .Y(n25) );
  OAI21BBX1 U562 ( .A(n369), .B(counter_st[2]), .C(n370), .Y(n276) );
  INVX1 U563 ( .A(N610), .Y(n355) );
  OAI21BBX1 U564 ( .A(counter_st[1]), .B(N610), .C(n369), .Y(n270) );
  NAND21X1 U565 ( .B(md3[5]), .A(n226), .Y(n308) );
  OAI31XL U566 ( .A(md3[7]), .B(n206), .C(n351), .D(n167), .Y(n347) );
  NAND5XL U567 ( .A(n286), .B(n285), .C(n284), .D(n283), .E(n282), .Y(n351) );
  INVX1 U568 ( .A(arcon[3]), .Y(n286) );
  INVX1 U569 ( .A(arcon[0]), .Y(n285) );
  INVX1 U570 ( .A(arcon[4]), .Y(n284) );
  NAND43X1 U571 ( .B(N610), .C(n453), .D(n346), .A(n236), .Y(n213) );
  NOR2X1 U572 ( .A(counter_st[3]), .B(counter_st[2]), .Y(n236) );
  NOR4XL U573 ( .A(n452), .B(N610), .C(counter_st[1]), .D(counter_st[3]), .Y(
        n228) );
  NAND2X1 U574 ( .A(counter_st[4]), .B(n228), .Y(n211) );
  INVX1 U575 ( .A(counter_st[4]), .Y(n453) );
  OAI31XL U576 ( .A(n220), .B(N610), .C(n346), .D(n281), .Y(n353) );
  NAND3X1 U577 ( .A(n454), .B(n453), .C(n452), .Y(n220) );
  INVX1 U578 ( .A(counter_st[3]), .Y(n454) );
  INVX1 U579 ( .A(counter_st[2]), .Y(n452) );
  OAI221X1 U580 ( .A(n167), .B(n353), .C(md3[7]), .D(n206), .E(n348), .Y(n287)
         );
  OAI22AX1 U581 ( .D(n209), .C(n210), .A(mdu_op[0]), .B(n208), .Y(n217) );
  INVX1 U582 ( .A(counter_st[1]), .Y(n346) );
  NAND3X1 U583 ( .A(n389), .B(oper_reg[3]), .C(oper_reg[2]), .Y(n223) );
  INVX1 U584 ( .A(arcon[1]), .Y(n283) );
  INVX1 U585 ( .A(arcon[2]), .Y(n282) );
  NAND31X1 U586 ( .C(n311), .A(n310), .B(n309), .Y(n312) );
  NAND31X1 U587 ( .C(md2[1]), .A(n303), .B(n301), .Y(n311) );
  NOR43XL U588 ( .B(n307), .C(n305), .D(n304), .A(md2[7]), .Y(n310) );
  NOR8XL U589 ( .A(md2[2]), .B(md2[4]), .C(md2[6]), .D(md3[0]), .E(md3[2]), 
        .F(md3[4]), .G(md3[7]), .H(n308), .Y(n309) );
  NAND3X1 U590 ( .A(n330), .B(n167), .C(arcon[6]), .Y(n324) );
  INVX1 U591 ( .A(md2[0]), .Y(n305) );
  INVX1 U592 ( .A(md0[1]), .Y(n97) );
  INVX1 U593 ( .A(md1[5]), .Y(n124) );
  INVX1 U594 ( .A(md1[4]), .Y(n120) );
  NAND42X1 U595 ( .C(n322), .D(n321), .A(n320), .B(n319), .Y(n323) );
  NOR32XL U596 ( .B(n316), .C(n315), .A(n314), .Y(n320) );
  NAND21X1 U597 ( .B(md4[3]), .A(n313), .Y(n322) );
  NOR8XL U598 ( .A(md5[6]), .B(md5[4]), .C(md4[2]), .D(md4[0]), .E(md4[6]), 
        .F(md4[4]), .G(md5[2]), .H(md5[0]), .Y(n319) );
  OR2X1 U599 ( .A(md5[3]), .B(md5[1]), .Y(n314) );
  OR2X1 U600 ( .A(md4[7]), .B(md4[5]), .Y(n321) );
  INVX1 U601 ( .A(md4[1]), .Y(n313) );
  INVX1 U602 ( .A(md0[0]), .Y(n95) );
  INVX1 U603 ( .A(set_div32), .Y(n397) );
  INVX1 U604 ( .A(md0[2]), .Y(n99) );
  INVX1 U605 ( .A(md0[3]), .Y(n101) );
  INVX1 U606 ( .A(md0[7]), .Y(n110) );
  INVX1 U607 ( .A(md0[6]), .Y(n108) );
  INVX1 U608 ( .A(md0[5]), .Y(n105) );
  INVX1 U609 ( .A(md0[4]), .Y(n103) );
  INVX1 U610 ( .A(md1[1]), .Y(n114) );
  INVX1 U611 ( .A(md1[3]), .Y(n118) );
  INVX1 U612 ( .A(md1[2]), .Y(n116) );
  INVX1 U613 ( .A(md1[0]), .Y(n112) );
  INVX1 U614 ( .A(md5[5]), .Y(n316) );
  INVX1 U615 ( .A(md5[7]), .Y(n315) );
  INVX1 U616 ( .A(arcon[5]), .Y(n293) );
  NOR43XL U617 ( .B(sfraddr[5]), .C(sfraddr[3]), .D(sfraddr[6]), .A(sfraddr[4]), .Y(n366) );
  XNOR2XL U618 ( .A(counter_st[4]), .B(r384_carry[4]), .Y(N614) );
  OR2X1 U619 ( .A(r384_carry[3]), .B(counter_st[3]), .Y(r384_carry[4]) );
  XNOR2XL U620 ( .A(r384_carry[3]), .B(counter_st[3]), .Y(N613) );
  OR2X1 U621 ( .A(counter_st[1]), .B(counter_st[2]), .Y(r384_carry[3]) );
  XNOR2XL U622 ( .A(counter_st[1]), .B(counter_st[2]), .Y(N612) );
  OR2X1 U623 ( .A(n369), .B(counter_st[2]), .Y(n370) );
endmodule


module mdu_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module mdu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module wakeupctrl_a0 ( irq, int0ff, int1ff, it0, it1, isreg, intprior0, 
        intprior1, eal, eint0, eint1, pmuintreq );
  input [3:0] isreg;
  input [1:0] intprior0;
  input [1:0] intprior1;
  input irq, int0ff, int1ff, it0, it1, eal, eint0, eint1;
  output pmuintreq;
  wire   n6, n7, n8, n9, n10, n11, n12, n1, n2, n3, n4, n5;

  OAI21BX1 U1 ( .C(eal), .B(n6), .A(n1), .Y(pmuintreq) );
  INVX1 U2 ( .A(irq), .Y(n1) );
  AOI33X1 U3 ( .A(eint0), .B(n7), .C(n8), .D(eint1), .E(n9), .F(n10), .Y(n6)
         );
  NOR3XL U4 ( .A(int1ff), .B(it1), .C(isreg[3]), .Y(n10) );
  NOR3XL U5 ( .A(int0ff), .B(it0), .C(isreg[3]), .Y(n8) );
  OAI21X1 U6 ( .B(n3), .C(n5), .A(n12), .Y(n7) );
  GEN2XL U7 ( .D(isreg[0]), .E(n3), .C(isreg[1]), .B(n5), .A(isreg[2]), .Y(n12) );
  INVX1 U8 ( .A(intprior1[0]), .Y(n5) );
  INVX1 U9 ( .A(intprior0[0]), .Y(n3) );
  OAI21X1 U10 ( .B(n2), .C(n4), .A(n11), .Y(n9) );
  GEN2XL U11 ( .D(isreg[0]), .E(n2), .C(isreg[1]), .B(n4), .A(isreg[2]), .Y(
        n11) );
  INVX1 U12 ( .A(intprior1[1]), .Y(n4) );
  INVX1 U13 ( .A(intprior0[1]), .Y(n2) );
endmodule


module pmurstctrl_a0 ( resetff, wdts, srst, pmuintreq, stop, idle, clkcpu_en, 
        clkper_en, cpu_resume, rsttowdt, rsttosrst, rst );
  input resetff, wdts, srst, pmuintreq, stop, idle;
  output clkcpu_en, clkper_en, cpu_resume, rsttowdt, rsttosrst, rst;
  wire   n2;

  OAI21X1 U1 ( .B(stop), .C(idle), .A(n2), .Y(clkcpu_en) );
  NAND2X1 U2 ( .A(stop), .B(n2), .Y(clkper_en) );
  INVX1 U3 ( .A(pmuintreq), .Y(n2) );
  OR2X1 U4 ( .A(srst), .B(resetff), .Y(rsttowdt) );
  OR2X1 U5 ( .A(wdts), .B(rsttowdt), .Y(rst) );
  OR2X1 U6 ( .A(resetff), .B(wdts), .Y(rsttosrst) );
  BUFX3 U7 ( .A(pmuintreq), .Y(cpu_resume) );
endmodule


module sfrmux_a0 ( isfrwait, sfraddr, c, ac, f0, rs, ov, f1, p, acc, b, dpl, 
        dph, dps, dpc, p2, sp, smod, pmw, p2sel, gf0, stop, idle, ckcon, port0, 
        port0ff, rmwinstr, arcon, md0, md1, md2, md3, md4, md5, t0_tmod, 
        t0_tf0, t0_tf1, t0_tr0, t0_tr1, tl0, th0, t1_tmod, t1_tf1, t1_tr1, tl1, 
        th1, wdtrel, ip0wdts, wdt_tm, t2con, s0con, s0buf, s0rell, s0relh, bd, 
        ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9, 
        iex10, iex11, iex12, ien0, ien1, ien2, ip0, ip1, isr_tm, i2c_int, 
        i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o, sfrdatai, tf1_gate, riti0_gate, 
        iex7_gate, iex2_gate, srstflag, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, ext_sfr_sel, sfrdatao );
  input [6:0] sfraddr;
  input [1:0] rs;
  input [7:0] acc;
  input [7:0] b;
  input [7:0] dpl;
  input [7:0] dph;
  input [3:0] dps;
  input [5:0] dpc;
  input [7:0] p2;
  input [7:0] sp;
  input [7:0] ckcon;
  input [7:0] port0;
  input [7:0] port0ff;
  input [7:0] arcon;
  input [7:0] md0;
  input [7:0] md1;
  input [7:0] md2;
  input [7:0] md3;
  input [7:0] md4;
  input [7:0] md5;
  input [3:0] t0_tmod;
  input [7:0] tl0;
  input [7:0] th0;
  input [3:0] t1_tmod;
  input [7:0] tl1;
  input [7:0] th1;
  input [7:0] wdtrel;
  input [7:0] t2con;
  input [7:0] s0con;
  input [7:0] s0buf;
  input [7:0] s0rell;
  input [7:0] s0relh;
  input [7:0] ien0;
  input [5:0] ien1;
  input [5:0] ien2;
  input [5:0] ip0;
  input [5:0] ip1;
  input [7:0] i2cdat_o;
  input [7:0] i2cadr_o;
  input [7:0] i2ccon_o;
  input [7:0] i2csta_o;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  input isfrwait, c, ac, f0, ov, f1, p, smod, pmw, p2sel, gf0, stop, idle,
         rmwinstr, t0_tf0, t0_tf1, t0_tr0, t0_tr1, t1_tf1, t1_tr1, ip0wdts,
         wdt_tm, bd, ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12, isr_tm, i2c_int, srstflag;
  output tf1_gate, riti0_gate, iex7_gate, iex2_gate, int_vect_8b, int_vect_93,
         int_vect_9b, int_vect_a3, ext_sfr_sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349;

  NAND32XL U2 ( .B(n31), .C(n79), .A(n14), .Y(n183) );
  OR3X1 U3 ( .A(n14), .B(n83), .C(n76), .Y(n139) );
  NAND32X4 U4 ( .B(sfraddr[2]), .C(n32), .A(n9), .Y(n79) );
  INVX3 U5 ( .A(sfraddr[2]), .Y(n34) );
  NAND31X2 U6 ( .C(sfraddr[0]), .A(sfraddr[1]), .B(n34), .Y(n77) );
  INVX3 U7 ( .A(n169), .Y(n342) );
  INVXL U8 ( .A(n168), .Y(n323) );
  INVX2 U9 ( .A(sfraddr[0]), .Y(n32) );
  INVX2 U10 ( .A(n160), .Y(n335) );
  NAND2X2 U11 ( .A(n6), .B(n7), .Y(sfrdatao[2]) );
  NAND43X2 U12 ( .B(n153), .C(n154), .D(n155), .A(n152), .Y(sfrdatao[0]) );
  NAND32X2 U13 ( .B(n37), .C(n35), .A(n36), .Y(n91) );
  NAND21X1 U14 ( .B(n11), .A(n104), .Y(n169) );
  INVX3 U15 ( .A(sfraddr[5]), .Y(n37) );
  NAND21X1 U16 ( .B(n18), .A(n85), .Y(n162) );
  INVX2 U17 ( .A(n48), .Y(n86) );
  NAND3XL U18 ( .A(sfraddr[4]), .B(sfraddr[3]), .C(n37), .Y(n76) );
  NAND21X1 U19 ( .B(n58), .A(n4), .Y(n95) );
  NAND32X1 U20 ( .B(n91), .C(n90), .A(n32), .Y(n164) );
  NAND3XL U21 ( .A(n82), .B(n89), .C(n32), .Y(n173) );
  INVX1 U22 ( .A(n38), .Y(n15) );
  NAND21X1 U23 ( .B(n37), .A(sfraddr[4]), .Y(n57) );
  INVX3 U24 ( .A(sfraddr[3]), .Y(n35) );
  NAND31X1 U25 ( .C(n147), .A(n146), .B(n145), .Y(n148) );
  NAND31XL U26 ( .C(n127), .A(n126), .B(n125), .Y(n147) );
  NOR43X1 U27 ( .B(n111), .C(n110), .D(n109), .A(n108), .Y(n151) );
  NOR43XL U28 ( .B(n122), .C(n121), .D(n120), .A(n119), .Y(n149) );
  AND3X1 U29 ( .A(n52), .B(n51), .C(n50), .Y(n53) );
  INVX2 U30 ( .A(n92), .Y(n309) );
  INVX2 U31 ( .A(n67), .Y(n312) );
  NAND21X1 U32 ( .B(n84), .A(n69), .Y(n160) );
  INVX1 U33 ( .A(n215), .Y(n7) );
  NAND32X1 U34 ( .B(n14), .C(n34), .A(n9), .Y(n90) );
  INVX2 U35 ( .A(n31), .Y(n82) );
  INVX1 U36 ( .A(n90), .Y(n89) );
  BUFX3 U37 ( .A(n33), .Y(n9) );
  INVX1 U38 ( .A(n175), .Y(n253) );
  INVX1 U39 ( .A(n113), .Y(n265) );
  INVX1 U40 ( .A(n348), .Y(n305) );
  INVX1 U41 ( .A(n163), .Y(n307) );
  INVX2 U42 ( .A(n118), .Y(n314) );
  INVX1 U43 ( .A(n185), .Y(n297) );
  INVX1 U44 ( .A(n159), .Y(n332) );
  INVX1 U45 ( .A(n162), .Y(n306) );
  INVX1 U46 ( .A(n165), .Y(n296) );
  INVX1 U47 ( .A(n166), .Y(n294) );
  INVX1 U48 ( .A(n112), .Y(n343) );
  INVX1 U49 ( .A(rmwinstr), .Y(n12) );
  NAND21X1 U50 ( .B(n71), .A(n4), .Y(n103) );
  INVX1 U51 ( .A(n138), .Y(n341) );
  NAND32X1 U52 ( .B(n35), .C(n60), .A(n36), .Y(n48) );
  INVX2 U53 ( .A(n62), .Y(n304) );
  NAND32X1 U54 ( .B(n71), .C(n31), .A(n39), .Y(n62) );
  NOR43XL U55 ( .B(n151), .C(n150), .D(n149), .A(n148), .Y(n152) );
  INVX1 U56 ( .A(n101), .Y(n344) );
  NOR5X1 U57 ( .A(n309), .B(n310), .C(n299), .D(n298), .E(n300), .Y(n97) );
  NOR5X1 U58 ( .A(n19), .B(n312), .C(n311), .D(n315), .E(n261), .Y(n74) );
  INVX1 U59 ( .A(n61), .Y(n347) );
  NAND21XL U60 ( .B(n77), .A(n78), .Y(n170) );
  NAND32XL U61 ( .B(n14), .C(n77), .A(n82), .Y(n171) );
  NAND21X2 U62 ( .B(sfraddr[6]), .A(n37), .Y(n60) );
  INVXL U63 ( .A(sfraddr[6]), .Y(n14) );
  INVX3 U64 ( .A(sfraddr[4]), .Y(n36) );
  NAND3X1 U65 ( .A(n47), .B(n46), .C(n45), .Y(n1) );
  NAND32X1 U66 ( .B(sfraddr[4]), .C(n60), .A(n35), .Y(n44) );
  INVX1 U67 ( .A(n183), .Y(n301) );
  INVXL U68 ( .A(sfraddr[6]), .Y(n38) );
  NAND21X2 U69 ( .B(n44), .A(n87), .Y(n68) );
  INVX1 U70 ( .A(n75), .Y(n345) );
  NOR21X2 U71 ( .B(n4), .A(n79), .Y(n19) );
  INVX2 U72 ( .A(n44), .Y(n4) );
  OR3X4 U73 ( .A(n71), .B(n39), .C(n13), .Y(n84) );
  BUFX1 U74 ( .A(sfraddr[3]), .Y(n13) );
  NAND21X1 U75 ( .B(n49), .A(sfraddr[0]), .Y(n58) );
  NAND32X2 U76 ( .B(n33), .C(n32), .A(n34), .Y(n83) );
  INVX3 U77 ( .A(sfraddr[1]), .Y(n33) );
  NAND43X2 U78 ( .B(n13), .C(n60), .D(n36), .A(n85), .Y(n113) );
  INVX3 U79 ( .A(n83), .Y(n85) );
  AND2XL U80 ( .A(md2[1]), .B(n306), .Y(n2) );
  AND2XL U81 ( .A(th0[1]), .B(n307), .Y(n3) );
  NOR3XL U82 ( .A(n2), .B(n3), .C(n167), .Y(n194) );
  NAND6X1 U83 ( .A(n213), .B(n212), .C(n214), .D(n211), .E(n210), .F(n209), 
        .Y(n215) );
  AOI222XL U84 ( .A(i2cdat_o[1]), .B(n324), .C(i2csta_o[1]), .D(n322), .E(
        i2ccon_o[1]), .F(n325), .Y(n176) );
  NAND6XL U85 ( .A(n131), .B(n160), .C(n165), .D(n157), .E(n182), .F(n113), 
        .Y(n61) );
  NAND21X1 U86 ( .B(n83), .A(n4), .Y(n67) );
  NAND21XL U87 ( .B(n71), .A(n4), .Y(n5) );
  NAND2X1 U88 ( .A(sfrdatai[2]), .B(n320), .Y(n6) );
  INVX2 U89 ( .A(n71), .Y(n81) );
  NAND32X1 U90 ( .B(n36), .C(n84), .A(n37), .Y(n138) );
  INVXL U91 ( .A(n156), .Y(n8) );
  NAND5X1 U92 ( .A(n347), .B(n349), .C(n102), .D(n345), .E(n344), .Y(n156) );
  INVX1 U93 ( .A(n17), .Y(n320) );
  NAND5X2 U94 ( .A(n81), .B(n20), .C(n39), .D(n36), .E(n35), .Y(n118) );
  NAND5X2 U95 ( .A(n13), .B(n15), .C(n81), .D(n37), .E(n36), .Y(n174) );
  INVXL U96 ( .A(n139), .Y(n326) );
  NAND31XL U97 ( .C(n32), .A(n82), .B(n89), .Y(n172) );
  NAND21X1 U98 ( .B(n175), .A(ip1[0]), .Y(n143) );
  NAND21X2 U99 ( .B(n79), .A(n78), .Y(n175) );
  INVX1 U100 ( .A(n173), .Y(n325) );
  BUFXL U101 ( .A(n315), .Y(n10) );
  BUFX8 U102 ( .A(n76), .Y(n31) );
  NAND43X1 U103 ( .B(n13), .C(n20), .D(n36), .A(n65), .Y(n112) );
  INVXL U104 ( .A(n11), .Y(n128) );
  INVX3 U105 ( .A(n93), .Y(n310) );
  NAND21X2 U106 ( .B(n48), .A(n85), .Y(n93) );
  NOR2X2 U107 ( .A(n103), .B(n12), .Y(n11) );
  NAND32X1 U108 ( .B(n32), .C(n91), .A(n89), .Y(n158) );
  INVXL U109 ( .A(n174), .Y(n331) );
  BUFXL U110 ( .A(n342), .Y(n16) );
  NAND21X1 U111 ( .B(n48), .A(n87), .Y(n94) );
  NAND5X1 U112 ( .A(n347), .B(n349), .C(n102), .D(n345), .E(n344), .Y(n17) );
  INVX3 U113 ( .A(n95), .Y(n298) );
  NAND5X1 U114 ( .A(n168), .B(n172), .C(n171), .D(n170), .E(n173), .Y(n100) );
  NOR21XL U115 ( .B(md1[0]), .A(n166), .Y(n127) );
  NAND32XL U116 ( .B(n91), .C(n79), .A(n39), .Y(n180) );
  OR2X1 U117 ( .A(n91), .B(n14), .Y(n18) );
  NAND21X2 U118 ( .B(n91), .A(n65), .Y(n73) );
  OR2X1 U119 ( .A(n91), .B(n14), .Y(n88) );
  NAND32X1 U120 ( .B(n37), .C(n84), .A(n36), .Y(n168) );
  NAND43X2 U121 ( .B(sfraddr[1]), .C(sfraddr[0]), .D(n34), .A(n86), .Y(n163)
         );
  NAND21X2 U122 ( .B(n88), .A(n80), .Y(n159) );
  NAND5X1 U123 ( .A(n140), .B(n159), .C(n174), .D(n139), .E(n175), .Y(n99) );
  INVX3 U124 ( .A(n72), .Y(n261) );
  NAND21X2 U125 ( .B(n71), .A(n78), .Y(n72) );
  OR2X2 U126 ( .A(n58), .B(n18), .Y(n157) );
  INVX1 U127 ( .A(n19), .Y(n66) );
  INVX2 U128 ( .A(n79), .Y(n80) );
  NAND32X1 U129 ( .B(n20), .C(n84), .A(n36), .Y(n140) );
  INVX3 U130 ( .A(n77), .Y(n87) );
  BUFXL U131 ( .A(sfraddr[5]), .Y(n20) );
  NAND21X2 U132 ( .B(n88), .A(n87), .Y(n166) );
  NAND21X1 U133 ( .B(n168), .A(acc[0]), .Y(n109) );
  INVX3 U134 ( .A(n70), .Y(n78) );
  AO222X1 U135 ( .A(port0[2]), .B(n11), .C(md0[2]), .D(n332), .E(b[2]), .F(
        n335), .Y(n197) );
  OAI21BBX1 U136 ( .A(sfrdatai[1]), .B(n320), .C(n23), .Y(sfrdatao[1]) );
  NAND21X1 U137 ( .B(n34), .A(sfraddr[1]), .Y(n49) );
  NAND21X2 U138 ( .B(n15), .A(n87), .Y(n43) );
  OR2X1 U139 ( .A(n18), .B(n59), .Y(n165) );
  AOI221X1 U140 ( .A(md2[2]), .B(n306), .C(th0[2]), .D(n307), .E(n198), .Y(
        n213) );
  AO222X1 U141 ( .A(md3[2]), .B(n293), .C(md5[2]), .D(n296), .E(md1[2]), .F(
        n294), .Y(n198) );
  INVX3 U142 ( .A(n96), .Y(n300) );
  NAND21X2 U143 ( .B(n71), .A(n86), .Y(n96) );
  INVX3 U144 ( .A(n73), .Y(n315) );
  INVX3 U145 ( .A(n43), .Y(n65) );
  INVX1 U146 ( .A(n170), .Y(n321) );
  INVX2 U147 ( .A(n94), .Y(n299) );
  NAND21XL U148 ( .B(n133), .A(n132), .Y(n134) );
  NOR5X1 U149 ( .A(n341), .B(n343), .C(n340), .D(n305), .E(n104), .Y(n102) );
  INVX3 U150 ( .A(n57), .Y(n69) );
  NAND43XL U151 ( .B(n55), .C(n54), .D(n1), .A(n53), .Y(n154) );
  NAND21XL U152 ( .B(n42), .A(n41), .Y(n155) );
  INVXL U153 ( .A(n134), .Y(n24) );
  AOI21BBXL U154 ( .B(n131), .C(n130), .A(n129), .Y(n132) );
  INVXL U155 ( .A(n182), .Y(n302) );
  INVX3 U156 ( .A(n68), .Y(n311) );
  INVXL U157 ( .A(n172), .Y(n322) );
  INVXL U158 ( .A(n140), .Y(n256) );
  INVXL U159 ( .A(n63), .Y(n349) );
  INVX1 U160 ( .A(n64), .Y(n340) );
  INVX1 U161 ( .A(n196), .Y(n23) );
  NOR43X1 U162 ( .B(n144), .C(n143), .D(n142), .A(n141), .Y(n145) );
  AND4X1 U163 ( .A(n177), .B(n176), .C(n21), .D(n22), .Y(n193) );
  AOI222XL U164 ( .A(iex2), .B(n256), .C(i2cadr_o[1]), .D(n326), .E(f1), .F(
        n341), .Y(n21) );
  AOI22X1 U165 ( .A(t2con[1]), .B(n331), .C(ip1[1]), .D(n253), .Y(n22) );
  AOI21BXL U166 ( .C(n165), .B(md5[0]), .A(n123), .Y(n126) );
  AOI21BXL U167 ( .C(n162), .B(md2[0]), .A(n124), .Y(n125) );
  NOR43X1 U168 ( .B(n117), .C(n116), .D(n115), .A(n114), .Y(n150) );
  AOI21BXL U169 ( .C(n348), .B(th1[0]), .A(n40), .Y(n41) );
  AOI21BXL U170 ( .C(n172), .B(i2csta_o[0]), .A(n105), .Y(n106) );
  INVX1 U171 ( .A(n158), .Y(n295) );
  INVX1 U172 ( .A(n157), .Y(n334) );
  INVX1 U173 ( .A(n180), .Y(n278) );
  INVXL U174 ( .A(n5), .Y(n104) );
  NAND21X1 U175 ( .B(n48), .A(n80), .Y(n92) );
  NAND21XL U176 ( .B(n59), .A(n4), .Y(n185) );
  NAND21XL U177 ( .B(n59), .A(n86), .Y(n182) );
  INVXL U178 ( .A(n178), .Y(n303) );
  INVX1 U179 ( .A(n171), .Y(n324) );
  INVX1 U180 ( .A(n164), .Y(n293) );
  INVX1 U181 ( .A(n179), .Y(n263) );
  NAND21XL U182 ( .B(n304), .A(n185), .Y(n63) );
  NAND43X1 U183 ( .B(n100), .C(n99), .D(n98), .A(n97), .Y(n101) );
  NAND21XL U184 ( .B(n31), .A(n65), .Y(n179) );
  OR2XL U185 ( .A(sfraddr[0]), .B(n49), .Y(n59) );
  NAND32XL U186 ( .B(n39), .C(n31), .A(n81), .Y(n64) );
  NAND6XL U187 ( .A(n349), .B(n348), .C(n347), .D(n346), .E(n345), .F(n344), 
        .Y(ext_sfr_sel) );
  INVXL U188 ( .A(n58), .Y(n56) );
  NAND43XL U189 ( .B(sfraddr[1]), .C(n48), .D(n34), .A(sfraddr[0]), .Y(n348)
         );
  NOR5XL U190 ( .A(n343), .B(n16), .C(n341), .D(n340), .E(n11), .Y(n346) );
  AND4X2 U191 ( .A(n137), .B(n136), .C(n135), .D(n24), .Y(n146) );
  AO21XL U192 ( .B(sfrdatai[3]), .C(n8), .A(n234), .Y(sfrdatao[3]) );
  NAND6XL U193 ( .A(n233), .B(n232), .C(n231), .D(n230), .E(n229), .F(n228), 
        .Y(n234) );
  AOI22XL U194 ( .A(dpl[1]), .B(n311), .C(s0rell[1]), .D(n315), .Y(n186) );
  AOI222XL U195 ( .A(t0_tmod[1]), .B(n309), .C(th1[1]), .D(n305), .E(tl1[1]), 
        .F(n310), .Y(n189) );
  AOI222XL U196 ( .A(sp[1]), .B(n19), .C(stop), .D(n298), .E(dph[1]), .F(n312), 
        .Y(n187) );
  AND4X1 U197 ( .A(n208), .B(n207), .C(n206), .D(n205), .Y(n209) );
  AOI22XL U198 ( .A(dpl[2]), .B(n311), .C(s0rell[2]), .D(n315), .Y(n205) );
  AOI222XL U199 ( .A(t0_tmod[2]), .B(n309), .C(th1[2]), .D(n305), .E(tl1[2]), 
        .F(n310), .Y(n208) );
  AOI222XL U200 ( .A(sp[2]), .B(n19), .C(gf0), .D(n298), .E(dph[2]), .F(n312), 
        .Y(n206) );
  AND4X1 U201 ( .A(n202), .B(n201), .C(n200), .D(n199), .Y(n212) );
  AOI22XL U202 ( .A(t2con[2]), .B(n331), .C(ip1[2]), .D(n253), .Y(n199) );
  AOI222XL U203 ( .A(i2cdat_o[2]), .B(n324), .C(i2csta_o[2]), .D(n322), .E(
        i2ccon_o[2]), .F(n325), .Y(n201) );
  AOI222XL U204 ( .A(iex3), .B(n256), .C(i2cadr_o[2]), .D(n326), .E(ov), .F(
        n341), .Y(n200) );
  AOI222XL U205 ( .A(wdtrel[1]), .B(n297), .C(tl0[1]), .D(n299), .E(ie0), .F(
        n300), .Y(n188) );
  AOI222XL U206 ( .A(acc[1]), .B(n323), .C(n342), .D(port0ff[1]), .E(s0relh[1]), .F(n321), .Y(n177) );
  AOI222XL U207 ( .A(acc[2]), .B(n323), .C(port0ff[2]), .D(n342), .E(s0relh[2]), .F(n321), .Y(n202) );
  AOI222XL U208 ( .A(wdtrel[2]), .B(n297), .C(tl0[2]), .D(n299), .E(it1), .F(
        n300), .Y(n207) );
  AOI221X1 U209 ( .A(ckcon[2]), .B(n302), .C(dps[2]), .D(n343), .E(n204), .Y(
        n210) );
  AOI221X1 U210 ( .A(ien0[1]), .B(n303), .C(ien2[1]), .D(n263), .E(n181), .Y(
        n192) );
  AOI221X1 U211 ( .A(arcon[1]), .B(n334), .C(md4[1]), .D(n295), .E(n161), .Y(
        n195) );
  AOI221X1 U212 ( .A(arcon[2]), .B(n334), .C(md4[2]), .D(n295), .E(n197), .Y(
        n214) );
  NOR21XL U213 ( .B(arcon[0]), .A(n157), .Y(n129) );
  NAND21XL U214 ( .B(n112), .A(dps[0]), .Y(n116) );
  NAND21XL U215 ( .B(n182), .A(ckcon[0]), .Y(n115) );
  NAND21XL U216 ( .B(n183), .A(s0buf[0]), .Y(n117) );
  NAND21XL U217 ( .B(n179), .A(ien2[0]), .Y(n121) );
  NAND21XL U218 ( .B(n180), .A(ip0[0]), .Y(n122) );
  NAND21X1 U219 ( .B(n107), .A(n106), .Y(n108) );
  NAND21XL U220 ( .B(n170), .A(s0relh[0]), .Y(n110) );
  NOR21XL U221 ( .B(tl1[0]), .A(n93), .Y(n40) );
  NOR21XL U222 ( .B(md3[0]), .A(n164), .Y(n123) );
  NOR21XL U223 ( .B(th0[0]), .A(n163), .Y(n124) );
  NOR21XL U224 ( .B(i2ccon_o[0]), .A(n173), .Y(n105) );
  NAND21XL U225 ( .B(n178), .A(ien0[0]), .Y(n120) );
  AO22XL U226 ( .A(i2cadr_o[0]), .B(n326), .C(iex7), .D(n256), .Y(n141) );
  NOR21XL U227 ( .B(md4[0]), .A(n158), .Y(n133) );
  INVX1 U228 ( .A(srstflag), .Y(n130) );
  NAND21XL U229 ( .B(n160), .A(b[0]), .Y(n135) );
  NAND21XL U230 ( .B(n159), .A(md0[0]), .Y(n137) );
  NAND21XL U231 ( .B(n138), .A(p), .Y(n144) );
  NAND21XL U232 ( .B(n66), .A(sp[0]), .Y(n46) );
  NAND21XL U233 ( .B(n95), .A(idle), .Y(n47) );
  NAND21XL U234 ( .B(n94), .A(tl0[0]), .Y(n52) );
  NAND21XL U235 ( .B(n185), .A(wdtrel[0]), .Y(n50) );
  NAND21XL U236 ( .B(n96), .A(it0), .Y(n51) );
  AOI221X1 U237 ( .A(ien0[2]), .B(n303), .C(ien2[2]), .D(n263), .E(n203), .Y(
        n211) );
  NOR21XL U238 ( .B(dpl[0]), .A(n68), .Y(n54) );
  NOR21XL U239 ( .B(i2cdat_o[0]), .A(n171), .Y(n107) );
  NOR21XL U240 ( .B(t0_tmod[0]), .A(n92), .Y(n42) );
  AOI221XL U241 ( .A(arcon[3]), .B(n334), .C(md4[3]), .D(n295), .E(n216), .Y(
        n233) );
  AO222XL U242 ( .A(port0[3]), .B(n11), .C(md0[3]), .D(n332), .E(b[3]), .F(
        n335), .Y(n216) );
  AND4X1 U243 ( .A(n227), .B(n226), .C(n225), .D(n224), .Y(n228) );
  AOI22XL U244 ( .A(dpl[3]), .B(n311), .C(s0rell[3]), .D(n10), .Y(n224) );
  AOI222XL U245 ( .A(t0_tmod[3]), .B(n309), .C(th1[3]), .D(n305), .E(tl1[3]), 
        .F(n310), .Y(n227) );
  AOI222XL U246 ( .A(sp[3]), .B(n19), .C(p2sel), .D(n298), .E(dph[3]), .F(n312), .Y(n225) );
  AND4X1 U247 ( .A(n221), .B(n220), .C(n219), .D(n218), .Y(n231) );
  AOI22XL U248 ( .A(t2con[3]), .B(n331), .C(ip1[3]), .D(n253), .Y(n218) );
  AOI222XL U249 ( .A(i2cdat_o[3]), .B(n324), .C(i2csta_o[3]), .D(n322), .E(
        i2ccon_o[3]), .F(n325), .Y(n220) );
  AOI222XL U250 ( .A(iex4), .B(n256), .C(i2cadr_o[3]), .D(n326), .E(rs[0]), 
        .F(n341), .Y(n219) );
  AOI222XL U251 ( .A(acc[3]), .B(n323), .C(port0ff[3]), .D(n16), .E(s0relh[3]), 
        .F(n321), .Y(n221) );
  AOI222XL U252 ( .A(wdtrel[3]), .B(n297), .C(tl0[3]), .D(n299), .E(ie1), .F(
        n300), .Y(n226) );
  AOI221XL U253 ( .A(ckcon[3]), .B(n302), .C(dps[3]), .D(n343), .E(n223), .Y(
        n229) );
  AO222XL U254 ( .A(s0buf[3]), .B(n301), .C(s0con[3]), .D(n304), .E(dpc[3]), 
        .F(n265), .Y(n223) );
  AOI221XL U255 ( .A(ien0[3]), .B(n303), .C(ien2[3]), .D(n263), .E(n222), .Y(
        n230) );
  AO222XL U256 ( .A(ip0[3]), .B(n278), .C(ien1[3]), .D(n261), .E(p2[3]), .F(
        n314), .Y(n222) );
  AOI221XL U257 ( .A(md2[3]), .B(n306), .C(th0[3]), .D(n307), .E(n217), .Y(
        n232) );
  AO222XL U258 ( .A(md3[3]), .B(n293), .C(md5[3]), .D(n296), .E(md1[3]), .F(
        n294), .Y(n217) );
  NAND6XL U259 ( .A(n275), .B(n274), .C(n273), .D(n272), .E(n271), .F(n270), 
        .Y(sfrdatao[5]) );
  AND4X1 U260 ( .A(n269), .B(n268), .C(n267), .D(n266), .Y(n270) );
  AOI221XL U261 ( .A(md1[5]), .B(n294), .C(md2[5]), .D(n306), .E(n255), .Y(
        n274) );
  AOI221XL U262 ( .A(b[5]), .B(n335), .C(arcon[5]), .D(n334), .E(n254), .Y(
        n275) );
  NAND6XL U263 ( .A(n252), .B(n251), .C(n250), .D(n249), .E(n248), .F(n247), 
        .Y(sfrdatao[4]) );
  AND4X1 U264 ( .A(n246), .B(n245), .C(n244), .D(n243), .Y(n247) );
  AOI221XL U265 ( .A(md1[4]), .B(n294), .C(md2[4]), .D(n306), .E(n236), .Y(
        n251) );
  AOI221XL U266 ( .A(b[4]), .B(n335), .C(arcon[4]), .D(n334), .E(n235), .Y(
        n252) );
  AND4X1 U267 ( .A(n260), .B(n259), .C(n258), .D(n257), .Y(n273) );
  AOI22XL U268 ( .A(iex6), .B(n256), .C(t2con[5]), .D(n331), .Y(n257) );
  AOI222XL U269 ( .A(i2ccon_o[5]), .B(n325), .C(acc[5]), .D(n323), .E(
        i2csta_o[5]), .F(n322), .Y(n259) );
  AOI222XL U270 ( .A(f0), .B(n341), .C(i2cdat_o[5]), .D(n324), .E(i2cadr_o[5]), 
        .F(n326), .Y(n258) );
  AND4X1 U271 ( .A(n240), .B(n239), .C(n238), .D(n237), .Y(n250) );
  AOI22XL U272 ( .A(iex5), .B(n256), .C(t2con[4]), .D(n331), .Y(n237) );
  AOI222XL U273 ( .A(i2ccon_o[4]), .B(n325), .C(acc[4]), .D(n323), .E(
        i2csta_o[4]), .F(n322), .Y(n239) );
  AOI222XL U274 ( .A(rs[1]), .B(n341), .C(i2cdat_o[4]), .D(n324), .E(
        i2cadr_o[4]), .F(n326), .Y(n238) );
  AOI222XL U275 ( .A(s0relh[5]), .B(n321), .C(port0ff[5]), .D(n16), .E(
        sfrdatai[5]), .F(n8), .Y(n260) );
  AOI222XL U276 ( .A(s0relh[4]), .B(n321), .C(port0ff[4]), .D(n16), .E(
        sfrdatai[4]), .F(n8), .Y(n240) );
  AO222XL U277 ( .A(md0[4]), .B(n332), .C(ip1[4]), .D(n253), .E(port0[4]), .F(
        n11), .Y(n235) );
  AO222XL U278 ( .A(md5[4]), .B(n296), .C(md4[4]), .D(n295), .E(md3[4]), .F(
        n293), .Y(n236) );
  AOI221XL U279 ( .A(dpc[4]), .B(n265), .C(ckcon[4]), .D(n302), .E(n242), .Y(
        n248) );
  AO222XL U280 ( .A(s0con[4]), .B(n304), .C(ien2[4]), .D(n263), .E(s0buf[4]), 
        .F(n301), .Y(n242) );
  AOI221XL U281 ( .A(p2[4]), .B(n314), .C(ien0[4]), .D(n303), .E(n241), .Y(
        n249) );
  AO222XL U282 ( .A(ien1[4]), .B(n261), .C(s0rell[4]), .D(n10), .E(ip0[4]), 
        .F(n278), .Y(n241) );
  NAND42X1 U283 ( .C(n339), .D(n338), .A(n337), .B(n336), .Y(sfrdatao[7]) );
  AO2222XL U284 ( .A(md5[7]), .B(n296), .C(md4[7]), .D(n295), .E(md1[7]), .F(
        n294), .G(md3[7]), .H(n293), .Y(n339) );
  AOI221XL U285 ( .A(b[7]), .B(n335), .C(arcon[7]), .D(n334), .E(n333), .Y(
        n336) );
  NAND42X1 U286 ( .C(n319), .D(n318), .A(n317), .B(n316), .Y(n338) );
  NAND42X1 U287 ( .C(n292), .D(n291), .A(n290), .B(n289), .Y(sfrdatao[6]) );
  AO2222XL U288 ( .A(md5[6]), .B(n296), .C(md4[6]), .D(n295), .E(md1[6]), .F(
        n294), .G(md3[6]), .H(n293), .Y(n292) );
  AOI221XL U289 ( .A(b[6]), .B(n335), .C(arcon[6]), .D(n334), .E(n288), .Y(
        n289) );
  NAND42X1 U290 ( .C(n282), .D(n281), .A(n280), .B(n279), .Y(n291) );
  AOI221XL U291 ( .A(tl1[6]), .B(n310), .C(t1_tmod[2]), .D(n309), .E(n276), 
        .Y(n280) );
  AO222XL U292 ( .A(th0[6]), .B(n307), .C(md2[6]), .D(n306), .E(th1[6]), .F(
        n305), .Y(n276) );
  AO222XL U293 ( .A(md0[5]), .B(n332), .C(ip1[5]), .D(n253), .E(port0[5]), .F(
        n11), .Y(n254) );
  AO222XL U294 ( .A(md5[5]), .B(n296), .C(md4[5]), .D(n295), .E(md3[5]), .F(
        n293), .Y(n255) );
  AND4X1 U295 ( .A(n287), .B(n286), .C(n285), .D(n284), .Y(n290) );
  AOI222XL U296 ( .A(i2cdat_o[6]), .B(n324), .C(i2csta_o[6]), .D(n322), .E(
        i2ccon_o[6]), .F(n325), .Y(n285) );
  AOI22XL U297 ( .A(s0relh[6]), .B(n321), .C(acc[6]), .D(n323), .Y(n286) );
  AOI22XL U298 ( .A(i2cadr_o[6]), .B(n326), .C(ac), .D(n341), .Y(n284) );
  AND4X1 U299 ( .A(n330), .B(n329), .C(n328), .D(n327), .Y(n337) );
  AOI222XL U300 ( .A(i2cadr_o[7]), .B(n326), .C(i2ccon_o[7]), .D(n325), .E(
        i2cdat_o[7]), .F(n324), .Y(n328) );
  AOI22XL U301 ( .A(acc[7]), .B(n323), .C(i2csta_o[7]), .D(n322), .Y(n329) );
  AOI22XL U302 ( .A(c), .B(n341), .C(bd), .D(n340), .Y(n327) );
  AOI221XL U303 ( .A(ip0wdts), .B(n278), .C(p2[6]), .D(n314), .E(n277), .Y(
        n279) );
  AO222XL U304 ( .A(dpl[6]), .B(n311), .C(sp[6]), .D(n19), .E(s0rell[6]), .F(
        n10), .Y(n277) );
  AOI222XL U305 ( .A(dph[5]), .B(n312), .C(wdtrel[5]), .D(n297), .E(isr_tm), 
        .F(n298), .Y(n267) );
  AOI222XL U306 ( .A(dph[4]), .B(n312), .C(wdtrel[4]), .D(n297), .E(pmw), .F(
        n298), .Y(n244) );
  AOI222XL U307 ( .A(tl1[4]), .B(n310), .C(th0[4]), .D(n307), .E(th1[4]), .F(
        n305), .Y(n246) );
  AOI222XL U308 ( .A(s0relh[7]), .B(n321), .C(port0ff[7]), .D(n16), .E(
        sfrdatai[7]), .F(n8), .Y(n330) );
  AOI222XL U309 ( .A(t0_tf0), .B(n300), .C(t1_tmod[1]), .D(n309), .E(tl0[5]), 
        .F(n299), .Y(n268) );
  AOI222XL U310 ( .A(t0_tr0), .B(n300), .C(t1_tmod[0]), .D(n309), .E(tl0[4]), 
        .F(n299), .Y(n245) );
  AOI221XL U311 ( .A(dpc[5]), .B(n265), .C(ckcon[5]), .D(n302), .E(n264), .Y(
        n271) );
  AO222XL U312 ( .A(s0con[5]), .B(n304), .C(ien2[5]), .D(n263), .E(s0buf[5]), 
        .F(n301), .Y(n264) );
  AOI221XL U313 ( .A(p2[5]), .B(n314), .C(ien0[5]), .D(n303), .E(n262), .Y(
        n272) );
  AO222XL U314 ( .A(ien1[5]), .B(n261), .C(s0rell[5]), .D(n10), .E(ip0[5]), 
        .F(n278), .Y(n262) );
  AOI221XL U315 ( .A(sfrdatai[6]), .B(n8), .C(port0ff[6]), .D(n16), .E(n283), 
        .Y(n287) );
  OA21XL U316 ( .B(t1_tr1), .C(t0_tr1), .A(n300), .Y(n283) );
  AOI22XL U317 ( .A(sp[4]), .B(n19), .C(dpl[4]), .D(n311), .Y(n243) );
  AO222XL U318 ( .A(md0[6]), .B(n332), .C(t2con[6]), .D(n331), .E(port0[6]), 
        .F(n11), .Y(n288) );
  AOI221XL U319 ( .A(s0rell[7]), .B(n10), .C(p2[7]), .D(n314), .E(n313), .Y(
        n316) );
  AO222XL U320 ( .A(sp[7]), .B(n19), .C(dph[7]), .D(n312), .E(dpl[7]), .F(n311), .Y(n313) );
  AOI221XL U321 ( .A(tl1[7]), .B(n310), .C(t1_tmod[3]), .D(n309), .E(n308), 
        .Y(n317) );
  AO222XL U322 ( .A(th0[7]), .B(n307), .C(md2[7]), .D(n306), .E(th1[7]), .F(
        n305), .Y(n308) );
  AO222XL U323 ( .A(md0[7]), .B(n332), .C(t2con[7]), .D(n331), .E(port0[7]), 
        .F(n11), .Y(n333) );
  AO2222XL U324 ( .A(s0con[6]), .B(n304), .C(ien0[6]), .D(n303), .E(ckcon[6]), 
        .F(n302), .G(s0buf[6]), .H(n301), .Y(n281) );
  AO2222XL U325 ( .A(s0con[7]), .B(n304), .C(ien0[7]), .D(n303), .E(ckcon[7]), 
        .F(n302), .G(s0buf[7]), .H(n301), .Y(n318) );
  AO2222XL U326 ( .A(n300), .B(tf1_gate), .C(tl0[7]), .D(n299), .E(smod), .F(
        n298), .G(wdtrel[7]), .H(n297), .Y(n319) );
  AO2222XL U327 ( .A(wdtrel[6]), .B(n297), .C(tl0[6]), .D(n299), .E(dph[6]), 
        .F(n312), .G(wdt_tm), .H(n298), .Y(n282) );
  AOI222XL U328 ( .A(tl1[5]), .B(n310), .C(th0[5]), .D(n307), .E(th1[5]), .F(
        n305), .Y(n269) );
  AOI22XL U329 ( .A(sp[5]), .B(n19), .C(dpl[5]), .D(n311), .Y(n266) );
  OR2X1 U330 ( .A(s0con[1]), .B(s0con[0]), .Y(riti0_gate) );
  OR2X1 U331 ( .A(t1_tf1), .B(t0_tf1), .Y(tf1_gate) );
  NAND21XL U332 ( .B(n174), .A(t2con[0]), .Y(n142) );
  BUFX3 U333 ( .A(iex2), .Y(iex2_gate) );
  BUFX3 U334 ( .A(iex7), .Y(iex7_gate) );
  BUFX3 U335 ( .A(iex8), .Y(int_vect_8b) );
  BUFX3 U336 ( .A(iex9), .Y(int_vect_93) );
  BUFX3 U337 ( .A(iex10), .Y(int_vect_9b) );
  BUFX3 U338 ( .A(iex11), .Y(int_vect_a3) );
  NAND32XL U339 ( .B(n71), .C(n91), .A(n14), .Y(n178) );
  NAND6X1 U340 ( .A(n74), .B(n179), .C(n178), .D(n180), .E(n118), .F(n183), 
        .Y(n75) );
  NAND21X1 U341 ( .B(n67), .A(dph[0]), .Y(n45) );
  NOR21XL U342 ( .B(s0rell[0]), .A(n73), .Y(n55) );
  AOI221X1 U343 ( .A(ckcon[1]), .B(n302), .C(dps[1]), .D(n343), .E(n184), .Y(
        n191) );
  NAND5XL U344 ( .A(n15), .B(n20), .C(sfraddr[4]), .D(n56), .E(n35), .Y(n131)
         );
  INVXL U345 ( .A(sfraddr[6]), .Y(n39) );
  AND4X1 U346 ( .A(n189), .B(n188), .C(n187), .D(n186), .Y(n190) );
  AO222X1 U347 ( .A(md3[1]), .B(n293), .C(md5[1]), .D(n296), .E(md1[1]), .F(
        n294), .Y(n167) );
  AO222X1 U348 ( .A(s0buf[1]), .B(n301), .C(s0con[1]), .D(n304), .E(dpc[1]), 
        .F(n265), .Y(n184) );
  AO222X1 U349 ( .A(s0buf[2]), .B(n301), .C(s0con[2]), .D(n304), .E(dpc[2]), 
        .F(n265), .Y(n204) );
  AO22X1 U350 ( .A(s0con[0]), .B(n304), .C(dpc[0]), .D(n265), .Y(n114) );
  NAND5X1 U351 ( .A(n162), .B(n166), .C(n163), .D(n158), .E(n164), .Y(n98) );
  NAND32X2 U352 ( .B(n15), .C(n35), .A(n69), .Y(n70) );
  NAND6X1 U353 ( .A(n193), .B(n194), .C(n195), .D(n192), .E(n191), .F(n190), 
        .Y(n196) );
  NAND21XL U354 ( .B(n128), .A(port0[0]), .Y(n136) );
  NAND21XL U355 ( .B(n169), .A(port0ff[0]), .Y(n111) );
  AO222X1 U356 ( .A(port0[1]), .B(n11), .C(md0[1]), .D(n332), .E(b[1]), .F(
        n335), .Y(n161) );
  NAND32X2 U357 ( .B(sfraddr[2]), .C(sfraddr[0]), .A(n33), .Y(n71) );
  AO222X1 U358 ( .A(ip0[1]), .B(n278), .C(ien1[1]), .D(n261), .E(p2[1]), .F(
        n314), .Y(n181) );
  AO222X1 U359 ( .A(ip0[2]), .B(n278), .C(ien1[2]), .D(n261), .E(p2[2]), .F(
        n314), .Y(n203) );
  AO22X1 U360 ( .A(ien1[0]), .B(n261), .C(p2[0]), .D(n314), .Y(n119) );
  NOR21X1 U361 ( .B(sfrdatai[0]), .A(n156), .Y(n153) );
endmodule


module syncneg_a0 ( clk, reset, rsttowdt, rsttosrst, rst, int0, int1, port0i, 
        rxd0i, sdai, int0ff, int1ff, port0ff, t0ff, t1ff, rxd0ff, sdaiff, 
        rsttowdtff, rsttosrstff, rstff, resetff );
  input [7:0] port0i;
  output [7:0] port0ff;
  input clk, reset, rsttowdt, rsttosrst, rst, int0, int1, rxd0i, sdai;
  output int0ff, int1ff, t0ff, t1ff, rxd0ff, sdaiff, rsttowdtff, rsttosrstff,
         rstff, resetff;
  wire   reset_ff1, int0_ff1, int1_ff1, rxd0_ff1, sdai_ff1;
  wire   [7:0] p0_ff1;

  DFFQX1 reset_ff2_reg ( .D(reset_ff1), .C(clk), .Q(resetff) );
  DFFQX1 rsttosrst_ff1_reg ( .D(rsttosrst), .C(clk), .Q(rsttosrstff) );
  DFFQX1 rsttowdt_ff1_reg ( .D(rsttowdt), .C(clk), .Q(rsttowdtff) );
  DFFQX1 int1_ff2_reg ( .D(int1_ff1), .C(clk), .Q(int1ff) );
  DFFQX1 int0_ff2_reg ( .D(int0_ff1), .C(clk), .Q(int0ff) );
  DFFQX1 p0_ff2_reg_6_ ( .D(p0_ff1[6]), .C(clk), .Q(port0ff[6]) );
  DFFQX1 p0_ff2_reg_7_ ( .D(p0_ff1[7]), .C(clk), .Q(port0ff[7]) );
  DFFQX1 p0_ff2_reg_5_ ( .D(p0_ff1[5]), .C(clk), .Q(port0ff[5]) );
  DFFQX1 p0_ff2_reg_4_ ( .D(p0_ff1[4]), .C(clk), .Q(port0ff[4]) );
  DFFQX1 rxd0_ff2_reg ( .D(rxd0_ff1), .C(clk), .Q(rxd0ff) );
  DFFQX1 sdai_ff2_reg ( .D(sdai_ff1), .C(clk), .Q(sdaiff) );
  DFFQX1 p0_ff2_reg_3_ ( .D(p0_ff1[3]), .C(clk), .Q(port0ff[3]) );
  DFFQX1 p0_ff2_reg_0_ ( .D(p0_ff1[0]), .C(clk), .Q(port0ff[0]) );
  DFFQX1 p0_ff2_reg_2_ ( .D(p0_ff1[2]), .C(clk), .Q(port0ff[2]) );
  DFFQX1 p0_ff2_reg_1_ ( .D(p0_ff1[1]), .C(clk), .Q(port0ff[1]) );
  DFFQX1 rst_ff1_reg ( .D(rst), .C(clk), .Q(rstff) );
  DFFQX1 int0_ff1_reg ( .D(int0), .C(clk), .Q(int0_ff1) );
  DFFQX1 int1_ff1_reg ( .D(int1), .C(clk), .Q(int1_ff1) );
  DFFQX1 p0_ff1_reg_6_ ( .D(port0i[6]), .C(clk), .Q(p0_ff1[6]) );
  DFFQX1 p0_ff1_reg_5_ ( .D(port0i[5]), .C(clk), .Q(p0_ff1[5]) );
  DFFQX1 p0_ff1_reg_4_ ( .D(port0i[4]), .C(clk), .Q(p0_ff1[4]) );
  DFFQX1 p0_ff1_reg_3_ ( .D(port0i[3]), .C(clk), .Q(p0_ff1[3]) );
  DFFQX1 p0_ff1_reg_2_ ( .D(port0i[2]), .C(clk), .Q(p0_ff1[2]) );
  DFFQX1 p0_ff1_reg_1_ ( .D(port0i[1]), .C(clk), .Q(p0_ff1[1]) );
  DFFQX1 p0_ff1_reg_0_ ( .D(port0i[0]), .C(clk), .Q(p0_ff1[0]) );
  DFFQX1 rxd0_ff1_reg ( .D(rxd0i), .C(clk), .Q(rxd0_ff1) );
  DFFQX1 p0_ff1_reg_7_ ( .D(port0i[7]), .C(clk), .Q(p0_ff1[7]) );
  DFFQX1 sdai_ff1_reg ( .D(sdai), .C(clk), .Q(sdai_ff1) );
  DFFQX1 reset_ff1_reg ( .D(reset), .C(clk), .Q(reset_ff1) );
  INVX1 U3 ( .A(1'b1), .Y(t1ff) );
  INVX1 U5 ( .A(1'b1), .Y(t0ff) );
endmodule


module mcu51_cpu_a0 ( clkcpu, rst, mempsack, memack, memdatai, memaddr, 
        mempsrd, mempswr, memrd, memwr, memaddr_comb, mempsrd_comb, 
        mempswr_comb, memrd_comb, memwr_comb, cpu_hold, cpu_resume, irq, 
        intvect, intcall, retiinstr, newinstr, rmwinstr, waitstaten, ramdatai, 
        sfrdatai, ramsfraddr, ramdatao, ramoe, ramwe, sfroe, sfrwe, sfroe_r, 
        sfrwe_r, sfroe_comb_s, sfrwe_comb_s, pc_o, pc_ini, cs_run, instr, 
        codefetch_s, sfrack, ramsfraddr_comb, ramdatao_comb, ramoe_comb, 
        ramwe_comb, ckcon, pmw, p2sel, gf0, stop, idle, acc, b, rs, c, ac, ov, 
        p, f0, f1, dph, dpl, dps, dpc, p2, sp );
  input [7:0] memdatai;
  output [15:0] memaddr;
  output [15:0] memaddr_comb;
  input [4:0] intvect;
  input [7:0] ramdatai;
  input [7:0] sfrdatai;
  output [7:0] ramsfraddr;
  output [7:0] ramdatao;
  output [15:0] pc_o;
  input [15:0] pc_ini;
  output [7:0] instr;
  output [7:0] ramsfraddr_comb;
  output [7:0] ramdatao_comb;
  output [7:0] ckcon;
  output [7:0] acc;
  output [7:0] b;
  output [1:0] rs;
  output [7:0] dph;
  output [7:0] dpl;
  output [3:0] dps;
  output [5:0] dpc;
  output [7:0] p2;
  output [7:0] sp;
  input clkcpu, rst, mempsack, memack, cpu_hold, cpu_resume, irq, sfrack;
  output mempsrd, mempswr, memrd, memwr, mempsrd_comb, mempswr_comb,
         memrd_comb, memwr_comb, intcall, retiinstr, newinstr, rmwinstr,
         waitstaten, ramoe, ramwe, sfroe, sfrwe, sfroe_r, sfrwe_r,
         sfroe_comb_s, sfrwe_comb_s, cs_run, codefetch_s, ramoe_comb,
         ramwe_comb, pmw, p2sel, gf0, stop, idle, c, ac, ov, p, f0, f1;
  wire   N343, N344, N345, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, finishmul, finishdiv, N370, N371, N372, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, d_hold, idle_r, cpu_resume_fff, stop_r, ramsfrwe,
         N512, N515, N520, pdmode, interrupt, N582, N583, N584, N585, N588,
         N589, N590, phase0_ff, newinstrlock, N670, N671, N672, N673, N674,
         N675, N676, N677, N679, N680, N681, N682, N683, N684, N685, N689,
         N690, accactv, N10562, N10563, N10564, N10565, N10566, N10567, N10568,
         N10569, N10570, N10571, N10572, N10573, N10574, N10575, N10576,
         N10577, N10578, N10581, N10582, N10583, N10584, N10585, N10586,
         N10587, N10588, N10589, N11478, N11479, N11480, N11481, N11482,
         N11483, N11484, N11485, N11486, N11487, N11488, N11489, N11491,
         N11498, N11499, N11500, N11501, N11502, N11503, N11504, N11505,
         N11787, N11788, N11789, N11790, N11791, N11792, N11793, N11804,
         N11805, N11806, N11807, N11808, N11809, N11810, N11821, N11822,
         N11823, N11824, N11825, N11826, N11827, dph_current_7_, N11845,
         N12469, N12470, N12472, N12477, N12478, N12479, N12480, N12481,
         N12482, N12483, N12484, N12485, N12486, N12487, N12488, N12489,
         N12490, N12491, N12492, N12493, N12494, N12495, N12496, N12497,
         N12498, N12499, N12500, N12501, N12502, N12503, N12504, N12505,
         N12506, N12507, N12508, N12509, N12510, N12511, N12512, N12513,
         N12514, N12515, N12516, N12517, N12518, N12519, N12520, N12521,
         N12522, N12523, N12524, N12525, N12526, N12527, N12528, N12529,
         N12530, N12531, N12532, N12533, N12534, N12535, N12536, N12537,
         N12538, N12539, N12540, N12541, N12542, N12543, N12544, N12545,
         N12546, N12547, N12548, N12549, N12550, N12551, N12552, N12553,
         N12554, N12555, N12556, N12557, N12558, N12559, N12560, N12561,
         N12562, N12563, N12564, N12566, N12567, N12568, N12569, N12570,
         N12571, N12572, N12573, N12575, N12576, N12577, N12578, N12579,
         N12580, N12581, N12582, N12584, N12585, N12586, N12587, N12588,
         N12589, N12590, N12591, N12593, N12594, N12595, N12596, N12597,
         N12598, N12599, N12600, N12602, N12603, N12604, N12605, N12606,
         N12607, N12608, N12609, N12611, N12612, N12613, N12614, N12615,
         N12616, N12617, N12618, N12620, N12621, N12622, N12623, N12624,
         N12625, N12626, N12627, N12629, N12630, N12631, N12632, N12633,
         N12634, N12635, N12636, N12637, N12644, N12651, N12658, N12665,
         N12672, N12679, N12686, N12690, N12691, N12692, N12693, N12694,
         N12695, N12697, N12698, N12699, N12700, N12701, N12702, N12703,
         N12704, N12705, N12706, N12709, N12710, N12711, N12713, N12714,
         N12715, N12716, N12717, N12718, N12719, N12720, N12721, N12722,
         N12723, N12724, N12725, N12726, N12727, N12728, N12729, N12730,
         N12770, N12776, N12801, N12802, N12803, N12804, N12805, N12806,
         N12807, N12808, N12824, N12825, N12826, N12827, N12828, N12829,
         N12830, N12831, N12841, N12842, N12843, N12844, N12845, N12846,
         N12847, N12848, N12849, N12850, N12851, N12852, N12853, N12854,
         N12855, N12856, N12905, israccess, N12912, N12965, N12966, N12967,
         N12968, N12969, N12970, N12971, N12972, N12974, N12975, N12976,
         N12977, N13014, N13023, N13032, N13041, N13050, N13059, N13068,
         N13077, N13086, N13095, N13104, N13113, N13122, N13131, N13140,
         N13149, N13158, N13167, N13176, N13185, N13194, N13203, N13212,
         N13221, N13230, N13239, N13248, N13257, N13266, N13275, N13284,
         N13293, rn_1_, multemp1_0_, N13324, N13325, N13326, N13327, N13328,
         N13329, N13330, N13331, N13332, N13336, N13337, N13338, N13339,
         N13340, N13341, N13342, N13343, divtemp1_0_, N13345, N13346, N13347,
         N13348, N13349, N13350, N13351, N13352, N13353, N13366, N13367,
         N13368, N13369, N13370, N13371, N13372, N13373, cpu_resume_ff1,
         N13379, N13380, net12372, net12378, net12383, net12388, net12393,
         net12398, net12403, net12408, net12413, net12418, net12423, net12428,
         net12433, net12438, net12443, net12448, net12453, net12458, net12463,
         net12468, net12473, net12478, net12483, net12488, net12493, net12498,
         net12503, net12508, net12513, net12518, net12523, net12528, net12533,
         net12538, net12543, net12548, net12553, net12558, net12563, net12568,
         net12573, net12578, net12583, net12588, net12593, net12598, net12603,
         net12608, net12613, net12618, net12623, net12628, net12633, net12638,
         net12643, n726, n1023, n1024, n1025, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, multemp1_8_, multemp1_7_, multemp1_6_,
         multemp1_5_, multemp1_4_, multemp1_3_, multemp1_2_, multemp1_1_,
         N14351, N14350, N14349, N14348, N14347, N14346, N14345, N14344,
         N14343, N14342, N14341, N14340, N14339, N14338, N14337, N14336,
         add_5280_3_carry_9_, add_5280_3_carry_10_, add_5280_3_carry_11_,
         add_5280_3_carry_12_, add_5280_3_carry_13_, add_5280_3_carry_14_,
         add_5280_3_carry_15_, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n34, n36, n38, n40, n42, n43, n44, n46, n47, n48,
         n50, n52, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n107,
         n108, n109, n111, n112, n113, n114, n116, n117, n118, n119, n122,
         n123, n124, n127, n128, n129, n130, n131, n132, n133, n135, n137,
         n138, n141, n142, n143, n144, n145, n147, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n543, n545, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         SYNOPSYS_UNCONNECTED_1;
  wire   [2:0] state;
  wire   [5:0] phase;
  wire   [15:0] alu_out;
  wire   [15:0] pc_i;
  wire   [7:0] temp;
  wire   [18:0] dec_accop;
  wire   [7:0] dec_cop;
  wire   [9:1] multemp2;
  wire   [7:0] temp2_comb;
  wire   [15:0] dptr_inc;
  wire   [63:0] dpl_reg;
  wire   [63:0] dph_reg;
  wire   [47:0] dpc_tab;
  wire   [2:0] waitcnt;
  wire   [255:0] rn_reg;
  wire   [7:0] multempreg;
  wire   [6:0] divtempreg;
  wire   [15:9] add_5280_4_carry;
  wire   [15:10] add_5280_2_carry;

  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 clk_gate_finishmul_reg ( .CLK(clkcpu), 
        .EN(N370), .ENCLK(net12372), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 clk_gate_instr_reg ( .CLK(clkcpu), .EN(
        N685), .ENCLK(net12378), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 clk_gate_bitno_reg ( .CLK(clkcpu), .EN(
        N11491), .ENCLK(net12383), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 clk_gate_dph_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N12556), .ENCLK(net12388), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 clk_gate_dph_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N12547), .ENCLK(net12393), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 clk_gate_dph_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N12538), .ENCLK(net12398), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 clk_gate_dph_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N12529), .ENCLK(net12403), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 clk_gate_dph_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N12520), .ENCLK(net12408), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 clk_gate_dph_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N12511), .ENCLK(net12413), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 clk_gate_dph_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N12502), .ENCLK(net12418), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 clk_gate_dph_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N12493), .ENCLK(net12423), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 clk_gate_dpc_tab_reg_7_ ( .CLK(clkcpu), 
        .EN(N12686), .ENCLK(net12428), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 clk_gate_dpc_tab_reg_6_ ( .CLK(clkcpu), 
        .EN(N12679), .ENCLK(net12433), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 clk_gate_dpc_tab_reg_5_ ( .CLK(clkcpu), 
        .EN(N12672), .ENCLK(net12438), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 clk_gate_dpc_tab_reg_4_ ( .CLK(clkcpu), 
        .EN(N12665), .ENCLK(net12443), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 clk_gate_dpc_tab_reg_3_ ( .CLK(clkcpu), 
        .EN(N12658), .ENCLK(net12448), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 clk_gate_dpc_tab_reg_2_ ( .CLK(clkcpu), 
        .EN(N12651), .ENCLK(net12453), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 clk_gate_dpc_tab_reg_1_ ( .CLK(clkcpu), 
        .EN(N12644), .ENCLK(net12458), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 clk_gate_dpc_tab_reg_0_ ( .CLK(clkcpu), 
        .EN(N12637), .ENCLK(net12463), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 clk_gate_temp_reg ( .CLK(clkcpu), .EN(
        N12722), .ENCLK(net12468), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 clk_gate_waitcnt_reg ( .CLK(clkcpu), 
        .EN(N12977), .ENCLK(net12473), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 clk_gate_rn_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N13293), .ENCLK(net12478), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 clk_gate_rn_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N13284), .ENCLK(net12483), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 clk_gate_rn_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N13275), .ENCLK(net12488), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 clk_gate_rn_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N13266), .ENCLK(net12493), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 clk_gate_rn_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N13257), .ENCLK(net12498), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 clk_gate_rn_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N13248), .ENCLK(net12503), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 clk_gate_rn_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N13239), .ENCLK(net12508), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 clk_gate_rn_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N13230), .ENCLK(net12513), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 clk_gate_rn_reg_reg_8_ ( .CLK(clkcpu), 
        .EN(N13221), .ENCLK(net12518), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 clk_gate_rn_reg_reg_9_ ( .CLK(clkcpu), 
        .EN(N13212), .ENCLK(net12523), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 clk_gate_rn_reg_reg_10_ ( .CLK(clkcpu), 
        .EN(N13203), .ENCLK(net12528), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 clk_gate_rn_reg_reg_11_ ( .CLK(clkcpu), 
        .EN(N13194), .ENCLK(net12533), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 clk_gate_rn_reg_reg_12_ ( .CLK(clkcpu), 
        .EN(N13185), .ENCLK(net12538), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 clk_gate_rn_reg_reg_13_ ( .CLK(clkcpu), 
        .EN(N13176), .ENCLK(net12543), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 clk_gate_rn_reg_reg_14_ ( .CLK(clkcpu), 
        .EN(N13167), .ENCLK(net12548), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 clk_gate_rn_reg_reg_15_ ( .CLK(clkcpu), 
        .EN(N13158), .ENCLK(net12553), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 clk_gate_rn_reg_reg_16_ ( .CLK(clkcpu), 
        .EN(N13149), .ENCLK(net12558), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 clk_gate_rn_reg_reg_17_ ( .CLK(clkcpu), 
        .EN(N13140), .ENCLK(net12563), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 clk_gate_rn_reg_reg_18_ ( .CLK(clkcpu), 
        .EN(N13131), .ENCLK(net12568), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 clk_gate_rn_reg_reg_19_ ( .CLK(clkcpu), 
        .EN(N13122), .ENCLK(net12573), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 clk_gate_rn_reg_reg_20_ ( .CLK(clkcpu), 
        .EN(N13113), .ENCLK(net12578), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 clk_gate_rn_reg_reg_21_ ( .CLK(clkcpu), 
        .EN(N13104), .ENCLK(net12583), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 clk_gate_rn_reg_reg_22_ ( .CLK(clkcpu), 
        .EN(N13095), .ENCLK(net12588), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 clk_gate_rn_reg_reg_23_ ( .CLK(clkcpu), 
        .EN(N13086), .ENCLK(net12593), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 clk_gate_rn_reg_reg_24_ ( .CLK(clkcpu), 
        .EN(N13077), .ENCLK(net12598), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 clk_gate_rn_reg_reg_25_ ( .CLK(clkcpu), 
        .EN(N13068), .ENCLK(net12603), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 clk_gate_rn_reg_reg_26_ ( .CLK(clkcpu), 
        .EN(N13059), .ENCLK(net12608), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 clk_gate_rn_reg_reg_27_ ( .CLK(clkcpu), 
        .EN(N13050), .ENCLK(net12613), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 clk_gate_rn_reg_reg_28_ ( .CLK(clkcpu), 
        .EN(N13041), .ENCLK(net12618), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 clk_gate_rn_reg_reg_29_ ( .CLK(clkcpu), 
        .EN(N13032), .ENCLK(net12623), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 clk_gate_rn_reg_reg_30_ ( .CLK(clkcpu), 
        .EN(N13023), .ENCLK(net12628), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 clk_gate_rn_reg_reg_31_ ( .CLK(clkcpu), 
        .EN(N13014), .ENCLK(net12633), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 clk_gate_multempreg_reg ( .CLK(clkcpu), 
        .EN(N13324), .ENCLK(net12638), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 clk_gate_divtempreg_reg ( .CLK(clkcpu), 
        .EN(N13366), .ENCLK(net12643), .TE(1'b0) );
  mcu51_cpu_a0_DW01_inc_0 add_5525 ( .A({N12776, n289, n290, n286, n285, n284, 
        N12770, n283}), .SUM({N12808, N12807, N12806, N12805, N12804, N12803, 
        N12802, N12801}) );
  mcu51_cpu_a0_DW01_inc_1 add_5286 ( .A({dph_current_7_, n24, n23, n22, n21, 
        n20, n18, n19, n17, n15, n14, n12, n13, n10, n8, n11}), .SUM(dptr_inc)
         );
  mcu51_cpu_a0_DW01_inc_2 r715 ( .A(pc_o), .SUM(pc_i) );
  mcu51_cpu_a0_DW01_add_8 add_5901_aco ( .A({1'b0, multempreg}), .B({1'b0, 
        N14343, N14342, N14341, N14340, N14339, N14338, N14337, N14336}), .CI(
        1'b0), .SUM({multemp1_8_, multemp1_7_, multemp1_6_, multemp1_5_, 
        multemp1_4_, multemp1_3_, multemp1_2_, multemp1_1_, multemp1_0_}), 
        .CO() );
  mcu51_cpu_a0_DW01_add_7 add_5907_aco ( .A({1'b0, multemp1_8_, multemp1_7_, 
        multemp1_6_, multemp1_5_, multemp1_4_, multemp1_3_, multemp1_2_, 
        multemp1_1_}), .B({1'b0, N14351, N14350, N14349, N14348, N14347, 
        N14346, N14345, N14344}), .CI(1'b0), .SUM(multemp2), .CO() );
  mcu51_cpu_a0_DW01_sub_2 sub_5969 ( .A({1'b0, n276, n275, n272, n273, n269, 
        n270, divtemp1_0_, acc[6]}), .B({1'b0, b}), .CI(1'b0), .DIFF({N13353, 
        N13352, N13351, N13350, N13349, N13348, N13347, N13346, N13345}), 
        .CO() );
  mcu51_cpu_a0_DW01_add_10 add_5586 ( .A({n2439, n2439, n2439, n2439, n2439, 
        n2439, n2439, n2439, N12831, N12830, N12829, N12828, N12827, N12826, 
        N12825, N12824}), .B({N12856, N12855, N12854, N12853, N12852, N12851, 
        N12850, N12849, N12848, N12847, N12846, N12845, N12844, N12843, N12842, 
        N12841}), .CI(1'b0), .SUM(alu_out), .CO() );
  mcu51_cpu_a0_DW01_sub_3 sub_5950 ( .A({1'b0, divtempreg, acc[7]}), .B({1'b0, 
        b}), .CI(1'b0), .DIFF({N13343, SYNOPSYS_UNCONNECTED_1, N13342, N13341, 
        N13340, N13339, N13338, N13337, N13336}), .CO() );
  DFFQX1 dec_accop_reg_9_ ( .D(N10572), .C(net12372), .Q(dec_accop[9]) );
  DFFQX1 dec_accop_reg_7_ ( .D(N10570), .C(net12372), .Q(dec_accop[7]) );
  DFFQX1 dec_accop_reg_18_ ( .D(N10581), .C(net12372), .Q(dec_accop[18]) );
  DFFQX1 dec_accop_reg_10_ ( .D(N10573), .C(net12372), .Q(dec_accop[10]) );
  DFFQX1 cpu_resume_ff1_reg ( .D(N13379), .C(clkcpu), .Q(cpu_resume_ff1) );
  DFFQX1 newinstrlock_reg ( .D(n1878), .C(net12372), .Q(newinstrlock) );
  DFFQX1 phase0_ff_reg ( .D(N689), .C(net12372), .Q(phase0_ff) );
  DFFQX1 finishmul_reg ( .D(N371), .C(net12372), .Q(finishmul) );
  DFFQX1 finishdiv_reg ( .D(N372), .C(net12372), .Q(finishdiv) );
  DFFQX1 multempreg_reg_7_ ( .D(N13332), .C(net12638), .Q(multempreg[7]) );
  DFFQX1 multempreg_reg_6_ ( .D(N13331), .C(net12638), .Q(multempreg[6]) );
  DFFQX1 multempreg_reg_5_ ( .D(N13330), .C(net12638), .Q(multempreg[5]) );
  DFFQX1 multempreg_reg_4_ ( .D(N13329), .C(net12638), .Q(multempreg[4]) );
  DFFQX1 multempreg_reg_3_ ( .D(N13328), .C(net12638), .Q(multempreg[3]) );
  DFFQX1 pdmode_reg ( .D(n2446), .C(net12372), .Q(pdmode) );
  DFFQX1 d_hold_reg ( .D(cpu_hold), .C(clkcpu), .Q(d_hold) );
  DFFQX1 cpu_resume_fff_reg ( .D(N13380), .C(clkcpu), .Q(cpu_resume_fff) );
  DFFQX1 multempreg_reg_2_ ( .D(N13327), .C(net12638), .Q(multempreg[2]) );
  DFFQX1 p2_reg_reg_7_ ( .D(N12492), .C(net12372), .Q(p2[7]) );
  DFFQX1 p2_reg_reg_6_ ( .D(N12491), .C(net12372), .Q(p2[6]) );
  DFFQX1 p2_reg_reg_5_ ( .D(N12490), .C(net12372), .Q(p2[5]) );
  DFFQX1 f0_reg ( .D(n1882), .C(net12372), .Q(f0) );
  DFFQX1 p2_reg_reg_4_ ( .D(N12489), .C(net12372), .Q(p2[4]) );
  DFFQX1 dpc_tab_reg_3__5_ ( .D(n2430), .C(net12448), .Q(dpc_tab[23]) );
  DFFQX1 dpc_tab_reg_3__4_ ( .D(N12691), .C(net12448), .Q(dpc_tab[22]) );
  DFFQX1 dpc_tab_reg_7__5_ ( .D(N12692), .C(net12428), .Q(dpc_tab[47]) );
  DFFQX1 dpc_tab_reg_7__4_ ( .D(N12691), .C(net12428), .Q(dpc_tab[46]) );
  DFFQX1 dpc_tab_reg_0__5_ ( .D(n521), .C(net12463), .Q(dpc_tab[5]) );
  DFFQX1 dpc_tab_reg_0__4_ ( .D(n2436), .C(net12463), .Q(dpc_tab[4]) );
  DFFQX1 dpc_tab_reg_4__5_ ( .D(N12692), .C(net12443), .Q(dpc_tab[29]) );
  DFFQX1 dpc_tab_reg_4__4_ ( .D(n2436), .C(net12443), .Q(dpc_tab[28]) );
  DFFQX1 dpc_tab_reg_1__5_ ( .D(n2430), .C(net12458), .Q(dpc_tab[11]) );
  DFFQX1 dpc_tab_reg_1__4_ ( .D(n2436), .C(net12458), .Q(dpc_tab[10]) );
  DFFQX1 dpc_tab_reg_5__5_ ( .D(N12692), .C(net12438), .Q(dpc_tab[35]) );
  DFFQX1 dpc_tab_reg_5__4_ ( .D(n2436), .C(net12438), .Q(dpc_tab[34]) );
  DFFQX1 dpc_tab_reg_2__5_ ( .D(n2430), .C(net12453), .Q(dpc_tab[17]) );
  DFFQX1 dpc_tab_reg_2__4_ ( .D(N12691), .C(net12453), .Q(dpc_tab[16]) );
  DFFQX1 dpc_tab_reg_6__5_ ( .D(N12692), .C(net12433), .Q(dpc_tab[41]) );
  DFFQX1 dpc_tab_reg_6__4_ ( .D(N12691), .C(net12433), .Q(dpc_tab[40]) );
  DFFQX1 dph_reg_reg_3__7_ ( .D(N12528), .C(net12408), .Q(dph_reg[31]) );
  DFFQX1 dph_reg_reg_3__6_ ( .D(N12527), .C(net12408), .Q(dph_reg[30]) );
  DFFQX1 dph_reg_reg_7__7_ ( .D(N12564), .C(net12388), .Q(dph_reg[63]) );
  DFFQX1 dph_reg_reg_7__6_ ( .D(N12563), .C(net12388), .Q(dph_reg[62]) );
  DFFQX1 dph_reg_reg_0__7_ ( .D(N12501), .C(net12423), .Q(dph_reg[7]) );
  DFFQX1 dph_reg_reg_0__6_ ( .D(N12500), .C(net12423), .Q(dph_reg[6]) );
  DFFQX1 dph_reg_reg_4__7_ ( .D(N12537), .C(net12403), .Q(dph_reg[39]) );
  DFFQX1 dph_reg_reg_4__6_ ( .D(N12536), .C(net12403), .Q(dph_reg[38]) );
  DFFQX1 dph_reg_reg_1__7_ ( .D(N12510), .C(net12418), .Q(dph_reg[15]) );
  DFFQX1 dph_reg_reg_1__6_ ( .D(N12509), .C(net12418), .Q(dph_reg[14]) );
  DFFQX1 dph_reg_reg_5__7_ ( .D(N12546), .C(net12398), .Q(dph_reg[47]) );
  DFFQX1 dph_reg_reg_5__6_ ( .D(N12545), .C(net12398), .Q(dph_reg[46]) );
  DFFQX1 dph_reg_reg_2__7_ ( .D(N12519), .C(net12413), .Q(dph_reg[23]) );
  DFFQX1 dph_reg_reg_2__6_ ( .D(N12518), .C(net12413), .Q(dph_reg[22]) );
  DFFQX1 dph_reg_reg_6__7_ ( .D(N12555), .C(net12393), .Q(dph_reg[55]) );
  DFFQX1 dph_reg_reg_6__6_ ( .D(N12554), .C(net12393), .Q(dph_reg[54]) );
  DFFQX1 dph_reg_reg_3__5_ ( .D(N12526), .C(net12408), .Q(dph_reg[29]) );
  DFFQX1 dph_reg_reg_3__4_ ( .D(N12525), .C(net12408), .Q(dph_reg[28]) );
  DFFQX1 dph_reg_reg_7__5_ ( .D(N12562), .C(net12388), .Q(dph_reg[61]) );
  DFFQX1 dph_reg_reg_7__4_ ( .D(N12561), .C(net12388), .Q(dph_reg[60]) );
  DFFQX1 dph_reg_reg_0__5_ ( .D(N12499), .C(net12423), .Q(dph_reg[5]) );
  DFFQX1 dph_reg_reg_0__4_ ( .D(N12498), .C(net12423), .Q(dph_reg[4]) );
  DFFQX1 dph_reg_reg_4__5_ ( .D(N12535), .C(net12403), .Q(dph_reg[37]) );
  DFFQX1 dph_reg_reg_4__4_ ( .D(N12534), .C(net12403), .Q(dph_reg[36]) );
  DFFQX1 dph_reg_reg_1__5_ ( .D(N12508), .C(net12418), .Q(dph_reg[13]) );
  DFFQX1 dph_reg_reg_1__4_ ( .D(N12507), .C(net12418), .Q(dph_reg[12]) );
  DFFQX1 dph_reg_reg_5__5_ ( .D(N12544), .C(net12398), .Q(dph_reg[45]) );
  DFFQX1 dph_reg_reg_5__4_ ( .D(N12543), .C(net12398), .Q(dph_reg[44]) );
  DFFQX1 dph_reg_reg_2__5_ ( .D(N12517), .C(net12413), .Q(dph_reg[21]) );
  DFFQX1 dph_reg_reg_2__4_ ( .D(N12516), .C(net12413), .Q(dph_reg[20]) );
  DFFQX1 dph_reg_reg_6__5_ ( .D(N12553), .C(net12393), .Q(dph_reg[53]) );
  DFFQX1 dph_reg_reg_6__4_ ( .D(N12552), .C(net12393), .Q(dph_reg[52]) );
  DFFQX1 p2sel_s_reg ( .D(N520), .C(net12372), .Q(p2sel) );
  DFFQX1 p2_reg_reg_3_ ( .D(N12488), .C(net12372), .Q(p2[3]) );
  DFFQX1 dph_reg_reg_3__3_ ( .D(N12524), .C(net12408), .Q(dph_reg[27]) );
  DFFQX1 dph_reg_reg_7__3_ ( .D(N12560), .C(net12388), .Q(dph_reg[59]) );
  DFFQX1 dph_reg_reg_0__3_ ( .D(N12497), .C(net12423), .Q(dph_reg[3]) );
  DFFQX1 dph_reg_reg_4__3_ ( .D(N12533), .C(net12403), .Q(dph_reg[35]) );
  DFFQX1 dph_reg_reg_1__3_ ( .D(N12506), .C(net12418), .Q(dph_reg[11]) );
  DFFQX1 dph_reg_reg_5__3_ ( .D(N12542), .C(net12398), .Q(dph_reg[43]) );
  DFFQX1 dph_reg_reg_2__3_ ( .D(N12515), .C(net12413), .Q(dph_reg[19]) );
  DFFQX1 dph_reg_reg_6__3_ ( .D(N12551), .C(net12393), .Q(dph_reg[51]) );
  DFFQX1 dpc_tab_reg_3__3_ ( .D(N12690), .C(net12448), .Q(dpc_tab[21]) );
  DFFQX1 dpc_tab_reg_7__3_ ( .D(N12690), .C(net12428), .Q(dpc_tab[45]) );
  DFFQX1 dpc_tab_reg_0__3_ ( .D(n532), .C(net12463), .Q(dpc_tab[3]) );
  DFFQX1 dpc_tab_reg_4__3_ ( .D(n532), .C(net12443), .Q(dpc_tab[27]) );
  DFFQX1 dpc_tab_reg_1__3_ ( .D(N12690), .C(net12458), .Q(dpc_tab[9]) );
  DFFQX1 dpc_tab_reg_5__3_ ( .D(N12690), .C(net12438), .Q(dpc_tab[33]) );
  DFFQX1 dpc_tab_reg_2__3_ ( .D(n532), .C(net12453), .Q(dpc_tab[15]) );
  DFFQX1 dpc_tab_reg_6__3_ ( .D(n532), .C(net12433), .Q(dpc_tab[39]) );
  DFFQX1 dpl_reg_reg_3__7_ ( .D(N12600), .C(net12408), .Q(dpl_reg[31]) );
  DFFQX1 dpl_reg_reg_7__7_ ( .D(N12636), .C(net12388), .Q(dpl_reg[63]) );
  DFFQX1 dpl_reg_reg_0__7_ ( .D(N12573), .C(net12423), .Q(dpl_reg[7]) );
  DFFQX1 dpl_reg_reg_4__7_ ( .D(N12609), .C(net12403), .Q(dpl_reg[39]) );
  DFFQX1 dpl_reg_reg_1__7_ ( .D(N12582), .C(net12418), .Q(dpl_reg[15]) );
  DFFQX1 dpl_reg_reg_5__7_ ( .D(N12618), .C(net12398), .Q(dpl_reg[47]) );
  DFFQX1 dpl_reg_reg_2__7_ ( .D(N12591), .C(net12413), .Q(dpl_reg[23]) );
  DFFQX1 dpl_reg_reg_6__7_ ( .D(N12627), .C(net12393), .Q(dpl_reg[55]) );
  DFFQX1 idle_r_reg ( .D(N512), .C(net12372), .Q(idle_r) );
  DFFQX1 israccess_reg ( .D(N12912), .C(net12372), .Q(israccess) );
  DFFQX1 stop_r_reg ( .D(N515), .C(net12372), .Q(stop_r) );
  DFFQX1 state_reg_2_ ( .D(N590), .C(net12372), .Q(state[2]) );
  DFFQX1 phase_reg_5_ ( .D(N684), .C(net12372), .Q(phase[5]) );
  DFFQX1 state_reg_1_ ( .D(N589), .C(net12372), .Q(state[1]) );
  DFFQX1 state_reg_0_ ( .D(N588), .C(net12372), .Q(state[0]) );
  DFFQX1 ramoe_r_reg ( .D(N11486), .C(net12372), .Q(ramoe) );
  DFFQX1 gf0_reg ( .D(n1881), .C(net12372), .Q(gf0) );
  DFFQX1 ov_reg_reg ( .D(N12711), .C(net12372), .Q(ov) );
  DFFQX1 p_reg ( .D(N12905), .C(net12372), .Q(p) );
  DFFQX1 p2_reg_reg_0_ ( .D(N12485), .C(net12372), .Q(p2[0]) );
  DFFQX1 phase_reg_4_ ( .D(N683), .C(net12372), .Q(phase[4]) );
  DFFQX1 phase_reg_3_ ( .D(N682), .C(net12372), .Q(phase[3]) );
  DFFQX1 idle_s_reg ( .D(n1879), .C(net12372), .Q(idle) );
  DFFQX1 pc_reg_5_ ( .D(N485), .C(net12372), .Q(pc_o[5]) );
  DFFQX1 dpl_reg_reg_3__6_ ( .D(N12599), .C(net12408), .Q(dpl_reg[30]) );
  DFFQX1 dpl_reg_reg_7__6_ ( .D(N12635), .C(net12388), .Q(dpl_reg[62]) );
  DFFQX1 dpl_reg_reg_0__6_ ( .D(N12572), .C(net12423), .Q(dpl_reg[6]) );
  DFFQX1 dpl_reg_reg_4__6_ ( .D(N12608), .C(net12403), .Q(dpl_reg[38]) );
  DFFQX1 dpl_reg_reg_1__6_ ( .D(N12581), .C(net12418), .Q(dpl_reg[14]) );
  DFFQX1 dpl_reg_reg_5__6_ ( .D(N12617), .C(net12398), .Q(dpl_reg[46]) );
  DFFQX1 dpl_reg_reg_2__6_ ( .D(N12590), .C(net12413), .Q(dpl_reg[22]) );
  DFFQX1 dpl_reg_reg_6__6_ ( .D(N12626), .C(net12393), .Q(dpl_reg[54]) );
  DFFQX1 dph_reg_reg_2__0_ ( .D(N12512), .C(net12413), .Q(dph_reg[16]) );
  DFFQX1 f1_reg ( .D(n1883), .C(net12372), .Q(f1) );
  DFFQX1 p2_reg_reg_2_ ( .D(N12487), .C(net12372), .Q(p2[2]) );
  DFFQX1 p2_reg_reg_1_ ( .D(N12486), .C(net12372), .Q(p2[1]) );
  DFFQX1 stop_s_reg ( .D(n1880), .C(net12372), .Q(stop) );
  DFFQX1 dpc_tab_reg_3__2_ ( .D(n519), .C(net12448), .Q(dpc_tab[20]) );
  DFFQX1 dpc_tab_reg_3__0_ ( .D(n538), .C(net12448), .Q(dpc_tab[18]) );
  DFFQX1 dpc_tab_reg_7__0_ ( .D(n538), .C(net12428), .Q(dpc_tab[42]) );
  DFFQX1 dpc_tab_reg_0__2_ ( .D(n2429), .C(net12463), .Q(dpc_tab[2]) );
  DFFQX1 dpc_tab_reg_0__0_ ( .D(n538), .C(net12463), .Q(dpc_tab[0]) );
  DFFQX1 dpc_tab_reg_4__0_ ( .D(n538), .C(net12443), .Q(dpc_tab[24]) );
  DFFQX1 dpc_tab_reg_1__2_ ( .D(n2429), .C(net12458), .Q(dpc_tab[8]) );
  DFFQX1 dpc_tab_reg_1__0_ ( .D(n538), .C(net12458), .Q(dpc_tab[6]) );
  DFFQX1 dpc_tab_reg_5__0_ ( .D(n538), .C(net12438), .Q(dpc_tab[30]) );
  DFFQX1 dpc_tab_reg_2__2_ ( .D(n519), .C(net12453), .Q(dpc_tab[14]) );
  DFFQX1 dpc_tab_reg_2__0_ ( .D(n538), .C(net12453), .Q(dpc_tab[12]) );
  DFFQX1 dpc_tab_reg_6__0_ ( .D(n538), .C(net12433), .Q(dpc_tab[36]) );
  DFFQX1 dph_reg_reg_3__2_ ( .D(N12523), .C(net12408), .Q(dph_reg[26]) );
  DFFQX1 dph_reg_reg_3__1_ ( .D(N12522), .C(net12408), .Q(dph_reg[25]) );
  DFFQX1 dpl_reg_reg_3__5_ ( .D(N12598), .C(net12408), .Q(dpl_reg[29]) );
  DFFQX1 dph_reg_reg_7__2_ ( .D(N12559), .C(net12388), .Q(dph_reg[58]) );
  DFFQX1 dph_reg_reg_7__1_ ( .D(N12558), .C(net12388), .Q(dph_reg[57]) );
  DFFQX1 dpl_reg_reg_7__5_ ( .D(N12634), .C(net12388), .Q(dpl_reg[61]) );
  DFFQX1 dph_reg_reg_7__0_ ( .D(N12557), .C(net12388), .Q(dph_reg[56]) );
  DFFQX1 dph_reg_reg_3__0_ ( .D(N12521), .C(net12408), .Q(dph_reg[24]) );
  DFFQX1 dph_reg_reg_0__2_ ( .D(N12496), .C(net12423), .Q(dph_reg[2]) );
  DFFQX1 dph_reg_reg_0__1_ ( .D(N12495), .C(net12423), .Q(dph_reg[1]) );
  DFFQX1 dpl_reg_reg_0__5_ ( .D(N12571), .C(net12423), .Q(dpl_reg[5]) );
  DFFQX1 dph_reg_reg_4__2_ ( .D(N12532), .C(net12403), .Q(dph_reg[34]) );
  DFFQX1 dph_reg_reg_4__1_ ( .D(N12531), .C(net12403), .Q(dph_reg[33]) );
  DFFQX1 dpl_reg_reg_4__5_ ( .D(N12607), .C(net12403), .Q(dpl_reg[37]) );
  DFFQX1 dph_reg_reg_4__0_ ( .D(N12530), .C(net12403), .Q(dph_reg[32]) );
  DFFQX1 dph_reg_reg_0__0_ ( .D(N12494), .C(net12423), .Q(dph_reg[0]) );
  DFFQX1 dph_reg_reg_1__2_ ( .D(N12505), .C(net12418), .Q(dph_reg[10]) );
  DFFQX1 dph_reg_reg_1__1_ ( .D(N12504), .C(net12418), .Q(dph_reg[9]) );
  DFFQX1 dpl_reg_reg_1__5_ ( .D(N12580), .C(net12418), .Q(dpl_reg[13]) );
  DFFQX1 dph_reg_reg_5__2_ ( .D(N12541), .C(net12398), .Q(dph_reg[42]) );
  DFFQX1 dph_reg_reg_5__1_ ( .D(N12540), .C(net12398), .Q(dph_reg[41]) );
  DFFQX1 dpl_reg_reg_5__5_ ( .D(N12616), .C(net12398), .Q(dpl_reg[45]) );
  DFFQX1 dph_reg_reg_5__0_ ( .D(N12539), .C(net12398), .Q(dph_reg[40]) );
  DFFQX1 dph_reg_reg_1__0_ ( .D(N12503), .C(net12418), .Q(dph_reg[8]) );
  DFFQX1 dph_reg_reg_2__2_ ( .D(N12514), .C(net12413), .Q(dph_reg[18]) );
  DFFQX1 dph_reg_reg_2__1_ ( .D(N12513), .C(net12413), .Q(dph_reg[17]) );
  DFFQX1 dpl_reg_reg_2__5_ ( .D(N12589), .C(net12413), .Q(dpl_reg[21]) );
  DFFQX1 dph_reg_reg_6__2_ ( .D(N12550), .C(net12393), .Q(dph_reg[50]) );
  DFFQX1 dph_reg_reg_6__1_ ( .D(N12549), .C(net12393), .Q(dph_reg[49]) );
  DFFQX1 dpl_reg_reg_6__5_ ( .D(N12625), .C(net12393), .Q(dpl_reg[53]) );
  DFFQX1 dph_reg_reg_6__0_ ( .D(N12548), .C(net12393), .Q(dph_reg[48]) );
  DFFQX1 rmwinstr_reg ( .D(N690), .C(net12372), .Q(rmwinstr) );
  DFFQX1 waitcnt_reg_2_ ( .D(N12976), .C(net12473), .Q(waitcnt[2]) );
  DFFQX1 sfrwe_r_reg ( .D(N11489), .C(net12372), .Q(sfrwe_r) );
  DFFQX1 sfroe_r_reg ( .D(N11488), .C(net12372), .Q(sfroe_r) );
  DFFQX1 rn_reg_reg_7__6_ ( .D(n527), .C(net12513), .Q(rn_reg[198]) );
  DFFQX1 rn_reg_reg_3__6_ ( .D(n527), .C(net12493), .Q(rn_reg[230]) );
  DFFQX1 rn_reg_reg_19__6_ ( .D(n526), .C(net12573), .Q(rn_reg[102]) );
  DFFQX1 rn_reg_reg_23__6_ ( .D(n2434), .C(net12593), .Q(rn_reg[70]) );
  DFFQX1 dpc_tab_reg_3__1_ ( .D(n515), .C(net12448), .Q(dpc_tab[19]) );
  DFFQX1 dpc_tab_reg_7__2_ ( .D(n519), .C(net12428), .Q(dpc_tab[44]) );
  DFFQX1 dpc_tab_reg_7__1_ ( .D(n515), .C(net12428), .Q(dpc_tab[43]) );
  DFFQX1 rn_reg_reg_27__6_ ( .D(n2434), .C(net12613), .Q(rn_reg[38]) );
  DFFQX1 rn_reg_reg_31__6_ ( .D(n528), .C(net12633), .Q(rn_reg[6]) );
  DFFQX1 rn_reg_reg_11__6_ ( .D(n527), .C(net12533), .Q(rn_reg[166]) );
  DFFQX1 rn_reg_reg_15__6_ ( .D(n526), .C(net12553), .Q(rn_reg[134]) );
  DFFQX1 rn_reg_reg_0__6_ ( .D(n528), .C(net12478), .Q(rn_reg[254]) );
  DFFQX1 rn_reg_reg_4__6_ ( .D(n527), .C(net12498), .Q(rn_reg[222]) );
  DFFQX1 rn_reg_reg_16__6_ ( .D(n526), .C(net12558), .Q(rn_reg[126]) );
  DFFQX1 rn_reg_reg_20__6_ ( .D(n526), .C(net12578), .Q(rn_reg[94]) );
  DFFQX1 dpc_tab_reg_0__1_ ( .D(n2428), .C(net12463), .Q(dpc_tab[1]) );
  DFFQX1 dpc_tab_reg_4__2_ ( .D(n519), .C(net12443), .Q(dpc_tab[26]) );
  DFFQX1 dpc_tab_reg_4__1_ ( .D(n515), .C(net12443), .Q(dpc_tab[25]) );
  DFFQX1 rn_reg_reg_24__6_ ( .D(n528), .C(net12598), .Q(rn_reg[62]) );
  DFFQX1 rn_reg_reg_28__6_ ( .D(n528), .C(net12618), .Q(rn_reg[30]) );
  DFFQX1 rn_reg_reg_8__6_ ( .D(n527), .C(net12518), .Q(rn_reg[190]) );
  DFFQX1 rn_reg_reg_12__6_ ( .D(n527), .C(net12538), .Q(rn_reg[158]) );
  DFFQX1 rn_reg_reg_5__6_ ( .D(n527), .C(net12503), .Q(rn_reg[214]) );
  DFFQX1 rn_reg_reg_1__6_ ( .D(n528), .C(net12483), .Q(rn_reg[246]) );
  DFFQX1 rn_reg_reg_17__6_ ( .D(n526), .C(net12563), .Q(rn_reg[118]) );
  DFFQX1 rn_reg_reg_21__6_ ( .D(n526), .C(net12583), .Q(rn_reg[86]) );
  DFFQX1 dpc_tab_reg_1__1_ ( .D(n515), .C(net12458), .Q(dpc_tab[7]) );
  DFFQX1 dpc_tab_reg_5__2_ ( .D(n519), .C(net12438), .Q(dpc_tab[32]) );
  DFFQX1 dpc_tab_reg_5__1_ ( .D(n515), .C(net12438), .Q(dpc_tab[31]) );
  DFFQX1 rn_reg_reg_25__6_ ( .D(n528), .C(net12603), .Q(rn_reg[54]) );
  DFFQX1 rn_reg_reg_29__6_ ( .D(n528), .C(net12623), .Q(rn_reg[22]) );
  DFFQX1 rn_reg_reg_9__6_ ( .D(n527), .C(net12523), .Q(rn_reg[182]) );
  DFFQX1 rn_reg_reg_13__6_ ( .D(n526), .C(net12543), .Q(rn_reg[150]) );
  DFFQX1 rn_reg_reg_2__6_ ( .D(n528), .C(net12488), .Q(rn_reg[238]) );
  DFFQX1 rn_reg_reg_6__6_ ( .D(n527), .C(net12508), .Q(rn_reg[206]) );
  DFFQX1 rn_reg_reg_18__6_ ( .D(n526), .C(net12568), .Q(rn_reg[110]) );
  DFFQX1 rn_reg_reg_22__6_ ( .D(n526), .C(net12588), .Q(rn_reg[78]) );
  DFFQX1 dpc_tab_reg_2__1_ ( .D(n515), .C(net12453), .Q(dpc_tab[13]) );
  DFFQX1 dpc_tab_reg_6__2_ ( .D(n519), .C(net12433), .Q(dpc_tab[38]) );
  DFFQX1 dpc_tab_reg_6__1_ ( .D(n515), .C(net12433), .Q(dpc_tab[37]) );
  DFFQX1 rn_reg_reg_26__6_ ( .D(n528), .C(net12608), .Q(rn_reg[46]) );
  DFFQX1 rn_reg_reg_30__6_ ( .D(n528), .C(net12628), .Q(rn_reg[14]) );
  DFFQX1 rn_reg_reg_10__6_ ( .D(n527), .C(net12528), .Q(rn_reg[174]) );
  DFFQX1 rn_reg_reg_14__6_ ( .D(n526), .C(net12548), .Q(rn_reg[142]) );
  DFFQX1 dec_cop_reg_0_ ( .D(N10582), .C(net12372), .Q(dec_cop[0]) );
  DFFQX1 dpl_reg_reg_3__4_ ( .D(N12597), .C(net12408), .Q(dpl_reg[28]) );
  DFFQX1 dpl_reg_reg_7__4_ ( .D(N12633), .C(net12388), .Q(dpl_reg[60]) );
  DFFQX1 dpl_reg_reg_0__4_ ( .D(N12570), .C(net12423), .Q(dpl_reg[4]) );
  DFFQX1 dpl_reg_reg_4__4_ ( .D(N12606), .C(net12403), .Q(dpl_reg[36]) );
  DFFQX1 dpl_reg_reg_1__4_ ( .D(N12579), .C(net12418), .Q(dpl_reg[12]) );
  DFFQX1 dpl_reg_reg_5__4_ ( .D(N12615), .C(net12398), .Q(dpl_reg[44]) );
  DFFQX1 dpl_reg_reg_2__4_ ( .D(N12588), .C(net12413), .Q(dpl_reg[20]) );
  DFFQX1 dpl_reg_reg_6__4_ ( .D(N12624), .C(net12393), .Q(dpl_reg[52]) );
  DFFQX1 waitcnt_reg_1_ ( .D(N12975), .C(net12473), .Q(waitcnt[1]) );
  DFFQX1 waitcnt_reg_0_ ( .D(N12974), .C(net12473), .Q(waitcnt[0]) );
  DFFQX1 ckcon_r_reg_5_ ( .D(N12970), .C(net12372), .Q(ckcon[5]) );
  DFFQX1 ckcon_r_reg_2_ ( .D(N12967), .C(net12372), .Q(ckcon[2]) );
  DFFQX1 ckcon_r_reg_6_ ( .D(N12971), .C(net12372), .Q(ckcon[6]) );
  DFFQX1 ckcon_r_reg_1_ ( .D(N12966), .C(net12372), .Q(ckcon[1]) );
  DFFQX1 mempsrd_r_reg ( .D(N582), .C(net12372), .Q(mempsrd) );
  DFFQX1 memwr_s_reg ( .D(N585), .C(net12372), .Q(memwr) );
  DFFQX1 mempswr_s_reg ( .D(N583), .C(net12372), .Q(mempswr) );
  DFFQX1 rn_reg_reg_3__2_ ( .D(n519), .C(net12493), .Q(rn_reg[226]) );
  DFFQX1 rn_reg_reg_7__2_ ( .D(n518), .C(net12513), .Q(rn_reg[194]) );
  DFFQX1 rn_reg_reg_7__5_ ( .D(n520), .C(net12513), .Q(rn_reg[197]) );
  DFFQX1 rn_reg_reg_3__5_ ( .D(n520), .C(net12493), .Q(rn_reg[229]) );
  DFFQX1 rn_reg_reg_19__5_ ( .D(n521), .C(net12573), .Q(rn_reg[101]) );
  DFFQX1 rn_reg_reg_19__2_ ( .D(n517), .C(net12573), .Q(rn_reg[98]) );
  DFFQX1 rn_reg_reg_23__5_ ( .D(n522), .C(net12593), .Q(rn_reg[69]) );
  DFFQX1 rn_reg_reg_23__2_ ( .D(n517), .C(net12593), .Q(rn_reg[66]) );
  DFFQX1 rn_reg_reg_27__5_ ( .D(n522), .C(net12613), .Q(rn_reg[37]) );
  DFFQX1 rn_reg_reg_27__2_ ( .D(n516), .C(net12613), .Q(rn_reg[34]) );
  DFFQX1 rn_reg_reg_31__5_ ( .D(n2430), .C(net12633), .Q(rn_reg[5]) );
  DFFQX1 rn_reg_reg_31__2_ ( .D(n516), .C(net12633), .Q(rn_reg[2]) );
  DFFQX1 rn_reg_reg_11__5_ ( .D(n520), .C(net12533), .Q(rn_reg[165]) );
  DFFQX1 rn_reg_reg_11__2_ ( .D(n518), .C(net12533), .Q(rn_reg[162]) );
  DFFQX1 rn_reg_reg_15__5_ ( .D(n521), .C(net12553), .Q(rn_reg[133]) );
  DFFQX1 rn_reg_reg_15__2_ ( .D(n517), .C(net12553), .Q(rn_reg[130]) );
  DFFQX1 rn_reg_reg_0__2_ ( .D(n2429), .C(net12478), .Q(rn_reg[250]) );
  DFFQX1 rn_reg_reg_4__2_ ( .D(n519), .C(net12498), .Q(rn_reg[218]) );
  DFFQX1 rn_reg_reg_0__5_ ( .D(n2430), .C(net12478), .Q(rn_reg[253]) );
  DFFQX1 rn_reg_reg_4__5_ ( .D(n520), .C(net12498), .Q(rn_reg[221]) );
  DFFQX1 rn_reg_reg_16__5_ ( .D(n521), .C(net12558), .Q(rn_reg[125]) );
  DFFQX1 rn_reg_reg_16__2_ ( .D(n517), .C(net12558), .Q(rn_reg[122]) );
  DFFQX1 rn_reg_reg_20__5_ ( .D(n521), .C(net12578), .Q(rn_reg[93]) );
  DFFQX1 rn_reg_reg_20__2_ ( .D(n517), .C(net12578), .Q(rn_reg[90]) );
  DFFQX1 rn_reg_reg_24__5_ ( .D(n522), .C(net12598), .Q(rn_reg[61]) );
  DFFQX1 rn_reg_reg_24__2_ ( .D(n517), .C(net12598), .Q(rn_reg[58]) );
  DFFQX1 rn_reg_reg_28__5_ ( .D(n522), .C(net12618), .Q(rn_reg[29]) );
  DFFQX1 rn_reg_reg_28__2_ ( .D(n516), .C(net12618), .Q(rn_reg[26]) );
  DFFQX1 rn_reg_reg_8__5_ ( .D(n520), .C(net12518), .Q(rn_reg[189]) );
  DFFQX1 rn_reg_reg_8__2_ ( .D(n518), .C(net12518), .Q(rn_reg[186]) );
  DFFQX1 rn_reg_reg_12__5_ ( .D(n520), .C(net12538), .Q(rn_reg[157]) );
  DFFQX1 rn_reg_reg_12__2_ ( .D(n518), .C(net12538), .Q(rn_reg[154]) );
  DFFQX1 rn_reg_reg_1__2_ ( .D(n519), .C(net12483), .Q(rn_reg[242]) );
  DFFQX1 rn_reg_reg_5__2_ ( .D(n518), .C(net12503), .Q(rn_reg[210]) );
  DFFQX1 rn_reg_reg_5__5_ ( .D(n520), .C(net12503), .Q(rn_reg[213]) );
  DFFQX1 rn_reg_reg_1__5_ ( .D(n2430), .C(net12483), .Q(rn_reg[245]) );
  DFFQX1 rn_reg_reg_17__5_ ( .D(n521), .C(net12563), .Q(rn_reg[117]) );
  DFFQX1 rn_reg_reg_17__2_ ( .D(n517), .C(net12563), .Q(rn_reg[114]) );
  DFFQX1 rn_reg_reg_21__5_ ( .D(n521), .C(net12583), .Q(rn_reg[85]) );
  DFFQX1 rn_reg_reg_21__2_ ( .D(n517), .C(net12583), .Q(rn_reg[82]) );
  DFFQX1 rn_reg_reg_25__5_ ( .D(n522), .C(net12603), .Q(rn_reg[53]) );
  DFFQX1 rn_reg_reg_25__2_ ( .D(n516), .C(net12603), .Q(rn_reg[50]) );
  DFFQX1 rn_reg_reg_29__5_ ( .D(n522), .C(net12623), .Q(rn_reg[21]) );
  DFFQX1 rn_reg_reg_29__2_ ( .D(n516), .C(net12623), .Q(rn_reg[18]) );
  DFFQX1 rn_reg_reg_9__5_ ( .D(n520), .C(net12523), .Q(rn_reg[181]) );
  DFFQX1 rn_reg_reg_9__2_ ( .D(n518), .C(net12523), .Q(rn_reg[178]) );
  DFFQX1 rn_reg_reg_13__5_ ( .D(n521), .C(net12543), .Q(rn_reg[149]) );
  DFFQX1 rn_reg_reg_13__2_ ( .D(n518), .C(net12543), .Q(rn_reg[146]) );
  DFFQX1 rn_reg_reg_2__2_ ( .D(n519), .C(net12488), .Q(rn_reg[234]) );
  DFFQX1 rn_reg_reg_6__2_ ( .D(n518), .C(net12508), .Q(rn_reg[202]) );
  DFFQX1 rn_reg_reg_2__5_ ( .D(n522), .C(net12488), .Q(rn_reg[237]) );
  DFFQX1 rn_reg_reg_6__5_ ( .D(n520), .C(net12508), .Q(rn_reg[205]) );
  DFFQX1 rn_reg_reg_18__5_ ( .D(n521), .C(net12568), .Q(rn_reg[109]) );
  DFFQX1 rn_reg_reg_18__2_ ( .D(n517), .C(net12568), .Q(rn_reg[106]) );
  DFFQX1 rn_reg_reg_22__5_ ( .D(n522), .C(net12588), .Q(rn_reg[77]) );
  DFFQX1 rn_reg_reg_22__2_ ( .D(n517), .C(net12588), .Q(rn_reg[74]) );
  DFFQX1 rn_reg_reg_26__5_ ( .D(n522), .C(net12608), .Q(rn_reg[45]) );
  DFFQX1 rn_reg_reg_26__2_ ( .D(n516), .C(net12608), .Q(rn_reg[42]) );
  DFFQX1 rn_reg_reg_30__5_ ( .D(n522), .C(net12628), .Q(rn_reg[13]) );
  DFFQX1 rn_reg_reg_30__2_ ( .D(n516), .C(net12628), .Q(rn_reg[10]) );
  DFFQX1 rn_reg_reg_10__5_ ( .D(n520), .C(net12528), .Q(rn_reg[173]) );
  DFFQX1 rn_reg_reg_10__2_ ( .D(n518), .C(net12528), .Q(rn_reg[170]) );
  DFFQX1 rn_reg_reg_14__5_ ( .D(n521), .C(net12548), .Q(rn_reg[141]) );
  DFFQX1 rn_reg_reg_14__2_ ( .D(n518), .C(net12548), .Q(rn_reg[138]) );
  DFFQX1 dpl_reg_reg_3__3_ ( .D(N12596), .C(net12408), .Q(dpl_reg[27]) );
  DFFQX1 dpl_reg_reg_3__2_ ( .D(N12595), .C(net12408), .Q(dpl_reg[26]) );
  DFFQX1 dpl_reg_reg_3__1_ ( .D(N12594), .C(net12408), .Q(dpl_reg[25]) );
  DFFQX1 dpl_reg_reg_7__3_ ( .D(N12632), .C(net12388), .Q(dpl_reg[59]) );
  DFFQX1 dpl_reg_reg_7__2_ ( .D(N12631), .C(net12388), .Q(dpl_reg[58]) );
  DFFQX1 dpl_reg_reg_0__3_ ( .D(N12569), .C(net12423), .Q(dpl_reg[3]) );
  DFFQX1 dpl_reg_reg_0__2_ ( .D(N12568), .C(net12423), .Q(dpl_reg[2]) );
  DFFQX1 dpl_reg_reg_4__3_ ( .D(N12605), .C(net12403), .Q(dpl_reg[35]) );
  DFFQX1 dpl_reg_reg_4__2_ ( .D(N12604), .C(net12403), .Q(dpl_reg[34]) );
  DFFQX1 dpl_reg_reg_1__3_ ( .D(N12578), .C(net12418), .Q(dpl_reg[11]) );
  DFFQX1 dpl_reg_reg_1__2_ ( .D(N12577), .C(net12418), .Q(dpl_reg[10]) );
  DFFQX1 dpl_reg_reg_5__3_ ( .D(N12614), .C(net12398), .Q(dpl_reg[43]) );
  DFFQX1 dpl_reg_reg_5__2_ ( .D(N12613), .C(net12398), .Q(dpl_reg[42]) );
  DFFQX1 dpl_reg_reg_2__3_ ( .D(N12587), .C(net12413), .Q(dpl_reg[19]) );
  DFFQX1 dpl_reg_reg_2__2_ ( .D(N12586), .C(net12413), .Q(dpl_reg[18]) );
  DFFQX1 dpl_reg_reg_2__1_ ( .D(N12585), .C(net12413), .Q(dpl_reg[17]) );
  DFFQX1 dpl_reg_reg_6__3_ ( .D(N12623), .C(net12393), .Q(dpl_reg[51]) );
  DFFQX1 dpl_reg_reg_6__2_ ( .D(N12622), .C(net12393), .Q(dpl_reg[50]) );
  DFFQX1 dec_cop_reg_5_ ( .D(N10587), .C(net12372), .Q(dec_cop[5]) );
  DFFQX1 multempreg_reg_1_ ( .D(N13326), .C(net12638), .Q(multempreg[1]) );
  DFFQX1 ramwe_r_reg ( .D(N11487), .C(net12372), .Q(ramwe) );
  DFFQX1 dec_cop_reg_2_ ( .D(N10584), .C(net12372), .Q(dec_cop[2]) );
  DFFQX1 dec_cop_reg_1_ ( .D(N10583), .C(net12372), .Q(dec_cop[1]) );
  DFFQX1 memrd_s_reg ( .D(N584), .C(net12372), .Q(memrd) );
  DFFQX1 sp_reg_reg_5_ ( .D(N12702), .C(net12372), .Q(sp[5]) );
  DFFQX1 ckcon_r_reg_4_ ( .D(N12969), .C(net12372), .Q(ckcon[4]) );
  DFFQX1 sp_reg_reg_6_ ( .D(N12703), .C(net12372), .Q(sp[6]) );
  DFFQX1 sp_reg_reg_7_ ( .D(N12704), .C(net12372), .Q(sp[7]) );
  DFFQX1 ckcon_r_reg_3_ ( .D(N12968), .C(net12372), .Q(ckcon[3]) );
  DFFQX1 temp2_reg_7_ ( .D(N12730), .C(net12372), .Q(temp2_comb[7]) );
  DFFQX1 ckcon_r_reg_7_ ( .D(N12972), .C(net12372), .Q(ckcon[7]) );
  DFFQX1 dec_cop_reg_7_ ( .D(N10589), .C(net12372), .Q(dec_cop[7]) );
  DFFQX1 ckcon_r_reg_0_ ( .D(N12965), .C(net12372), .Q(ckcon[0]) );
  DFFQX1 phase_reg_2_ ( .D(N681), .C(net12372), .Q(phase[2]) );
  DFFQX1 dec_accop_reg_17_ ( .D(n217), .C(net12372), .Q(dec_accop[17]) );
  DFFQX1 ramdatao_r_reg_7_ ( .D(N11505), .C(net12372), .Q(ramdatao[7]) );
  DFFQX1 ramdatao_r_reg_6_ ( .D(N11504), .C(net12372), .Q(ramdatao[6]) );
  DFFQX1 ramdatao_r_reg_5_ ( .D(N11503), .C(net12372), .Q(ramdatao[5]) );
  DFFQX1 rn_reg_reg_3__7_ ( .D(n525), .C(net12493), .Q(rn_reg[231]) );
  DFFQX1 rn_reg_reg_3__3_ ( .D(n532), .C(net12493), .Q(rn_reg[227]) );
  DFFQX1 rn_reg_reg_3__1_ ( .D(n515), .C(net12493), .Q(rn_reg[225]) );
  DFFQX1 rn_reg_reg_3__0_ ( .D(n537), .C(net12493), .Q(rn_reg[224]) );
  DFFQX1 rn_reg_reg_7__7_ ( .D(n525), .C(net12513), .Q(rn_reg[199]) );
  DFFQX1 rn_reg_reg_7__3_ ( .D(n533), .C(net12513), .Q(rn_reg[195]) );
  DFFQX1 rn_reg_reg_7__1_ ( .D(n514), .C(net12513), .Q(rn_reg[193]) );
  DFFQX1 rn_reg_reg_7__0_ ( .D(n537), .C(net12513), .Q(rn_reg[192]) );
  DFFQX1 rn_reg_reg_7__4_ ( .D(n529), .C(net12513), .Q(rn_reg[196]) );
  DFFQX1 rn_reg_reg_3__4_ ( .D(n2436), .C(net12493), .Q(rn_reg[228]) );
  DFFQX1 rn_reg_reg_19__7_ ( .D(n524), .C(net12573), .Q(rn_reg[103]) );
  DFFQX1 rn_reg_reg_19__4_ ( .D(n530), .C(net12573), .Q(rn_reg[100]) );
  DFFQX1 rn_reg_reg_19__3_ ( .D(n534), .C(net12573), .Q(rn_reg[99]) );
  DFFQX1 rn_reg_reg_19__1_ ( .D(n513), .C(net12573), .Q(rn_reg[97]) );
  DFFQX1 rn_reg_reg_19__0_ ( .D(n536), .C(net12573), .Q(rn_reg[96]) );
  DFFQX1 rn_reg_reg_23__7_ ( .D(n523), .C(net12593), .Q(rn_reg[71]) );
  DFFQX1 rn_reg_reg_23__4_ ( .D(n531), .C(net12593), .Q(rn_reg[68]) );
  DFFQX1 rn_reg_reg_23__3_ ( .D(n2438), .C(net12593), .Q(rn_reg[67]) );
  DFFQX1 rn_reg_reg_23__1_ ( .D(n513), .C(net12593), .Q(rn_reg[65]) );
  DFFQX1 rn_reg_reg_23__0_ ( .D(n535), .C(net12593), .Q(rn_reg[64]) );
  DFFQX1 rn_reg_reg_27__7_ ( .D(n523), .C(net12613), .Q(rn_reg[39]) );
  DFFQX1 rn_reg_reg_27__4_ ( .D(n531), .C(net12613), .Q(rn_reg[36]) );
  DFFQX1 rn_reg_reg_27__3_ ( .D(n2438), .C(net12613), .Q(rn_reg[35]) );
  DFFQX1 rn_reg_reg_27__1_ ( .D(n512), .C(net12613), .Q(rn_reg[33]) );
  DFFQX1 rn_reg_reg_27__0_ ( .D(n535), .C(net12613), .Q(rn_reg[32]) );
  DFFQX1 rn_reg_reg_31__7_ ( .D(n523), .C(net12633), .Q(rn_reg[7]) );
  DFFQX1 rn_reg_reg_31__4_ ( .D(n2436), .C(net12633), .Q(rn_reg[4]) );
  DFFQX1 rn_reg_reg_31__3_ ( .D(n532), .C(net12633), .Q(rn_reg[3]) );
  DFFQX1 rn_reg_reg_31__1_ ( .D(n512), .C(net12633), .Q(rn_reg[1]) );
  DFFQX1 rn_reg_reg_31__0_ ( .D(n535), .C(net12633), .Q(rn_reg[0]) );
  DFFQX1 rn_reg_reg_11__7_ ( .D(n525), .C(net12533), .Q(rn_reg[167]) );
  DFFQX1 rn_reg_reg_11__4_ ( .D(n529), .C(net12533), .Q(rn_reg[164]) );
  DFFQX1 rn_reg_reg_11__3_ ( .D(n533), .C(net12533), .Q(rn_reg[163]) );
  DFFQX1 rn_reg_reg_11__1_ ( .D(n514), .C(net12533), .Q(rn_reg[161]) );
  DFFQX1 rn_reg_reg_11__0_ ( .D(n537), .C(net12533), .Q(rn_reg[160]) );
  DFFQX1 rn_reg_reg_15__7_ ( .D(n524), .C(net12553), .Q(rn_reg[135]) );
  DFFQX1 rn_reg_reg_15__4_ ( .D(n530), .C(net12553), .Q(rn_reg[132]) );
  DFFQX1 rn_reg_reg_15__3_ ( .D(n534), .C(net12553), .Q(rn_reg[131]) );
  DFFQX1 rn_reg_reg_15__1_ ( .D(n513), .C(net12553), .Q(rn_reg[129]) );
  DFFQX1 rn_reg_reg_15__0_ ( .D(n536), .C(net12553), .Q(rn_reg[128]) );
  DFFQX1 rn_reg_reg_0__7_ ( .D(n2431), .C(net12478), .Q(rn_reg[255]) );
  DFFQX1 rn_reg_reg_0__3_ ( .D(n534), .C(net12478), .Q(rn_reg[251]) );
  DFFQX1 rn_reg_reg_0__1_ ( .D(n2428), .C(net12478), .Q(rn_reg[249]) );
  DFFQX1 rn_reg_reg_0__0_ ( .D(n2440), .C(net12478), .Q(rn_reg[248]) );
  DFFQX1 rn_reg_reg_4__7_ ( .D(n525), .C(net12498), .Q(rn_reg[223]) );
  DFFQX1 rn_reg_reg_4__3_ ( .D(n533), .C(net12498), .Q(rn_reg[219]) );
  DFFQX1 rn_reg_reg_4__1_ ( .D(n514), .C(net12498), .Q(rn_reg[217]) );
  DFFQX1 rn_reg_reg_4__0_ ( .D(n537), .C(net12498), .Q(rn_reg[216]) );
  DFFQX1 rn_reg_reg_0__4_ ( .D(n530), .C(net12478), .Q(rn_reg[252]) );
  DFFQX1 rn_reg_reg_4__4_ ( .D(n529), .C(net12498), .Q(rn_reg[220]) );
  DFFQX1 rn_reg_reg_16__7_ ( .D(n524), .C(net12558), .Q(rn_reg[127]) );
  DFFQX1 rn_reg_reg_16__4_ ( .D(n530), .C(net12558), .Q(rn_reg[124]) );
  DFFQX1 rn_reg_reg_16__3_ ( .D(n534), .C(net12558), .Q(rn_reg[123]) );
  DFFQX1 rn_reg_reg_16__1_ ( .D(n513), .C(net12558), .Q(rn_reg[121]) );
  DFFQX1 rn_reg_reg_16__0_ ( .D(n536), .C(net12558), .Q(rn_reg[120]) );
  DFFQX1 rn_reg_reg_20__7_ ( .D(n524), .C(net12578), .Q(rn_reg[95]) );
  DFFQX1 rn_reg_reg_20__4_ ( .D(n530), .C(net12578), .Q(rn_reg[92]) );
  DFFQX1 rn_reg_reg_20__3_ ( .D(n534), .C(net12578), .Q(rn_reg[91]) );
  DFFQX1 rn_reg_reg_20__1_ ( .D(n513), .C(net12578), .Q(rn_reg[89]) );
  DFFQX1 rn_reg_reg_20__0_ ( .D(n536), .C(net12578), .Q(rn_reg[88]) );
  DFFQX1 rn_reg_reg_24__7_ ( .D(n523), .C(net12598), .Q(rn_reg[63]) );
  DFFQX1 rn_reg_reg_24__4_ ( .D(n531), .C(net12598), .Q(rn_reg[60]) );
  DFFQX1 rn_reg_reg_24__3_ ( .D(n2438), .C(net12598), .Q(rn_reg[59]) );
  DFFQX1 rn_reg_reg_24__1_ ( .D(n512), .C(net12598), .Q(rn_reg[57]) );
  DFFQX1 rn_reg_reg_24__0_ ( .D(n535), .C(net12598), .Q(rn_reg[56]) );
  DFFQX1 rn_reg_reg_28__7_ ( .D(n523), .C(net12618), .Q(rn_reg[31]) );
  DFFQX1 rn_reg_reg_28__4_ ( .D(n531), .C(net12618), .Q(rn_reg[28]) );
  DFFQX1 rn_reg_reg_28__3_ ( .D(n2438), .C(net12618), .Q(rn_reg[27]) );
  DFFQX1 rn_reg_reg_28__1_ ( .D(n512), .C(net12618), .Q(rn_reg[25]) );
  DFFQX1 rn_reg_reg_28__0_ ( .D(n535), .C(net12618), .Q(rn_reg[24]) );
  DFFQX1 rn_reg_reg_8__7_ ( .D(n525), .C(net12518), .Q(rn_reg[191]) );
  DFFQX1 rn_reg_reg_8__4_ ( .D(n529), .C(net12518), .Q(rn_reg[188]) );
  DFFQX1 rn_reg_reg_8__3_ ( .D(n533), .C(net12518), .Q(rn_reg[187]) );
  DFFQX1 rn_reg_reg_8__1_ ( .D(n514), .C(net12518), .Q(rn_reg[185]) );
  DFFQX1 rn_reg_reg_8__0_ ( .D(n537), .C(net12518), .Q(rn_reg[184]) );
  DFFQX1 rn_reg_reg_12__7_ ( .D(n524), .C(net12538), .Q(rn_reg[159]) );
  DFFQX1 rn_reg_reg_12__4_ ( .D(n529), .C(net12538), .Q(rn_reg[156]) );
  DFFQX1 rn_reg_reg_12__3_ ( .D(n533), .C(net12538), .Q(rn_reg[155]) );
  DFFQX1 rn_reg_reg_12__1_ ( .D(n514), .C(net12538), .Q(rn_reg[153]) );
  DFFQX1 rn_reg_reg_12__0_ ( .D(n537), .C(net12538), .Q(rn_reg[152]) );
  DFFQX1 rn_reg_reg_1__7_ ( .D(n2431), .C(net12483), .Q(rn_reg[247]) );
  DFFQX1 rn_reg_reg_1__3_ ( .D(n532), .C(net12483), .Q(rn_reg[243]) );
  DFFQX1 rn_reg_reg_1__1_ ( .D(n515), .C(net12483), .Q(rn_reg[241]) );
  DFFQX1 rn_reg_reg_1__0_ ( .D(n538), .C(net12483), .Q(rn_reg[240]) );
  DFFQX1 rn_reg_reg_5__7_ ( .D(n525), .C(net12503), .Q(rn_reg[215]) );
  DFFQX1 rn_reg_reg_5__3_ ( .D(n533), .C(net12503), .Q(rn_reg[211]) );
  DFFQX1 rn_reg_reg_5__1_ ( .D(n514), .C(net12503), .Q(rn_reg[209]) );
  DFFQX1 rn_reg_reg_5__0_ ( .D(n537), .C(net12503), .Q(rn_reg[208]) );
  DFFQX1 rn_reg_reg_5__4_ ( .D(n529), .C(net12503), .Q(rn_reg[212]) );
  DFFQX1 rn_reg_reg_1__4_ ( .D(n531), .C(net12483), .Q(rn_reg[244]) );
  DFFQX1 rn_reg_reg_17__7_ ( .D(n524), .C(net12563), .Q(rn_reg[119]) );
  DFFQX1 rn_reg_reg_17__4_ ( .D(n530), .C(net12563), .Q(rn_reg[116]) );
  DFFQX1 rn_reg_reg_17__3_ ( .D(n534), .C(net12563), .Q(rn_reg[115]) );
  DFFQX1 rn_reg_reg_17__1_ ( .D(n513), .C(net12563), .Q(rn_reg[113]) );
  DFFQX1 rn_reg_reg_17__0_ ( .D(n536), .C(net12563), .Q(rn_reg[112]) );
  DFFQX1 rn_reg_reg_21__7_ ( .D(n524), .C(net12583), .Q(rn_reg[87]) );
  DFFQX1 rn_reg_reg_21__4_ ( .D(n530), .C(net12583), .Q(rn_reg[84]) );
  DFFQX1 rn_reg_reg_21__3_ ( .D(n534), .C(net12583), .Q(rn_reg[83]) );
  DFFQX1 rn_reg_reg_21__1_ ( .D(n513), .C(net12583), .Q(rn_reg[81]) );
  DFFQX1 rn_reg_reg_21__0_ ( .D(n536), .C(net12583), .Q(rn_reg[80]) );
  DFFQX1 rn_reg_reg_25__7_ ( .D(n523), .C(net12603), .Q(rn_reg[55]) );
  DFFQX1 rn_reg_reg_25__4_ ( .D(n531), .C(net12603), .Q(rn_reg[52]) );
  DFFQX1 rn_reg_reg_25__3_ ( .D(n2438), .C(net12603), .Q(rn_reg[51]) );
  DFFQX1 rn_reg_reg_25__1_ ( .D(n512), .C(net12603), .Q(rn_reg[49]) );
  DFFQX1 rn_reg_reg_25__0_ ( .D(n535), .C(net12603), .Q(rn_reg[48]) );
  DFFQX1 rn_reg_reg_29__7_ ( .D(n523), .C(net12623), .Q(rn_reg[23]) );
  DFFQX1 rn_reg_reg_29__4_ ( .D(n531), .C(net12623), .Q(rn_reg[20]) );
  DFFQX1 rn_reg_reg_29__3_ ( .D(n2438), .C(net12623), .Q(rn_reg[19]) );
  DFFQX1 rn_reg_reg_29__1_ ( .D(n512), .C(net12623), .Q(rn_reg[17]) );
  DFFQX1 rn_reg_reg_29__0_ ( .D(n535), .C(net12623), .Q(rn_reg[16]) );
  DFFQX1 rn_reg_reg_9__7_ ( .D(n525), .C(net12523), .Q(rn_reg[183]) );
  DFFQX1 rn_reg_reg_9__4_ ( .D(n529), .C(net12523), .Q(rn_reg[180]) );
  DFFQX1 rn_reg_reg_9__3_ ( .D(n533), .C(net12523), .Q(rn_reg[179]) );
  DFFQX1 rn_reg_reg_9__1_ ( .D(n514), .C(net12523), .Q(rn_reg[177]) );
  DFFQX1 rn_reg_reg_9__0_ ( .D(n537), .C(net12523), .Q(rn_reg[176]) );
  DFFQX1 rn_reg_reg_13__7_ ( .D(n524), .C(net12543), .Q(rn_reg[151]) );
  DFFQX1 rn_reg_reg_13__4_ ( .D(n529), .C(net12543), .Q(rn_reg[148]) );
  DFFQX1 rn_reg_reg_13__3_ ( .D(n533), .C(net12543), .Q(rn_reg[147]) );
  DFFQX1 rn_reg_reg_13__1_ ( .D(n514), .C(net12543), .Q(rn_reg[145]) );
  DFFQX1 rn_reg_reg_13__0_ ( .D(n536), .C(net12543), .Q(rn_reg[144]) );
  DFFQX1 rn_reg_reg_2__7_ ( .D(n525), .C(net12488), .Q(rn_reg[239]) );
  DFFQX1 rn_reg_reg_2__3_ ( .D(n532), .C(net12488), .Q(rn_reg[235]) );
  DFFQX1 rn_reg_reg_2__1_ ( .D(n515), .C(net12488), .Q(rn_reg[233]) );
  DFFQX1 rn_reg_reg_2__0_ ( .D(n538), .C(net12488), .Q(rn_reg[232]) );
  DFFQX1 rn_reg_reg_6__7_ ( .D(n525), .C(net12508), .Q(rn_reg[207]) );
  DFFQX1 rn_reg_reg_6__3_ ( .D(n533), .C(net12508), .Q(rn_reg[203]) );
  DFFQX1 rn_reg_reg_6__1_ ( .D(n514), .C(net12508), .Q(rn_reg[201]) );
  DFFQX1 rn_reg_reg_6__0_ ( .D(n537), .C(net12508), .Q(rn_reg[200]) );
  DFFQX1 rn_reg_reg_2__4_ ( .D(n531), .C(net12488), .Q(rn_reg[236]) );
  DFFQX1 rn_reg_reg_6__4_ ( .D(n529), .C(net12508), .Q(rn_reg[204]) );
  DFFQX1 rn_reg_reg_18__7_ ( .D(n524), .C(net12568), .Q(rn_reg[111]) );
  DFFQX1 rn_reg_reg_18__4_ ( .D(n530), .C(net12568), .Q(rn_reg[108]) );
  DFFQX1 rn_reg_reg_18__3_ ( .D(n534), .C(net12568), .Q(rn_reg[107]) );
  DFFQX1 rn_reg_reg_18__1_ ( .D(n513), .C(net12568), .Q(rn_reg[105]) );
  DFFQX1 rn_reg_reg_18__0_ ( .D(n536), .C(net12568), .Q(rn_reg[104]) );
  DFFQX1 rn_reg_reg_22__7_ ( .D(n523), .C(net12588), .Q(rn_reg[79]) );
  DFFQX1 rn_reg_reg_22__4_ ( .D(n530), .C(net12588), .Q(rn_reg[76]) );
  DFFQX1 rn_reg_reg_22__3_ ( .D(n534), .C(net12588), .Q(rn_reg[75]) );
  DFFQX1 rn_reg_reg_22__1_ ( .D(n513), .C(net12588), .Q(rn_reg[73]) );
  DFFQX1 rn_reg_reg_22__0_ ( .D(n536), .C(net12588), .Q(rn_reg[72]) );
  DFFQX1 rn_reg_reg_26__7_ ( .D(n523), .C(net12608), .Q(rn_reg[47]) );
  DFFQX1 rn_reg_reg_26__4_ ( .D(n531), .C(net12608), .Q(rn_reg[44]) );
  DFFQX1 rn_reg_reg_26__3_ ( .D(n2438), .C(net12608), .Q(rn_reg[43]) );
  DFFQX1 rn_reg_reg_26__1_ ( .D(n512), .C(net12608), .Q(rn_reg[41]) );
  DFFQX1 rn_reg_reg_26__0_ ( .D(n535), .C(net12608), .Q(rn_reg[40]) );
  DFFQX1 rn_reg_reg_30__7_ ( .D(n523), .C(net12628), .Q(rn_reg[15]) );
  DFFQX1 rn_reg_reg_30__4_ ( .D(n531), .C(net12628), .Q(rn_reg[12]) );
  DFFQX1 rn_reg_reg_30__3_ ( .D(n2438), .C(net12628), .Q(rn_reg[11]) );
  DFFQX1 rn_reg_reg_30__1_ ( .D(n512), .C(net12628), .Q(rn_reg[9]) );
  DFFQX1 rn_reg_reg_30__0_ ( .D(n535), .C(net12628), .Q(rn_reg[8]) );
  DFFQX1 rn_reg_reg_10__7_ ( .D(n525), .C(net12528), .Q(rn_reg[175]) );
  DFFQX1 rn_reg_reg_10__4_ ( .D(n529), .C(net12528), .Q(rn_reg[172]) );
  DFFQX1 rn_reg_reg_10__3_ ( .D(n533), .C(net12528), .Q(rn_reg[171]) );
  DFFQX1 rn_reg_reg_10__1_ ( .D(n514), .C(net12528), .Q(rn_reg[169]) );
  DFFQX1 rn_reg_reg_10__0_ ( .D(n537), .C(net12528), .Q(rn_reg[168]) );
  DFFQX1 rn_reg_reg_14__7_ ( .D(n524), .C(net12548), .Q(rn_reg[143]) );
  DFFQX1 rn_reg_reg_14__4_ ( .D(n530), .C(net12548), .Q(rn_reg[140]) );
  DFFQX1 rn_reg_reg_14__3_ ( .D(n534), .C(net12548), .Q(rn_reg[139]) );
  DFFQX1 rn_reg_reg_14__1_ ( .D(n513), .C(net12548), .Q(rn_reg[137]) );
  DFFQX1 rn_reg_reg_14__0_ ( .D(n536), .C(net12548), .Q(rn_reg[136]) );
  DFFQX1 dpl_reg_reg_3__0_ ( .D(N12593), .C(net12408), .Q(dpl_reg[24]) );
  DFFQX1 dpl_reg_reg_7__1_ ( .D(N12630), .C(net12388), .Q(dpl_reg[57]) );
  DFFQX1 dpl_reg_reg_7__0_ ( .D(N12629), .C(net12388), .Q(dpl_reg[56]) );
  DFFQX1 dpl_reg_reg_0__1_ ( .D(N12567), .C(net12423), .Q(dpl_reg[1]) );
  DFFQX1 dpl_reg_reg_0__0_ ( .D(N12566), .C(net12423), .Q(dpl_reg[0]) );
  DFFQX1 dpl_reg_reg_4__1_ ( .D(N12603), .C(net12403), .Q(dpl_reg[33]) );
  DFFQX1 dpl_reg_reg_4__0_ ( .D(N12602), .C(net12403), .Q(dpl_reg[32]) );
  DFFQX1 dpl_reg_reg_1__1_ ( .D(N12576), .C(net12418), .Q(dpl_reg[9]) );
  DFFQX1 dpl_reg_reg_1__0_ ( .D(N12575), .C(net12418), .Q(dpl_reg[8]) );
  DFFQX1 dpl_reg_reg_5__1_ ( .D(N12612), .C(net12398), .Q(dpl_reg[41]) );
  DFFQX1 dpl_reg_reg_5__0_ ( .D(N12611), .C(net12398), .Q(dpl_reg[40]) );
  DFFQX1 dpl_reg_reg_2__0_ ( .D(N12584), .C(net12413), .Q(dpl_reg[16]) );
  DFFQX1 dpl_reg_reg_6__1_ ( .D(N12621), .C(net12393), .Q(dpl_reg[49]) );
  DFFQX1 dpl_reg_reg_6__0_ ( .D(N12620), .C(net12393), .Q(dpl_reg[48]) );
  DFFQX1 multempreg_reg_0_ ( .D(N13325), .C(net12638), .Q(multempreg[0]) );
  DFFQX1 dec_accop_reg_15_ ( .D(N10578), .C(net12372), .Q(dec_accop[15]) );
  DFFQX1 dec_cop_reg_3_ ( .D(N10585), .C(net12372), .Q(dec_cop[3]) );
  DFFQX1 dec_cop_reg_4_ ( .D(N10586), .C(net12372), .Q(dec_cop[4]) );
  DFFQX1 sp_reg_reg_4_ ( .D(N12701), .C(net12372), .Q(sp[4]) );
  DFFQX1 pmw_reg_reg ( .D(N12713), .C(net12372), .Q(pmw) );
  DFFQX1 sp_reg_reg_3_ ( .D(N12700), .C(net12372), .Q(sp[3]) );
  DFFQX1 dec_cop_reg_6_ ( .D(N10588), .C(net12372), .Q(dec_cop[6]) );
  DFFQX1 bitno_reg_2_ ( .D(n2442), .C(net12383), .Q(N345) );
  DFFQX1 pc_reg_14_ ( .D(N494), .C(net12372), .Q(memaddr[14]) );
  DFFQX1 dps_reg_reg_2_ ( .D(N12695), .C(net12372), .Q(N351) );
  DFFQX1 dec_accop_reg_13_ ( .D(N10576), .C(net12372), .Q(dec_accop[13]) );
  DFFQX1 dec_accop_reg_14_ ( .D(N10577), .C(net12372), .Q(dec_accop[14]) );
  DFFQX1 dec_accop_reg_12_ ( .D(N10575), .C(net12372), .Q(dec_accop[12]) );
  DFFQX1 dec_accop_reg_2_ ( .D(N10565), .C(net12372), .Q(dec_accop[2]) );
  DFFQX1 sp_reg_reg_1_ ( .D(N12698), .C(net12372), .Q(sp[1]) );
  DFFQX1 sp_reg_reg_2_ ( .D(N12699), .C(net12372), .Q(sp[2]) );
  DFFQX1 rs_reg_reg_1_ ( .D(N12710), .C(net12372), .Q(rs[1]) );
  DFFQX1 temp2_reg_6_ ( .D(N12729), .C(net12372), .Q(temp2_comb[6]) );
  DFFQX1 sp_reg_reg_0_ ( .D(N12697), .C(net12372), .Q(sp[0]) );
  DFFQX1 temp_reg_2_ ( .D(N12716), .C(net12468), .Q(temp[2]) );
  DFFQX1 temp_reg_1_ ( .D(N12715), .C(net12468), .Q(temp[1]) );
  DFFQX1 temp_reg_0_ ( .D(N12714), .C(net12468), .Q(temp[0]) );
  DFFQX1 temp_reg_4_ ( .D(N12718), .C(net12468), .Q(temp[4]) );
  DFFQX1 temp_reg_3_ ( .D(N12717), .C(net12468), .Q(temp[3]) );
  DFFQX1 temp_reg_7_ ( .D(N12721), .C(net12468), .Q(temp[7]) );
  DFFQX1 temp_reg_6_ ( .D(N12720), .C(net12468), .Q(temp[6]) );
  DFFQX1 temp_reg_5_ ( .D(N12719), .C(net12468), .Q(temp[5]) );
  DFFQX1 ramdatao_r_reg_4_ ( .D(N11502), .C(net12372), .Q(ramdatao[4]) );
  DFFQX1 interrupt_reg ( .D(n2445), .C(net12378), .Q(interrupt) );
  DFFQX1 ramdatao_r_reg_2_ ( .D(N11500), .C(net12372), .Q(ramdatao[2]) );
  DFFQX1 pc_reg_15_ ( .D(N495), .C(net12372), .Q(pc_o[15]) );
  DFFQX1 pc_reg_4_ ( .D(N484), .C(net12372), .Q(pc_o[4]) );
  DFFQX1 pc_reg_12_ ( .D(N492), .C(net12372), .Q(memaddr[12]) );
  DFFQX1 pc_reg_7_ ( .D(N487), .C(net12372), .Q(pc_o[7]) );
  DFFQX1 pc_reg_11_ ( .D(N491), .C(net12372), .Q(pc_o[11]) );
  DFFQX1 pc_reg_13_ ( .D(N493), .C(net12372), .Q(memaddr[13]) );
  DFFQX1 pc_reg_10_ ( .D(N490), .C(net12372), .Q(memaddr[10]) );
  DFFQX1 dec_accop_reg_11_ ( .D(N10574), .C(net12372), .Q(dec_accop[11]) );
  DFFQX1 dec_accop_reg_3_ ( .D(N10566), .C(net12372), .Q(dec_accop[3]) );
  DFFQX1 dec_accop_reg_0_ ( .D(N10563), .C(net12372), .Q(dec_accop[0]) );
  DFFQX1 dps_reg_reg_3_ ( .D(n1884), .C(net12372), .Q(dps[3]) );
  DFFQX1 bitno_reg_0_ ( .D(n2443), .C(net12383), .Q(N343) );
  DFFQX1 rs_reg_reg_0_ ( .D(N12709), .C(net12372), .Q(rs[0]) );
  DFFQX1 temp2_reg_5_ ( .D(N12728), .C(net12372), .Q(temp2_comb[5]) );
  DFFQX1 bitno_reg_1_ ( .D(n2444), .C(net12383), .Q(N344) );
  DFFQX1 dec_accop_reg_4_ ( .D(N10567), .C(net12372), .Q(dec_accop[4]) );
  DFFQX1 ramdatao_r_reg_1_ ( .D(N11499), .C(net12372), .Q(ramdatao[1]) );
  DFFQX1 phase_reg_1_ ( .D(N680), .C(net12372), .Q(phase[1]) );
  DFFQX1 pc_reg_3_ ( .D(N483), .C(net12372), .Q(pc_o[3]) );
  DFFQX1 pc_reg_8_ ( .D(N488), .C(net12372), .Q(pc_o[8]) );
  DFFQX1 pc_reg_9_ ( .D(N489), .C(net12372), .Q(pc_o[9]) );
  DFFQX1 temp2_reg_4_ ( .D(N12727), .C(net12372), .Q(temp2_comb[4]) );
  DFFQX1 dps_reg_reg_1_ ( .D(N12694), .C(net12372), .Q(N350) );
  DFFQX1 dps_reg_reg_0_ ( .D(N12693), .C(net12372), .Q(N349) );
  DFFQX1 accactv_reg ( .D(N10562), .C(net12372), .Q(accactv) );
  DFFQX1 temp2_reg_1_ ( .D(N12724), .C(net12372), .Q(temp2_comb[1]) );
  DFFQX1 divtempreg_reg_6_ ( .D(N13373), .C(net12643), .Q(divtempreg[6]) );
  DFFQX1 dec_accop_reg_1_ ( .D(N10564), .C(net12372), .Q(dec_accop[1]) );
  DFFQX1 temp2_reg_3_ ( .D(N12726), .C(net12372), .Q(temp2_comb[3]) );
  DFFQX1 temp2_reg_2_ ( .D(N12725), .C(net12372), .Q(temp2_comb[2]) );
  DFFQX1 ramdatao_r_reg_3_ ( .D(N11501), .C(net12372), .Q(ramdatao[3]) );
  DFFQX1 phase_reg_0_ ( .D(N679), .C(net12372), .Q(phase[0]) );
  DFFQX1 instr_reg_1_ ( .D(N671), .C(net12378), .Q(n2457) );
  DFFQX1 instr_reg_0_ ( .D(N670), .C(net12378), .Q(N352) );
  DFFQX1 pc_reg_6_ ( .D(N486), .C(net12372), .Q(pc_o[6]) );
  DFFQX1 ac_reg_reg ( .D(N12706), .C(net12372), .Q(ac) );
  DFFQX1 divtempreg_reg_0_ ( .D(N13367), .C(net12643), .Q(divtempreg[0]) );
  DFFQX1 ramsfraddr_s_reg_6_ ( .D(N11484), .C(net12372), .Q(ramsfraddr[6]) );
  DFFQX1 dec_accop_reg_8_ ( .D(N10571), .C(net12372), .Q(dec_accop[8]) );
  DFFQX1 divtempreg_reg_1_ ( .D(N13368), .C(net12643), .Q(divtempreg[1]) );
  DFFQX1 ramsfrwe_reg ( .D(n2441), .C(net12372), .Q(ramsfrwe) );
  DFFQX1 pc_reg_2_ ( .D(N482), .C(net12372), .Q(pc_o[2]) );
  DFFQX1 instr_reg_7_ ( .D(N677), .C(net12378), .Q(n2451) );
  DFFQX1 instr_reg_4_ ( .D(N674), .C(net12378), .Q(n2454) );
  DFFQX1 pc_reg_0_ ( .D(N480), .C(net12372), .Q(memaddr[0]) );
  DFFQX1 acc_reg_reg_0_ ( .D(N12469), .C(net12372), .Q(n2459) );
  DFFQX1 instr_reg_5_ ( .D(N675), .C(net12378), .Q(n2453) );
  DFFQX1 pc_reg_1_ ( .D(N481), .C(net12372), .Q(memaddr[1]) );
  DFFQX1 instr_reg_6_ ( .D(N676), .C(net12378), .Q(n2452) );
  DFFQX1 instr_reg_3_ ( .D(N673), .C(net12378), .Q(n2455) );
  DFFQX1 instr_reg_2_ ( .D(N672), .C(net12378), .Q(n2456) );
  DFFQX2 b_reg_reg_1_ ( .D(N12478), .C(net12372), .Q(b[1]) );
  DFFQX2 b_reg_reg_0_ ( .D(N12477), .C(net12372), .Q(b[0]) );
  DFFQX2 acc_reg_reg_7_ ( .D(n2427), .C(net12372), .Q(acc[7]) );
  DFFQX1 dec_accop_reg_5_ ( .D(N10568), .C(net12372), .Q(dec_accop[5]) );
  DFFQX1 dec_accop_reg_16_ ( .D(n206), .C(net12372), .Q(dec_accop[16]) );
  DFFQX1 dec_accop_reg_6_ ( .D(N10569), .C(net12372), .Q(dec_accop[6]) );
  DFFQX1 ramsfraddr_s_reg_0_ ( .D(N11478), .C(net12372), .Q(ramsfraddr[0]) );
  DFFQX1 ramsfraddr_s_reg_1_ ( .D(N11479), .C(net12372), .Q(ramsfraddr[1]) );
  DFFQX1 ramsfraddr_s_reg_4_ ( .D(N11482), .C(net12372), .Q(ramsfraddr[4]) );
  DFFQX1 ramsfraddr_s_reg_7_ ( .D(N11485), .C(net12372), .Q(ramsfraddr[7]) );
  DFFQX1 ramsfraddr_s_reg_3_ ( .D(N11481), .C(net12372), .Q(ramsfraddr[3]) );
  DFFQX1 ramsfraddr_s_reg_5_ ( .D(N11483), .C(net12372), .Q(ramsfraddr[5]) );
  DFFQX1 divtempreg_reg_5_ ( .D(N13372), .C(net12643), .Q(divtempreg[5]) );
  DFFQX1 divtempreg_reg_4_ ( .D(N13371), .C(net12643), .Q(divtempreg[4]) );
  DFFQX1 divtempreg_reg_3_ ( .D(N13370), .C(net12643), .Q(divtempreg[3]) );
  DFFQX1 divtempreg_reg_2_ ( .D(N13369), .C(net12643), .Q(divtempreg[2]) );
  DFFQX1 ramsfraddr_s_reg_2_ ( .D(N11480), .C(net12372), .Q(ramsfraddr[2]) );
  DFFQX1 b_reg_reg_7_ ( .D(N12484), .C(net12372), .Q(b[7]) );
  DFFQX1 temp2_reg_0_ ( .D(N12723), .C(net12372), .Q(temp2_comb[0]) );
  DFFQX1 c_reg_reg ( .D(N12705), .C(net12372), .Q(c) );
  DFFQX1 acc_reg_reg_1_ ( .D(N12470), .C(net12372), .Q(n2458) );
  DFFQX1 b_reg_reg_5_ ( .D(N12482), .C(net12372), .Q(b[5]) );
  DFFQX1 b_reg_reg_6_ ( .D(N12483), .C(net12372), .Q(b[6]) );
  DFFQX1 b_reg_reg_4_ ( .D(N12481), .C(net12372), .Q(b[4]) );
  DFFQX1 b_reg_reg_3_ ( .D(N12480), .C(net12372), .Q(b[3]) );
  DFFQX1 b_reg_reg_2_ ( .D(N12479), .C(net12372), .Q(b[2]) );
  DFFQX1 acc_reg_reg_2_ ( .D(n2437), .C(net12372), .Q(acc[2]) );
  DFFQX1 acc_reg_reg_3_ ( .D(N12472), .C(net12372), .Q(acc[3]) );
  DFFQX1 acc_reg_reg_5_ ( .D(n2432), .C(net12372), .Q(acc[5]) );
  DFFQX1 acc_reg_reg_4_ ( .D(n2435), .C(net12372), .Q(acc[4]) );
  DFFQX1 ramdatao_r_reg_0_ ( .D(N11498), .C(net12372), .Q(ramdatao[0]) );
  DFFQX1 acc_reg_reg_6_ ( .D(n2433), .C(net12372), .Q(acc[6]) );
  INVX2 U3 ( .A(memdatai[0]), .Y(n1855) );
  INVX3 U4 ( .A(memdatai[3]), .Y(n1550) );
  INVX2 U5 ( .A(n2398), .Y(n2387) );
  NOR21X4 U6 ( .B(n2395), .A(n2394), .Y(n2397) );
  NAND21X2 U7 ( .B(n2274), .A(n2331), .Y(n2395) );
  NAND42X2 U8 ( .C(n2399), .D(n2398), .A(n2397), .B(n2396), .Y(n2400) );
  INVX1 U9 ( .A(n76), .Y(n70) );
  MUX2IX1 U10 ( .D0(n1854), .D1(n62), .S(n76), .Y(memaddr_comb[0]) );
  NOR32X1 U11 ( .B(n2406), .C(n2405), .A(n2404), .Y(n76) );
  NAND32X2 U12 ( .B(n2380), .C(n2394), .A(n2379), .Y(n2406) );
  NOR21X2 U13 ( .B(n2395), .A(n2378), .Y(n2379) );
  MUX2IX2 U14 ( .D0(n54), .D1(n63), .S(n491), .Y(memaddr_comb[3]) );
  INVX2 U15 ( .A(n945), .Y(n946) );
  MUX2XL U16 ( .D0(n2061), .D1(n2062), .S(n230), .Y(n1899) );
  MUX2IX2 U17 ( .D0(n92), .D1(n34), .S(n490), .Y(memaddr_comb[4]) );
  AND2X2 U18 ( .A(n78), .B(n97), .Y(n940) );
  INVX1 U19 ( .A(dec_accop[6]), .Y(n744) );
  NOR2X1 U20 ( .A(dec_accop[18]), .B(dec_accop[5]), .Y(n266) );
  NAND21X1 U21 ( .B(n266), .A(n743), .Y(n997) );
  MUX2X1 U22 ( .D0(n1321), .D1(n1320), .S(codefetch_s), .Y(n1445) );
  INVX1 U23 ( .A(n1322), .Y(n1323) );
  INVX1 U24 ( .A(n2391), .Y(n2376) );
  INVX1 U28 ( .A(acc[6]), .Y(n1921) );
  NAND21X2 U29 ( .B(n2376), .A(n1978), .Y(n2192) );
  OR3XL U30 ( .A(n714), .B(n2206), .C(n713), .Y(n2040) );
  AND2XL U31 ( .A(n2391), .B(codefetch_s), .Y(n160) );
  GEN2XL U32 ( .D(acc[3]), .E(n989), .C(ac), .B(n994), .A(n992), .Y(n985) );
  NAND21X1 U33 ( .B(n753), .A(n1567), .Y(n921) );
  AO21X1 U34 ( .B(n1131), .C(n1029), .A(n988), .Y(n1143) );
  INVX1 U35 ( .A(dec_accop[16]), .Y(n740) );
  NOR2X1 U36 ( .A(n261), .B(n998), .Y(n225) );
  OAI221X1 U37 ( .A(n636), .B(n1458), .C(n635), .D(n477), .E(n634), .Y(n638)
         );
  INVX1 U38 ( .A(n2040), .Y(n87) );
  INVX1 U39 ( .A(n2410), .Y(n63) );
  AO21X1 U40 ( .B(mempsack), .C(n2235), .A(n578), .Y(n579) );
  MUX2X1 U41 ( .D0(n2328), .D1(ramoe), .S(n552), .Y(ramoe_comb) );
  OAI222X1 U42 ( .A(n683), .B(n26), .C(n688), .D(n1550), .E(n1579), .F(n1855), 
        .Y(n2348) );
  AO2222XL U43 ( .A(n1992), .B(n2193), .C(alu_out[1]), .D(n2192), .E(n2046), 
        .F(ramdatai[1]), .G(n2048), .H(n1474), .Y(n1478) );
  AO2222XL U44 ( .A(n1994), .B(n2193), .C(alu_out[0]), .D(n2192), .E(n2046), 
        .F(ramdatai[0]), .G(n2048), .H(n1853), .Y(n1857) );
  NAND42X1 U45 ( .C(n1008), .D(n1007), .A(n178), .B(n1005), .Y(n2073) );
  NAND5XL U46 ( .A(n1910), .B(n2062), .C(n2061), .D(n1926), .E(n1770), .Y(n888) );
  INVX1 U47 ( .A(n928), .Y(n994) );
  NOR2X1 U48 ( .A(dec_accop[10]), .B(dec_accop[8]), .Y(n265) );
  NAND21X1 U49 ( .B(n2383), .A(n160), .Y(n2385) );
  XNOR2XL U50 ( .A(n1036), .B(n2459), .Y(n264) );
  XNOR2XL U51 ( .A(n1036), .B(n2458), .Y(n268) );
  MUX2BXL U52 ( .D0(n2148), .D1(n1213), .S(n1848), .Y(n1217) );
  INVX1 U53 ( .A(n929), .Y(n992) );
  NAND32X1 U54 ( .B(n920), .C(n921), .A(n763), .Y(n749) );
  NAND3X1 U55 ( .A(n7), .B(n2382), .C(n2381), .Y(n2405) );
  NAND21X1 U56 ( .B(n1948), .A(n1598), .Y(n1594) );
  NOR2X1 U57 ( .A(n2192), .B(n203), .Y(n202) );
  INVX1 U58 ( .A(n1768), .Y(n83) );
  OA222X1 U59 ( .A(n122), .B(n79), .C(n1485), .D(n2080), .E(n2082), .F(n1483), 
        .Y(n1064) );
  OA222X1 U60 ( .A(n122), .B(n1575), .C(n1421), .D(n2080), .E(n2082), .F(n1574), .Y(n249) );
  INVX1 U61 ( .A(acc[2]), .Y(n1898) );
  INVX1 U62 ( .A(acc[5]), .Y(n1777) );
  MUX2X1 U63 ( .D0(n1310), .D1(n1309), .S(instr[6]), .Y(n1311) );
  NAND43X1 U64 ( .B(n748), .C(n751), .D(n750), .A(n731), .Y(n747) );
  INVX1 U65 ( .A(n749), .Y(n731) );
  OAI221X1 U66 ( .A(n636), .B(n1809), .C(n1596), .D(n635), .E(n629), .Y(n639)
         );
  INVX1 U67 ( .A(n894), .Y(n86) );
  NAND21X1 U68 ( .B(n2206), .A(ramsfrwe), .Y(n597) );
  INVX1 U69 ( .A(memack), .Y(n2240) );
  NAND21X1 U70 ( .B(ramsfraddr[3]), .A(n2218), .Y(n2224) );
  INVX1 U71 ( .A(ramsfraddr[1]), .Y(n2211) );
  OA22X1 U72 ( .A(n1482), .B(n1499), .C(n1418), .D(n1483), .Y(n941) );
  MUX2X1 U73 ( .D0(N13337), .D1(divtempreg[0]), .S(N13343), .Y(n270) );
  INVX1 U74 ( .A(n639), .Y(n684) );
  ENOX1 U75 ( .A(n267), .B(N13343), .C(N13343), .D(acc[7]), .Y(divtemp1_0_) );
  INVX1 U76 ( .A(n1583), .Y(n1598) );
  OAI21X1 U77 ( .B(n1228), .C(n909), .A(n2387), .Y(n1914) );
  NAND6XL U78 ( .A(n1969), .B(n1972), .C(n768), .D(n1973), .E(n1967), .F(n767), 
        .Y(n1155) );
  MUX2BXL U79 ( .D0(sp[0]), .D1(n2178), .S(n235), .Y(n283) );
  NAND21X1 U80 ( .B(n2154), .A(n2314), .Y(n2156) );
  AO21X1 U81 ( .B(waitcnt[1]), .C(n2177), .A(n573), .Y(n574) );
  OAI21X1 U82 ( .B(n1143), .C(n1144), .A(n995), .Y(n262) );
  NAND21X1 U83 ( .B(n746), .A(n732), .Y(n761) );
  INVX1 U84 ( .A(n747), .Y(n732) );
  NAND21X1 U85 ( .B(n2224), .A(n1580), .Y(n1442) );
  INVX1 U86 ( .A(ramsfraddr[6]), .Y(n2205) );
  INVX1 U87 ( .A(n2409), .Y(n61) );
  INVX1 U88 ( .A(n2408), .Y(n94) );
  MUX2IX1 U89 ( .D0(n258), .D1(n259), .S(n551), .Y(ramwe_comb) );
  OA222X1 U90 ( .A(n2041), .B(n1550), .C(n2044), .D(n1555), .E(n2040), .F(
        n1791), .Y(n1079) );
  INVX1 U91 ( .A(temp2_comb[0]), .Y(n1872) );
  MUX2AXL U92 ( .D0(rn_1_), .D1(n2176), .S(n655), .Y(n1485) );
  AO2222XL U93 ( .A(n1990), .B(n2193), .C(alu_out[3]), .D(n2192), .E(n2046), 
        .F(ramdatai[3]), .G(n2048), .H(n1553), .Y(n1552) );
  NAND32X1 U94 ( .B(n2250), .C(n1581), .A(n1580), .Y(n1583) );
  AO2222XL U95 ( .A(n1989), .B(n2193), .C(alu_out[4]), .D(n2192), .E(
        ramdatai[4]), .F(n2046), .G(n2048), .H(n1542), .Y(n1540) );
  INVX1 U96 ( .A(memdatai[5]), .Y(n1956) );
  INVX1 U97 ( .A(memdatai[1]), .Y(n1476) );
  INVX1 U98 ( .A(sfrdatai[2]), .Y(n1575) );
  OA2222XL U99 ( .A(n2050), .B(n44), .C(n2051), .D(n1788), .E(n1935), .F(n2001), .G(n2000), .H(n1957), .Y(n1761) );
  OA222X1 U100 ( .A(n2041), .B(n2016), .C(n2040), .D(n2021), .E(n218), .F(
        n2018), .Y(n1503) );
  OA222X1 U101 ( .A(n2041), .B(n1573), .C(n2044), .D(n1904), .E(n2040), .F(
        n1575), .Y(n1419) );
  OA222X1 U102 ( .A(n2041), .B(n2052), .C(n2040), .D(n2078), .E(n218), .F(
        n2099), .Y(n2042) );
  MUX2BXL U103 ( .D0(n646), .D1(n645), .S(n685), .Y(n647) );
  OAI31XL U104 ( .A(n2125), .B(n958), .C(n1505), .D(mempsrd), .Y(n2389) );
  MUX2X1 U105 ( .D0(n1849), .D1(n1090), .S(n1082), .Y(n955) );
  INVX2 U106 ( .A(n553), .Y(n550) );
  OAI222X1 U107 ( .A(n1579), .B(n1476), .C(n688), .D(n1546), .E(n680), .F(n26), 
        .Y(n2349) );
  NOR2X1 U108 ( .A(n2046), .B(n1760), .Y(n4) );
  NOR2X1 U109 ( .A(n1444), .B(n5), .Y(n207) );
  INVX1 U110 ( .A(n4), .Y(n5) );
  NAND21X1 U111 ( .B(n2048), .A(n202), .Y(n1444) );
  NAND21X1 U112 ( .B(n1449), .A(n207), .Y(n1322) );
  OR3XL U113 ( .A(n944), .B(n943), .C(n1912), .Y(n6) );
  NAND2X1 U114 ( .A(n6), .B(n60), .Y(n948) );
  INVX1 U115 ( .A(n2412), .Y(n71) );
  AOI32X1 U116 ( .A(n946), .B(n241), .C(n2068), .D(n241), .E(n2067), .Y(n947)
         );
  MUX2AXL U117 ( .D0(N349), .D1(n2178), .S(n1598), .Y(n2266) );
  INVX1 U118 ( .A(n43), .Y(n541) );
  INVX1 U119 ( .A(N352), .Y(n549) );
  XOR3X1 U120 ( .A(n1063), .B(n914), .C(n2084), .Y(n7) );
  MUX2IX1 U121 ( .D0(n179), .D1(n2176), .S(n1660), .Y(n8) );
  AOI21X1 U122 ( .B(temp2_comb[6]), .C(n997), .A(n1026), .Y(n9) );
  INVX1 U123 ( .A(n540), .Y(n539) );
  INVX1 U124 ( .A(n552), .Y(n551) );
  INVX1 U125 ( .A(n2388), .Y(n2450) );
  OAI31X1 U126 ( .A(n1243), .B(n1242), .C(n1241), .D(n1240), .Y(n2391) );
  INVX1 U127 ( .A(dec_accop[8]), .Y(n741) );
  INVX1 U128 ( .A(dec_accop[5]), .Y(n926) );
  MUX2IX1 U129 ( .D0(n185), .D1(n2333), .S(n1660), .Y(n10) );
  MUX2IX1 U130 ( .D0(n186), .D1(n2178), .S(n1660), .Y(n11) );
  MUX2IX1 U131 ( .D0(n180), .D1(n2336), .S(n1660), .Y(n12) );
  MUX2IX1 U132 ( .D0(n184), .D1(n1948), .S(n1660), .Y(n13) );
  MUX2IX1 U133 ( .D0(n188), .D1(n2339), .S(n1660), .Y(n14) );
  MUX2IX1 U134 ( .D0(n189), .D1(n2342), .S(n1660), .Y(n15) );
  OA22X1 U135 ( .A(n2452), .B(n2315), .C(n1371), .D(n1333), .Y(n16) );
  INVX1 U136 ( .A(n2377), .Y(n2378) );
  MUX2IX1 U137 ( .D0(n192), .D1(n2344), .S(n1660), .Y(n17) );
  MUX2IX1 U138 ( .D0(n194), .D1(n2176), .S(n1679), .Y(n18) );
  MUX2IX1 U139 ( .D0(n193), .D1(n2178), .S(n1679), .Y(n19) );
  MUX2IX1 U140 ( .D0(n195), .D1(n2333), .S(n1679), .Y(n20) );
  MUX2IX1 U141 ( .D0(n196), .D1(n1948), .S(n1679), .Y(n21) );
  MUX2IX1 U142 ( .D0(n197), .D1(n2336), .S(n1679), .Y(n22) );
  MUX2IX1 U143 ( .D0(n198), .D1(n2339), .S(n1679), .Y(n23) );
  MUX2IX1 U144 ( .D0(n199), .D1(n2342), .S(n1679), .Y(n24) );
  OAI31XL U145 ( .A(n1999), .B(n43), .C(n2262), .D(n502), .Y(n1711) );
  INVX1 U146 ( .A(n2355), .Y(n2327) );
  INVX1 U147 ( .A(n1865), .Y(n91) );
  INVXL U148 ( .A(n690), .Y(n25) );
  INVXL U149 ( .A(n25), .Y(n26) );
  INVXL U150 ( .A(n1245), .Y(n27) );
  INVXL U151 ( .A(n1244), .Y(n28) );
  INVXL U152 ( .A(n1244), .Y(n29) );
  INVXL U153 ( .A(n1342), .Y(n30) );
  INVXL U154 ( .A(n30), .Y(n31) );
  INVXL U155 ( .A(pc_o[2]), .Y(n32) );
  INVXL U156 ( .A(n32), .Y(memaddr[2]) );
  INVXL U157 ( .A(pc_o[4]), .Y(n34) );
  INVXL U158 ( .A(n34), .Y(memaddr[4]) );
  INVXL U159 ( .A(pc_o[6]), .Y(n36) );
  INVXL U160 ( .A(n36), .Y(memaddr[6]) );
  INVXL U161 ( .A(pc_o[15]), .Y(n38) );
  INVXL U162 ( .A(n38), .Y(memaddr[15]) );
  INVXL U163 ( .A(pc_o[8]), .Y(n40) );
  INVXL U164 ( .A(n40), .Y(memaddr[8]) );
  INVXL U165 ( .A(n2266), .Y(n42) );
  INVXL U166 ( .A(n42), .Y(n43) );
  INVXL U167 ( .A(pc_o[5]), .Y(n44) );
  INVXL U168 ( .A(n44), .Y(memaddr[5]) );
  INVXL U169 ( .A(n1711), .Y(n46) );
  INVXL U170 ( .A(n46), .Y(n47) );
  INVXL U171 ( .A(pc_o[9]), .Y(n48) );
  INVXL U172 ( .A(n48), .Y(memaddr[9]) );
  INVXL U173 ( .A(pc_o[7]), .Y(n50) );
  INVXL U174 ( .A(n50), .Y(memaddr[7]) );
  INVXL U175 ( .A(pc_o[11]), .Y(n52) );
  INVXL U176 ( .A(n52), .Y(memaddr[11]) );
  INVXL U177 ( .A(pc_o[3]), .Y(n54) );
  INVXL U178 ( .A(n54), .Y(memaddr[3]) );
  OAI21BBXL U179 ( .A(n895), .B(n1926), .C(n86), .Y(n56) );
  AND2XL U180 ( .A(n508), .B(n2351), .Y(N11481) );
  AO22AX1 U181 ( .A(n57), .B(n59), .C(n644), .D(n690), .Y(n2354) );
  AOI21AXL U182 ( .B(n1579), .C(n2052), .A(n26), .Y(n57) );
  INVX2 U183 ( .A(memdatai[6]), .Y(n2016) );
  BUFXL U184 ( .A(memdatai[3]), .Y(n58) );
  BUFXL U185 ( .A(memdatai[6]), .Y(n59) );
  ENOXL U186 ( .A(n1767), .B(n1472), .C(n83), .D(ramdatai[1]), .Y(n60) );
  MUX2IX1 U187 ( .D0(n1479), .D1(n94), .S(n491), .Y(memaddr_comb[1]) );
  INVX2 U188 ( .A(sfrdatai[1]), .Y(n1472) );
  NAND31X1 U189 ( .C(n2062), .A(n893), .B(n892), .Y(n895) );
  INVX2 U190 ( .A(n2351), .Y(n693) );
  INVX3 U191 ( .A(N13353), .Y(n766) );
  INVX1 U192 ( .A(n2407), .Y(n62) );
  INVX2 U193 ( .A(memdatai[7]), .Y(n2052) );
  NAND21X1 U194 ( .B(n61), .A(n491), .Y(n157) );
  INVX1 U195 ( .A(n2327), .Y(n65) );
  INVX3 U196 ( .A(n490), .Y(n491) );
  NAND2X1 U197 ( .A(n491), .B(n2413), .Y(n159) );
  NAND21X1 U198 ( .B(n32), .A(n70), .Y(n156) );
  MUX2IX1 U199 ( .D0(n71), .D1(n44), .S(n490), .Y(memaddr_comb[5]) );
  INVX2 U200 ( .A(n867), .Y(n260) );
  NAND21X1 U201 ( .B(n2390), .A(n128), .Y(n865) );
  OR2XL U202 ( .A(n88), .B(n85), .Y(n64) );
  NAND2X1 U203 ( .A(n1449), .B(n207), .Y(n2054) );
  INVXL U204 ( .A(n2354), .Y(n694) );
  OAI22X1 U205 ( .A(n67), .B(n1546), .C(n684), .D(n690), .Y(n2352) );
  INVX1 U206 ( .A(memdatai[4]), .Y(n1546) );
  OAI22AX1 U207 ( .D(n681), .C(n26), .A(n1956), .B(n688), .Y(n1577) );
  INVX1 U208 ( .A(n2411), .Y(n92) );
  BUFXL U209 ( .A(n65), .Y(n66) );
  OAI21BBX1 U210 ( .A(n1579), .B(n2052), .C(n690), .Y(n67) );
  OAI22AX1 U211 ( .D(n2140), .C(n26), .A(n689), .B(n2052), .Y(n2355) );
  NAND21X1 U212 ( .B(n2136), .A(n2390), .Y(n864) );
  AOI22AX1 U213 ( .A(sfrdatai[2]), .B(n1066), .D(n1574), .C(n83), .Y(n230) );
  INVX1 U214 ( .A(n1456), .Y(n68) );
  INVXL U215 ( .A(n692), .Y(n69) );
  OAI221X1 U216 ( .A(n691), .B(n690), .C(n67), .D(n1956), .E(n688), .Y(n2353)
         );
  NAND2X2 U217 ( .A(sfrdatai[0]), .B(n1066), .Y(n893) );
  BUFXL U218 ( .A(n2349), .Y(n72) );
  OAI211XL U219 ( .C(n1485), .D(n2038), .A(n941), .B(n940), .Y(n73) );
  BUFXL U220 ( .A(n69), .Y(n74) );
  NAND8X2 U221 ( .A(n2349), .B(n2350), .C(n2348), .D(n695), .E(n694), .F(n693), 
        .G(sfrwe_comb_s), .H(n692), .Y(n2390) );
  INVXL U222 ( .A(n2052), .Y(n75) );
  NAND6X1 U223 ( .A(n896), .B(n899), .C(n897), .D(n1869), .E(n2137), .F(n898), 
        .Y(n2384) );
  NAND42X2 U224 ( .C(n2403), .D(n2402), .A(n2401), .B(n2400), .Y(n2404) );
  AOI22CXL U225 ( .C(n87), .D(sfrdatai[0]), .A(n1418), .B(n1460), .Y(n774) );
  NAND21X2 U226 ( .B(n2383), .A(n160), .Y(n77) );
  AND2X2 U227 ( .A(n868), .B(n260), .Y(n2383) );
  AND2X1 U228 ( .A(n96), .B(n95), .Y(n78) );
  AND2XL U229 ( .A(n511), .B(n74), .Y(N11483) );
  BUFXL U230 ( .A(n1472), .Y(n79) );
  NAND32X1 U231 ( .B(n80), .C(n81), .A(n200), .Y(n914) );
  NOR2X4 U232 ( .A(n2082), .B(n1483), .Y(n80) );
  NOR2X4 U233 ( .A(n1485), .B(n2080), .Y(n81) );
  NOR32X2 U234 ( .B(n2406), .C(n2405), .A(n2404), .Y(n2417) );
  BUFXL U235 ( .A(n491), .Y(n82) );
  OAI222X1 U236 ( .A(n686), .B(n690), .C(n688), .D(n2016), .E(n67), .F(n1550), 
        .Y(n2351) );
  OAI22CX1 U237 ( .C(n1767), .D(n1472), .A(n83), .B(ramdatai[1]), .Y(n945) );
  BUFXL U238 ( .A(n2275), .Y(n84) );
  AND2X2 U239 ( .A(n893), .B(n892), .Y(n85) );
  OAI21BBX1 U240 ( .A(n895), .B(n1926), .C(n86), .Y(n1867) );
  NAND21X1 U241 ( .B(n98), .A(n917), .Y(n1859) );
  BUFX1 U242 ( .A(n1456), .Y(n98) );
  INVXL U243 ( .A(sfrdatai[0]), .Y(n1456) );
  AND2XL U244 ( .A(n509), .B(n2328), .Y(N11486) );
  NOR3XL U245 ( .A(n891), .B(n890), .C(n1912), .Y(n88) );
  OR2X1 U246 ( .A(n85), .B(n88), .Y(n1866) );
  BUFXL U247 ( .A(n2383), .Y(n89) );
  OR2X1 U248 ( .A(n1472), .B(n2079), .Y(n200) );
  BUFXL U249 ( .A(n82), .Y(n90) );
  NAND21X1 U250 ( .B(n2390), .A(n2275), .Y(n868) );
  OAI221X1 U251 ( .A(n917), .B(n916), .C(n916), .D(n68), .E(n915), .Y(n1063)
         );
  INVX3 U252 ( .A(n2417), .Y(n490) );
  NAND21X1 U253 ( .B(n36), .A(n70), .Y(n158) );
  OAI21BBX1 U254 ( .A(n1866), .B(n1867), .C(n91), .Y(n896) );
  NOR32X4 U255 ( .B(n2387), .C(n2386), .A(n77), .Y(n2402) );
  BUFXL U256 ( .A(n2384), .Y(n93) );
  NAND2X1 U257 ( .A(n157), .B(n156), .Y(memaddr_comb[2]) );
  NAND2X1 U258 ( .A(n158), .B(n159), .Y(memaddr_comb[6]) );
  NAND32X1 U259 ( .B(n908), .C(N345), .A(n907), .Y(n2398) );
  OR2XL U260 ( .A(n2041), .B(n1476), .Y(n95) );
  OR2X1 U261 ( .A(n2044), .B(n1480), .Y(n96) );
  OR2X1 U262 ( .A(n2040), .B(n1472), .Y(n97) );
  BUFX3 U263 ( .A(n1706), .Y(n99) );
  OAI31XL U264 ( .A(n1999), .B(n2266), .C(n2259), .D(n502), .Y(n1706) );
  INVX1 U265 ( .A(n2157), .Y(n100) );
  INVX1 U266 ( .A(n1656), .Y(n101) );
  BUFX3 U267 ( .A(n1751), .Y(n102) );
  OAI31XL U268 ( .A(n540), .B(n43), .C(n1722), .D(n502), .Y(n1751) );
  BUFX3 U269 ( .A(n2315), .Y(n103) );
  INVX1 U270 ( .A(n1700), .Y(n104) );
  BUFX3 U271 ( .A(n1718), .Y(n105) );
  INVX1 U272 ( .A(n703), .Y(instr[2]) );
  BUFX3 U273 ( .A(n1715), .Y(n107) );
  BUFX3 U274 ( .A(n1704), .Y(n108) );
  INVX1 U275 ( .A(n1980), .Y(n109) );
  INVX1 U276 ( .A(n129), .Y(instr[1]) );
  NAND21X1 U277 ( .B(n2457), .A(n548), .Y(n1278) );
  INVX1 U278 ( .A(n2454), .Y(n111) );
  BUFX3 U279 ( .A(n1708), .Y(n112) );
  OAI31XL U280 ( .A(n541), .B(n1999), .C(n2262), .D(n502), .Y(n1708) );
  BUFX3 U281 ( .A(n1712), .Y(n113) );
  NAND21XL U282 ( .B(n2376), .A(n1978), .Y(n114) );
  INVX1 U283 ( .A(n1901), .Y(pc_o[10]) );
  INVX1 U284 ( .A(n1841), .Y(n116) );
  NAND21X1 U285 ( .B(n2315), .A(n2157), .Y(n1392) );
  INVX1 U286 ( .A(n873), .Y(n117) );
  BUFX3 U287 ( .A(n1756), .Y(n118) );
  OAI31XL U288 ( .A(n541), .B(n1999), .C(n2259), .D(n502), .Y(n1756) );
  BUFX3 U289 ( .A(n1709), .Y(n119) );
  BUFX3 U290 ( .A(n2455), .Y(instr[3]) );
  INVX1 U291 ( .A(n2015), .Y(pc_o[14]) );
  OR2X1 U292 ( .A(n2206), .B(n874), .Y(n122) );
  INVX1 U293 ( .A(ramsfraddr[7]), .Y(n2206) );
  BUFX3 U294 ( .A(n1719), .Y(n123) );
  OAI31XL U295 ( .A(n541), .B(n540), .C(n1722), .D(n502), .Y(n1719) );
  BUFX3 U296 ( .A(n1707), .Y(n124) );
  INVX1 U297 ( .A(n708), .Y(instr[6]) );
  NAND21X1 U298 ( .B(n2315), .A(n2452), .Y(n2146) );
  INVX1 U299 ( .A(n1827), .Y(pc_o[12]) );
  INVX1 U300 ( .A(n2163), .Y(n127) );
  GEN2XL U301 ( .D(n1260), .E(n2167), .C(n2128), .B(n127), .A(n1259), .Y(n1449) );
  INVX1 U302 ( .A(n2331), .Y(n128) );
  AND3X1 U303 ( .A(n1862), .B(n875), .C(n2332), .Y(n897) );
  NAND6X1 U304 ( .A(n951), .B(n2332), .C(n950), .D(n949), .E(n948), .F(n947), 
        .Y(n2377) );
  BUFX3 U305 ( .A(n2316), .Y(n129) );
  INVX1 U306 ( .A(n871), .Y(n130) );
  BUFX3 U307 ( .A(n1716), .Y(n131) );
  BUFX3 U308 ( .A(n1752), .Y(n132) );
  INVX1 U309 ( .A(n1807), .Y(n133) );
  BUFX3 U310 ( .A(memaddr[1]), .Y(pc_o[1]) );
  MUX2X1 U311 ( .D0(n1658), .D1(n1657), .S(pc_o[1]), .Y(n1659) );
  INVX1 U312 ( .A(n1701), .Y(n135) );
  BUFX3 U313 ( .A(n2453), .Y(instr[5]) );
  BUFX3 U314 ( .A(n653), .Y(n137) );
  INVX1 U315 ( .A(n2246), .Y(n138) );
  NAND5XL U316 ( .A(n861), .B(n2094), .C(n2097), .D(n1258), .E(n2086), .Y(n853) );
  INVX1 U317 ( .A(n1226), .Y(acc[0]) );
  INVX1 U318 ( .A(n1225), .Y(acc[1]) );
  AOI21X1 U319 ( .B(n220), .C(n42), .A(n505), .Y(n1717) );
  INVX1 U320 ( .A(n1717), .Y(n141) );
  INVX1 U321 ( .A(n1717), .Y(n142) );
  BUFX3 U322 ( .A(n1758), .Y(n143) );
  BUFX3 U323 ( .A(n1720), .Y(n144) );
  INVX1 U324 ( .A(n1588), .Y(n145) );
  MUX2X1 U325 ( .D0(n1587), .D1(n1948), .S(n2307), .Y(n1588) );
  BUFX3 U326 ( .A(memaddr[0]), .Y(pc_o[0]) );
  INVX1 U327 ( .A(n1248), .Y(n147) );
  BUFX3 U328 ( .A(n2454), .Y(instr[4]) );
  INVX1 U329 ( .A(n1955), .Y(pc_o[13]) );
  INVX1 U330 ( .A(n1361), .Y(instr[7]) );
  BUFX3 U331 ( .A(N348), .Y(n151) );
  BUFX3 U332 ( .A(N348), .Y(n152) );
  BUFX3 U333 ( .A(N348), .Y(n153) );
  OAI221X1 U334 ( .A(n1596), .B(n1595), .C(n1594), .D(n1593), .E(n1592), .Y(
        N348) );
  INVX1 U335 ( .A(accactv), .Y(n154) );
  INVX1 U336 ( .A(accactv), .Y(n155) );
  INVX1 U337 ( .A(accactv), .Y(n1190) );
  NAND21XL U338 ( .B(n597), .A(n598), .Y(n2249) );
  INVX1 U339 ( .A(n43), .Y(n391) );
  INVX1 U340 ( .A(n393), .Y(n395) );
  AND3XL U341 ( .A(n683), .B(n691), .C(n639), .Y(n641) );
  MUX2BXL U342 ( .D0(n2336), .D1(pmw), .S(n2309), .Y(n2181) );
  NAND5X1 U343 ( .A(n266), .B(n741), .C(n744), .D(n740), .E(n739), .Y(n1036)
         );
  NOR8X1 U344 ( .A(n1964), .B(n1155), .C(n1962), .D(n1963), .E(n1933), .F(
        n2073), .G(n1961), .H(n1960), .Y(n1222) );
  NAND32X1 U345 ( .B(n1392), .C(n2371), .A(n1266), .Y(n2086) );
  INVX1 U346 ( .A(n624), .Y(n686) );
  OAI221XL U347 ( .A(n636), .B(n1554), .C(n1588), .D(n635), .E(n623), .Y(n624)
         );
  NAND21XL U348 ( .B(n283), .A(n613), .Y(n595) );
  NAND21XL U349 ( .B(n265), .A(c), .Y(n742) );
  NAND21X1 U350 ( .B(n2455), .A(n1094), .Y(n2154) );
  INVXL U351 ( .A(n593), .Y(n598) );
  NAND21X1 U352 ( .B(ramsfraddr[5]), .A(n2205), .Y(n593) );
  INVXL U353 ( .A(n2352), .Y(n695) );
  INVXL U354 ( .A(n2353), .Y(n692) );
  INVX1 U355 ( .A(n687), .Y(sfrwe_comb_s) );
  AOI21BX1 U356 ( .C(n594), .B(n2000), .A(n653), .Y(n208) );
  NAND32XL U357 ( .B(n2370), .C(n653), .A(n161), .Y(n657) );
  OR2X1 U358 ( .A(n761), .B(n736), .Y(n755) );
  OR2X1 U359 ( .A(n887), .B(n591), .Y(n633) );
  NAND21X1 U360 ( .B(n591), .A(n887), .Y(n636) );
  XOR2X1 U361 ( .A(n686), .B(n684), .Y(n637) );
  INVX1 U362 ( .A(n1277), .Y(n1840) );
  INVX1 U363 ( .A(n792), .Y(n793) );
  INVX1 U364 ( .A(n638), .Y(n683) );
  NOR2X1 U365 ( .A(n2214), .B(n1442), .Y(n235) );
  OR2XL U366 ( .A(n2316), .B(n234), .Y(n1806) );
  INVX1 U367 ( .A(n1363), .Y(n2148) );
  INVX1 U368 ( .A(n497), .Y(n495) );
  OAI221X1 U369 ( .A(n636), .B(n1897), .C(n635), .D(n703), .E(n608), .Y(n681)
         );
  INVXL U370 ( .A(n1113), .Y(n607) );
  INVX1 U371 ( .A(n580), .Y(n1261) );
  INVX1 U372 ( .A(n581), .Y(n582) );
  INVX1 U373 ( .A(n2319), .Y(n2147) );
  INVXL U374 ( .A(n1371), .Y(n842) );
  NAND5XL U375 ( .A(n876), .B(n2088), .C(n1865), .D(n2097), .E(n863), .Y(n2332) );
  OR3XL U376 ( .A(n2382), .B(n857), .C(n856), .Y(n1908) );
  AO222XL U377 ( .A(n1305), .B(n804), .C(n803), .D(n2316), .E(n802), .F(n801), 
        .Y(n807) );
  INVXL U378 ( .A(n1963), .Y(n1909) );
  INVX1 U379 ( .A(n2325), .Y(n177) );
  INVX1 U380 ( .A(n1006), .Y(n178) );
  OAI221X1 U381 ( .A(n237), .B(n1810), .C(n1150), .D(n1052), .E(n1051), .Y(
        n1053) );
  OAI221X1 U382 ( .A(n237), .B(n1227), .C(n1150), .D(n1121), .E(n1120), .Y(
        n1122) );
  NAND21X1 U383 ( .B(n2454), .A(n2456), .Y(n1092) );
  INVX1 U384 ( .A(n2453), .Y(n2315) );
  MUX2XL U385 ( .D0(n1963), .D1(temp[2]), .S(n1978), .Y(N12826) );
  INVXL U386 ( .A(n2454), .Y(n1333) );
  INVX1 U387 ( .A(n2456), .Y(n703) );
  INVX1 U388 ( .A(ramdatao[3]), .Y(n1948) );
  AOI31XL U389 ( .A(n976), .B(n2457), .C(n1267), .D(n673), .Y(n674) );
  INVXL U390 ( .A(n2266), .Y(n390) );
  INVXL U391 ( .A(n393), .Y(n394) );
  NAND21XL U392 ( .B(n554), .A(n550), .Y(n2359) );
  NAND21XL U393 ( .B(n2390), .A(n160), .Y(n2394) );
  INVX1 U394 ( .A(n1999), .Y(n203) );
  NAND21XL U395 ( .B(n1459), .A(n936), .Y(n1862) );
  INVXL U396 ( .A(n999), .Y(n1150) );
  INVXL U397 ( .A(n2152), .Y(n715) );
  INVXL U398 ( .A(n2322), .Y(n2370) );
  NAND21XL U399 ( .B(n852), .A(n845), .Y(n856) );
  NAND21XL U400 ( .B(n2331), .A(n550), .Y(n2347) );
  AND2XL U401 ( .A(n510), .B(n72), .Y(N11479) );
  AND2XL U402 ( .A(n510), .B(n2348), .Y(N11478) );
  AND2XL U403 ( .A(n511), .B(n145), .Y(N12709) );
  AND2XL U404 ( .A(n1494), .B(n1846), .Y(N10581) );
  AND2XL U405 ( .A(n1847), .B(n1846), .Y(N10582) );
  NAND21XL U406 ( .B(n1045), .A(n65), .Y(n687) );
  NAND21X2 U407 ( .B(n1448), .A(n1323), .Y(n2050) );
  AO21XL U408 ( .B(n589), .C(n585), .A(n2323), .Y(n161) );
  INVXL U409 ( .A(n548), .Y(n477) );
  OAI211XL U410 ( .C(n1392), .D(n1382), .A(n1107), .B(n846), .Y(n1288) );
  AOI21XL U411 ( .B(n1364), .C(n842), .A(n1059), .Y(n209) );
  NAND21XL U412 ( .B(n2321), .A(n812), .Y(n1409) );
  NAND43XL U413 ( .B(n1234), .C(n884), .D(n902), .A(n1771), .Y(n1780) );
  NAND21XL U414 ( .B(n792), .A(n1840), .Y(n882) );
  NAND21XL U415 ( .B(n849), .A(n978), .Y(n1247) );
  INVXL U416 ( .A(n1171), .Y(n1125) );
  INVXL U417 ( .A(memdatai[2]), .Y(n1573) );
  NAND21XL U418 ( .B(n2321), .A(n715), .Y(n589) );
  NAND21XL U419 ( .B(n495), .A(n583), .Y(n844) );
  INVXL U420 ( .A(n1047), .Y(n1049) );
  INVXL U421 ( .A(n1130), .Y(n1563) );
  INVXL U422 ( .A(n1282), .Y(n2358) );
  AO21XL U423 ( .B(n800), .C(n1253), .A(n799), .Y(n803) );
  INVXL U424 ( .A(n1143), .Y(n1146) );
  AND4XL U425 ( .A(n691), .B(n680), .C(n637), .D(n638), .Y(n646) );
  NAND21XL U426 ( .B(n2321), .A(n793), .Y(n1770) );
  NAND21XL U427 ( .B(n1852), .A(n871), .Y(n1860) );
  INVXL U428 ( .A(n1116), .Y(n1118) );
  NAND21XL U429 ( .B(n495), .A(n969), .Y(n1356) );
  NAND32XL U430 ( .B(n969), .C(n1215), .A(n1214), .Y(n970) );
  NAND32XL U431 ( .B(n1316), .C(n1315), .A(n1314), .Y(n1317) );
  AO21XL U432 ( .B(n2072), .C(n2071), .A(n2070), .Y(n2075) );
  NAND21XL U433 ( .B(n1448), .A(n212), .Y(n1894) );
  OAI32XL U434 ( .A(n2269), .B(codefetch_s), .C(n2270), .D(n2145), .E(n2268), 
        .Y(N679) );
  NAND3XL U435 ( .A(n1860), .B(n1859), .C(n1858), .Y(n213) );
  AND3XL U436 ( .A(n2444), .B(n959), .C(codefetch_s), .Y(N671) );
  AND2XL U437 ( .A(n2138), .B(n58), .Y(N673) );
  AND2XL U438 ( .A(n2138), .B(n59), .Y(N676) );
  NAND21XL U439 ( .B(n2332), .A(n550), .Y(n2345) );
  AND2XL U440 ( .A(n509), .B(n84), .Y(N12469) );
  NAND21XL U441 ( .B(n1855), .A(n498), .Y(n1464) );
  AO21XL U442 ( .B(n2234), .C(n2226), .A(n558), .Y(N13230) );
  AO21XL U443 ( .B(n2222), .C(n2226), .A(n559), .Y(N13158) );
  AO21XL U444 ( .B(n2217), .C(n2226), .A(n560), .Y(N13086) );
  AO21XL U445 ( .B(n2215), .C(n2226), .A(n561), .Y(N13014) );
  OAI22AXL U446 ( .D(n1577), .C(n2359), .A(n1579), .B(n1578), .Y(N11480) );
  NAND21XL U447 ( .B(n1476), .A(n498), .Y(n1489) );
  AOI21XL U448 ( .B(n1432), .C(n1431), .A(n1430), .Y(n216) );
  AO21XL U449 ( .B(n509), .C(n1885), .A(n561), .Y(N12697) );
  AO21XL U450 ( .B(n507), .C(n1113), .A(n561), .Y(N12699) );
  AO21XL U451 ( .B(n509), .C(n1091), .A(n561), .Y(N12698) );
  AND2XL U452 ( .A(n509), .B(n2354), .Y(N11484) );
  AND2XL U453 ( .A(n508), .B(n66), .Y(N11485) );
  AND2XL U454 ( .A(n511), .B(n1834), .Y(N12701) );
  AND2XL U455 ( .A(n511), .B(n1886), .Y(N12700) );
  AND2XL U456 ( .A(n1842), .B(n1432), .Y(N10567) );
  AND2XL U457 ( .A(n507), .B(n2171), .Y(N12713) );
  AND2XL U458 ( .A(n508), .B(n1945), .Y(N12702) );
  AND2XL U459 ( .A(n510), .B(n1944), .Y(N12703) );
  AND2XL U460 ( .A(n510), .B(n2103), .Y(N12704) );
  AOI31XL U461 ( .A(n1409), .B(n1408), .C(n1407), .D(n505), .Y(N10569) );
  NAND21XL U462 ( .B(n1425), .A(n1432), .Y(n1426) );
  AOI21BBXL U463 ( .B(n1062), .C(n2323), .A(n162), .Y(n2077) );
  AOI21X1 U464 ( .B(n2357), .C(n1061), .A(n2163), .Y(n162) );
  INVXL U465 ( .A(n2124), .Y(n2144) );
  OA22XL U466 ( .A(n1393), .B(n116), .C(n2143), .D(n1391), .Y(n1394) );
  OA21XL U467 ( .B(n1840), .C(n1846), .A(n240), .Y(n1387) );
  MUX2XL U468 ( .D0(mempswr), .D1(n2374), .S(n550), .Y(mempswr_comb) );
  MUX2X1 U469 ( .D0(n942), .D1(n2068), .S(n894), .Y(n891) );
  AOI31XL U470 ( .A(n1861), .B(n2382), .C(n916), .D(n2390), .Y(n899) );
  INVXL U471 ( .A(n261), .Y(n229) );
  INVXL U472 ( .A(n1117), .Y(n226) );
  XOR2XL U473 ( .A(n231), .B(n300), .Y(n1209) );
  AO21X1 U474 ( .B(n1143), .C(n1144), .A(n1145), .Y(n995) );
  OA21X1 U475 ( .B(n1131), .C(n1029), .A(n1130), .Y(n988) );
  AOI31XL U476 ( .A(n201), .B(n1237), .C(n1299), .D(n1222), .Y(n1242) );
  OA2222XL U477 ( .A(n1872), .B(n2054), .C(n2053), .D(n1855), .E(n2051), .F(
        n1871), .G(n1854), .H(n2050), .Y(n1856) );
  NAND32X1 U478 ( .B(n1511), .C(n2207), .A(n1439), .Y(n757) );
  INVXL U479 ( .A(n1031), .Y(n1131) );
  NAND32X1 U480 ( .B(n1180), .C(n1564), .A(n1179), .Y(n1508) );
  NAND21X1 U481 ( .B(n1142), .A(n1003), .Y(n1180) );
  NAND21X1 U482 ( .B(n755), .A(n754), .Y(n918) );
  XNOR3XL U483 ( .A(n268), .B(n986), .C(n987), .Y(n932) );
  NAND21XL U484 ( .B(n548), .A(n2316), .Y(n1342) );
  INVXL U485 ( .A(n1367), .Y(n1257) );
  AND4XL U486 ( .A(n1379), .B(n2321), .C(n1220), .D(n1277), .Y(n586) );
  MUX2X1 U487 ( .D0(n163), .D1(n2333), .S(n655), .Y(n1421) );
  MUX2IX1 U488 ( .D0(n426), .D1(n421), .S(N356), .Y(n163) );
  INVXL U489 ( .A(n1379), .Y(n1406) );
  MUX2X1 U490 ( .D0(n164), .D1(n2178), .S(n655), .Y(n1852) );
  MUX2IX1 U491 ( .D0(n406), .D1(n401), .S(N356), .Y(n164) );
  MUX2X1 U492 ( .D0(n165), .D1(n1948), .S(n655), .Y(n1792) );
  MUX2IX1 U493 ( .D0(n436), .D1(n431), .S(N356), .Y(n165) );
  AO21XL U494 ( .B(n1329), .C(n877), .A(n1432), .Y(n804) );
  NAND21XL U495 ( .B(n1365), .A(n1257), .Y(n2155) );
  MUX2X1 U496 ( .D0(n166), .D1(n2336), .S(n655), .Y(n1820) );
  MUX2IX1 U497 ( .D0(n446), .D1(n441), .S(N356), .Y(n166) );
  MUX2X1 U498 ( .D0(n167), .D1(n2339), .S(n655), .Y(n1935) );
  MUX2IX1 U499 ( .D0(n456), .D1(n451), .S(N356), .Y(n167) );
  MUX2X1 U500 ( .D0(n168), .D1(n2342), .S(n655), .Y(n2002) );
  MUX2IX1 U501 ( .D0(n466), .D1(n461), .S(N356), .Y(n168) );
  AO21XL U502 ( .B(N12770), .C(n283), .A(n614), .Y(n615) );
  AO21XL U503 ( .B(n284), .C(n595), .A(n609), .Y(n596) );
  XOR2XL U504 ( .A(n649), .B(n289), .Y(n643) );
  NAND21XL U505 ( .B(n759), .A(n1169), .Y(n1174) );
  NAND21XL U506 ( .B(n2118), .A(n1316), .Y(n2000) );
  INVXL U507 ( .A(n1032), .Y(n1145) );
  MUX2X1 U508 ( .D0(n169), .D1(n2344), .S(n655), .Y(n2081) );
  MUX2IX1 U509 ( .D0(n476), .D1(n471), .S(N356), .Y(n169) );
  NAND21XL U510 ( .B(n1379), .A(n1266), .Y(n2362) );
  INVXL U511 ( .A(n1327), .Y(n800) );
  NAND32XL U512 ( .B(n2211), .C(n2212), .A(n2209), .Y(n1946) );
  NAND21XL U513 ( .B(n1101), .A(n2148), .Y(n660) );
  NAND32XL U514 ( .B(n1511), .C(n2250), .A(n2207), .Y(n2271) );
  NAND21XL U515 ( .B(n1371), .A(n2148), .Y(n843) );
  NAND32XL U516 ( .B(n100), .C(n1363), .A(n1362), .Y(n670) );
  NAND32XL U517 ( .B(n849), .C(n1363), .A(n976), .Y(n885) );
  NAND21XL U518 ( .B(n1363), .A(n2147), .Y(n1269) );
  NAND21XL U519 ( .B(n1150), .A(n745), .Y(n1972) );
  MUX2X1 U520 ( .D0(n641), .D1(n640), .S(n680), .Y(n642) );
  OA21XL U521 ( .B(n1132), .C(n1031), .A(n1030), .Y(n1033) );
  AO21XL U522 ( .B(n1132), .C(n1031), .A(n1563), .Y(n1030) );
  MUX4XL U523 ( .D0(n415), .D1(n413), .D2(n414), .D3(n412), .S0(N355), .S1(
        N354), .Y(n416) );
  MUX4XL U524 ( .D0(n410), .D1(n408), .D2(n409), .D3(n407), .S0(N355), .S1(
        N354), .Y(n411) );
  NAND32XL U525 ( .B(n2313), .C(n2319), .A(n111), .Y(n809) );
  INVXL U526 ( .A(n1204), .Y(n1196) );
  NAND21XL U527 ( .B(n1835), .A(n1102), .Y(n666) );
  INVX1 U528 ( .A(n2146), .Y(n1100) );
  AO21XL U529 ( .B(n825), .C(n1266), .A(n794), .Y(n667) );
  NAND21XL U530 ( .B(n2316), .A(n548), .Y(n849) );
  NAND32XL U531 ( .B(n2382), .C(n856), .A(n857), .Y(n1865) );
  NAND32XL U532 ( .B(n1333), .C(n2152), .A(n1406), .Y(n2356) );
  NAND21XL U533 ( .B(n848), .A(n2314), .Y(n1382) );
  INVXL U534 ( .A(n1308), .Y(n1309) );
  INVXL U535 ( .A(n1029), .Y(n1132) );
  NAND21XL U536 ( .B(n1379), .A(n1372), .Y(n1061) );
  NAND21XL U537 ( .B(n708), .A(n1843), .Y(n1220) );
  NAND32XL U538 ( .B(n2316), .C(n1392), .A(n2314), .Y(n2161) );
  OAI222XL U539 ( .A(n672), .B(n496), .C(n671), .D(n2163), .E(n2118), .F(n2361), .Y(n2311) );
  OA21XL U540 ( .B(n663), .C(n1327), .A(n1291), .Y(n669) );
  NAND21XL U541 ( .B(n871), .A(n872), .Y(n874) );
  INVXL U542 ( .A(n1026), .Y(n1027) );
  NOR2XL U543 ( .A(n1367), .B(n849), .Y(n240) );
  OAI31XL U544 ( .A(n1255), .B(n496), .C(n31), .D(n1600), .Y(n2193) );
  NAND21XL U545 ( .B(n2315), .A(n548), .Y(n877) );
  NAND32XL U546 ( .B(n1302), .C(n31), .A(n1101), .Y(n1378) );
  NAND32XL U547 ( .B(n31), .C(n1092), .A(n1101), .Y(n1265) );
  OAI21BBX1 U548 ( .A(n702), .B(n701), .C(n1356), .Y(n772) );
  NAND21XL U549 ( .B(n1371), .A(n715), .Y(n1332) );
  AND3XL U550 ( .A(n1432), .B(n1257), .C(n477), .Y(n817) );
  OA21XL U551 ( .B(n1361), .C(n1333), .A(n1367), .Y(n824) );
  NAND21XL U552 ( .B(n2313), .A(n1364), .Y(n661) );
  INVXL U553 ( .A(n497), .Y(n496) );
  OA22XL U554 ( .A(n1417), .B(n1273), .C(n1272), .D(n1835), .Y(n1274) );
  AND3XL U555 ( .A(n1415), .B(n2318), .C(n1385), .Y(n1273) );
  OR2XL U556 ( .A(n2246), .B(n1258), .Y(n2085) );
  NAND32XL U557 ( .B(n2152), .C(n2318), .A(n1333), .Y(n1233) );
  NAND21XL U558 ( .B(n1278), .A(n1257), .Y(n1292) );
  NAND32XL U559 ( .B(n1432), .C(n1338), .A(n1385), .Y(n1263) );
  NAND21XL U560 ( .B(n854), .A(n1379), .Y(n1105) );
  NAND21XL U561 ( .B(n1261), .A(n973), .Y(n1287) );
  NAND32XL U562 ( .B(n1342), .C(n1835), .A(n2148), .Y(n968) );
  AND3XL U563 ( .A(n2155), .B(n1363), .C(n1237), .Y(n1238) );
  AO21XL U564 ( .B(n1268), .C(n1267), .A(n1342), .Y(n1271) );
  OAI221XL U565 ( .A(n709), .B(n111), .C(n1843), .D(n708), .E(n2318), .Y(n710)
         );
  AND3XL U566 ( .A(n1085), .B(n2125), .C(n2124), .Y(n2131) );
  AOI22AXL U567 ( .A(n1085), .B(n2389), .D(n170), .C(n2365), .Y(n1087) );
  AOI21X1 U568 ( .B(codefetch_s), .C(n2113), .A(n1085), .Y(n170) );
  XNOR3X1 U569 ( .A(n2084), .B(n2083), .C(n171), .Y(n2087) );
  OAI222XL U570 ( .A(n117), .B(n2099), .C(n2081), .D(n130), .E(n122), .F(n2078), .Y(n171) );
  AOI22XL U571 ( .A(n91), .B(n1934), .C(n2074), .D(n1933), .Y(n244) );
  XNOR3X1 U572 ( .A(n2084), .B(n1936), .C(n1797), .Y(n1801) );
  NAND43X1 U573 ( .B(n1803), .C(n172), .D(n173), .A(n1802), .Y(n1804) );
  OAI222XL U574 ( .A(n2097), .B(n1789), .C(n2093), .D(n1788), .E(n2091), .F(
        n1787), .Y(n172) );
  OAI222XL U575 ( .A(n2094), .B(n1790), .C(n2085), .D(n1955), .E(n44), .F(
        n2086), .Y(n173) );
  XNOR3X1 U576 ( .A(n2084), .B(n1823), .C(n1822), .Y(n1826) );
  OA21XL U577 ( .B(n1772), .C(n1771), .A(n1770), .Y(n1774) );
  NAND42X1 U578 ( .C(n1831), .D(n174), .A(n1830), .B(n1829), .Y(n1832) );
  OAI222XL U579 ( .A(n2097), .B(n1819), .C(n2093), .D(n1818), .E(n2091), .F(
        n1817), .Y(n174) );
  OAI221XL U580 ( .A(n1909), .B(n1908), .C(n2088), .D(n1907), .E(n1906), .Y(
        n1917) );
  AO21XL U581 ( .B(n1864), .C(n2382), .A(n1863), .Y(n1876) );
  NOR3XL U582 ( .A(n1918), .B(n1917), .C(n176), .Y(n175) );
  OAI222XL U583 ( .A(n2091), .B(n1916), .C(n230), .D(n1915), .E(n1929), .F(
        n1914), .Y(n176) );
  OAI211XL U584 ( .C(n1421), .D(n2038), .A(n1420), .B(n1419), .Y(n1422) );
  NAND32XL U585 ( .B(n540), .C(n1710), .A(n2266), .Y(n1709) );
  NAND21XL U586 ( .B(n43), .A(n204), .Y(n1718) );
  NAND21XL U587 ( .B(n2266), .A(n214), .Y(n1707) );
  NAND21XL U588 ( .B(n2266), .A(n500), .Y(n2260) );
  AO22AXL U589 ( .A(n2307), .B(n516), .C(n2308), .D(n2285), .Y(N12711) );
  AO21XL U590 ( .B(n205), .C(n43), .A(n557), .Y(N12529) );
  OAI21BBXL U591 ( .A(n220), .B(n2266), .C(n507), .Y(n1715) );
  OAI211XL U592 ( .C(n292), .D(n493), .A(n2143), .B(n2389), .Y(n2123) );
  OA21XL U593 ( .B(n1854), .C(n2031), .A(n138), .Y(n1463) );
  OA22XL U594 ( .A(n1458), .B(n2030), .C(n1872), .D(n2032), .Y(n1462) );
  NAND32XL U595 ( .B(n2125), .C(n506), .A(n2389), .Y(n963) );
  OA21XL U596 ( .B(n1479), .C(n2031), .A(n138), .Y(n1488) );
  NAND21XL U597 ( .B(n1835), .A(n500), .Y(n1836) );
  NAND21XL U598 ( .B(n2327), .A(n2326), .Y(n2164) );
  AND2XL U599 ( .A(n206), .B(n1505), .Y(N371) );
  AND2XL U600 ( .A(n217), .B(n1505), .Y(N372) );
  NAND32XL U601 ( .B(n2241), .C(n2240), .A(n2239), .Y(n2424) );
  INVXL U602 ( .A(n1960), .Y(n1954) );
  INVXL U603 ( .A(n1961), .Y(n1824) );
  INVXL U604 ( .A(n1798), .Y(n1799) );
  INVXL U605 ( .A(n1933), .Y(n2013) );
  MUX2IXL U606 ( .D0(n2060), .D1(n2059), .S(n295), .Y(n254) );
  NAND21XL U607 ( .B(n1910), .A(n1228), .Y(n2064) );
  MUX2XL U608 ( .D0(n1898), .D1(n1897), .S(n295), .Y(n1913) );
  INVXL U609 ( .A(n1990), .Y(n1730) );
  INVXL U610 ( .A(n1989), .Y(n1728) );
  NAND21XL U611 ( .B(n1500), .A(n1846), .Y(n2098) );
  AOI31XL U612 ( .A(n972), .B(n971), .C(n1301), .D(n495), .Y(n974) );
  AO21XL U613 ( .B(n1328), .C(n1386), .A(n1327), .Y(n1331) );
  INVXL U614 ( .A(n2371), .Y(intcall) );
  NAND21XL U615 ( .B(n1365), .A(n1364), .Y(n1400) );
  OAI211XL U616 ( .C(n1423), .D(n2321), .A(n1407), .B(n1380), .Y(n1381) );
  AO21XL U617 ( .B(n1379), .C(n2318), .A(n1403), .Y(n1380) );
  NAND21XL U618 ( .B(n2171), .A(n2180), .Y(n2172) );
  OAI22XL U619 ( .A(n1369), .B(n2318), .C(n2318), .D(n1382), .Y(n1430) );
  NAND32XL U620 ( .B(n1365), .C(n1363), .A(n1362), .Y(n1399) );
  NAND21XL U621 ( .B(n2318), .A(n1372), .Y(n1427) );
  NAND21XL U622 ( .B(n1371), .A(n1370), .Y(n1428) );
  INVXL U623 ( .A(n2214), .Y(n2232) );
  NAND32XL U624 ( .B(n2209), .C(n2212), .A(n2211), .Y(n2210) );
  OR2X1 U625 ( .A(n2206), .B(n874), .Y(n2079) );
  OA33X1 U626 ( .A(n905), .B(n230), .C(n1929), .D(n946), .E(n905), .F(n2399), 
        .Y(n907) );
  INVXL U627 ( .A(n875), .Y(n866) );
  INVX1 U628 ( .A(ramwe), .Y(n258) );
  OAI21BBX1 U629 ( .A(n2327), .B(n2326), .C(n177), .Y(n2328) );
  OAI21AX1 U630 ( .B(sfroe_r), .C(sfrwe_r), .A(sfrack), .Y(n2239) );
  OAI221XL U631 ( .A(n1979), .B(n1777), .C(n1194), .D(n1566), .E(n1002), .Y(
        n1006) );
  NAND21XL U632 ( .B(instr[5]), .A(instr[4]), .Y(n1213) );
  INVX1 U633 ( .A(n1212), .Y(n1848) );
  OAI221XL U634 ( .A(n1226), .B(n1566), .C(n2060), .D(n1211), .E(n1210), .Y(
        n1212) );
  NAND21X1 U635 ( .B(dec_accop[9]), .A(n265), .Y(n927) );
  NAND31XL U636 ( .C(n927), .A(dec_accop[18]), .B(n926), .Y(n928) );
  INVX1 U637 ( .A(N13336), .Y(n267) );
  MUX2XL U638 ( .D0(n1960), .D1(temp[5]), .S(n1978), .Y(N12829) );
  MUX2XL U639 ( .D0(n1961), .D1(temp[4]), .S(n1978), .Y(N12828) );
  NAND32X1 U640 ( .B(ramsfraddr[0]), .C(ramsfraddr[2]), .A(n2211), .Y(n1437)
         );
  NAND21X1 U641 ( .B(n2452), .A(n2451), .Y(n2313) );
  OAI211XL U642 ( .C(instr[5]), .D(instr[7]), .A(n775), .B(n1371), .Y(n783) );
  INVXL U643 ( .A(n2457), .Y(n2316) );
  XOR3XL U644 ( .A(n1146), .B(n1145), .C(n1144), .Y(n1149) );
  NAND21X1 U645 ( .B(dps[3]), .A(dps[1]), .Y(n1585) );
  NAND21XL U646 ( .B(n2455), .A(n2457), .Y(n848) );
  AOI33XL U647 ( .A(n1370), .B(phase[0]), .C(n855), .D(n854), .E(phase[1]), 
        .F(n1362), .Y(n858) );
  NAND21XL U648 ( .B(N344), .A(N343), .Y(n2399) );
  NAND21XL U649 ( .B(N343), .A(N344), .Y(n1929) );
  MUX2X1 U650 ( .D0(pc_o[0]), .D1(n1994), .S(n1993), .Y(N12841) );
  NAND21XL U651 ( .B(n2165), .A(instr[4]), .Y(n820) );
  NAND21XL U652 ( .B(n2456), .A(n2454), .Y(n1097) );
  NAND21XL U653 ( .B(n1304), .A(n2456), .Y(n1807) );
  NAND21XL U654 ( .B(n2316), .A(n2454), .Y(n665) );
  MUX2IX1 U655 ( .D0(n377), .D1(n376), .S(n151), .Y(n179) );
  AOI22XL U656 ( .A(multemp1_0_), .B(n1522), .C(acc[4]), .D(n2294), .Y(n1041)
         );
  MUX4XL U657 ( .D0(dpl_reg[32]), .D1(dpl_reg[40]), .D2(dpl_reg[48]), .D3(
        dpl_reg[56]), .S0(n391), .S1(n395), .Y(n374) );
  AO22AXL U658 ( .A(phase[0]), .B(n675), .C(phase[1]), .D(n846), .Y(n682) );
  NAND21XL U659 ( .B(n1333), .A(n2455), .Y(n1386) );
  NAND21X1 U660 ( .B(n2209), .A(ramsfraddr[1]), .Y(n784) );
  MUX2IX1 U661 ( .D0(n383), .D1(n382), .S(n152), .Y(n180) );
  OR4X1 U662 ( .A(n935), .B(n934), .C(n933), .D(n181), .Y(n1964) );
  OAI22XL U663 ( .A(n2305), .B(n1227), .C(N13343), .D(n1979), .Y(n181) );
  OA22XL U664 ( .A(n2060), .B(n2305), .C(n1979), .D(n1227), .Y(n1151) );
  OR4X1 U665 ( .A(n1124), .B(n1123), .C(n1122), .D(n182), .Y(n1963) );
  OAI22X1 U666 ( .A(n2305), .B(n1810), .C(n1979), .D(n1226), .Y(n182) );
  OR4X1 U667 ( .A(n1055), .B(n1054), .C(n1053), .D(n183), .Y(n1962) );
  OAI22XL U668 ( .A(n2305), .B(n1777), .C(n1225), .D(n1979), .Y(n183) );
  NAND32XL U669 ( .B(ramsfraddr[2]), .C(n2211), .A(n2209), .Y(n1581) );
  NAND21XL U670 ( .B(ramsfraddr[3]), .A(ramsfraddr[4]), .Y(n2250) );
  INVXL U671 ( .A(n644), .Y(n685) );
  OA21X1 U672 ( .B(dec_cop[0]), .C(n1200), .A(accactv), .Y(n1201) );
  MUX2X1 U673 ( .D0(pc_o[1]), .D1(n1992), .S(n1993), .Y(N12842) );
  NAND21X1 U674 ( .B(n1190), .A(dec_accop[0]), .Y(n1003) );
  MUX2X1 U675 ( .D0(memaddr[2]), .D1(n1991), .S(n1993), .Y(N12843) );
  INVXL U676 ( .A(n2451), .Y(n1361) );
  NAND21XL U677 ( .B(n1204), .A(dec_cop[6]), .Y(n1188) );
  INVX1 U678 ( .A(ramdatao[0]), .Y(n2178) );
  INVX1 U679 ( .A(N350), .Y(n545) );
  MUX2IX1 U680 ( .D0(n381), .D1(n380), .S(n153), .Y(n184) );
  MUX2IX1 U681 ( .D0(n379), .D1(n378), .S(n152), .Y(n185) );
  MUX2IX1 U682 ( .D0(n375), .D1(n374), .S(n151), .Y(n186) );
  AOI21XL U683 ( .B(phase[1]), .C(n1288), .A(n888), .Y(n298) );
  INVX1 U684 ( .A(n730), .Y(n753) );
  AND3XL U685 ( .A(n849), .B(n1101), .C(n31), .Y(n829) );
  INVXL U686 ( .A(n2455), .Y(n1101) );
  AND4XL U687 ( .A(n1108), .B(n1107), .C(n2160), .D(n1106), .Y(n1109) );
  NAND21XL U688 ( .B(n703), .A(n2454), .Y(n1302) );
  AOI32XL U689 ( .A(n1257), .B(n2457), .C(n825), .D(n1338), .E(n1101), .Y(n826) );
  NAND21XL U690 ( .B(n2455), .A(n2456), .Y(n1360) );
  NAND21XL U691 ( .B(n848), .A(n2456), .Y(n1500) );
  NAND21XL U692 ( .B(n2454), .A(n2457), .Y(n1366) );
  AOI21XL U693 ( .B(n1312), .C(n1392), .A(n1311), .Y(n293) );
  OAI32XL U694 ( .A(n820), .B(n1342), .C(n1255), .D(n787), .E(n848), .Y(n788)
         );
  NAND21XL U695 ( .B(n2456), .A(n30), .Y(n2320) );
  NAND31XL U696 ( .C(n496), .A(n187), .B(n1257), .Y(n679) );
  AOI21X1 U697 ( .B(n678), .C(n805), .A(N352), .Y(n187) );
  MUX2IX1 U698 ( .D0(n385), .D1(n384), .S(n153), .Y(n188) );
  NAND21XL U699 ( .B(n2455), .A(n1841), .Y(n717) );
  AO21XL U700 ( .B(instr[3]), .C(n1105), .A(n1098), .Y(n1099) );
  OAI211XL U701 ( .C(n1295), .D(n1338), .A(n1020), .B(phase[0]), .Y(n1980) );
  OAI211XL U702 ( .C(n2457), .D(n814), .A(n813), .B(n1409), .Y(n815) );
  AND3XL U703 ( .A(n1408), .B(n813), .C(n1291), .Y(n723) );
  NAND21XL U704 ( .B(n1254), .A(n1253), .Y(n1600) );
  MUX2IX1 U705 ( .D0(n387), .D1(n386), .S(n152), .Y(n189) );
  NAND21XL U706 ( .B(n495), .A(n2455), .Y(n859) );
  NAND21XL U707 ( .B(n2454), .A(n2455), .Y(n1369) );
  NAND21XL U708 ( .B(n1267), .A(instr[3]), .Y(n697) );
  OR4XL U709 ( .A(instr[3]), .B(n492), .C(instr[1]), .D(n190), .Y(n713) );
  MUX2IXL U710 ( .D0(n707), .D1(n706), .S(n548), .Y(n190) );
  AOI31XL U711 ( .A(n1253), .B(instr[4]), .C(n477), .D(n793), .Y(n663) );
  OAI21BBXL U712 ( .A(phase[0]), .B(n1059), .C(n191), .Y(n913) );
  OAI21X1 U713 ( .B(n869), .C(n1060), .A(n127), .Y(n191) );
  NAND4XL U714 ( .A(n1493), .B(n1257), .C(n2169), .D(n239), .Y(n299) );
  NAND21XL U715 ( .B(n2316), .A(phase[0]), .Y(n1010) );
  OAI211XL U716 ( .C(n1480), .D(n2097), .A(n938), .B(n937), .Y(n939) );
  NAND32XL U717 ( .B(phase[2]), .C(phase[0]), .A(n492), .Y(n956) );
  AO21XL U718 ( .B(n1316), .C(instr[4]), .A(israccess), .Y(n2139) );
  MUX2XL U719 ( .D0(n1303), .D1(n1302), .S(instr[1]), .Y(n1307) );
  NAND21XL U720 ( .B(instr[4]), .A(interrupt), .Y(n1303) );
  AND2XL U721 ( .A(n2370), .B(instr[4]), .Y(retiinstr) );
  MUX2AXL U722 ( .D0(state[0]), .D1(n1087), .S(n1086), .Y(n1088) );
  OAI22XL U723 ( .A(n2093), .B(n1647), .C(n1557), .D(n1908), .Y(n1078) );
  AOI211XL U724 ( .C(n2114), .D(n2389), .A(n555), .B(n2145), .Y(n2115) );
  MUX2IX1 U725 ( .D0(n389), .D1(n388), .S(n153), .Y(n192) );
  MUX2IX1 U726 ( .D0(n359), .D1(n358), .S(n152), .Y(n193) );
  MUX2IX1 U727 ( .D0(n361), .D1(n360), .S(n153), .Y(n194) );
  MUX2IX1 U728 ( .D0(n363), .D1(n362), .S(n152), .Y(n195) );
  MUX2IX1 U729 ( .D0(n365), .D1(n364), .S(n153), .Y(n196) );
  MUX2IX1 U730 ( .D0(n367), .D1(n366), .S(n152), .Y(n197) );
  MUX2IX1 U731 ( .D0(n369), .D1(n368), .S(n153), .Y(n198) );
  MUX2IX1 U732 ( .D0(n371), .D1(n370), .S(n152), .Y(n199) );
  NAND2XL U733 ( .A(n2309), .B(n563), .Y(n302) );
  AND2XL U734 ( .A(n2134), .B(n497), .Y(N680) );
  MUX2XL U735 ( .D0(n1639), .D1(n1638), .S(memaddr[3]), .Y(n1646) );
  NAND21XL U736 ( .B(pc_o[3]), .A(n1602), .Y(n1631) );
  MUX2XL U737 ( .D0(n1336), .D1(n1335), .S(instr[3]), .Y(n1344) );
  OAI211XL U738 ( .C(n111), .D(n1332), .A(n1331), .B(n1330), .Y(n1345) );
  NAND32XL U739 ( .B(pc_o[3]), .C(n1650), .A(n34), .Y(n1619) );
  OA21XL U740 ( .B(instr[3]), .C(n1339), .A(n1338), .Y(n1340) );
  AND2XL U741 ( .A(cs_run), .B(phase[0]), .Y(n2127) );
  XOR2XL U742 ( .A(n1649), .B(pc_o[3]), .Y(n1642) );
  AO21XL U743 ( .B(n2128), .C(n497), .A(n2048), .Y(n1352) );
  MUX2XL U744 ( .D0(n127), .D1(n497), .S(n2165), .Y(n2166) );
  NAND21XL U745 ( .B(instr[4]), .A(n1450), .Y(n1490) );
  AO21XL U746 ( .B(memaddr[3]), .C(n1641), .A(n1640), .Y(n1644) );
  NOR43XL U747 ( .B(n2288), .C(n2287), .D(n2286), .A(b[0]), .Y(n2289) );
  INVX1 U748 ( .A(n504), .Y(n499) );
  INVX1 U749 ( .A(n505), .Y(n498) );
  INVX1 U750 ( .A(n504), .Y(n500) );
  INVX1 U751 ( .A(n503), .Y(n501) );
  INVX1 U752 ( .A(n510), .Y(n504) );
  INVX1 U753 ( .A(n510), .Y(n505) );
  INVX1 U754 ( .A(n503), .Y(n502) );
  INVX1 U755 ( .A(n508), .Y(n506) );
  INVX1 U756 ( .A(n2359), .Y(n510) );
  INVX1 U757 ( .A(n511), .Y(n503) );
  INVX1 U758 ( .A(n2359), .Y(n511) );
  INVX1 U759 ( .A(n2359), .Y(n508) );
  INVX1 U760 ( .A(n2359), .Y(n507) );
  INVX1 U761 ( .A(n2359), .Y(n509) );
  NAND21X1 U762 ( .B(n551), .A(n569), .Y(N370) );
  INVX1 U763 ( .A(n566), .Y(n554) );
  INVX1 U764 ( .A(n566), .Y(n555) );
  INVX1 U765 ( .A(n564), .Y(n561) );
  INVX1 U766 ( .A(n565), .Y(n556) );
  INVX1 U767 ( .A(n565), .Y(n557) );
  INVX1 U768 ( .A(n566), .Y(n558) );
  INVX1 U769 ( .A(n565), .Y(n559) );
  INVX1 U770 ( .A(n564), .Y(n560) );
  INVX1 U771 ( .A(n2394), .Y(n2381) );
  INVX1 U772 ( .A(n1806), .Y(n485) );
  INVX1 U773 ( .A(n1806), .Y(n488) );
  INVX1 U774 ( .A(n1806), .Y(n486) );
  INVX1 U775 ( .A(n1806), .Y(n487) );
  INVX1 U776 ( .A(n1806), .Y(n489) );
  INVX1 U777 ( .A(n1806), .Y(n484) );
  NOR2X1 U778 ( .A(n1219), .B(n1466), .Y(n201) );
  INVX1 U779 ( .A(n1760), .Y(n2053) );
  INVX1 U780 ( .A(n1833), .Y(n2435) );
  INVX1 U781 ( .A(n1887), .Y(n516) );
  INVX1 U782 ( .A(n1468), .Y(n512) );
  INVX1 U783 ( .A(n1440), .Y(n535) );
  INVX1 U784 ( .A(n1862), .Y(n1863) );
  INVX1 U785 ( .A(n1943), .Y(n2433) );
  NAND21X1 U786 ( .B(n2430), .A(n562), .Y(N12692) );
  NAND21X1 U787 ( .B(n532), .A(n562), .Y(N12690) );
  NAND21X1 U788 ( .B(n2436), .A(n568), .Y(N12691) );
  INVX1 U789 ( .A(n1440), .Y(n536) );
  INVX1 U790 ( .A(n1468), .Y(n513) );
  INVX1 U791 ( .A(n1887), .Y(n517) );
  INVX1 U792 ( .A(n1951), .Y(n521) );
  INVX1 U793 ( .A(n2023), .Y(n526) );
  INVX1 U794 ( .A(n2188), .Y(n524) );
  INVX1 U795 ( .A(n1951), .Y(n520) );
  INVX1 U796 ( .A(n2023), .Y(n527) );
  INVX1 U797 ( .A(n1535), .Y(n529) );
  INVX1 U798 ( .A(n1535), .Y(n530) );
  INVX1 U799 ( .A(n1887), .Y(n518) );
  INVX1 U800 ( .A(n1468), .Y(n514) );
  INVX1 U801 ( .A(n1582), .Y(n533) );
  INVX1 U802 ( .A(n1440), .Y(n537) );
  INVX1 U803 ( .A(n2188), .Y(n525) );
  INVX1 U804 ( .A(n1440), .Y(n538) );
  INVX1 U805 ( .A(n1468), .Y(n515) );
  INVX1 U806 ( .A(n1887), .Y(n519) );
  INVX1 U807 ( .A(n1582), .Y(n534) );
  INVX1 U808 ( .A(n1951), .Y(n522) );
  INVX1 U809 ( .A(n1535), .Y(n531) );
  INVX1 U810 ( .A(n2023), .Y(n528) );
  INVX1 U811 ( .A(n1578), .Y(n2442) );
  INVX1 U812 ( .A(n1111), .Y(n2441) );
  OA21X1 U813 ( .B(n1467), .C(n1466), .A(n511), .Y(N10572) );
  AND2X1 U814 ( .A(n510), .B(n2352), .Y(N11482) );
  INVX1 U815 ( .A(n1060), .Y(n2357) );
  INVX1 U816 ( .A(n2091), .Y(n1058) );
  INVX1 U817 ( .A(n570), .Y(n566) );
  INVX1 U818 ( .A(n571), .Y(n564) );
  INVX1 U819 ( .A(n571), .Y(n563) );
  INVX1 U820 ( .A(n571), .Y(n562) );
  INVX1 U821 ( .A(n570), .Y(n565) );
  INVX1 U822 ( .A(n570), .Y(n567) );
  INVX1 U823 ( .A(n2450), .Y(n553) );
  INVX1 U824 ( .A(n2450), .Y(n552) );
  INVX1 U825 ( .A(n2050), .Y(n1995) );
  INVX1 U826 ( .A(n539), .Y(n393) );
  INVX1 U827 ( .A(n540), .Y(n396) );
  INVX1 U828 ( .A(n2266), .Y(n392) );
  INVX1 U829 ( .A(n549), .Y(n480) );
  INVX1 U830 ( .A(n549), .Y(n481) );
  INVX1 U831 ( .A(n549), .Y(n479) );
  INVX1 U832 ( .A(n549), .Y(n478) );
  INVX1 U833 ( .A(n585), .Y(n1316) );
  INVX1 U834 ( .A(n657), .Y(n632) );
  INVX1 U835 ( .A(n633), .Y(n658) );
  INVX1 U836 ( .A(n636), .Y(n659) );
  NAND21X1 U837 ( .B(n2152), .A(n1840), .Y(n1107) );
  INVX1 U838 ( .A(n549), .Y(n482) );
  INVX1 U839 ( .A(n923), .Y(n1569) );
  NAND21X1 U840 ( .B(n922), .A(n1181), .Y(n923) );
  AO21X1 U841 ( .B(n1841), .C(n1264), .A(n1347), .Y(n1466) );
  INVX1 U842 ( .A(n543), .Y(n357) );
  INVX1 U843 ( .A(n1286), .Y(n971) );
  INVX1 U844 ( .A(n1771), .Y(n904) );
  NAND21X1 U845 ( .B(n1219), .A(n838), .Y(n1060) );
  INVX1 U846 ( .A(n2068), .Y(n2062) );
  INVX1 U847 ( .A(n2080), .Y(n871) );
  INVX1 U848 ( .A(n543), .Y(n356) );
  INVX1 U849 ( .A(n543), .Y(n355) );
  INVX1 U850 ( .A(n543), .Y(n354) );
  INVX1 U851 ( .A(n1780), .Y(n1910) );
  INVX1 U852 ( .A(n545), .Y(n353) );
  INVX1 U853 ( .A(n545), .Y(n352) );
  INVX1 U854 ( .A(n545), .Y(n350) );
  INVX1 U855 ( .A(n1264), .Y(n1425) );
  INVX1 U856 ( .A(n1431), .Y(n1417) );
  INVX1 U857 ( .A(n1409), .Y(n1219) );
  INVX1 U858 ( .A(n850), .Y(n879) );
  INVX1 U859 ( .A(n2067), .Y(n1926) );
  INVX1 U860 ( .A(n547), .Y(n349) );
  INVX1 U861 ( .A(n1484), .Y(n2028) );
  INVX1 U862 ( .A(n545), .Y(n351) );
  INVX1 U863 ( .A(n942), .Y(n2061) );
  INVX1 U864 ( .A(n1315), .Y(n1239) );
  INVX1 U865 ( .A(n964), .Y(n716) );
  OR2X1 U866 ( .A(n862), .B(n861), .Y(n2091) );
  INVX1 U867 ( .A(n1279), .Y(n1359) );
  INVX1 U868 ( .A(n844), .Y(n852) );
  INVX1 U869 ( .A(n1770), .Y(n903) );
  INVX1 U870 ( .A(n862), .Y(n876) );
  NAND21X1 U871 ( .B(n1450), .A(n1326), .Y(n1760) );
  NAND21X1 U872 ( .B(n1533), .A(n1894), .Y(n2197) );
  INVXL U873 ( .A(n2390), .Y(n1082) );
  OA21X1 U874 ( .B(n2062), .C(n1069), .A(n1926), .Y(n1070) );
  INVX1 U875 ( .A(n1245), .Y(n2057) );
  NAND21X1 U876 ( .B(n1533), .A(n498), .Y(n1245) );
  MUX2X1 U877 ( .D0(n2061), .D1(n2062), .S(n1931), .Y(n1925) );
  INVX1 U878 ( .A(n1069), .Y(n1073) );
  AO21X1 U879 ( .B(n2442), .C(n959), .A(n2445), .Y(N672) );
  AO21X1 U880 ( .B(n2443), .C(n959), .A(n2445), .Y(N670) );
  NAND21X1 U881 ( .B(n506), .A(n1533), .Y(n1244) );
  NAND21X1 U882 ( .B(n2337), .A(n500), .Y(n1833) );
  AND2X1 U883 ( .A(n2330), .B(n501), .Y(N11499) );
  NAND21X1 U884 ( .B(n2343), .A(n500), .Y(n1943) );
  INVX1 U885 ( .A(n2101), .Y(n2427) );
  INVX1 U886 ( .A(n1805), .Y(n2432) );
  NAND21X1 U887 ( .B(n541), .A(n204), .Y(n1716) );
  NAND21X1 U888 ( .B(n541), .A(n214), .Y(n1758) );
  INVX1 U889 ( .A(n1446), .Y(n1684) );
  INVX1 U890 ( .A(n1447), .Y(n1682) );
  NAND21X1 U891 ( .B(n1683), .A(n1446), .Y(n1447) );
  INVX1 U892 ( .A(n1611), .Y(n1713) );
  NAND21X1 U893 ( .B(n1999), .A(n499), .Y(n1611) );
  NOR2X1 U894 ( .A(n539), .B(n1721), .Y(n204) );
  INVX1 U895 ( .A(n1582), .Y(n532) );
  INVX1 U896 ( .A(n1919), .Y(n2437) );
  NAND21X1 U897 ( .B(n1520), .A(n499), .Y(n1527) );
  NAND21X1 U898 ( .B(n2307), .A(n500), .Y(n2285) );
  NAND21X1 U899 ( .B(n1045), .A(n498), .Y(n1111) );
  NAND21X1 U900 ( .B(n1573), .A(n498), .Y(n1578) );
  NAND21X1 U901 ( .B(n2331), .A(n500), .Y(n2102) );
  NAND21X1 U902 ( .B(n505), .A(n2144), .Y(n2269) );
  AO21X1 U903 ( .B(n205), .C(n42), .A(n557), .Y(N12538) );
  AND2X1 U904 ( .A(n1494), .B(n1840), .Y(N10565) );
  AND2X1 U905 ( .A(n1842), .B(n1841), .Y(N10589) );
  INVX1 U906 ( .A(n2188), .Y(n523) );
  INVX1 U907 ( .A(n1489), .Y(n2444) );
  INVX1 U908 ( .A(n1464), .Y(n2443) );
  NOR2X1 U909 ( .A(n539), .B(n2265), .Y(n205) );
  AND3X1 U910 ( .A(n508), .B(n1493), .C(n1492), .Y(N10577) );
  AND2X1 U911 ( .A(n508), .B(N356), .Y(N12710) );
  AND2X1 U912 ( .A(n511), .B(sfrwe_comb_s), .Y(N11489) );
  AND2X1 U913 ( .A(n1847), .B(n1840), .Y(N10583) );
  AND2X1 U914 ( .A(n1838), .B(n501), .Y(N10585) );
  NOR2X1 U915 ( .A(n2359), .B(n1429), .Y(n206) );
  INVX1 U916 ( .A(n1326), .Y(n1888) );
  INVX1 U917 ( .A(n1701), .Y(n1693) );
  INVX1 U918 ( .A(n1656), .Y(n1695) );
  INVX1 U919 ( .A(n1700), .Y(n1697) );
  NAND21X1 U920 ( .B(n1697), .A(n1656), .Y(n1662) );
  INVX1 U921 ( .A(n2295), .Y(n2296) );
  INVX1 U922 ( .A(n2097), .Y(n1056) );
  INVX1 U923 ( .A(n1564), .Y(n1568) );
  NAND21X1 U924 ( .B(n2370), .A(n2017), .Y(n1011) );
  INVX1 U925 ( .A(n1299), .Y(n1467) );
  INVX1 U926 ( .A(n572), .Y(n570) );
  INVX1 U927 ( .A(n572), .Y(n571) );
  INVX1 U928 ( .A(n1541), .Y(n2027) );
  INVX1 U929 ( .A(n571), .Y(n568) );
  INVX1 U930 ( .A(n571), .Y(n569) );
  OAI21BBX1 U931 ( .A(n1579), .B(n2052), .C(n690), .Y(n689) );
  INVX1 U932 ( .A(n997), .Y(n1028) );
  INVX1 U933 ( .A(n2054), .Y(n1996) );
  INVX1 U934 ( .A(n1155), .Y(n1459) );
  INVX1 U935 ( .A(n2271), .Y(n2307) );
  INVX1 U936 ( .A(n1594), .Y(n1589) );
  NAND43X1 U937 ( .B(n1178), .C(n1177), .D(n1176), .A(n1175), .Y(n1564) );
  INVX1 U938 ( .A(n1166), .Y(n1178) );
  AND4X1 U939 ( .A(n1174), .B(n1173), .C(n1172), .D(n1171), .Y(n1175) );
  INVX1 U940 ( .A(n1167), .Y(n1177) );
  INVX1 U941 ( .A(n757), .Y(n1142) );
  INVX1 U942 ( .A(n2249), .Y(n1580) );
  INVX1 U943 ( .A(n918), .Y(n1168) );
  INVX1 U944 ( .A(n1180), .Y(n1567) );
  NAND21X1 U945 ( .B(n492), .A(n583), .Y(n2097) );
  NAND21X1 U946 ( .B(n495), .A(n582), .Y(n2094) );
  NAND21X1 U947 ( .B(n984), .A(n1185), .Y(n1139) );
  NAND21X1 U948 ( .B(n492), .A(n1316), .Y(n2322) );
  INVX1 U949 ( .A(n1588), .Y(N355) );
  NAND21X1 U950 ( .B(n1442), .A(n2226), .Y(n2309) );
  NAND21X1 U951 ( .B(n492), .A(n582), .Y(n861) );
  NAND21X1 U952 ( .B(n792), .A(n1432), .Y(n585) );
  NAND32X1 U953 ( .B(n738), .C(n1208), .A(n1166), .Y(n999) );
  INVX1 U954 ( .A(n1172), .Y(n738) );
  OAI211X1 U955 ( .C(n493), .D(n1107), .A(n844), .B(n845), .Y(n653) );
  OAI31XL U956 ( .A(n2321), .B(n493), .C(n2152), .D(n2322), .Y(n594) );
  INVX1 U957 ( .A(n2305), .Y(n1522) );
  INVX1 U958 ( .A(n1174), .Y(n1140) );
  INVX1 U959 ( .A(n2156), .Y(n1266) );
  INVX1 U960 ( .A(n477), .Y(instr[0]) );
  INVX1 U961 ( .A(n592), .Y(n654) );
  NAND32XL U962 ( .B(n653), .C(n594), .A(n2000), .Y(n592) );
  INVXL U963 ( .A(n761), .Y(n1169) );
  INVX1 U964 ( .A(n1173), .Y(n984) );
  INVX1 U965 ( .A(n1096), .Y(n583) );
  INVX1 U966 ( .A(n595), .Y(n614) );
  INVX1 U967 ( .A(n853), .Y(n845) );
  INVX1 U968 ( .A(n2081), .Y(n2047) );
  INVX1 U969 ( .A(n1935), .Y(n1763) );
  INVX1 U970 ( .A(n620), .Y(n609) );
  INVX1 U971 ( .A(n626), .Y(n619) );
  INVX1 U972 ( .A(n612), .Y(n625) );
  INVX1 U973 ( .A(n1806), .Y(N353) );
  NAND21X1 U974 ( .B(n2267), .A(n1579), .Y(n690) );
  NAND21X1 U975 ( .B(n31), .A(n1257), .Y(n2152) );
  NAND21X1 U976 ( .B(n921), .A(n920), .Y(n1181) );
  INVX1 U977 ( .A(n1596), .Y(N356) );
  INVX1 U978 ( .A(n1185), .Y(n2299) );
  INVX1 U979 ( .A(n1211), .Y(n922) );
  INVX1 U980 ( .A(n2002), .Y(n2005) );
  INVX1 U981 ( .A(n1566), .Y(n2297) );
  INVX1 U982 ( .A(n2161), .Y(n1104) );
  NAND21X1 U983 ( .B(n977), .A(n799), .Y(n1771) );
  NAND21X1 U984 ( .B(n1392), .A(n1383), .Y(n2160) );
  NAND43X1 U985 ( .B(n1236), .C(n1235), .D(n1234), .A(n201), .Y(n1315) );
  INVX1 U986 ( .A(n1233), .Y(n1236) );
  NAND21X1 U987 ( .B(n2156), .A(n1338), .Y(n846) );
  NAND2X1 U988 ( .A(n670), .B(n589), .Y(n1286) );
  NAND21X1 U989 ( .B(n1218), .A(n1358), .Y(n1264) );
  INVX1 U990 ( .A(n1114), .Y(n1660) );
  NAND21X1 U991 ( .B(n1442), .A(n2231), .Y(n1114) );
  NAND2X1 U992 ( .A(n1860), .B(n1858), .Y(n916) );
  INVX1 U993 ( .A(n1248), .Y(n1683) );
  NAND21X1 U994 ( .B(n1247), .A(n1845), .Y(n1248) );
  INVX1 U995 ( .A(n2155), .Y(n976) );
  INVX1 U996 ( .A(n1392), .Y(n1841) );
  INVX1 U997 ( .A(n2150), .Y(n1253) );
  INVX1 U998 ( .A(n1250), .Y(n1665) );
  NAND21X1 U999 ( .B(n1683), .A(n1249), .Y(n1250) );
  INVX1 U1000 ( .A(n1280), .Y(n1493) );
  INVX1 U1001 ( .A(n1946), .Y(n2227) );
  INVX1 U1002 ( .A(n977), .Y(n1102) );
  INVX1 U1003 ( .A(n590), .Y(n635) );
  INVX1 U1004 ( .A(n2149), .Y(n812) );
  INVX1 U1005 ( .A(n630), .Y(n656) );
  INVX1 U1006 ( .A(n1382), .Y(n1294) );
  INVX1 U1007 ( .A(n1378), .Y(n1218) );
  OR2X1 U1008 ( .A(n495), .B(n209), .Y(n2080) );
  AO21X1 U1009 ( .B(n880), .C(n879), .A(n878), .Y(n2068) );
  INVX1 U1010 ( .A(n877), .Y(n880) );
  NAND21X1 U1011 ( .B(n2155), .A(n1839), .Y(n886) );
  NAND21X1 U1012 ( .B(n1358), .A(n1406), .Y(n838) );
  OR2X1 U1013 ( .A(n1460), .B(n1768), .Y(n892) );
  INVX1 U1014 ( .A(n882), .Y(n884) );
  AO21X1 U1015 ( .B(n1410), .C(n1406), .A(n969), .Y(n1059) );
  AO21X1 U1016 ( .B(n1493), .C(n662), .A(n719), .Y(n1283) );
  NAND21X1 U1017 ( .B(n2155), .A(n1260), .Y(n850) );
  NAND21X1 U1018 ( .B(n1266), .A(n1265), .Y(n1431) );
  NAND21X1 U1019 ( .B(n1482), .A(n936), .Y(n950) );
  INVX1 U1020 ( .A(n1974), .Y(n1978) );
  INVX1 U1021 ( .A(n2193), .Y(n1999) );
  INVX1 U1022 ( .A(n2321), .Y(n1846) );
  INVX1 U1023 ( .A(n2332), .Y(n2331) );
  INVX1 U1024 ( .A(n1249), .Y(n1666) );
  AND3X1 U1025 ( .A(n1301), .B(n1300), .C(n1299), .Y(n1318) );
  INVX1 U1026 ( .A(n1298), .Y(n1300) );
  INVX1 U1027 ( .A(n1358), .Y(n662) );
  INVX1 U1028 ( .A(n2356), .Y(n1234) );
  INVX1 U1029 ( .A(n1332), .Y(n1223) );
  INVX1 U1030 ( .A(n1408), .Y(n969) );
  INVX1 U1031 ( .A(n1270), .Y(n1837) );
  INVX1 U1032 ( .A(n813), .Y(n1347) );
  INVX1 U1033 ( .A(n1269), .Y(n1839) );
  NAND3X1 U1034 ( .A(n789), .B(n838), .C(n2362), .Y(n1284) );
  INVX1 U1035 ( .A(n2396), .Y(n2380) );
  INVX1 U1036 ( .A(n790), .Y(n878) );
  NAND21X1 U1037 ( .B(n2155), .A(n1837), .Y(n790) );
  INVX1 U1038 ( .A(n2311), .Y(n1045) );
  NAND21X1 U1039 ( .B(n495), .A(n1347), .Y(n1484) );
  NAND2X1 U1040 ( .A(n885), .B(n886), .Y(n2067) );
  OR2X1 U1041 ( .A(n31), .B(n1220), .Y(n1279) );
  NAND21X1 U1042 ( .B(n1020), .A(n881), .Y(n942) );
  NAND21X1 U1043 ( .B(n1392), .A(n1339), .Y(n814) );
  NAND21X1 U1044 ( .B(n2148), .A(n1223), .Y(n964) );
  INVX1 U1045 ( .A(n712), .Y(n1418) );
  NAND21X1 U1046 ( .B(n1502), .A(n1501), .Y(n712) );
  NAND2X1 U1047 ( .A(n772), .B(n2041), .Y(n2038) );
  NAND43X1 U1048 ( .B(n887), .C(n1288), .D(n903), .A(n1926), .Y(n1778) );
  INVX1 U1049 ( .A(n1265), .Y(n1492) );
  INVX1 U1050 ( .A(n1435), .Y(n1372) );
  OR2X1 U1051 ( .A(n719), .B(n718), .Y(n720) );
  NAND21X1 U1052 ( .B(n1234), .A(n1233), .Y(n1232) );
  INVX1 U1053 ( .A(n714), .Y(n2041) );
  AND2X1 U1054 ( .A(n1372), .B(n855), .Y(n778) );
  INVX1 U1055 ( .A(n1403), .Y(n1020) );
  INVX1 U1056 ( .A(n1820), .Y(n1542) );
  INVX1 U1057 ( .A(n1423), .Y(n696) );
  INVX1 U1058 ( .A(n711), .Y(n1502) );
  NAND21X1 U1059 ( .B(n770), .A(n771), .Y(n711) );
  INVX1 U1060 ( .A(n797), .Y(n798) );
  NAND21X1 U1061 ( .B(n31), .A(n976), .Y(n1214) );
  NAND21X1 U1062 ( .B(n1392), .A(n1372), .Y(n1299) );
  NAND21X1 U1063 ( .B(n853), .A(n852), .Y(n2093) );
  INVX1 U1064 ( .A(n910), .Y(n2386) );
  NAND21X1 U1065 ( .B(n1865), .A(n1816), .Y(n910) );
  INVX1 U1066 ( .A(n1317), .Y(n2119) );
  MUX2X1 U1067 ( .D0(n2068), .D1(n942), .S(n241), .Y(n944) );
  INVX1 U1068 ( .A(n2086), .Y(n2246) );
  INVX1 U1069 ( .A(n2382), .Y(n2088) );
  INVX1 U1070 ( .A(n1908), .Y(n936) );
  INVX1 U1071 ( .A(n2079), .Y(n917) );
  INVX1 U1072 ( .A(n915), .Y(n1861) );
  NAND2X1 U1073 ( .A(n2094), .B(n2086), .Y(n862) );
  INVX1 U1074 ( .A(n1792), .Y(n1553) );
  INVX1 U1075 ( .A(n724), .Y(n771) );
  INVX1 U1076 ( .A(n970), .Y(n1301) );
  INVX1 U1077 ( .A(n1262), .Y(n1450) );
  NAND21X1 U1078 ( .B(n492), .A(n1261), .Y(n1262) );
  INVX1 U1079 ( .A(n2198), .Y(n1533) );
  INVX1 U1080 ( .A(n2001), .Y(n2048) );
  INVX1 U1081 ( .A(n2368), .Y(n2365) );
  INVX1 U1082 ( .A(n1255), .Y(n2167) );
  NOR2X1 U1083 ( .A(n1533), .B(n1892), .Y(n210) );
  NOR2X1 U1084 ( .A(n1533), .B(n1891), .Y(n211) );
  INVX1 U1085 ( .A(n2000), .Y(n2046) );
  OR2X1 U1086 ( .A(n495), .B(n1292), .Y(n1326) );
  NOR2XL U1087 ( .A(n1444), .B(n1451), .Y(n212) );
  INVX1 U1088 ( .A(n1532), .Y(n1889) );
  NAND21X1 U1089 ( .B(n1888), .A(n1532), .Y(n2196) );
  INVX1 U1090 ( .A(n1893), .Y(n2195) );
  INVX1 U1091 ( .A(sfrdatai[3]), .Y(n1791) );
  AO21X1 U1092 ( .B(n2072), .C(n1816), .A(n1815), .Y(n1831) );
  GEN2XL U1093 ( .D(n1814), .E(n2068), .C(n2067), .B(n255), .A(n1813), .Y(
        n1815) );
  AOI31X1 U1094 ( .A(n2065), .B(n1812), .C(n1811), .D(n1814), .Y(n1813) );
  MUX2X1 U1095 ( .D0(n2062), .D1(n2061), .S(n255), .Y(n1811) );
  AO21X1 U1096 ( .B(n2072), .C(n1786), .A(n1785), .Y(n1803) );
  GEN2XL U1097 ( .D(n1784), .E(n2068), .C(n2067), .B(n256), .A(n1783), .Y(
        n1785) );
  AOI31X1 U1098 ( .A(n2065), .B(n1782), .C(n1781), .D(n1784), .Y(n1783) );
  MUX2X1 U1099 ( .D0(n2062), .D1(n2061), .S(n256), .Y(n1781) );
  INVX1 U1100 ( .A(n1928), .Y(n2072) );
  AO21X1 U1101 ( .B(sfrdatai[3]), .C(n1066), .A(n1065), .Y(n1069) );
  GEN2XL U1102 ( .D(n2069), .E(n2068), .C(n2067), .B(n254), .A(n2066), .Y(
        n2070) );
  AOI31X1 U1103 ( .A(n2065), .B(n2064), .C(n2063), .D(n2069), .Y(n2066) );
  MUX2X1 U1104 ( .D0(n2062), .D1(n2061), .S(n254), .Y(n2063) );
  OAI22X1 U1105 ( .A(n246), .B(n2102), .C(n2332), .D(n2101), .Y(N11505) );
  INVX1 U1106 ( .A(n1775), .Y(n1784) );
  INVX1 U1107 ( .A(n2058), .Y(n2069) );
  INVX1 U1108 ( .A(n1808), .Y(n1814) );
  AO21X1 U1109 ( .B(n1926), .C(n1899), .A(n1913), .Y(n1900) );
  XNOR2XL U1110 ( .A(n1861), .B(n213), .Y(n1864) );
  AND2X1 U1111 ( .A(n2107), .B(n563), .Y(N512) );
  OAI22XL U1112 ( .A(n2106), .B(n2390), .C(n2105), .D(n2104), .Y(n2107) );
  INVX1 U1113 ( .A(n2329), .Y(n2106) );
  OAI22X1 U1114 ( .A(n243), .B(n2102), .C(n2332), .D(n1943), .Y(N11504) );
  INVX1 U1115 ( .A(n1090), .Y(n2330) );
  INVX1 U1116 ( .A(n2278), .Y(n2337) );
  INVX1 U1117 ( .A(n1920), .Y(n1931) );
  NAND21X1 U1118 ( .B(n2144), .A(n2145), .Y(n2110) );
  AND2X1 U1119 ( .A(n511), .B(n2375), .Y(N582) );
  OAI22X1 U1120 ( .A(n2341), .B(n2102), .C(n2332), .D(n1805), .Y(N11503) );
  OAI31XL U1121 ( .A(n962), .B(n1956), .C(n506), .D(n961), .Y(N675) );
  OAI31XL U1122 ( .A(n962), .B(n2052), .C(n506), .D(n961), .Y(N677) );
  INVX1 U1123 ( .A(n961), .Y(n2445) );
  INVX1 U1124 ( .A(n2276), .Y(n2343) );
  INVX1 U1125 ( .A(n960), .Y(n2138) );
  NAND21X1 U1126 ( .B(n2268), .A(n959), .Y(n960) );
  NOR21XL U1127 ( .B(n507), .A(n2284), .Y(N12905) );
  XOR2X1 U1128 ( .A(n2283), .B(n2282), .Y(n2284) );
  XNOR3X1 U1129 ( .A(n2277), .B(n2346), .C(n2276), .Y(n2283) );
  XOR3X1 U1130 ( .A(n2281), .B(n2334), .C(n2280), .Y(n2282) );
  XOR2X1 U1131 ( .A(n2278), .B(n2340), .Y(n2281) );
  INVX1 U1132 ( .A(n962), .Y(n959) );
  AND2XL U1133 ( .A(n2138), .B(memdatai[4]), .Y(N674) );
  OAI22X1 U1134 ( .A(n2338), .B(n2102), .C(n2332), .D(n1833), .Y(N11502) );
  NAND21X1 U1135 ( .B(n2340), .A(n500), .Y(n1805) );
  AND2X1 U1136 ( .A(n510), .B(n2329), .Y(N11498) );
  OAI22X1 U1137 ( .A(n175), .B(n2102), .C(n2332), .D(n1919), .Y(N11500) );
  INVX1 U1138 ( .A(n2279), .Y(n2280) );
  NAND21X1 U1139 ( .B(n2346), .A(n499), .Y(n2101) );
  NAND21X1 U1140 ( .B(n2334), .A(n499), .Y(n1919) );
  XOR2XL U1141 ( .A(n84), .B(n73), .Y(n2277) );
  NAND21X1 U1142 ( .B(n492), .A(n1246), .Y(n1446) );
  NAND21X1 U1143 ( .B(n1714), .A(n1713), .Y(n1721) );
  INVX1 U1144 ( .A(n1443), .Y(n1679) );
  NAND21X1 U1145 ( .B(n1442), .A(n2230), .Y(n1443) );
  AO21X1 U1146 ( .B(n2234), .C(n2233), .A(n558), .Y(N13293) );
  AO21X1 U1147 ( .B(n2234), .C(n2232), .A(n558), .Y(N13284) );
  AO21X1 U1148 ( .B(n2234), .C(n2231), .A(n558), .Y(N13275) );
  AO21X1 U1149 ( .B(n2234), .C(n2230), .A(n558), .Y(N13266) );
  AO21X1 U1150 ( .B(n2228), .C(n2234), .A(n558), .Y(N13248) );
  AO21X1 U1151 ( .B(n2234), .C(n2227), .A(n558), .Y(N13239) );
  AO21X1 U1152 ( .B(n2222), .C(n2233), .A(n559), .Y(N13221) );
  AO21X1 U1153 ( .B(n2222), .C(n2232), .A(n559), .Y(N13212) );
  AO21X1 U1154 ( .B(n2222), .C(n2231), .A(n559), .Y(N13203) );
  AO21X1 U1155 ( .B(n2222), .C(n2230), .A(n559), .Y(N13194) );
  AO21X1 U1156 ( .B(n2222), .C(n2228), .A(n559), .Y(N13176) );
  AO21X1 U1157 ( .B(n2222), .C(n2227), .A(n559), .Y(N13167) );
  AO21X1 U1158 ( .B(n2217), .C(n2233), .A(n559), .Y(N13149) );
  AO21X1 U1159 ( .B(n2217), .C(n2232), .A(n560), .Y(N13140) );
  AO21X1 U1160 ( .B(n2217), .C(n2231), .A(n560), .Y(N13131) );
  AO21X1 U1161 ( .B(n2217), .C(n2230), .A(n560), .Y(N13122) );
  AO21X1 U1162 ( .B(n2217), .C(n2228), .A(n560), .Y(N13104) );
  AO21X1 U1163 ( .B(n2217), .C(n2227), .A(n560), .Y(N13095) );
  AO21X1 U1164 ( .B(n2215), .C(n2233), .A(n560), .Y(N13077) );
  AO21X1 U1165 ( .B(n2215), .C(n2232), .A(n560), .Y(N13068) );
  AO21X1 U1166 ( .B(n2215), .C(n2231), .A(n560), .Y(N13059) );
  AO21X1 U1167 ( .B(n2215), .C(n2230), .A(n561), .Y(N13050) );
  AO21X1 U1168 ( .B(n2215), .C(n2228), .A(n561), .Y(N13032) );
  AO21X1 U1169 ( .B(n2215), .C(n2227), .A(n561), .Y(N13023) );
  AND2XL U1170 ( .A(n508), .B(n73), .Y(N12470) );
  AND2X1 U1171 ( .A(n511), .B(n2279), .Y(N12472) );
  NOR2XL U1172 ( .A(n539), .B(n1710), .Y(n214) );
  OAI22X1 U1173 ( .A(n1733), .B(n1716), .C(n1732), .D(n1715), .Y(N12604) );
  OAI22X1 U1174 ( .A(n1733), .B(n1718), .C(n1732), .D(n141), .Y(N12613) );
  OAI22X1 U1175 ( .A(n1733), .B(n1720), .C(n1732), .D(n1719), .Y(N12622) );
  OAI22X1 U1176 ( .A(n1733), .B(n1752), .C(n1732), .D(n1751), .Y(N12631) );
  OAI22X1 U1177 ( .A(n1733), .B(n1758), .C(n1732), .D(n1756), .Y(N12568) );
  OAI22X1 U1178 ( .A(n1733), .B(n1707), .C(n1732), .D(n1706), .Y(N12577) );
  OAI22X1 U1179 ( .A(n1733), .B(n1709), .C(n1732), .D(n1708), .Y(N12586) );
  OAI22X1 U1180 ( .A(n1733), .B(n1712), .C(n1732), .D(n1711), .Y(N12595) );
  INVX1 U1181 ( .A(n2023), .Y(n2434) );
  INVX1 U1182 ( .A(n1582), .Y(n2438) );
  INVX1 U1183 ( .A(n1951), .Y(n2430) );
  INVX1 U1184 ( .A(n1535), .Y(n2436) );
  INVX1 U1185 ( .A(n1440), .Y(n2440) );
  INVX1 U1186 ( .A(n1468), .Y(n2428) );
  INVX1 U1187 ( .A(n1887), .Y(n2429) );
  NAND21X1 U1188 ( .B(n1714), .A(n499), .Y(n2265) );
  NAND21X1 U1189 ( .B(dps[2]), .A(n2255), .Y(n2252) );
  INVX1 U1190 ( .A(n1424), .Y(n1494) );
  NAND21X1 U1191 ( .B(n1423), .A(n498), .Y(n1424) );
  NAND21X1 U1192 ( .B(n1452), .A(n498), .Y(n2190) );
  NAND21X1 U1193 ( .B(n503), .A(n1755), .Y(n1754) );
  AO21X1 U1194 ( .B(n509), .C(n2267), .A(n557), .Y(N11491) );
  AO21X1 U1195 ( .B(n2264), .C(n2263), .A(n557), .Y(N12520) );
  INVX1 U1196 ( .A(n2262), .Y(n2264) );
  AO21X1 U1197 ( .B(n2261), .C(n2263), .A(n557), .Y(N12502) );
  INVX1 U1198 ( .A(n2259), .Y(n2261) );
  AO21X1 U1199 ( .B(n2258), .C(n2257), .A(n558), .Y(N12686) );
  INVX1 U1200 ( .A(n2256), .Y(n2257) );
  AO21X1 U1201 ( .B(n2254), .C(n2258), .A(n558), .Y(N12658) );
  INVX1 U1202 ( .A(n2252), .Y(n2254) );
  AND3X1 U1203 ( .A(n1845), .B(n30), .C(n1844), .Y(N10587) );
  AND3X1 U1204 ( .A(n1844), .B(n30), .C(n1843), .Y(N10588) );
  AND2X1 U1205 ( .A(n1842), .B(n1406), .Y(N10564) );
  AND2X1 U1206 ( .A(n1844), .B(n1839), .Y(N10586) );
  AND2X1 U1207 ( .A(n1844), .B(n1837), .Y(N10584) );
  NOR2X1 U1208 ( .A(n1525), .B(n1527), .Y(n215) );
  OAI31XL U1209 ( .A(n541), .B(n540), .C(n2265), .D(n562), .Y(N12547) );
  OAI31XL U1210 ( .A(dps[1]), .B(dps[0]), .C(n2256), .D(n564), .Y(N12665) );
  OAI31XL U1211 ( .A(dps[1]), .B(dps[0]), .C(n2252), .D(n567), .Y(N12637) );
  INVX1 U1212 ( .A(n2188), .Y(n2431) );
  INVX1 U1213 ( .A(n1404), .Y(n1842) );
  NAND21X1 U1214 ( .B(n1403), .A(n499), .Y(n1404) );
  INVX1 U1215 ( .A(n2260), .Y(n2263) );
  OAI211X1 U1216 ( .C(n2270), .D(n2269), .A(n2268), .B(n568), .Y(N685) );
  INVX1 U1217 ( .A(n1401), .Y(n1847) );
  NAND21X1 U1218 ( .B(n505), .A(n240), .Y(n1401) );
  INVX1 U1219 ( .A(n2203), .Y(n1507) );
  AND3X1 U1220 ( .A(n508), .B(n1406), .C(n1492), .Y(N10568) );
  AND2X1 U1221 ( .A(n2372), .B(n501), .Y(N585) );
  AND2X1 U1222 ( .A(n2374), .B(n501), .Y(N583) );
  AND2X1 U1223 ( .A(n2373), .B(n501), .Y(N584) );
  AND2X1 U1224 ( .A(n1530), .B(n1514), .Y(N13372) );
  AND2X1 U1225 ( .A(n1530), .B(n1516), .Y(N13370) );
  AND2X1 U1226 ( .A(n1530), .B(n1518), .Y(N13368) );
  AND2X1 U1227 ( .A(n1530), .B(n1529), .Y(N13373) );
  AND2X1 U1228 ( .A(n1530), .B(n1515), .Y(N13371) );
  AND2X1 U1229 ( .A(n1530), .B(n1517), .Y(N13369) );
  AND2X1 U1230 ( .A(n1496), .B(n501), .Y(N10578) );
  INVX1 U1231 ( .A(n1495), .Y(n1496) );
  AND2X1 U1232 ( .A(n1847), .B(n1402), .Y(N10563) );
  AND2X1 U1233 ( .A(n1405), .B(n501), .Y(N10566) );
  AND2X1 U1234 ( .A(n508), .B(n1414), .Y(N10575) );
  AO21X1 U1235 ( .B(n1413), .C(n1433), .A(n1412), .Y(n1414) );
  INVX1 U1236 ( .A(n1411), .Y(n1412) );
  NOR21XL U1237 ( .B(n509), .A(n216), .Y(N10570) );
  OAI31XL U1238 ( .A(n541), .B(n504), .C(n2262), .D(n562), .Y(N12511) );
  OAI31XL U1239 ( .A(n541), .B(n503), .C(n2259), .D(n567), .Y(N12493) );
  AOI31X1 U1240 ( .A(n2362), .B(n2361), .C(n2360), .D(n505), .Y(N690) );
  AND3X1 U1241 ( .A(n2358), .B(n2357), .C(n2356), .Y(n2360) );
  AOI31X1 U1242 ( .A(n1428), .B(n1427), .C(n1426), .D(n504), .Y(N10571) );
  AOI31X1 U1243 ( .A(n1400), .B(n1399), .C(n1398), .D(n503), .Y(N10574) );
  NAND21X1 U1244 ( .B(n1417), .A(n1413), .Y(n1398) );
  NOR2X1 U1245 ( .A(n505), .B(n1497), .Y(n217) );
  INVX1 U1246 ( .A(n1059), .Y(n1062) );
  NAND32X1 U1247 ( .B(n1661), .C(n1603), .A(n1604), .Y(n1701) );
  MUX2X1 U1248 ( .D0(n2061), .D1(n2062), .S(n1071), .Y(n1067) );
  INVX1 U1249 ( .A(n1922), .Y(n2065) );
  AOI21AX1 U1250 ( .B(n1502), .C(n2098), .A(n1501), .Y(n218) );
  AND2X1 U1251 ( .A(n1499), .B(n2098), .Y(n219) );
  INVX1 U1252 ( .A(n1932), .Y(n2074) );
  OA22X1 U1253 ( .A(n496), .B(n1378), .C(n493), .D(n1358), .Y(n1393) );
  NOR5X1 U1254 ( .A(n1390), .B(n1389), .C(n1388), .D(n1492), .E(n1387), .Y(
        n1391) );
  NAND32X1 U1255 ( .B(n1661), .C(n1604), .A(n1603), .Y(n1656) );
  NAND32X1 U1256 ( .B(n1603), .C(n1604), .A(n1687), .Y(n1700) );
  NAND21X1 U1257 ( .B(n1508), .A(n1569), .Y(n2295) );
  INVX1 U1258 ( .A(n1661), .Y(n1687) );
  NAND21X1 U1259 ( .B(n2200), .A(n1695), .Y(n1699) );
  INVX1 U1260 ( .A(n2085), .Y(n1057) );
  INVX1 U1261 ( .A(n1637), .Y(n1638) );
  INVX1 U1262 ( .A(n1620), .Y(n1621) );
  INVX1 U1263 ( .A(n1692), .Y(n1601) );
  NOR2XL U1264 ( .A(n539), .B(n1722), .Y(n220) );
  INVX1 U1265 ( .A(n1014), .Y(n2017) );
  INVX1 U1266 ( .A(n1612), .Y(n1691) );
  INVX1 U1267 ( .A(n1630), .Y(n1623) );
  OR2X1 U1268 ( .A(n2243), .B(n1351), .Y(n2031) );
  INVX1 U1269 ( .A(n2012), .Y(n1015) );
  INVX1 U1270 ( .A(n2014), .Y(n1013) );
  INVX1 U1271 ( .A(rst), .Y(n572) );
  INVX1 U1272 ( .A(n2270), .Y(n2112) );
  NAND21X1 U1273 ( .B(n492), .A(n1467), .Y(n1541) );
  NAND21X1 U1274 ( .B(n1378), .A(n1406), .Y(n1407) );
  INVX1 U1275 ( .A(n1275), .Y(n1838) );
  INVX1 U1276 ( .A(n1384), .Y(n1416) );
  NAND21X1 U1277 ( .B(n1383), .A(n1382), .Y(n1384) );
  INVX1 U1278 ( .A(n1427), .Y(n1374) );
  NAND21X1 U1279 ( .B(n1435), .A(n1413), .Y(n1411) );
  NAND21X1 U1280 ( .B(n1410), .A(n1425), .Y(n1433) );
  INVX1 U1281 ( .A(n2272), .Y(n2273) );
  NAND21X1 U1282 ( .B(n554), .A(n2271), .Y(n2272) );
  NAND21X1 U1283 ( .B(n116), .A(n1492), .Y(n1429) );
  INVX1 U1284 ( .A(n1526), .Y(n1520) );
  MUX2X1 U1285 ( .D0(memwr), .D1(n2372), .S(n2450), .Y(memwr_comb) );
  NAND3X1 U1286 ( .A(n2239), .B(n221), .C(n579), .Y(n2388) );
  OAI21X1 U1287 ( .B(n296), .C(n2240), .A(n2236), .Y(n221) );
  NAND21X1 U1288 ( .B(n1445), .A(n1323), .Y(n2051) );
  NAND21X1 U1289 ( .B(n1478), .A(n1477), .Y(n2408) );
  OA2222XL U1290 ( .A(n1480), .B(n2054), .C(n2053), .D(n1476), .E(n1475), .F(
        n2051), .G(n2050), .H(n1479), .Y(n1477) );
  INVX1 U1291 ( .A(n1485), .Y(n1474) );
  NAND21X1 U1292 ( .B(n1857), .A(n1856), .Y(n2407) );
  INVX1 U1293 ( .A(n1852), .Y(n1853) );
  OAI21BBX1 U1294 ( .A(n274), .B(n1048), .C(n222), .Y(n1130) );
  OAI21X1 U1295 ( .B(n274), .C(n1048), .A(n1047), .Y(n222) );
  OAI21BBX1 U1296 ( .A(n264), .B(n925), .C(n223), .Y(n986) );
  OAI21X1 U1297 ( .B(n264), .C(n925), .A(n924), .Y(n223) );
  OAI21BBX1 U1298 ( .A(n268), .B(n987), .C(n224), .Y(n1116) );
  OAI21X1 U1299 ( .B(n268), .C(n987), .A(n986), .Y(n224) );
  MUX2X1 U1300 ( .D0(n1232), .D1(n1235), .S(n1231), .Y(n1241) );
  OAI222XL U1301 ( .A(n1239), .B(n2118), .C(n1238), .D(n2163), .E(n2120), .F(
        n1299), .Y(n1240) );
  NAND32X1 U1302 ( .B(n744), .C(n927), .A(n926), .Y(n929) );
  OAI211X1 U1303 ( .C(n2041), .D(n1855), .A(n774), .B(n773), .Y(n2275) );
  OA222X1 U1304 ( .A(n1872), .B(n2044), .C(n1459), .D(n1499), .E(n1852), .F(
        n2038), .Y(n773) );
  NAND43X1 U1305 ( .B(n2088), .C(n1861), .D(n916), .A(n1859), .Y(n898) );
  NAND21X1 U1306 ( .B(n1540), .A(n1539), .Y(n2411) );
  OA2222XL U1307 ( .A(n1819), .B(n2054), .C(n2053), .D(n1546), .E(n2051), .F(
        n1818), .G(n2050), .H(n34), .Y(n1539) );
  NAND21X1 U1308 ( .B(n1552), .A(n1551), .Y(n2410) );
  OA2222XL U1309 ( .A(n1555), .B(n2054), .C(n2053), .D(n1550), .E(n2051), .F(
        n1647), .G(n2050), .H(n54), .Y(n1551) );
  NAND21X1 U1310 ( .B(n1325), .A(n1324), .Y(n2409) );
  AO2222XL U1311 ( .A(n1991), .B(n2193), .C(alu_out[2]), .D(n2192), .E(n2046), 
        .F(ramdatai[2]), .G(n2048), .H(n1256), .Y(n1325) );
  OA2222XL U1312 ( .A(n1904), .B(n2054), .C(n2053), .D(n1573), .E(n2051), .F(
        n1905), .G(n2050), .H(n32), .Y(n1324) );
  INVX1 U1313 ( .A(n1421), .Y(n1256) );
  XOR2X1 U1314 ( .A(n1156), .B(n228), .Y(n1000) );
  OAI21BX1 U1315 ( .C(n271), .B(n226), .A(n227), .Y(n1047) );
  OAI21X1 U1316 ( .B(n271), .C(n1117), .A(n1116), .Y(n227) );
  OAI221X1 U1317 ( .A(n1028), .B(n1872), .C(n926), .D(n927), .E(n929), .Y(n925) );
  INVX1 U1318 ( .A(n1812), .Y(n890) );
  INVX1 U1319 ( .A(n927), .Y(n743) );
  INVX1 U1320 ( .A(n1782), .Y(n943) );
  AOI21BX1 U1321 ( .C(n229), .B(n998), .A(n225), .Y(n228) );
  AND3X1 U1322 ( .A(n1971), .B(n1968), .C(n1965), .Y(n768) );
  AOI211X1 U1323 ( .C(n2294), .D(n766), .A(n765), .B(n764), .Y(n767) );
  INVX1 U1324 ( .A(n1966), .Y(n764) );
  AOI21XL U1325 ( .B(n228), .C(n1156), .A(n225), .Y(n231) );
  NAND32XL U1326 ( .B(n682), .C(n679), .A(n2052), .Y(n688) );
  AO21X1 U1327 ( .B(memdatai[2]), .C(n682), .A(n1577), .Y(n2350) );
  INVX1 U1328 ( .A(n1035), .Y(n1037) );
  OA21XL U1329 ( .B(n1028), .C(n1789), .A(n1027), .Y(n1034) );
  NAND32X1 U1330 ( .B(n1437), .C(n2205), .A(n1438), .Y(n1511) );
  INVX1 U1331 ( .A(N347), .Y(n540) );
  AO21X1 U1332 ( .B(n1170), .C(n1169), .A(n1168), .Y(n1176) );
  INVX1 U1333 ( .A(n597), .Y(n1438) );
  OAI211X1 U1334 ( .C(n1184), .D(n1183), .A(n1182), .B(n1181), .Y(n1207) );
  OAI221X1 U1335 ( .A(n1190), .B(n1162), .C(n1161), .D(n155), .E(n1202), .Y(
        n1184) );
  NAND43X1 U1336 ( .B(n1205), .C(n1192), .D(n1165), .A(n288), .Y(n1183) );
  INVX1 U1337 ( .A(n1508), .Y(n1182) );
  NAND43X1 U1338 ( .B(n751), .C(n750), .D(n749), .A(n748), .Y(n1173) );
  NAND32XL U1339 ( .B(n761), .C(n760), .A(n759), .Y(n1167) );
  NAND21XL U1340 ( .B(n747), .A(n746), .Y(n1171) );
  NAND32XL U1341 ( .B(n761), .C(n1506), .A(n288), .Y(n2305) );
  AO222XL U1342 ( .A(n654), .B(n285), .C(n208), .D(n621), .E(N12804), .F(n653), 
        .Y(n1886) );
  AO21X1 U1343 ( .B(n285), .C(n620), .A(n619), .Y(n621) );
  AO222XL U1344 ( .A(n654), .B(n286), .C(n208), .D(n627), .E(N12805), .F(n653), 
        .Y(n1834) );
  AO21X1 U1345 ( .B(n286), .C(n626), .A(n625), .Y(n627) );
  AO222XL U1346 ( .A(n654), .B(N12770), .C(n208), .D(n615), .E(N12802), .F(
        n653), .Y(n1091) );
  AO222XL U1347 ( .A(n654), .B(n284), .C(n208), .D(n596), .E(N12803), .F(n653), 
        .Y(n1113) );
  NAND31X1 U1348 ( .C(n2139), .A(n232), .B(irq), .Y(n2124) );
  NAND3X1 U1349 ( .A(n2141), .B(n2140), .C(n2311), .Y(n232) );
  MUX2XL U1350 ( .D0(n1593), .D1(n2336), .S(n2307), .Y(n1596) );
  NAND43X1 U1351 ( .B(n1165), .C(n1498), .D(n761), .A(n288), .Y(n1185) );
  NAND21XL U1352 ( .B(n749), .A(n751), .Y(n1166) );
  MUX2X1 U1353 ( .D0(n416), .D1(n411), .S(N356), .Y(rn_1_) );
  NAND21X1 U1354 ( .B(n1367), .A(n2147), .Y(n792) );
  MUX4X1 U1355 ( .D0(n405), .D1(n403), .D2(n404), .D3(n402), .S0(N355), .S1(
        N354), .Y(n406) );
  MUX4X1 U1356 ( .D0(n400), .D1(n398), .D2(n399), .D3(n397), .S0(N355), .S1(
        N354), .Y(n401) );
  GEN2XL U1357 ( .D(n290), .E(n612), .C(n649), .B(n208), .A(n611), .Y(n1945)
         );
  AO22XL U1358 ( .A(n654), .B(n290), .C(N12806), .D(n653), .Y(n611) );
  MUX4X1 U1359 ( .D0(n445), .D1(n443), .D2(n444), .D3(n442), .S0(N355), .S1(
        N354), .Y(n446) );
  MUX4X1 U1360 ( .D0(n440), .D1(n438), .D2(n439), .D3(n437), .S0(N355), .S1(
        N354), .Y(n441) );
  MUX4X1 U1361 ( .D0(n435), .D1(n433), .D2(n434), .D3(n432), .S0(N355), .S1(
        N354), .Y(n436) );
  MUX4X1 U1362 ( .D0(n430), .D1(n428), .D2(n429), .D3(n427), .S0(N355), .S1(
        N354), .Y(n431) );
  MUX4X1 U1363 ( .D0(n425), .D1(n423), .D2(n424), .D3(n422), .S0(n145), .S1(
        n133), .Y(n426) );
  MUX4X1 U1364 ( .D0(n420), .D1(n418), .D2(n419), .D3(n417), .S0(n145), .S1(
        n133), .Y(n421) );
  MUX4X1 U1365 ( .D0(n455), .D1(n453), .D2(n454), .D3(n452), .S0(n145), .S1(
        n133), .Y(n456) );
  MUX4X1 U1366 ( .D0(n450), .D1(n448), .D2(n449), .D3(n447), .S0(n145), .S1(
        n133), .Y(n451) );
  NAND21X1 U1367 ( .B(n1361), .A(n1100), .Y(n1280) );
  OAI21BBXL U1368 ( .A(N12801), .B(n137), .C(n233), .Y(n1885) );
  MUX2IXL U1369 ( .D0(n208), .D1(n654), .S(n283), .Y(n233) );
  AOI21XL U1370 ( .B(n1280), .C(n703), .A(n848), .Y(n234) );
  NAND21XL U1371 ( .B(n749), .A(n750), .Y(n1172) );
  NAND32X1 U1372 ( .B(n657), .C(n590), .A(n606), .Y(n591) );
  NAND21X1 U1373 ( .B(n2154), .A(n847), .Y(n1096) );
  NAND21X1 U1374 ( .B(n284), .A(n614), .Y(n620) );
  NAND21X1 U1375 ( .B(n285), .A(n609), .Y(n626) );
  NAND21X1 U1376 ( .B(n286), .A(n619), .Y(n612) );
  MUX4X1 U1377 ( .D0(n470), .D1(n468), .D2(n469), .D3(n467), .S0(N355), .S1(
        N354), .Y(n471) );
  MUX4X1 U1378 ( .D0(n475), .D1(n473), .D2(n474), .D3(n472), .S0(N355), .S1(
        N354), .Y(n476) );
  AO222XL U1379 ( .A(n654), .B(N12776), .C(N12808), .D(n653), .E(n208), .F(
        n652), .Y(n2103) );
  XOR2X1 U1380 ( .A(n651), .B(n650), .Y(n652) );
  NAND21X1 U1381 ( .B(n289), .A(n649), .Y(n650) );
  OA222X1 U1382 ( .A(n2218), .B(n633), .C(n632), .D(n628), .E(n1820), .F(n630), 
        .Y(n629) );
  INVX1 U1383 ( .A(n1834), .Y(n628) );
  OA222X1 U1384 ( .A(n633), .B(n2209), .C(n632), .D(n631), .E(n1852), .F(n630), 
        .Y(n634) );
  INVX1 U1385 ( .A(n1885), .Y(n631) );
  OA222X1 U1386 ( .A(n633), .B(n2220), .C(n632), .D(n622), .E(n1792), .F(n630), 
        .Y(n623) );
  INVX1 U1387 ( .A(n1886), .Y(n622) );
  INVX1 U1388 ( .A(n618), .Y(n680) );
  OAI221X1 U1389 ( .A(n636), .B(n1481), .C(n635), .D(n129), .E(n617), .Y(n618)
         );
  OA222X1 U1390 ( .A(n633), .B(n2211), .C(n632), .D(n616), .E(n1485), .F(n630), 
        .Y(n617) );
  INVX1 U1391 ( .A(n1091), .Y(n616) );
  OA222X1 U1392 ( .A(n633), .B(n2212), .C(n632), .D(n607), .E(n1421), .F(n630), 
        .Y(n608) );
  INVX1 U1393 ( .A(n2399), .Y(n1786) );
  INVX1 U1394 ( .A(n1929), .Y(n1769) );
  INVX1 U1395 ( .A(n1092), .Y(n2314) );
  INVX1 U1396 ( .A(n2313), .Y(n2157) );
  XOR3XL U1397 ( .A(n264), .B(n924), .C(n925), .Y(n745) );
  NAND32XL U1398 ( .B(n1190), .C(n1565), .A(n1169), .Y(n758) );
  INVX1 U1399 ( .A(n1278), .Y(n1094) );
  NAND21X1 U1400 ( .B(n236), .A(n1179), .Y(n1208) );
  AO21X1 U1401 ( .B(n1196), .C(n1194), .A(n1193), .Y(n1199) );
  AO21X1 U1402 ( .B(n1140), .C(n2096), .A(n1139), .Y(n982) );
  INVX1 U1403 ( .A(n786), .Y(n2165) );
  INVX1 U1404 ( .A(n2389), .Y(codefetch_s) );
  INVX1 U1405 ( .A(n2181), .Y(n2171) );
  INVX1 U1406 ( .A(n1868), .Y(n1816) );
  INVX1 U1407 ( .A(n613), .Y(N12770) );
  INVX1 U1408 ( .A(n762), .Y(n920) );
  INVX1 U1409 ( .A(n549), .Y(n548) );
  INVX1 U1410 ( .A(n640), .Y(n691) );
  INVX1 U1411 ( .A(n1228), .Y(n2071) );
  NAND21X1 U1412 ( .B(n1379), .A(n793), .Y(n580) );
  INVX1 U1413 ( .A(n1445), .Y(n1448) );
  INVX1 U1414 ( .A(n545), .Y(dps[1]) );
  NAND21X1 U1415 ( .B(n1333), .A(n1261), .Y(n581) );
  INVX1 U1416 ( .A(n1036), .Y(n996) );
  INVX1 U1417 ( .A(n494), .Y(n493) );
  OAI221X1 U1418 ( .A(n237), .B(n1898), .C(n1150), .D(n932), .E(n931), .Y(n933) );
  AO21XL U1419 ( .B(n930), .C(n1173), .A(n1480), .Y(n931) );
  INVX1 U1420 ( .A(n2224), .Y(n1439) );
  NOR3XL U1421 ( .A(n754), .B(n737), .C(n755), .Y(n236) );
  INVX1 U1422 ( .A(n610), .Y(n649) );
  NAND21X1 U1423 ( .B(n290), .A(n625), .Y(n610) );
  NAND32X1 U1424 ( .B(n735), .C(n1170), .A(n760), .Y(n736) );
  INVX1 U1425 ( .A(n759), .Y(n735) );
  INVX1 U1426 ( .A(n648), .Y(n2141) );
  NAND21X1 U1427 ( .B(n681), .A(n647), .Y(n648) );
  NAND21XL U1428 ( .B(n686), .A(n642), .Y(n645) );
  NAND21X1 U1429 ( .B(n1333), .A(n854), .Y(n2321) );
  NAND21XL U1430 ( .B(n1180), .A(n753), .Y(n1566) );
  NAND21X1 U1431 ( .B(n776), .A(n2148), .Y(n1277) );
  NAND21X1 U1432 ( .B(n2143), .A(cpu_hold), .Y(n875) );
  MUX4X1 U1433 ( .D0(n465), .D1(n463), .D2(n464), .D3(n462), .S0(n145), .S1(
        n133), .Y(n466) );
  MUX4X1 U1434 ( .D0(n460), .D1(n458), .D2(n459), .D3(n457), .S0(n145), .S1(
        n133), .Y(n461) );
  NAND32XL U1435 ( .B(n921), .C(n763), .A(n762), .Y(n1211) );
  AO222XL U1436 ( .A(n654), .B(n289), .C(N12807), .D(n137), .E(n208), .F(n643), 
        .Y(n1944) );
  AO21XL U1437 ( .B(n743), .C(n739), .A(n155), .Y(n737) );
  INVX1 U1438 ( .A(n2318), .Y(n1432) );
  AOI21BBXL U1439 ( .B(cpu_resume), .C(irq), .A(n554), .Y(N13379) );
  NAND32X1 U1440 ( .B(n754), .C(n736), .A(n737), .Y(n1565) );
  INVX1 U1441 ( .A(n1979), .Y(n2294) );
  AO21X1 U1442 ( .B(n812), .C(n2313), .A(n1104), .Y(n673) );
  INVX1 U1443 ( .A(n1987), .Y(n1998) );
  INVX1 U1444 ( .A(n1097), .Y(n847) );
  AOI21BXL U1445 ( .C(n1003), .B(n757), .A(n2297), .Y(n237) );
  INVX1 U1446 ( .A(n682), .Y(n1579) );
  INVX1 U1447 ( .A(n494), .Y(n492) );
  INVX1 U1448 ( .A(n785), .Y(n2226) );
  NAND21X1 U1449 ( .B(n2212), .A(n1441), .Y(n785) );
  INVX1 U1450 ( .A(n584), .Y(n854) );
  NAND21X1 U1451 ( .B(n1361), .A(n800), .Y(n584) );
  INVX1 U1452 ( .A(n547), .Y(dps[2]) );
  INVX1 U1453 ( .A(n1970), .Y(n765) );
  INVX1 U1454 ( .A(n1505), .Y(n2143) );
  NAND21X1 U1455 ( .B(n1302), .A(n802), .Y(n1358) );
  NAND21X1 U1456 ( .B(n606), .A(n635), .Y(n630) );
  AND4X1 U1457 ( .A(n2085), .B(n2093), .C(n1798), .D(n2091), .Y(n863) );
  NAND43X1 U1458 ( .B(n796), .C(n878), .D(n904), .A(n795), .Y(n1282) );
  INVX1 U1459 ( .A(n886), .Y(n796) );
  AND4X1 U1460 ( .A(n882), .B(n1770), .C(n881), .D(n883), .Y(n795) );
  NAND21X1 U1461 ( .B(n2118), .A(n1246), .Y(n1249) );
  NAND21X1 U1462 ( .B(n548), .A(n2169), .Y(n977) );
  NAND21X1 U1463 ( .B(n1194), .A(n922), .Y(n1966) );
  NAND21X1 U1464 ( .B(n1360), .A(n1094), .Y(n2149) );
  NAND21X1 U1465 ( .B(n1415), .A(n2169), .Y(n805) );
  NAND21X1 U1466 ( .B(n1361), .A(n1257), .Y(n2150) );
  INVX1 U1467 ( .A(n967), .Y(n2168) );
  NAND21X1 U1468 ( .B(n1333), .A(n30), .Y(n967) );
  INVX1 U1469 ( .A(n791), .Y(n799) );
  NAND21X1 U1470 ( .B(n2315), .A(n978), .Y(n791) );
  INVX1 U1471 ( .A(n1283), .Y(n672) );
  AND4X1 U1472 ( .A(n670), .B(n2356), .C(n669), .D(n668), .Y(n671) );
  INVX1 U1473 ( .A(n1807), .Y(N354) );
  OAI22X1 U1474 ( .A(n493), .B(n2160), .C(n586), .D(n859), .Y(n590) );
  NAND6XL U1475 ( .A(n1293), .B(n1292), .C(n2160), .D(n1291), .E(n1290), .F(
        n1289), .Y(n1298) );
  OA222X1 U1476 ( .A(n1281), .B(n1360), .C(n2156), .D(n1280), .E(n1415), .F(
        n1435), .Y(n1290) );
  INVX1 U1477 ( .A(n1373), .Y(n1293) );
  NOR8XL U1478 ( .A(n1288), .B(n1287), .C(n1286), .D(n1285), .E(n1284), .F(
        n1283), .G(n1282), .H(n1315), .Y(n1289) );
  INVX1 U1479 ( .A(n1500), .Y(n1362) );
  INVX1 U1480 ( .A(n1267), .Y(n1843) );
  INVX1 U1481 ( .A(n1369), .Y(n1383) );
  INVX1 U1482 ( .A(n973), .Y(n1246) );
  INVX1 U1483 ( .A(n1835), .Y(n978) );
  NAND6XL U1484 ( .A(n811), .B(n2358), .C(n1292), .D(n810), .E(n809), .F(n808), 
        .Y(n835) );
  AOI31X1 U1485 ( .A(n1338), .B(n1339), .C(n1101), .D(n798), .Y(n810) );
  INVX1 U1486 ( .A(n1284), .Y(n811) );
  INVX1 U1487 ( .A(n848), .Y(n1304) );
  INVX1 U1488 ( .A(n1964), .Y(n1482) );
  INVX1 U1489 ( .A(n889), .Y(n887) );
  INVX1 U1490 ( .A(n1581), .Y(n2231) );
  INVX1 U1491 ( .A(n651), .Y(N12776) );
  INVX1 U1492 ( .A(n543), .Y(dps[0]) );
  INVX1 U1493 ( .A(n2154), .Y(n802) );
  INVX1 U1494 ( .A(n1195), .Y(n1192) );
  INVX1 U1495 ( .A(n709), .Y(n676) );
  AOI221XL U1496 ( .A(n812), .B(n1105), .C(n879), .D(n477), .E(n667), .Y(n668)
         );
  AOI211X1 U1497 ( .C(n1362), .D(n1267), .A(n807), .B(n806), .Y(n808) );
  INVX1 U1498 ( .A(n805), .Y(n806) );
  INVX1 U1499 ( .A(n666), .Y(n794) );
  INVX1 U1500 ( .A(n679), .Y(n2267) );
  AO21X1 U1501 ( .B(n298), .C(n889), .A(n1066), .Y(n1768) );
  OR3XL U1502 ( .A(n872), .B(n871), .C(n238), .Y(n2382) );
  AOI21X1 U1503 ( .B(n1061), .C(n870), .A(n2163), .Y(n238) );
  NAND32X1 U1504 ( .B(n848), .C(n477), .A(n847), .Y(n1403) );
  NAND21X1 U1505 ( .B(n1101), .A(n1846), .Y(n1408) );
  NAND21X1 U1506 ( .B(n2313), .A(n1370), .Y(n813) );
  NAND21X1 U1507 ( .B(n2313), .A(n1383), .Y(n797) );
  NAND32X1 U1508 ( .B(n2315), .C(n1366), .A(n477), .Y(n1270) );
  INVX1 U1509 ( .A(n1224), .Y(n1235) );
  NAND21X1 U1510 ( .B(n1267), .A(n1223), .Y(n1224) );
  OAI31XL U1511 ( .A(n1247), .B(n496), .C(n1363), .D(n1980), .Y(n1974) );
  NAND5XL U1512 ( .A(n950), .B(n2332), .C(n951), .D(n1865), .E(n949), .Y(n2396) );
  NAND21X1 U1513 ( .B(n2082), .A(ramdatai[0]), .Y(n1858) );
  OAI221X1 U1514 ( .A(n850), .B(n877), .C(n1403), .D(n1385), .E(n885), .Y(
        n1285) );
  OAI211X1 U1515 ( .C(n1276), .D(n1425), .A(n1275), .B(n1274), .Y(n1373) );
  INVX1 U1516 ( .A(n1263), .Y(n1276) );
  NAND32X1 U1517 ( .B(n2155), .C(n977), .A(n2315), .Y(n881) );
  NAND21X1 U1518 ( .B(n1415), .A(n662), .Y(n1291) );
  NAND43X1 U1519 ( .B(n817), .C(n816), .D(n1234), .A(n965), .Y(n834) );
  INVX1 U1520 ( .A(n1314), .Y(n816) );
  NAND32XL U1521 ( .B(n921), .C(n2060), .A(n920), .Y(n1968) );
  NAND21X1 U1522 ( .B(n1302), .A(n1094), .Y(n1328) );
  INVX1 U1523 ( .A(ramdatai[0]), .Y(n1460) );
  INVX1 U1524 ( .A(n697), .Y(n1370) );
  INVX1 U1525 ( .A(n1365), .Y(n1329) );
  INVX1 U1526 ( .A(ramdatai[1]), .Y(n1483) );
  INVX1 U1527 ( .A(ramdatai[2]), .Y(n1574) );
  INVX1 U1528 ( .A(n1434), .Y(n1338) );
  INVX1 U1529 ( .A(n1268), .Y(n1845) );
  INVX1 U1530 ( .A(n1767), .Y(n1066) );
  AND3X1 U1531 ( .A(n1271), .B(n1270), .C(n1269), .Y(n1272) );
  AND3X1 U1532 ( .A(n1102), .B(n1406), .C(n1101), .Y(n1103) );
  INVX1 U1533 ( .A(n1366), .Y(n1260) );
  MUX2IX1 U1534 ( .D0(n2120), .D1(n2163), .S(n2165), .Y(n239) );
  INVX1 U1535 ( .A(n1415), .Y(n1295) );
  INVX1 U1536 ( .A(n883), .Y(n902) );
  INVX1 U1537 ( .A(n1506), .Y(n1165) );
  NAND21X1 U1538 ( .B(n848), .A(n1339), .Y(n1435) );
  OAI21AX1 U1539 ( .B(n1010), .C(n814), .A(n2028), .Y(n2244) );
  NAND21X1 U1540 ( .B(n2313), .A(n1492), .Y(n1314) );
  NAND32X1 U1541 ( .B(n771), .C(n770), .A(n769), .Y(n1499) );
  NAND32X1 U1542 ( .B(n714), .C(n713), .A(n2206), .Y(n1501) );
  NAND21XL U1543 ( .B(n2146), .A(n1253), .Y(n1255) );
  NAND21X1 U1544 ( .B(n1360), .A(n30), .Y(n1423) );
  NAND21X1 U1545 ( .B(n697), .A(n1329), .Y(n789) );
  NAND32X1 U1546 ( .B(n103), .C(n977), .A(n976), .Y(n1275) );
  OAI221X1 U1547 ( .A(n700), .B(n496), .C(n699), .D(n2163), .E(n698), .Y(n714)
         );
  AND3X1 U1548 ( .A(n2173), .B(n1291), .C(n1009), .Y(n699) );
  INVX1 U1549 ( .A(n2244), .Y(n698) );
  AOI221XL U1550 ( .A(n1218), .B(n2157), .C(n696), .D(n1335), .E(n718), .Y(
        n700) );
  NAND32X1 U1551 ( .B(n770), .C(n769), .A(n724), .Y(n2044) );
  OAI31XL U1552 ( .A(n1415), .B(n2316), .C(n1302), .D(n789), .Y(n718) );
  NAND32X1 U1553 ( .B(n849), .C(n2155), .A(n1267), .Y(n2361) );
  INVX1 U1554 ( .A(n1980), .Y(n1993) );
  INVX1 U1555 ( .A(n1302), .Y(n1339) );
  NAND32X1 U1556 ( .B(n772), .C(n714), .A(n713), .Y(n770) );
  NAND21X1 U1557 ( .B(n1500), .A(n1402), .Y(n870) );
  INVX1 U1558 ( .A(n859), .Y(n702) );
  NAND32X1 U1559 ( .B(n1840), .C(n1263), .A(n1251), .Y(n701) );
  INVX1 U1560 ( .A(n1360), .Y(n1305) );
  AND3XL U1561 ( .A(n1434), .B(n2146), .C(n1365), .Y(n777) );
  INVX1 U1562 ( .A(n660), .Y(n1364) );
  INVX1 U1563 ( .A(n1386), .Y(n1410) );
  INVX1 U1564 ( .A(n2153), .Y(n2312) );
  INVX1 U1565 ( .A(n801), .Y(n775) );
  INVX1 U1566 ( .A(n661), .Y(n719) );
  NAND21X1 U1567 ( .B(n1910), .A(n2399), .Y(n1782) );
  MUX2X1 U1568 ( .D0(n1226), .D1(n1458), .S(n295), .Y(n894) );
  MUX2IX1 U1569 ( .D0(n1225), .D1(n1481), .S(n295), .Y(n241) );
  NAND21X1 U1570 ( .B(n1910), .A(n1868), .Y(n1812) );
  OR3XL U1571 ( .A(n1364), .B(n913), .C(n242), .Y(n915) );
  AOI21X1 U1572 ( .B(n2362), .C(n870), .A(n2163), .Y(n242) );
  INVX1 U1573 ( .A(ramdatai[5]), .Y(n1957) );
  NAND21X1 U1574 ( .B(n1329), .A(n1337), .Y(n1335) );
  INVX1 U1575 ( .A(ramdatai[6]), .Y(n2018) );
  INVX1 U1576 ( .A(n776), .Y(n855) );
  INVX1 U1577 ( .A(n843), .Y(n1402) );
  INVX1 U1578 ( .A(n2174), .Y(n2373) );
  NAND32X1 U1579 ( .B(n496), .C(n2173), .A(n2181), .Y(n2174) );
  INVX1 U1580 ( .A(n968), .Y(n1215) );
  INVX1 U1581 ( .A(n704), .Y(n1334) );
  NAND21X1 U1582 ( .B(n103), .A(n2312), .Y(n704) );
  INVX1 U1583 ( .A(n2238), .Y(n578) );
  NAND32X1 U1584 ( .B(n1500), .C(n493), .A(n710), .Y(n724) );
  NAND21X1 U1585 ( .B(n2091), .A(pc_i[9]), .Y(n951) );
  INVX1 U1586 ( .A(n913), .Y(n2084) );
  NAND2X1 U1587 ( .A(n2104), .B(n955), .Y(n2368) );
  NAND32XL U1588 ( .B(n2365), .C(n2389), .A(n2391), .Y(n2198) );
  NAND21X1 U1589 ( .B(n1010), .A(n2167), .Y(n2001) );
  OAI211XL U1590 ( .C(n954), .D(n2396), .A(n2395), .B(n953), .Y(n1090) );
  INVX1 U1591 ( .A(n952), .Y(n954) );
  OAI211X1 U1592 ( .C(n2399), .D(n1914), .A(n952), .B(n2378), .Y(n953) );
  NAND21X1 U1593 ( .B(n2088), .A(n7), .Y(n952) );
  NAND21X1 U1594 ( .B(n1194), .A(n902), .Y(n1773) );
  OAI221X1 U1595 ( .A(n1066), .B(n1065), .C(sfrdatai[3]), .D(n1065), .E(n906), 
        .Y(n909) );
  INVX1 U1596 ( .A(n905), .Y(n906) );
  INVX1 U1597 ( .A(pc_i[1]), .Y(n1475) );
  INVX1 U1598 ( .A(n1009), .Y(n2128) );
  NAND21X1 U1599 ( .B(n1914), .A(n2386), .Y(n911) );
  NAND21X1 U1600 ( .B(n2056), .A(n2055), .Y(n2414) );
  AO2222XL U1601 ( .A(n2049), .B(n2193), .C(alu_out[7]), .D(n114), .E(n2048), 
        .F(n2047), .G(ramdatai[7]), .H(n2046), .Y(n2056) );
  OA2222XL U1602 ( .A(n2096), .B(n2054), .C(n2053), .D(n2052), .E(n2051), .F(
        n2092), .G(n2050), .H(n50), .Y(n2055) );
  INVX1 U1603 ( .A(pc_i[4]), .Y(n1818) );
  INVX1 U1604 ( .A(pc_i[5]), .Y(n1788) );
  INVX1 U1605 ( .A(n2109), .Y(n2125) );
  INVX1 U1606 ( .A(n2364), .Y(n1086) );
  INVX1 U1607 ( .A(pc_i[3]), .Y(n1647) );
  INVX1 U1608 ( .A(pc_i[2]), .Y(n1905) );
  NAND21X1 U1609 ( .B(n1445), .A(n212), .Y(n1532) );
  OAI31XL U1610 ( .A(n1450), .B(n2046), .C(n1449), .D(n202), .Y(n1893) );
  OA222X1 U1611 ( .A(n2082), .B(n1957), .C(n1935), .D(n2080), .E(n122), .F(
        n1958), .Y(n1937) );
  OA222X1 U1612 ( .A(n2082), .B(n1793), .C(n1792), .D(n2080), .E(n122), .F(
        n1791), .Y(n1795) );
  OA222X1 U1613 ( .A(n2082), .B(n1825), .C(n1820), .D(n2080), .E(n122), .F(
        n1821), .Y(n1796) );
  GEN2XL U1614 ( .D(cs_run), .E(n2132), .C(n2131), .B(n2133), .A(n2130), .Y(
        n2375) );
  NAND21X1 U1615 ( .B(n2123), .A(n2122), .Y(n2132) );
  GEN2XL U1616 ( .D(n2129), .E(n2171), .C(n2128), .B(n2127), .A(n2126), .Y(
        n2130) );
  OAI221X1 U1617 ( .A(n2093), .B(n1940), .C(n2091), .D(n2009), .E(n1939), .Y(
        n1942) );
  OA222X1 U1618 ( .A(n2088), .B(n1938), .C(n2085), .D(n2015), .E(n36), .F(
        n2086), .Y(n1939) );
  XOR3X1 U1619 ( .A(n2084), .B(n250), .C(n2076), .Y(n1938) );
  OAI222XL U1620 ( .A(n243), .B(n2347), .C(n2343), .D(n2345), .E(n551), .F(
        n2342), .Y(ramdatao_comb[6]) );
  OAI222XL U1621 ( .A(n246), .B(n2347), .C(n2346), .D(n2345), .E(waitstaten), 
        .F(n2344), .Y(ramdatao_comb[7]) );
  OAI221X1 U1622 ( .A(n2093), .B(n2092), .C(n2091), .D(n2090), .E(n2089), .Y(
        n2100) );
  OA222X1 U1623 ( .A(n2088), .B(n2087), .C(n50), .D(n2086), .E(n2085), .F(n38), 
        .Y(n2089) );
  NOR31X1 U1624 ( .C(n244), .A(n1942), .B(n245), .Y(n243) );
  OAI222XL U1625 ( .A(n2018), .B(n2098), .C(n2097), .D(n2007), .E(n2094), .F(
        n1941), .Y(n245) );
  NOR31X1 U1626 ( .C(n247), .A(n2100), .B(n248), .Y(n246) );
  AOI22X1 U1627 ( .A(n91), .B(n2075), .C(n2074), .D(n2073), .Y(n247) );
  OAI222XL U1628 ( .A(n2099), .B(n2098), .C(n2097), .D(n2096), .E(n2095), .F(
        n2094), .Y(n248) );
  INVX1 U1629 ( .A(n726), .Y(n1085) );
  INVX1 U1630 ( .A(sfrdatai[5]), .Y(n1958) );
  INVX1 U1631 ( .A(sfrdatai[4]), .Y(n1821) );
  OA222X1 U1632 ( .A(n2088), .B(n1801), .C(n1957), .D(n2098), .E(n1954), .F(
        n1932), .Y(n1802) );
  OAI222XL U1633 ( .A(n122), .B(n1958), .C(n1935), .D(n2080), .E(n2082), .F(
        n1957), .Y(n1797) );
  OAI22X1 U1634 ( .A(n1768), .B(n1957), .C(n1767), .D(n1958), .Y(n1775) );
  OAI22X1 U1635 ( .A(n1768), .B(n1825), .C(n1767), .D(n1821), .Y(n1808) );
  OA222X1 U1636 ( .A(n2088), .B(n1826), .C(n1825), .D(n2098), .E(n1824), .F(
        n1932), .Y(n1830) );
  OAI222XL U1637 ( .A(n122), .B(n1821), .C(n1820), .D(n2080), .E(n2082), .F(
        n1825), .Y(n1822) );
  INVX1 U1638 ( .A(n1832), .Y(n2338) );
  OA222X1 U1639 ( .A(n2094), .B(n1828), .C(n2085), .D(n1827), .E(n34), .F(
        n2086), .Y(n1829) );
  INVX1 U1640 ( .A(n1804), .Y(n2341) );
  AO21X1 U1641 ( .B(n1774), .C(n1773), .A(n1779), .Y(n1928) );
  AO2222XL U1642 ( .A(n1786), .B(n1775), .C(n1816), .D(n1808), .E(n1769), .F(
        n1920), .G(n2071), .H(n2058), .Y(n1772) );
  OAI222XL U1643 ( .A(n2338), .B(n2347), .C(n2337), .D(n2345), .E(waitstaten), 
        .F(n2336), .Y(ramdatao_comb[4]) );
  OAI222XL U1644 ( .A(n2341), .B(n2347), .C(n2340), .D(n2345), .E(waitstaten), 
        .F(n2339), .Y(ramdatao_comb[5]) );
  OAI221X1 U1645 ( .A(n1931), .B(n1930), .C(n1929), .D(n1928), .E(n1927), .Y(
        n1934) );
  AOI211X1 U1646 ( .C(n1924), .D(n2068), .A(n1923), .B(n1922), .Y(n1930) );
  AO21X1 U1647 ( .B(n1926), .C(n1925), .A(n1924), .Y(n1927) );
  MUX2X1 U1648 ( .D0(n1921), .D1(n2006), .S(n295), .Y(n1924) );
  MUX2XL U1649 ( .D0(n1877), .D1(n2275), .S(n2331), .Y(n2329) );
  NAND32X1 U1650 ( .B(n1876), .C(n1875), .A(n1874), .Y(n1877) );
  OA2222XL U1651 ( .A(n2091), .B(n1873), .C(n1872), .D(n2097), .E(n2093), .F(
        n1871), .G(n2085), .H(n40), .Y(n1874) );
  OA222X1 U1652 ( .A(n2088), .B(n1075), .C(n2094), .D(n1642), .E(n1074), .F(
        n1865), .Y(n1076) );
  OA222X1 U1653 ( .A(n1073), .B(n1072), .C(n1071), .D(n1070), .E(n1228), .F(
        n1914), .Y(n1074) );
  XOR3X1 U1654 ( .A(n2084), .B(n1794), .C(n251), .Y(n1075) );
  AND3X1 U1655 ( .A(n1068), .B(n2064), .C(n1067), .Y(n1072) );
  OAI22X1 U1656 ( .A(n1768), .B(n2018), .C(n1767), .D(n2021), .Y(n1920) );
  OAI22X1 U1657 ( .A(n1768), .B(n2099), .C(n1767), .D(n2078), .Y(n2058) );
  OAI222XL U1658 ( .A(n175), .B(n2347), .C(n2334), .D(n2345), .E(waitstaten), 
        .F(n2333), .Y(ramdatao_comb[2]) );
  OAI21BBX1 U1659 ( .A(n91), .B(n1870), .C(n1869), .Y(n1875) );
  INVX1 U1660 ( .A(sfrdatai[6]), .Y(n2021) );
  INVX1 U1661 ( .A(sfrdatai[7]), .Y(n2078) );
  OA222X1 U1662 ( .A(n2093), .B(n1905), .C(n2097), .D(n1904), .E(n1903), .F(
        n2094), .Y(n1906) );
  XOR3X1 U1663 ( .A(n2084), .B(n249), .C(n1902), .Y(n1907) );
  OAI221X1 U1664 ( .A(n2085), .B(n1901), .C(n32), .D(n2086), .E(n1900), .Y(
        n1918) );
  OA222X1 U1665 ( .A(n122), .B(n2021), .C(n2002), .D(n2080), .E(n2082), .F(
        n2018), .Y(n250) );
  OA222X1 U1666 ( .A(n122), .B(n1791), .C(n1792), .D(n130), .E(n117), .F(n1793), .Y(n251) );
  OAI211X1 U1667 ( .C(n2044), .D(n1819), .A(n1548), .B(n1547), .Y(n2278) );
  OA22XL U1668 ( .A(n1824), .B(n219), .C(n1820), .D(n2038), .Y(n1548) );
  OA222X1 U1669 ( .A(n2041), .B(n1546), .C(n2040), .D(n1821), .E(n218), .F(
        n1825), .Y(n1547) );
  OAI211XL U1670 ( .C(n1792), .D(n2038), .A(n1080), .B(n1079), .Y(n2279) );
  OA22X1 U1671 ( .A(n1557), .B(n1499), .C(n1418), .D(n1793), .Y(n1080) );
  INVX1 U1672 ( .A(n1562), .Y(n2340) );
  OAI211X1 U1673 ( .C(n2044), .D(n1789), .A(n1561), .B(n1560), .Y(n1562) );
  OA22X1 U1674 ( .A(n1954), .B(n219), .C(n1935), .D(n2038), .Y(n1561) );
  OA222X1 U1675 ( .A(n2041), .B(n1956), .C(n2040), .D(n1958), .E(n218), .F(
        n1957), .Y(n1560) );
  OR2X1 U1676 ( .A(n554), .B(n252), .Y(n2135) );
  AOI21X1 U1677 ( .B(cs_run), .C(n2133), .A(n2364), .Y(n252) );
  OAI31XL U1678 ( .A(n2366), .B(cs_run), .C(n2364), .D(n2390), .Y(n2105) );
  INVX1 U1679 ( .A(n2133), .Y(n2366) );
  OAI22X1 U1680 ( .A(n2363), .B(n2113), .C(n1849), .D(n2135), .Y(n1880) );
  OAI22X1 U1681 ( .A(n2363), .B(n2137), .C(n2136), .D(n2135), .Y(n1879) );
  AOI21X1 U1682 ( .B(n1851), .C(n1850), .A(n557), .Y(N515) );
  NAND21XL U1683 ( .B(n2390), .A(n2330), .Y(n1851) );
  AO21X1 U1684 ( .B(n2113), .C(n1849), .A(n2105), .Y(n1850) );
  OR2X1 U1685 ( .A(n505), .B(n253), .Y(n961) );
  AOI21X1 U1686 ( .B(n2144), .C(n2108), .A(n2389), .Y(n253) );
  NAND32X1 U1687 ( .B(n2364), .C(n506), .A(n2366), .Y(n2363) );
  OAI211X1 U1688 ( .C(n2013), .D(n219), .A(n1504), .B(n1503), .Y(n2276) );
  OA22X1 U1689 ( .A(n2002), .B(n2038), .C(n2044), .D(n2007), .Y(n1504) );
  NAND21X1 U1690 ( .B(n2365), .A(n726), .Y(n2111) );
  INVX1 U1691 ( .A(n2108), .Y(n2145) );
  AND2X1 U1692 ( .A(n510), .B(n2133), .Y(N588) );
  INVX1 U1693 ( .A(n2045), .Y(n2346) );
  OAI211X1 U1694 ( .C(n2044), .D(n2096), .A(n2043), .B(n2042), .Y(n2045) );
  OA22XL U1695 ( .A(n2039), .B(n219), .C(n2081), .D(n2038), .Y(n2043) );
  INVX1 U1696 ( .A(n1422), .Y(n2334) );
  OA22X1 U1697 ( .A(n1909), .B(n1499), .C(n1418), .D(n1574), .Y(n1420) );
  NAND21X1 U1698 ( .B(n2144), .A(n2108), .Y(n962) );
  AND2X1 U1699 ( .A(n511), .B(n2335), .Y(N11501) );
  INVX1 U1700 ( .A(n901), .Y(n1065) );
  NAND21X1 U1701 ( .B(n1768), .A(ramdatai[3]), .Y(n901) );
  NAND21X1 U1702 ( .B(n1452), .A(n301), .Y(n1891) );
  NAND21X1 U1703 ( .B(n2189), .A(n301), .Y(n1892) );
  NAND32X1 U1704 ( .B(n1449), .C(n1760), .A(n2000), .Y(n1451) );
  INVX1 U1705 ( .A(n2073), .Y(n2039) );
  NAND32XL U1706 ( .B(n540), .C(n1721), .A(n43), .Y(n1720) );
  NAND32XL U1707 ( .B(n2266), .C(n1721), .A(n539), .Y(n1752) );
  NAND32XL U1708 ( .B(n43), .C(n1710), .A(n539), .Y(n1712) );
  NAND21X1 U1709 ( .B(n153), .A(n1713), .Y(n1710) );
  NAND21X1 U1710 ( .B(n2342), .A(n500), .Y(n2023) );
  NAND21X1 U1711 ( .B(n1948), .A(n499), .Y(n1582) );
  NAND21X1 U1712 ( .B(n2339), .A(n500), .Y(n1951) );
  NAND21X1 U1713 ( .B(n2336), .A(n499), .Y(n1535) );
  NAND21X1 U1714 ( .B(n2178), .A(n498), .Y(n1440) );
  NAND21X1 U1715 ( .B(n2176), .A(n498), .Y(n1468) );
  NAND21X1 U1716 ( .B(n2333), .A(n499), .Y(n1887) );
  INVX1 U1717 ( .A(n1021), .Y(n2439) );
  NAND21X1 U1718 ( .B(n2059), .A(n1978), .Y(n1021) );
  AO21X1 U1719 ( .B(n2229), .C(n2234), .A(n559), .Y(N13257) );
  AO21X1 U1720 ( .B(n2222), .C(n2229), .A(n559), .Y(N13185) );
  AO21X1 U1721 ( .B(n2217), .C(n2229), .A(n560), .Y(N13113) );
  AO21X1 U1722 ( .B(n2215), .C(n2229), .A(n561), .Y(N13041) );
  OAI211X1 U1723 ( .C(n2306), .D(n2305), .A(n2304), .B(n2303), .Y(n2308) );
  NAND6XL U1724 ( .A(n2294), .B(n2293), .C(n2292), .D(n2291), .E(n2290), .F(
        n2289), .Y(n2304) );
  INVX1 U1725 ( .A(n2219), .Y(n2223) );
  INVX1 U1726 ( .A(n2221), .Y(n2222) );
  NAND32X1 U1727 ( .B(n2220), .C(n2219), .A(n2218), .Y(n2221) );
  INVX1 U1728 ( .A(n2208), .Y(n2215) );
  NAND32X1 U1729 ( .B(n2218), .C(n2220), .A(n2223), .Y(n2208) );
  INVX1 U1730 ( .A(n2248), .Y(n2230) );
  INVX1 U1731 ( .A(n2216), .Y(n2217) );
  NAND21X1 U1732 ( .B(n2250), .A(n2223), .Y(n2216) );
  INVX1 U1733 ( .A(n2225), .Y(n2234) );
  NAND21X1 U1734 ( .B(n2224), .A(n2223), .Y(n2225) );
  OAI22X1 U1735 ( .A(n1759), .B(n1716), .C(n1757), .D(n1715), .Y(N12530) );
  OAI22X1 U1736 ( .A(n1759), .B(n1718), .C(n1757), .D(n141), .Y(N12539) );
  OAI22X1 U1737 ( .A(n1736), .B(n1716), .C(n1735), .D(n1715), .Y(N12602) );
  OAI22X1 U1738 ( .A(n304), .B(n1716), .C(n1734), .D(n1715), .Y(N12603) );
  OAI22X1 U1739 ( .A(n1731), .B(n1716), .C(n1730), .D(n1715), .Y(N12605) );
  OAI22X1 U1740 ( .A(n1729), .B(n1716), .C(n1728), .D(n1715), .Y(N12606) );
  OAI22X1 U1741 ( .A(n1727), .B(n1716), .C(n1726), .D(n1715), .Y(N12607) );
  OAI22X1 U1742 ( .A(n1725), .B(n1716), .C(n1998), .D(n1715), .Y(N12608) );
  OAI22X1 U1743 ( .A(n1724), .B(n1716), .C(n1723), .D(n1715), .Y(N12609) );
  OAI22X1 U1744 ( .A(n1750), .B(n131), .C(n1749), .D(n107), .Y(N12531) );
  OAI22X1 U1745 ( .A(n1748), .B(n131), .C(n1747), .D(n107), .Y(N12532) );
  OAI22X1 U1746 ( .A(n1746), .B(n131), .C(n1745), .D(n107), .Y(N12533) );
  OAI22X1 U1747 ( .A(n1744), .B(n131), .C(n1743), .D(n107), .Y(N12534) );
  OAI22X1 U1748 ( .A(n1742), .B(n131), .C(n1741), .D(n107), .Y(N12535) );
  OAI22X1 U1749 ( .A(n1740), .B(n131), .C(n1739), .D(n107), .Y(N12536) );
  OAI22X1 U1750 ( .A(n1738), .B(n131), .C(n1737), .D(n107), .Y(N12537) );
  OAI22X1 U1751 ( .A(n1736), .B(n1718), .C(n1735), .D(n141), .Y(N12611) );
  OAI22X1 U1752 ( .A(n304), .B(n1718), .C(n1734), .D(n141), .Y(N12612) );
  OAI22X1 U1753 ( .A(n1731), .B(n1718), .C(n1730), .D(n141), .Y(N12614) );
  OAI22X1 U1754 ( .A(n1729), .B(n1718), .C(n1728), .D(n141), .Y(N12615) );
  OAI22X1 U1755 ( .A(n1727), .B(n1718), .C(n1726), .D(n142), .Y(N12616) );
  OAI22X1 U1756 ( .A(n1725), .B(n1718), .C(n1998), .D(n142), .Y(N12617) );
  OAI22X1 U1757 ( .A(n1724), .B(n1718), .C(n1723), .D(n142), .Y(N12618) );
  OAI22X1 U1758 ( .A(n1750), .B(n105), .C(n1749), .D(n142), .Y(N12540) );
  OAI22X1 U1759 ( .A(n1748), .B(n105), .C(n1747), .D(n142), .Y(N12541) );
  OAI22X1 U1760 ( .A(n1746), .B(n105), .C(n1745), .D(n142), .Y(N12542) );
  OAI22X1 U1761 ( .A(n1744), .B(n105), .C(n1743), .D(n142), .Y(N12543) );
  OAI22X1 U1762 ( .A(n1742), .B(n105), .C(n1741), .D(n142), .Y(N12544) );
  OAI22X1 U1763 ( .A(n1740), .B(n105), .C(n1739), .D(n142), .Y(N12545) );
  OAI22X1 U1764 ( .A(n1738), .B(n105), .C(n1737), .D(n142), .Y(N12546) );
  OAI22X1 U1765 ( .A(n555), .B(n1959), .C(n1958), .D(n2020), .Y(N12719) );
  OA2222XL U1766 ( .A(n2019), .B(n1957), .C(n2017), .D(n1956), .E(n1955), .F(
        n2014), .G(n1954), .H(n2012), .Y(n1959) );
  OAI22X1 U1767 ( .A(n555), .B(n1538), .C(n1821), .D(n2020), .Y(N12718) );
  OA2222XL U1768 ( .A(n2019), .B(n1825), .C(n2017), .D(n1546), .E(n1827), .F(
        n2014), .G(n1824), .H(n2012), .Y(n1538) );
  OAI22X1 U1769 ( .A(n1759), .B(n1758), .C(n1757), .D(n1756), .Y(N12494) );
  OAI22X1 U1770 ( .A(n1759), .B(n1707), .C(n1757), .D(n1706), .Y(N12503) );
  OAI22X1 U1771 ( .A(n1759), .B(n1709), .C(n1757), .D(n1708), .Y(N12512) );
  OAI22X1 U1772 ( .A(n1759), .B(n1712), .C(n1757), .D(n47), .Y(N12521) );
  OAI22X1 U1773 ( .A(n1759), .B(n1720), .C(n1757), .D(n1719), .Y(N12548) );
  OAI22X1 U1774 ( .A(n1759), .B(n1752), .C(n1757), .D(n1751), .Y(N12557) );
  OAI22X1 U1775 ( .A(n1736), .B(n1720), .C(n1735), .D(n1719), .Y(N12620) );
  OAI22X1 U1776 ( .A(n304), .B(n1720), .C(n1734), .D(n1719), .Y(N12621) );
  OAI22X1 U1777 ( .A(n1731), .B(n1720), .C(n1730), .D(n1719), .Y(N12623) );
  OAI22X1 U1778 ( .A(n1729), .B(n1720), .C(n1728), .D(n1719), .Y(N12624) );
  OAI22X1 U1779 ( .A(n1727), .B(n1720), .C(n1726), .D(n1719), .Y(N12625) );
  OAI22X1 U1780 ( .A(n1725), .B(n1720), .C(n1998), .D(n1719), .Y(N12626) );
  OAI22X1 U1781 ( .A(n1724), .B(n1720), .C(n1723), .D(n1719), .Y(N12627) );
  OAI22X1 U1782 ( .A(n1750), .B(n144), .C(n1749), .D(n123), .Y(N12549) );
  OAI22X1 U1783 ( .A(n1748), .B(n144), .C(n1747), .D(n123), .Y(N12550) );
  OAI22X1 U1784 ( .A(n1746), .B(n144), .C(n1745), .D(n123), .Y(N12551) );
  OAI22X1 U1785 ( .A(n1744), .B(n144), .C(n1743), .D(n123), .Y(N12552) );
  OAI22X1 U1786 ( .A(n1742), .B(n144), .C(n1741), .D(n123), .Y(N12553) );
  OAI22X1 U1787 ( .A(n1740), .B(n144), .C(n1739), .D(n123), .Y(N12554) );
  OAI22X1 U1788 ( .A(n1738), .B(n144), .C(n1737), .D(n123), .Y(N12555) );
  OAI22X1 U1789 ( .A(n1736), .B(n1752), .C(n1735), .D(n1751), .Y(N12629) );
  OAI22X1 U1790 ( .A(n304), .B(n1752), .C(n1734), .D(n1751), .Y(N12630) );
  OAI22X1 U1791 ( .A(n1731), .B(n1752), .C(n1730), .D(n1751), .Y(N12632) );
  OAI22X1 U1792 ( .A(n1729), .B(n1752), .C(n1728), .D(n1751), .Y(N12633) );
  OAI22X1 U1793 ( .A(n1727), .B(n1752), .C(n1726), .D(n1751), .Y(N12634) );
  OAI22X1 U1794 ( .A(n1725), .B(n1752), .C(n1998), .D(n1751), .Y(N12635) );
  OAI22X1 U1795 ( .A(n1724), .B(n1752), .C(n1723), .D(n1751), .Y(N12636) );
  OAI22X1 U1796 ( .A(n1750), .B(n132), .C(n1749), .D(n102), .Y(N12558) );
  OAI22X1 U1797 ( .A(n1748), .B(n132), .C(n1747), .D(n102), .Y(N12559) );
  OAI22X1 U1798 ( .A(n1746), .B(n132), .C(n1745), .D(n102), .Y(N12560) );
  OAI22X1 U1799 ( .A(n1744), .B(n132), .C(n1743), .D(n102), .Y(N12561) );
  OAI22X1 U1800 ( .A(n1742), .B(n132), .C(n1741), .D(n102), .Y(N12562) );
  OAI22X1 U1801 ( .A(n1740), .B(n132), .C(n1739), .D(n102), .Y(N12563) );
  OAI22X1 U1802 ( .A(n1738), .B(n132), .C(n1737), .D(n102), .Y(N12564) );
  OAI22X1 U1803 ( .A(n1736), .B(n1758), .C(n1735), .D(n1756), .Y(N12566) );
  OAI22X1 U1804 ( .A(n304), .B(n1758), .C(n1734), .D(n1756), .Y(N12567) );
  OAI22X1 U1805 ( .A(n1731), .B(n1758), .C(n1730), .D(n1756), .Y(N12569) );
  OAI22X1 U1806 ( .A(n1729), .B(n1758), .C(n1728), .D(n1756), .Y(N12570) );
  OAI22X1 U1807 ( .A(n1727), .B(n1758), .C(n1726), .D(n1756), .Y(N12571) );
  OAI22X1 U1808 ( .A(n1725), .B(n1758), .C(n1998), .D(n1756), .Y(N12572) );
  OAI22X1 U1809 ( .A(n1724), .B(n1758), .C(n1723), .D(n1756), .Y(N12573) );
  OAI22X1 U1810 ( .A(n1750), .B(n143), .C(n1749), .D(n118), .Y(N12495) );
  OAI22X1 U1811 ( .A(n1748), .B(n143), .C(n1747), .D(n118), .Y(N12496) );
  OAI22X1 U1812 ( .A(n1746), .B(n143), .C(n1745), .D(n118), .Y(N12497) );
  OAI22X1 U1813 ( .A(n1744), .B(n143), .C(n1743), .D(n118), .Y(N12498) );
  OAI22X1 U1814 ( .A(n1742), .B(n143), .C(n1741), .D(n118), .Y(N12499) );
  OAI22X1 U1815 ( .A(n1740), .B(n143), .C(n1739), .D(n118), .Y(N12500) );
  OAI22X1 U1816 ( .A(n1738), .B(n143), .C(n1737), .D(n118), .Y(N12501) );
  OAI22X1 U1817 ( .A(n1736), .B(n1707), .C(n1735), .D(n1706), .Y(N12575) );
  OAI22X1 U1818 ( .A(n304), .B(n1707), .C(n1734), .D(n1706), .Y(N12576) );
  OAI22X1 U1819 ( .A(n1731), .B(n1707), .C(n1730), .D(n1706), .Y(N12578) );
  OAI22X1 U1820 ( .A(n1729), .B(n1707), .C(n1728), .D(n1706), .Y(N12579) );
  OAI22X1 U1821 ( .A(n1727), .B(n1707), .C(n1726), .D(n1706), .Y(N12580) );
  OAI22X1 U1822 ( .A(n1725), .B(n1707), .C(n1998), .D(n1706), .Y(N12581) );
  OAI22X1 U1823 ( .A(n1724), .B(n1707), .C(n1723), .D(n1706), .Y(N12582) );
  OAI22X1 U1824 ( .A(n1750), .B(n124), .C(n1749), .D(n99), .Y(N12504) );
  OAI22X1 U1825 ( .A(n1748), .B(n124), .C(n1747), .D(n99), .Y(N12505) );
  OAI22X1 U1826 ( .A(n1746), .B(n124), .C(n1745), .D(n99), .Y(N12506) );
  OAI22X1 U1827 ( .A(n1744), .B(n124), .C(n1743), .D(n99), .Y(N12507) );
  OAI22X1 U1828 ( .A(n1742), .B(n124), .C(n1741), .D(n99), .Y(N12508) );
  OAI22X1 U1829 ( .A(n1740), .B(n124), .C(n1739), .D(n99), .Y(N12509) );
  OAI22X1 U1830 ( .A(n1738), .B(n124), .C(n1737), .D(n99), .Y(N12510) );
  OAI22X1 U1831 ( .A(n1736), .B(n1709), .C(n1735), .D(n1708), .Y(N12584) );
  OAI22X1 U1832 ( .A(n304), .B(n1709), .C(n1734), .D(n1708), .Y(N12585) );
  OAI22X1 U1833 ( .A(n1731), .B(n1709), .C(n1730), .D(n1708), .Y(N12587) );
  OAI22X1 U1834 ( .A(n1729), .B(n1709), .C(n1728), .D(n1708), .Y(N12588) );
  OAI22X1 U1835 ( .A(n1727), .B(n1709), .C(n1726), .D(n1708), .Y(N12589) );
  OAI22X1 U1836 ( .A(n1725), .B(n1709), .C(n1998), .D(n1708), .Y(N12590) );
  OAI22X1 U1837 ( .A(n1724), .B(n1709), .C(n1723), .D(n1708), .Y(N12591) );
  OAI22X1 U1838 ( .A(n1750), .B(n119), .C(n1749), .D(n112), .Y(N12513) );
  OAI22X1 U1839 ( .A(n1748), .B(n119), .C(n1747), .D(n112), .Y(N12514) );
  OAI22X1 U1840 ( .A(n1746), .B(n119), .C(n1745), .D(n112), .Y(N12515) );
  OAI22X1 U1841 ( .A(n1744), .B(n119), .C(n1743), .D(n112), .Y(N12516) );
  OAI22X1 U1842 ( .A(n1742), .B(n119), .C(n1741), .D(n112), .Y(N12517) );
  OAI22X1 U1843 ( .A(n1740), .B(n119), .C(n1739), .D(n112), .Y(N12518) );
  OAI22X1 U1844 ( .A(n1738), .B(n119), .C(n1737), .D(n112), .Y(N12519) );
  OAI22X1 U1845 ( .A(n1736), .B(n1712), .C(n1735), .D(n47), .Y(N12593) );
  OAI22X1 U1846 ( .A(n304), .B(n1712), .C(n1734), .D(n1711), .Y(N12594) );
  OAI22X1 U1847 ( .A(n1731), .B(n1712), .C(n1730), .D(n47), .Y(N12596) );
  OAI22X1 U1848 ( .A(n1729), .B(n1712), .C(n1728), .D(n1711), .Y(N12597) );
  OAI22X1 U1849 ( .A(n1727), .B(n1712), .C(n1726), .D(n47), .Y(N12598) );
  OAI22X1 U1850 ( .A(n1725), .B(n1712), .C(n1998), .D(n1711), .Y(N12599) );
  OAI22X1 U1851 ( .A(n1724), .B(n1712), .C(n1723), .D(n47), .Y(N12600) );
  OAI22X1 U1852 ( .A(n1750), .B(n113), .C(n1749), .D(n1711), .Y(N12522) );
  OAI22X1 U1853 ( .A(n1748), .B(n113), .C(n1747), .D(n47), .Y(N12523) );
  OAI22X1 U1854 ( .A(n1746), .B(n113), .C(n1745), .D(n1711), .Y(N12524) );
  OAI22X1 U1855 ( .A(n1744), .B(n113), .C(n1743), .D(n47), .Y(N12525) );
  OAI22X1 U1856 ( .A(n1742), .B(n113), .C(n1741), .D(n1711), .Y(N12526) );
  OAI22X1 U1857 ( .A(n1740), .B(n113), .C(n1739), .D(n47), .Y(N12527) );
  OAI22X1 U1858 ( .A(n1738), .B(n113), .C(n1737), .D(n1711), .Y(N12528) );
  NAND21X1 U1859 ( .B(n2344), .A(n499), .Y(n2188) );
  NAND21X1 U1860 ( .B(n547), .A(n2255), .Y(n2256) );
  NAND32X1 U1861 ( .B(n1506), .C(n506), .A(n2204), .Y(n2203) );
  INVX1 U1862 ( .A(n1513), .Y(n1519) );
  NAND32X1 U1863 ( .B(n2204), .C(n1527), .A(n1522), .Y(n1513) );
  NAND21X1 U1864 ( .B(n2389), .A(n498), .Y(n2268) );
  AO21X1 U1865 ( .B(n2442), .C(n2029), .A(n1355), .Y(N12725) );
  AOI21X1 U1866 ( .B(n1354), .C(n1353), .A(n506), .Y(n1355) );
  OA2222XL U1867 ( .A(n1904), .B(n2032), .C(n1916), .D(n2035), .E(n32), .F(
        n2031), .G(n1897), .H(n2030), .Y(n1354) );
  OA222X1 U1868 ( .A(n1574), .B(n1541), .C(n1909), .D(n2034), .E(n1421), .F(
        n1484), .Y(n1353) );
  AO21X1 U1869 ( .B(n509), .C(n2247), .A(n558), .Y(N12722) );
  NAND43X1 U1870 ( .B(n2246), .C(n2245), .D(n2244), .A(n2243), .Y(n2247) );
  NOR21XL U1871 ( .B(n2143), .A(n2142), .Y(N12912) );
  AOI32XL U1872 ( .A(n2441), .B(n2141), .C(n2140), .D(n502), .E(n2139), .Y(
        n2142) );
  INVX1 U1873 ( .A(n2251), .Y(n2255) );
  NAND43X1 U1874 ( .B(n2250), .C(n2249), .D(n2248), .A(n500), .Y(n2251) );
  INVX1 U1875 ( .A(n1512), .Y(n1521) );
  NAND32X1 U1876 ( .B(n2202), .C(n1527), .A(n2294), .Y(n1512) );
  OAI32X1 U1877 ( .A(n1755), .B(n540), .C(n2359), .D(n1754), .E(n1753), .Y(
        N12694) );
  INVX1 U1878 ( .A(dpc[4]), .Y(n1753) );
  OAI221X1 U1879 ( .A(n1453), .B(n2190), .C(n2189), .D(n1440), .E(n562), .Y(
        N12485) );
  OAI221X1 U1880 ( .A(n1469), .B(n2190), .C(n2189), .D(n1468), .E(n569), .Y(
        N12486) );
  OAI221X1 U1881 ( .A(n1890), .B(n2190), .C(n2189), .D(n1887), .E(n569), .Y(
        N12487) );
  OAI22XL U1882 ( .A(n1848), .B(n2285), .C(n2271), .D(n2188), .Y(N12705) );
  OAI22X1 U1883 ( .A(n1491), .B(n505), .C(n1490), .D(n1489), .Y(N12724) );
  AND3X1 U1884 ( .A(n1488), .B(n1487), .C(n1486), .Y(n1491) );
  OA22X1 U1885 ( .A(n1481), .B(n2030), .C(n1480), .D(n2032), .Y(n1487) );
  OAI22X1 U1886 ( .A(n1465), .B(n503), .C(n1490), .D(n1464), .Y(N12723) );
  AND3X1 U1887 ( .A(n1463), .B(n1462), .C(n1461), .Y(n1465) );
  OAI22XL U1888 ( .A(n1583), .B(n1582), .C(n556), .D(n1595), .Y(n1884) );
  OAI22XL U1889 ( .A(n1112), .B(n505), .C(n66), .D(n1111), .Y(N11487) );
  INVX1 U1890 ( .A(n2310), .Y(n1112) );
  OAI22X1 U1891 ( .A(n1754), .B(n1597), .C(n1755), .D(n2265), .Y(N12695) );
  INVX1 U1892 ( .A(dpc[5]), .Y(n1597) );
  OAI22X1 U1893 ( .A(n1754), .B(n1599), .C(n1755), .D(n2260), .Y(N12693) );
  INVX1 U1894 ( .A(dpc[3]), .Y(n1599) );
  OAI22X1 U1895 ( .A(n554), .B(n2022), .C(n2021), .D(n2020), .Y(N12720) );
  OA2222XL U1896 ( .A(n2019), .B(n2018), .C(n2017), .D(n2016), .E(n2015), .F(
        n2014), .G(n2013), .H(n2012), .Y(n2022) );
  OAI22X1 U1897 ( .A(n555), .B(n1549), .C(n1791), .D(n2020), .Y(N12717) );
  OA2222XL U1898 ( .A(n2019), .B(n1793), .C(n2017), .D(n1550), .E(n52), .F(
        n2014), .G(n1557), .H(n2012), .Y(n1549) );
  OAI22XL U1899 ( .A(n555), .B(n1576), .C(n1575), .D(n2020), .Y(N12716) );
  OA2222XL U1900 ( .A(n2019), .B(n1574), .C(n2017), .D(n1573), .E(n1901), .F(
        n2014), .G(n1909), .H(n2012), .Y(n1576) );
  INVX1 U1901 ( .A(n1836), .Y(n1844) );
  OAI31XL U1902 ( .A(n540), .B(n2266), .C(n2265), .D(n569), .Y(N12556) );
  OAI31XL U1903 ( .A(dps[1]), .B(n543), .C(n2256), .D(n563), .Y(N12672) );
  OAI31XL U1904 ( .A(dps[0]), .B(n545), .C(n2252), .D(n565), .Y(N12651) );
  OAI31XL U1905 ( .A(dps[1]), .B(n543), .C(n2252), .D(n566), .Y(N12644) );
  OAI211X1 U1906 ( .C(n506), .D(n2204), .A(n2203), .B(n567), .Y(N13324) );
  OAI211X1 U1907 ( .C(n506), .D(n2202), .A(n2201), .B(n567), .Y(N13366) );
  OA2222XL U1908 ( .A(n2019), .B(n1460), .C(n2017), .D(n1855), .E(n40), .F(
        n2014), .G(n1459), .H(n2012), .Y(n1457) );
  INVX1 U1909 ( .A(n2201), .Y(n1530) );
  INVX1 U1910 ( .A(n963), .Y(n2134) );
  AND2X1 U1911 ( .A(n1507), .B(multemp2[2]), .Y(N13325) );
  AND2X1 U1912 ( .A(n1507), .B(multemp2[3]), .Y(N13326) );
  AND2X1 U1913 ( .A(n1507), .B(multemp2[4]), .Y(N13327) );
  AND2X1 U1914 ( .A(n1507), .B(multemp2[5]), .Y(N13328) );
  AND2X1 U1915 ( .A(n1507), .B(multemp2[6]), .Y(N13329) );
  AND2X1 U1916 ( .A(n1507), .B(multemp2[7]), .Y(N13330) );
  AND2X1 U1917 ( .A(n1507), .B(multemp2[8]), .Y(N13331) );
  AND2X1 U1918 ( .A(n1507), .B(multemp2[9]), .Y(N13332) );
  AND2X1 U1919 ( .A(sfroe_comb_s), .B(n501), .Y(N11488) );
  INVX1 U1920 ( .A(n2164), .Y(sfroe_comb_s) );
  AND2X1 U1921 ( .A(n1530), .B(n303), .Y(N13367) );
  OAI22XL U1922 ( .A(n554), .B(n1473), .C(n79), .D(n2020), .Y(N12715) );
  OA2222XL U1923 ( .A(n2019), .B(n1483), .C(n2017), .D(n1476), .E(n48), .F(
        n2014), .G(n1482), .H(n2012), .Y(n1473) );
  AOI211X1 U1924 ( .C(n1417), .D(n1416), .A(n1415), .B(n2359), .Y(N10576) );
  AOI211X1 U1925 ( .C(n1436), .D(n1435), .A(n1434), .B(n504), .Y(N10573) );
  INVX1 U1926 ( .A(n1433), .Y(n1436) );
  AOI31X1 U1927 ( .A(n1397), .B(n1396), .C(n1395), .D(n2359), .Y(N10562) );
  OA21X1 U1928 ( .B(n493), .C(n1409), .A(n1356), .Y(n1397) );
  AO21X1 U1929 ( .B(n1497), .C(n1429), .A(n1357), .Y(n1396) );
  AND3X1 U1930 ( .A(n1541), .B(n1484), .C(n1394), .Y(n1395) );
  INVX1 U1931 ( .A(ramdatai[4]), .Y(n1825) );
  INVX1 U1932 ( .A(pc_i[7]), .Y(n2092) );
  INVX1 U1933 ( .A(ramdatai[3]), .Y(n1793) );
  OA2222XL U1934 ( .A(n1852), .B(n1484), .C(n1460), .D(n1541), .E(n1873), .F(
        n2035), .G(n1459), .H(n2034), .Y(n1461) );
  OA222X1 U1935 ( .A(n2121), .B(n2120), .C(n2119), .D(n2118), .E(n2117), .F(
        n495), .Y(n2122) );
  OAI221X1 U1936 ( .A(n2426), .B(n2425), .C(n296), .D(n2424), .E(n567), .Y(
        n1024) );
  INVX1 U1937 ( .A(n2194), .Y(n1737) );
  INVXL U1938 ( .A(ramdatai[7]), .Y(n2099) );
  INVX1 U1939 ( .A(n1962), .Y(n1557) );
  INVX1 U1940 ( .A(n1983), .Y(n1745) );
  INVX1 U1941 ( .A(n1982), .Y(n1743) );
  INVX1 U1942 ( .A(n1981), .Y(n1741) );
  INVX1 U1943 ( .A(n2025), .Y(n1739) );
  NAND32X1 U1944 ( .B(n555), .C(n2242), .A(n2424), .Y(N12977) );
  GEN2XL U1945 ( .D(mempsack), .E(n2239), .C(n2426), .B(n2238), .A(n2425), .Y(
        n2242) );
  INVX1 U1946 ( .A(n1437), .Y(n2233) );
  INVX1 U1947 ( .A(n2189), .Y(n1452) );
  NAND21X1 U1948 ( .B(n1800), .A(n1799), .Y(n1932) );
  INVX1 U1949 ( .A(n2098), .Y(n1800) );
  MUX2XL U1950 ( .D0(N13350), .D1(n272), .S(N13353), .Y(n1514) );
  MUX2XL U1951 ( .D0(N13346), .D1(divtemp1_0_), .S(N13353), .Y(n1518) );
  MUX2XL U1952 ( .D0(N13348), .D1(n269), .S(N13353), .Y(n1516) );
  MUX2XL U1953 ( .D0(N13351), .D1(n275), .S(N13353), .Y(n1529) );
  MUX2XL U1954 ( .D0(N13349), .D1(n273), .S(N13353), .Y(n1515) );
  MUX2XL U1955 ( .D0(N13347), .D1(n270), .S(N13353), .Y(n1517) );
  INVX1 U1956 ( .A(n1986), .Y(n1757) );
  INVX1 U1957 ( .A(n1985), .Y(n1749) );
  INVX1 U1958 ( .A(n1984), .Y(n1747) );
  NAND21X1 U1959 ( .B(n1600), .A(dpc[0]), .Y(n1661) );
  MUX2X1 U1960 ( .D0(n1227), .D1(n1554), .S(n295), .Y(n1071) );
  AO21X1 U1961 ( .B(n1780), .C(n1779), .A(n1778), .Y(n1922) );
  AO21X1 U1962 ( .B(n1693), .C(n1650), .A(n1661), .Y(n1637) );
  AO21X1 U1963 ( .B(n1693), .C(n1619), .A(n1661), .Y(n1620) );
  AO21X1 U1964 ( .B(n1693), .C(n1689), .A(n1661), .Y(n1692) );
  INVX1 U1965 ( .A(pc_i[15]), .Y(n2090) );
  INVX1 U1966 ( .A(pc_i[13]), .Y(n1787) );
  INVX1 U1967 ( .A(pc_i[14]), .Y(n2009) );
  INVX1 U1968 ( .A(n1988), .Y(n1726) );
  INVX1 U1969 ( .A(n2049), .Y(n1723) );
  MUX2IX1 U1970 ( .D0(n1810), .D1(n1809), .S(n295), .Y(n255) );
  MUX2IX1 U1971 ( .D0(n1777), .D1(n1776), .S(n295), .Y(n256) );
  INVX1 U1972 ( .A(n1912), .Y(n1068) );
  AOI211X1 U1973 ( .C(n1913), .D(n2068), .A(n1923), .B(n1912), .Y(n1915) );
  INVX1 U1974 ( .A(pc_i[10]), .Y(n1916) );
  INVX1 U1975 ( .A(pc_i[12]), .Y(n1817) );
  INVX1 U1976 ( .A(n1991), .Y(n1732) );
  INVX1 U1977 ( .A(n1911), .Y(n1923) );
  NAND21X1 U1978 ( .B(n1910), .A(n1929), .Y(n1911) );
  NAND32X1 U1979 ( .B(dpc[2]), .C(n1661), .A(n1603), .Y(n1704) );
  NAND21X1 U1980 ( .B(n1999), .A(n152), .Y(n1722) );
  NOR8XL U1981 ( .A(multemp2[8]), .B(multemp2[9]), .C(multemp2[6]), .D(
        multemp2[7]), .E(multemp2[4]), .F(multemp2[5]), .G(multemp2[2]), .H(
        multemp2[3]), .Y(n2306) );
  MUX2X1 U1982 ( .D0(n1656), .D1(n1700), .S(n1903), .Y(n1651) );
  NAND21X1 U1983 ( .B(n1619), .A(n135), .Y(n1635) );
  NAND21X1 U1984 ( .B(n1689), .A(n135), .Y(n1617) );
  INVX1 U1985 ( .A(pc_i[8]), .Y(n1873) );
  AO21X1 U1986 ( .B(n135), .C(n1854), .A(n1662), .Y(n1658) );
  INVX1 U1987 ( .A(n1994), .Y(n1735) );
  INVX1 U1988 ( .A(n1992), .Y(n1734) );
  NAND21X1 U1989 ( .B(n1650), .A(n135), .Y(n1639) );
  INVX1 U1990 ( .A(n1510), .Y(n1525) );
  NAND43X1 U1991 ( .B(n2297), .C(n236), .D(n2295), .A(n1509), .Y(n1510) );
  AOI221XL U1992 ( .A(n2294), .B(n2202), .C(n1522), .D(n2204), .E(n2299), .Y(
        n1509) );
  INVX1 U1993 ( .A(n1655), .Y(n1733) );
  OAI211X1 U1994 ( .C(n1654), .D(n32), .A(n1653), .B(n1652), .Y(n1655) );
  AO21X1 U1995 ( .B(n1650), .C(n1649), .A(n1701), .Y(n1653) );
  OA21X1 U1996 ( .B(n1905), .C(n1704), .A(n1651), .Y(n1652) );
  INVX1 U1997 ( .A(n1657), .Y(n1654) );
  INVX1 U1998 ( .A(n2173), .Y(n2129) );
  OA2222XL U1999 ( .A(n1485), .B(n1484), .C(n1483), .D(n1541), .E(n1686), .F(
        n2035), .G(n1482), .H(n2034), .Y(n1486) );
  INVX1 U2000 ( .A(pc_i[6]), .Y(n1940) );
  INVX1 U2001 ( .A(dpc[1]), .Y(n1603) );
  INVX1 U2002 ( .A(n1641), .Y(n1602) );
  INVX1 U2003 ( .A(n1696), .Y(n1690) );
  INVX1 U2004 ( .A(n1631), .Y(n1640) );
  INVX1 U2005 ( .A(n1613), .Y(n1622) );
  OR2X1 U2006 ( .A(n2243), .B(n2245), .Y(n2014) );
  NAND43X1 U2007 ( .B(n975), .C(n1346), .D(n974), .A(n1446), .Y(n1014) );
  AOI31X1 U2008 ( .A(n965), .B(n964), .C(n2361), .D(n492), .Y(n975) );
  INVX1 U2009 ( .A(n1287), .Y(n972) );
  NAND43X1 U2010 ( .B(n1349), .C(n1351), .D(n1352), .A(n1348), .Y(n2032) );
  INVX1 U2011 ( .A(n1350), .Y(n1348) );
  INVX1 U2012 ( .A(n2035), .Y(n1349) );
  NAND32X1 U2013 ( .B(n44), .C(n34), .A(n1623), .Y(n1612) );
  NAND32X1 U2014 ( .B(n1352), .C(n1351), .A(n1350), .Y(n2030) );
  NAND5XL U2015 ( .A(n2086), .B(n1484), .C(n1541), .D(n1490), .E(n2034), .Y(
        n1351) );
  INVX1 U2016 ( .A(dpc[2]), .Y(n1604) );
  OR2X1 U2017 ( .A(n54), .B(n1649), .Y(n1630) );
  NAND6XL U2018 ( .A(n1411), .B(n1495), .C(n1399), .D(n1377), .E(n1400), .F(
        n1376), .Y(n1390) );
  AO21X1 U2019 ( .B(n1386), .C(n1435), .A(n1434), .Y(n1377) );
  NOR5X1 U2020 ( .A(n1405), .B(n1430), .C(n1375), .D(n1374), .E(n1373), .Y(
        n1376) );
  INVX1 U2021 ( .A(n1428), .Y(n1375) );
  NAND32X1 U2022 ( .B(n1352), .C(n1014), .A(n2244), .Y(n2012) );
  NAND21X1 U2023 ( .B(n153), .A(n540), .Y(n2259) );
  NAND21XL U2024 ( .B(n152), .A(n539), .Y(n2262) );
  NAND21X1 U2025 ( .B(n726), .A(n2125), .Y(n2270) );
  NAND32X1 U2026 ( .B(n50), .C(n36), .A(n1691), .Y(n2200) );
  INVX1 U2027 ( .A(pc_i[11]), .Y(n1677) );
  INVX1 U2028 ( .A(n2019), .Y(n1016) );
  INVX1 U2029 ( .A(n1352), .Y(n2243) );
  AND2X1 U2030 ( .A(n1334), .B(n129), .Y(n1336) );
  INVX1 U2031 ( .A(n1600), .Y(n1755) );
  NOR2X1 U2032 ( .A(n40), .B(n2200), .Y(n257) );
  INVX1 U2033 ( .A(n2182), .Y(n2374) );
  NAND21X1 U2034 ( .B(n2181), .A(n2180), .Y(n2182) );
  INVX1 U2035 ( .A(n2172), .Y(n2372) );
  INVX1 U2036 ( .A(n966), .Y(n1346) );
  NAND21X1 U2037 ( .B(n2118), .A(n1467), .Y(n966) );
  NAND21X1 U2038 ( .B(n111), .A(n1888), .Y(n2035) );
  NAND32X1 U2039 ( .B(n1361), .C(n1360), .A(n1359), .Y(n1495) );
  INVX1 U2040 ( .A(pc_i[9]), .Y(n1686) );
  AO21X1 U2041 ( .B(n240), .C(n1402), .A(n1381), .Y(n1389) );
  INVX1 U2042 ( .A(n152), .Y(n1714) );
  OAI222XL U2043 ( .A(n1392), .B(n1403), .C(n1416), .D(n1415), .E(n1386), .F(
        n1385), .Y(n1388) );
  INVX1 U2044 ( .A(n1337), .Y(n1341) );
  INVX1 U2045 ( .A(n1368), .Y(n1405) );
  NAND43X1 U2046 ( .B(n1367), .C(n1366), .D(n477), .A(n1432), .Y(n1368) );
  NAND21X1 U2047 ( .B(n554), .A(n1947), .Y(n2186) );
  OR2X1 U2048 ( .A(n554), .B(n1947), .Y(n2185) );
  INVX1 U2049 ( .A(n1385), .Y(n1413) );
  INVX1 U2050 ( .A(n1490), .Y(n2029) );
  OAI22X1 U2051 ( .A(n2184), .B(n2186), .C(n2339), .D(n2185), .Y(N12970) );
  OAI22X1 U2052 ( .A(n2183), .B(n2186), .C(n2342), .D(n2185), .Y(N12971) );
  OAI22X1 U2053 ( .A(n2187), .B(n2186), .C(n2336), .D(n2185), .Y(N12969) );
  OAI22X1 U2054 ( .A(n2179), .B(n2186), .C(n2178), .D(n2185), .Y(N12965) );
  OAI22X1 U2055 ( .A(n2177), .B(n2186), .C(n2176), .D(n2185), .Y(N12966) );
  OAI22X1 U2056 ( .A(n2175), .B(n2186), .C(n2333), .D(n2185), .Y(N12967) );
  INVX1 U2057 ( .A(n2095), .Y(n1606) );
  INVX1 U2058 ( .A(n1642), .Y(n1643) );
  INVX1 U2059 ( .A(n1790), .Y(n1625) );
  INVX1 U2060 ( .A(n2237), .Y(n2425) );
  NAND21X1 U2061 ( .B(n2241), .A(n296), .Y(n2237) );
  NAND21X1 U2062 ( .B(n1434), .A(n1492), .Y(n1497) );
  OR3XL U2063 ( .A(n2207), .B(n2250), .C(n1511), .Y(n1526) );
  INVX1 U2064 ( .A(n2235), .Y(n2426) );
  INVX1 U2065 ( .A(n2236), .Y(n2241) );
  INVX1 U2066 ( .A(n2253), .Y(n2258) );
  NAND21X1 U2067 ( .B(n545), .A(dps[0]), .Y(n2253) );
  INVX1 U2068 ( .A(n2210), .Y(n2228) );
  MUX2X2 U2069 ( .D0(memrd), .D1(n2373), .S(n550), .Y(memrd_comb) );
  MUX2XL U2070 ( .D0(n1004), .D1(n2344), .S(n1142), .Y(n1005) );
  OAI22XL U2071 ( .A(n1167), .B(n1227), .C(n1569), .D(n1921), .Y(n1007) );
  MUX2XL U2072 ( .D0(n1168), .D1(n982), .S(acc[7]), .Y(n1008) );
  NAND21X1 U2073 ( .B(n1762), .A(n1761), .Y(n2412) );
  AO2222XL U2074 ( .A(n1996), .B(temp2_comb[5]), .C(alu_out[5]), .D(n2192), 
        .E(n1988), .F(n2193), .G(memdatai[5]), .H(n1760), .Y(n1762) );
  AOI21X1 U2075 ( .B(n2327), .C(n2311), .A(n2310), .Y(n259) );
  INVX1 U2076 ( .A(n1214), .Y(n1216) );
  XOR2X1 U2077 ( .A(n742), .B(n1036), .Y(n924) );
  OAI31XL U2078 ( .A(n2324), .B(instr[3]), .C(n2323), .D(n2322), .Y(n2325) );
  OA222X1 U2079 ( .A(n2321), .B(n2320), .C(n2319), .D(n2318), .E(n2317), .F(
        n129), .Y(n2324) );
  AOI221XL U2080 ( .A(instr[2]), .B(n103), .C(n2314), .D(n2313), .E(n2312), 
        .Y(n2317) );
  MAJ3X1 U2081 ( .A(n262), .B(n263), .C(n9), .Y(n261) );
  XNOR2XL U2082 ( .A(acc[6]), .B(n996), .Y(n263) );
  NAND21X1 U2083 ( .B(n2004), .A(n2003), .Y(n2413) );
  OA2222XL U2084 ( .A(n2002), .B(n2001), .C(n2000), .D(n2018), .E(n2053), .F(
        n2016), .G(n1999), .H(n1998), .Y(n2003) );
  AO2222XL U2085 ( .A(pc_i[6]), .B(n1997), .C(alu_out[6]), .D(n114), .E(n1996), 
        .F(temp2_comb[6]), .G(pc_o[6]), .H(n1995), .Y(n2004) );
  INVXL U2086 ( .A(n2051), .Y(n1997) );
  AOI222XL U2087 ( .A(multemp2[1]), .B(n1522), .C(temp2_comb[7]), .D(n1001), 
        .E(n1000), .F(n999), .Y(n1002) );
  NAND21X1 U2088 ( .B(n984), .A(n983), .Y(n1001) );
  AOI222XL U2089 ( .A(n1209), .B(n1208), .C(c), .D(n1207), .E(n2299), .F(n1206), .Y(n1210) );
  GEN3XL U2090 ( .F(dec_cop[4]), .G(c), .E(n1205), .D(n1204), .C(n1203), .B(
        n1202), .A(n1201), .Y(n1206) );
  AO21XL U2091 ( .B(temp2_comb[1]), .C(n997), .A(n985), .Y(n987) );
  INVX1 U2092 ( .A(dec_accop[7]), .Y(n739) );
  NOR21X2 U2093 ( .B(waitstaten), .A(n2392), .Y(n2401) );
  INVXL U2094 ( .A(n2388), .Y(waitstaten) );
  NOR43XL U2095 ( .B(n2391), .C(n2390), .D(stop), .A(n2389), .Y(n2392) );
  MUX2X1 U2096 ( .D0(n320), .D1(n319), .S(N351), .Y(dpl[0]) );
  MUX4X1 U2097 ( .D0(dpl_reg[0]), .D1(dpl_reg[8]), .D2(dpl_reg[16]), .D3(
        dpl_reg[24]), .S0(n355), .S1(n351), .Y(n320) );
  MUX4X1 U2098 ( .D0(dpl_reg[32]), .D1(dpl_reg[40]), .D2(dpl_reg[48]), .D3(
        dpl_reg[56]), .S0(n355), .S1(n351), .Y(n319) );
  AO21XL U2099 ( .B(temp2_comb[2]), .C(n997), .A(n985), .Y(n1117) );
  NAND21X1 U2100 ( .B(n2458), .A(n1898), .Y(n989) );
  MUX2XL U2101 ( .D0(N13338), .D1(divtempreg[1]), .S(N13343), .Y(n269) );
  XNOR2XL U2102 ( .A(n1036), .B(acc[2]), .Y(n271) );
  MUX2X1 U2103 ( .D0(memaddr[4]), .D1(n1989), .S(n1993), .Y(N12845) );
  MUX2X1 U2104 ( .D0(memaddr[5]), .D1(n1988), .S(n1993), .Y(N12846) );
  NAND43X1 U2105 ( .B(n1044), .C(n1043), .D(n1042), .A(n1041), .Y(n1933) );
  OAI22XL U2106 ( .A(n1898), .B(n1167), .C(n1569), .D(n1777), .Y(n1043) );
  AO21XL U2107 ( .B(ramdatao[6]), .C(n1142), .A(n1022), .Y(n1044) );
  AND2XL U2108 ( .A(sfrwe_r), .B(n551), .Y(sfrwe) );
  MUX2X1 U2109 ( .D0(memaddr[6]), .D1(n1987), .S(n1993), .Y(N12847) );
  MUX2XL U2110 ( .D0(n1933), .D1(temp[6]), .S(n1978), .Y(N12830) );
  AO21XL U2111 ( .B(temp2_comb[3]), .C(n997), .A(n992), .Y(n1048) );
  OAI31XL U2112 ( .A(n1979), .B(N13353), .C(n1978), .D(n1977), .Y(N12824) );
  OAI22X1 U2113 ( .A(n1976), .B(n1975), .C(temp[0]), .D(n1974), .Y(n1977) );
  NAND5XL U2114 ( .A(n1974), .B(n1968), .C(n1967), .D(n1966), .E(n1965), .Y(
        n1976) );
  NAND5XL U2115 ( .A(n1973), .B(n1972), .C(n1971), .D(n1970), .E(n1969), .Y(
        n1975) );
  MUX2XL U2116 ( .D0(N13340), .D1(divtempreg[3]), .S(N13343), .Y(n272) );
  MUX2XL U2117 ( .D0(N13339), .D1(divtempreg[2]), .S(N13343), .Y(n273) );
  XNOR2XL U2118 ( .A(n1036), .B(acc[3]), .Y(n274) );
  OAI221X1 U2119 ( .A(n237), .B(n2060), .C(n1150), .D(n1040), .E(n1039), .Y(
        n1042) );
  AO21XL U2120 ( .B(n1038), .C(n1173), .A(n2007), .Y(n1039) );
  XOR3X1 U2121 ( .A(n1037), .B(n291), .C(n9), .Y(n1040) );
  MUX2XL U2122 ( .D0(n1174), .D1(n1171), .S(acc[6]), .Y(n1038) );
  AO222X1 U2123 ( .A(n1666), .B(temp[1]), .C(dptr_inc[1]), .D(n1683), .E(n1665), .F(n8), .Y(n1992) );
  NAND43X1 U2124 ( .B(n1154), .C(n1153), .D(n1152), .A(n1151), .Y(n1960) );
  OAI22XL U2125 ( .A(n1225), .B(n1167), .C(n1569), .D(n1810), .Y(n1153) );
  AO21XL U2126 ( .B(ramdatao[5]), .C(n1142), .A(n1141), .Y(n1154) );
  AO21XL U2127 ( .B(temp2_comb[4]), .C(n997), .A(n992), .Y(n1029) );
  XOR2XL U2128 ( .A(n1036), .B(acc[4]), .Y(n1031) );
  OAI221X1 U2129 ( .A(n1588), .B(n1595), .C(n1594), .D(n1587), .E(n1586), .Y(
        N347) );
  MUX2X1 U2130 ( .D0(n1585), .D1(n1584), .S(n1598), .Y(n1586) );
  NAND21X1 U2131 ( .B(n1589), .A(ramdatao[1]), .Y(n1584) );
  OAI221X1 U2132 ( .A(n1150), .B(n1149), .C(n237), .D(n1921), .E(n1148), .Y(
        n1152) );
  AO21XL U2133 ( .B(n1147), .C(n1173), .A(n1789), .Y(n1148) );
  MUX2XL U2134 ( .D0(n1174), .D1(n1171), .S(acc[5]), .Y(n1147) );
  MUX2XL U2135 ( .D0(N13341), .D1(divtempreg[4]), .S(N13343), .Y(n275) );
  MUX4XL U2136 ( .D0(dpl_reg[0]), .D1(dpl_reg[8]), .D2(dpl_reg[16]), .D3(
        dpl_reg[24]), .S0(n391), .S1(n395), .Y(n375) );
  AO222X1 U2137 ( .A(n1666), .B(temp[3]), .C(dptr_inc[3]), .D(n1683), .E(n1665), .F(n13), .Y(n1990) );
  AO222X1 U2138 ( .A(n1666), .B(temp[2]), .C(dptr_inc[2]), .D(n1683), .E(n1665), .F(n10), .Y(n1991) );
  AO222XL U2139 ( .A(n1666), .B(temp[0]), .C(dptr_inc[0]), .D(n1683), .E(n1665), .F(n11), .Y(n1994) );
  MUX4XL U2140 ( .D0(dpl_reg[33]), .D1(dpl_reg[41]), .D2(dpl_reg[49]), .D3(
        dpl_reg[57]), .S0(n391), .S1(n395), .Y(n376) );
  MUX4XL U2141 ( .D0(dpl_reg[34]), .D1(dpl_reg[42]), .D2(dpl_reg[50]), .D3(
        dpl_reg[58]), .S0(n391), .S1(n395), .Y(n378) );
  MUX4X1 U2142 ( .D0(dpl_reg[35]), .D1(dpl_reg[43]), .D2(dpl_reg[51]), .D3(
        dpl_reg[59]), .S0(n392), .S1(n396), .Y(n380) );
  NAND43X1 U2143 ( .B(n1138), .C(n1137), .D(n1136), .A(n1135), .Y(n1961) );
  OAI22XL U2144 ( .A(n1167), .B(n1226), .C(n1569), .D(n1227), .Y(n1137) );
  OAI22XL U2145 ( .A(n1898), .B(n1979), .C(n2305), .D(n1921), .Y(n1136) );
  AO21XL U2146 ( .B(ramdatao[4]), .C(n1142), .A(n1129), .Y(n1138) );
  AO21XL U2147 ( .B(n994), .C(n993), .A(n992), .Y(n1026) );
  NAND32XL U2148 ( .B(n991), .C(c), .A(n990), .Y(n993) );
  AO21X1 U2149 ( .B(n1921), .C(n1777), .A(n2060), .Y(n990) );
  AND4XL U2150 ( .A(acc[3]), .B(acc[4]), .C(acc[7]), .D(n989), .Y(n991) );
  XOR2XL U2151 ( .A(n1036), .B(acc[5]), .Y(n1032) );
  OA222X1 U2152 ( .A(n237), .B(n1777), .C(n1134), .D(n1819), .E(n1150), .F(
        n1133), .Y(n1135) );
  OA21XL U2153 ( .B(acc[4]), .C(n1174), .A(n1173), .Y(n1134) );
  XOR3XL U2154 ( .A(n1132), .B(n1131), .C(n1130), .Y(n1133) );
  MUX2X1 U2155 ( .D0(pc_o[3]), .D1(n1990), .S(n1993), .Y(N12844) );
  AO21XL U2156 ( .B(temp2_comb[5]), .C(n997), .A(n1026), .Y(n1144) );
  NAND21XL U2157 ( .B(n1598), .A(dps[3]), .Y(n1595) );
  INVXL U2158 ( .A(ramsfraddr[0]), .Y(n2209) );
  MUX2XL U2159 ( .D0(N13342), .D1(divtempreg[5]), .S(N13343), .Y(n276) );
  MUX4XL U2160 ( .D0(dpl_reg[1]), .D1(dpl_reg[9]), .D2(dpl_reg[17]), .D3(
        dpl_reg[25]), .S0(n391), .S1(n395), .Y(n377) );
  MUX4XL U2161 ( .D0(dpl_reg[2]), .D1(dpl_reg[10]), .D2(dpl_reg[18]), .D3(
        dpl_reg[26]), .S0(n391), .S1(n395), .Y(n379) );
  MUX4XL U2162 ( .D0(dpl_reg[3]), .D1(dpl_reg[11]), .D2(dpl_reg[19]), .D3(
        dpl_reg[27]), .S0(n392), .S1(n396), .Y(n381) );
  MUX2XL U2163 ( .D0(n1591), .D1(n1590), .S(n1598), .Y(n1592) );
  NAND21XL U2164 ( .B(dps[3]), .A(dps[2]), .Y(n1591) );
  NAND21XL U2165 ( .B(n1589), .A(ramdatao[2]), .Y(n1590) );
  MUX4X1 U2166 ( .D0(ramdatao[3]), .D1(ramdatao[7]), .D2(ckcon[3]), .D3(
        ckcon[7]), .S0(n2171), .S1(n277), .Y(n786) );
  NAND4XL U2167 ( .A(ramsfraddr[3]), .B(n1580), .C(n2227), .D(n2218), .Y(n277)
         );
  NOR43XL U2168 ( .B(n2120), .C(n957), .D(n1357), .A(phase[5]), .Y(n958) );
  NAND21X1 U2169 ( .B(n2453), .A(n842), .Y(n1379) );
  NAND21X1 U2170 ( .B(n2451), .A(n708), .Y(n1371) );
  NAND21X1 U2171 ( .B(n900), .A(N343), .Y(n1228) );
  NAND21X1 U2172 ( .B(N343), .A(n900), .Y(n1868) );
  AO222X1 U2173 ( .A(n1666), .B(temp[5]), .C(dptr_inc[5]), .D(n1683), .E(n1665), .F(n14), .Y(n1988) );
  AO222X1 U2174 ( .A(n1666), .B(temp[4]), .C(dptr_inc[4]), .D(n1683), .E(n1665), .F(n12), .Y(n1989) );
  NAND43X1 U2175 ( .B(n1392), .C(n2156), .D(n493), .A(interrupt), .Y(n1258) );
  AO222X1 U2176 ( .A(n1666), .B(temp[6]), .C(dptr_inc[6]), .D(n1683), .E(n1665), .F(n15), .Y(n1987) );
  MUX2AXL U2177 ( .D0(sp[1]), .D1(n2176), .S(n235), .Y(n613) );
  NAND21X1 U2178 ( .B(n2455), .A(n703), .Y(n1367) );
  NAND21XL U2179 ( .B(n758), .A(dec_accop[18]), .Y(n1179) );
  AO2222XL U2180 ( .A(temp[7]), .B(n659), .C(n658), .D(ramsfraddr[7]), .E(
        n2103), .F(n657), .G(n656), .H(n2047), .Y(n2140) );
  NAND21X1 U2181 ( .B(n155), .A(dec_accop[13]), .Y(n759) );
  MUX4X1 U2182 ( .D0(rn_reg[89]), .D1(rn_reg[81]), .D2(rn_reg[73]), .D3(
        rn_reg[65]), .S0(n478), .S1(n485), .Y(n409) );
  MUX4X1 U2183 ( .D0(rn_reg[217]), .D1(rn_reg[209]), .D2(rn_reg[201]), .D3(
        rn_reg[193]), .S0(n479), .S1(n486), .Y(n414) );
  MUX4XL U2184 ( .D0(rn_reg[216]), .D1(rn_reg[208]), .D2(rn_reg[200]), .D3(
        rn_reg[192]), .S0(n478), .S1(n485), .Y(n404) );
  MUX4XL U2185 ( .D0(rn_reg[92]), .D1(rn_reg[84]), .D2(rn_reg[76]), .D3(
        rn_reg[68]), .S0(n481), .S1(n488), .Y(n439) );
  MUX4XL U2186 ( .D0(rn_reg[220]), .D1(rn_reg[212]), .D2(rn_reg[204]), .D3(
        rn_reg[196]), .S0(n481), .S1(n488), .Y(n444) );
  MUX4XL U2187 ( .D0(rn_reg[91]), .D1(rn_reg[83]), .D2(rn_reg[75]), .D3(
        rn_reg[67]), .S0(n480), .S1(n487), .Y(n429) );
  MUX4XL U2188 ( .D0(rn_reg[219]), .D1(rn_reg[211]), .D2(rn_reg[203]), .D3(
        rn_reg[195]), .S0(n480), .S1(n487), .Y(n434) );
  MUX4X1 U2189 ( .D0(rn_reg[223]), .D1(rn_reg[215]), .D2(rn_reg[207]), .D3(
        rn_reg[199]), .S0(instr[0]), .S1(N353), .Y(n474) );
  MUX4X1 U2190 ( .D0(rn_reg[95]), .D1(rn_reg[87]), .D2(rn_reg[79]), .D3(
        rn_reg[71]), .S0(instr[0]), .S1(N353), .Y(n469) );
  MUX4XL U2191 ( .D0(rn_reg[93]), .D1(rn_reg[85]), .D2(rn_reg[77]), .D3(
        rn_reg[69]), .S0(n481), .S1(n488), .Y(n449) );
  MUX4X1 U2192 ( .D0(rn_reg[221]), .D1(rn_reg[213]), .D2(rn_reg[205]), .D3(
        rn_reg[197]), .S0(n482), .S1(n489), .Y(n454) );
  MUX4XL U2193 ( .D0(rn_reg[90]), .D1(rn_reg[82]), .D2(rn_reg[74]), .D3(
        rn_reg[66]), .S0(n479), .S1(n486), .Y(n419) );
  MUX4XL U2194 ( .D0(rn_reg[218]), .D1(rn_reg[210]), .D2(rn_reg[202]), .D3(
        rn_reg[194]), .S0(n479), .S1(n486), .Y(n424) );
  MUX4XL U2195 ( .D0(rn_reg[88]), .D1(rn_reg[80]), .D2(rn_reg[72]), .D3(
        rn_reg[64]), .S0(N352), .S1(n484), .Y(n399) );
  MUX4XL U2196 ( .D0(rn_reg[57]), .D1(rn_reg[49]), .D2(rn_reg[41]), .D3(
        rn_reg[33]), .S0(n478), .S1(n485), .Y(n408) );
  MUX4XL U2197 ( .D0(rn_reg[185]), .D1(rn_reg[177]), .D2(rn_reg[169]), .D3(
        rn_reg[161]), .S0(n478), .S1(n485), .Y(n413) );
  MUX4XL U2198 ( .D0(rn_reg[184]), .D1(rn_reg[176]), .D2(rn_reg[168]), .D3(
        rn_reg[160]), .S0(n478), .S1(n485), .Y(n403) );
  MUX4XL U2199 ( .D0(rn_reg[60]), .D1(rn_reg[52]), .D2(rn_reg[44]), .D3(
        rn_reg[36]), .S0(n480), .S1(n487), .Y(n438) );
  MUX4XL U2200 ( .D0(rn_reg[188]), .D1(rn_reg[180]), .D2(rn_reg[172]), .D3(
        rn_reg[164]), .S0(n481), .S1(n488), .Y(n443) );
  MUX4XL U2201 ( .D0(rn_reg[59]), .D1(rn_reg[51]), .D2(rn_reg[43]), .D3(
        rn_reg[35]), .S0(n480), .S1(n487), .Y(n428) );
  MUX4XL U2202 ( .D0(rn_reg[187]), .D1(rn_reg[179]), .D2(rn_reg[171]), .D3(
        rn_reg[163]), .S0(n480), .S1(n487), .Y(n433) );
  MUX4X1 U2203 ( .D0(rn_reg[191]), .D1(rn_reg[183]), .D2(rn_reg[175]), .D3(
        rn_reg[167]), .S0(instr[0]), .S1(n484), .Y(n473) );
  MUX4XL U2204 ( .D0(rn_reg[63]), .D1(rn_reg[55]), .D2(rn_reg[47]), .D3(
        rn_reg[39]), .S0(instr[0]), .S1(n484), .Y(n468) );
  MUX4XL U2205 ( .D0(rn_reg[61]), .D1(rn_reg[53]), .D2(rn_reg[45]), .D3(
        rn_reg[37]), .S0(n481), .S1(n488), .Y(n448) );
  MUX4X1 U2206 ( .D0(rn_reg[189]), .D1(rn_reg[181]), .D2(rn_reg[173]), .D3(
        rn_reg[165]), .S0(n482), .S1(n489), .Y(n453) );
  MUX4XL U2207 ( .D0(rn_reg[58]), .D1(rn_reg[50]), .D2(rn_reg[42]), .D3(
        rn_reg[34]), .S0(n479), .S1(n486), .Y(n418) );
  MUX4XL U2208 ( .D0(rn_reg[186]), .D1(rn_reg[178]), .D2(rn_reg[170]), .D3(
        rn_reg[162]), .S0(n479), .S1(n486), .Y(n423) );
  MUX4XL U2209 ( .D0(rn_reg[56]), .D1(rn_reg[48]), .D2(rn_reg[40]), .D3(
        rn_reg[32]), .S0(N352), .S1(n484), .Y(n398) );
  MUX4XL U2210 ( .D0(rn_reg[121]), .D1(rn_reg[113]), .D2(rn_reg[105]), .D3(
        rn_reg[97]), .S0(n478), .S1(n485), .Y(n410) );
  MUX4XL U2211 ( .D0(rn_reg[249]), .D1(rn_reg[241]), .D2(rn_reg[233]), .D3(
        rn_reg[225]), .S0(n479), .S1(n486), .Y(n415) );
  MUX4XL U2212 ( .D0(rn_reg[248]), .D1(rn_reg[240]), .D2(rn_reg[232]), .D3(
        rn_reg[224]), .S0(n478), .S1(n485), .Y(n405) );
  MUX4XL U2213 ( .D0(rn_reg[124]), .D1(rn_reg[116]), .D2(rn_reg[108]), .D3(
        rn_reg[100]), .S0(n481), .S1(n488), .Y(n440) );
  MUX4XL U2214 ( .D0(rn_reg[252]), .D1(rn_reg[244]), .D2(rn_reg[236]), .D3(
        rn_reg[228]), .S0(n481), .S1(n488), .Y(n445) );
  MUX4XL U2215 ( .D0(rn_reg[123]), .D1(rn_reg[115]), .D2(rn_reg[107]), .D3(
        rn_reg[99]), .S0(n480), .S1(n487), .Y(n430) );
  MUX4XL U2216 ( .D0(rn_reg[251]), .D1(rn_reg[243]), .D2(rn_reg[235]), .D3(
        rn_reg[227]), .S0(n480), .S1(n487), .Y(n435) );
  MUX4XL U2217 ( .D0(rn_reg[255]), .D1(rn_reg[247]), .D2(rn_reg[239]), .D3(
        rn_reg[231]), .S0(instr[0]), .S1(n484), .Y(n475) );
  MUX4XL U2218 ( .D0(rn_reg[127]), .D1(rn_reg[119]), .D2(rn_reg[111]), .D3(
        rn_reg[103]), .S0(instr[0]), .S1(n484), .Y(n470) );
  MUX4XL U2219 ( .D0(rn_reg[125]), .D1(rn_reg[117]), .D2(rn_reg[109]), .D3(
        rn_reg[101]), .S0(n481), .S1(n488), .Y(n450) );
  MUX4X1 U2220 ( .D0(rn_reg[253]), .D1(rn_reg[245]), .D2(rn_reg[237]), .D3(
        rn_reg[229]), .S0(n482), .S1(n489), .Y(n455) );
  MUX4XL U2221 ( .D0(rn_reg[122]), .D1(rn_reg[114]), .D2(rn_reg[106]), .D3(
        rn_reg[98]), .S0(n479), .S1(n486), .Y(n420) );
  MUX4XL U2222 ( .D0(rn_reg[250]), .D1(rn_reg[242]), .D2(rn_reg[234]), .D3(
        rn_reg[226]), .S0(n479), .S1(n486), .Y(n425) );
  MUX4XL U2223 ( .D0(rn_reg[120]), .D1(rn_reg[112]), .D2(rn_reg[104]), .D3(
        rn_reg[96]), .S0(N352), .S1(n484), .Y(n400) );
  MUX4XL U2224 ( .D0(dpl_reg[36]), .D1(dpl_reg[44]), .D2(dpl_reg[52]), .D3(
        dpl_reg[60]), .S0(n392), .S1(n396), .Y(n382) );
  MUX4XL U2225 ( .D0(dpl_reg[37]), .D1(dpl_reg[45]), .D2(dpl_reg[53]), .D3(
        dpl_reg[61]), .S0(n392), .S1(n396), .Y(n384) );
  MUX4XL U2226 ( .D0(rn_reg[25]), .D1(rn_reg[17]), .D2(rn_reg[9]), .D3(
        rn_reg[1]), .S0(n478), .S1(n485), .Y(n407) );
  MUX4XL U2227 ( .D0(rn_reg[153]), .D1(rn_reg[145]), .D2(rn_reg[137]), .D3(
        rn_reg[129]), .S0(n478), .S1(n485), .Y(n412) );
  MUX4XL U2228 ( .D0(rn_reg[152]), .D1(rn_reg[144]), .D2(rn_reg[136]), .D3(
        rn_reg[128]), .S0(n478), .S1(n485), .Y(n402) );
  MUX4XL U2229 ( .D0(rn_reg[28]), .D1(rn_reg[20]), .D2(rn_reg[12]), .D3(
        rn_reg[4]), .S0(n480), .S1(n487), .Y(n437) );
  MUX4XL U2230 ( .D0(rn_reg[156]), .D1(rn_reg[148]), .D2(rn_reg[140]), .D3(
        rn_reg[132]), .S0(n481), .S1(n488), .Y(n442) );
  MUX4XL U2231 ( .D0(rn_reg[27]), .D1(rn_reg[19]), .D2(rn_reg[11]), .D3(
        rn_reg[3]), .S0(n480), .S1(n487), .Y(n427) );
  MUX4XL U2232 ( .D0(rn_reg[155]), .D1(rn_reg[147]), .D2(rn_reg[139]), .D3(
        rn_reg[131]), .S0(n480), .S1(n487), .Y(n432) );
  MUX4XL U2233 ( .D0(rn_reg[159]), .D1(rn_reg[151]), .D2(rn_reg[143]), .D3(
        rn_reg[135]), .S0(instr[0]), .S1(n484), .Y(n472) );
  MUX4XL U2234 ( .D0(rn_reg[31]), .D1(rn_reg[23]), .D2(rn_reg[15]), .D3(
        rn_reg[7]), .S0(instr[0]), .S1(n484), .Y(n467) );
  MUX4XL U2235 ( .D0(rn_reg[29]), .D1(rn_reg[21]), .D2(rn_reg[13]), .D3(
        rn_reg[5]), .S0(n481), .S1(n488), .Y(n447) );
  MUX4X1 U2236 ( .D0(rn_reg[157]), .D1(rn_reg[149]), .D2(rn_reg[141]), .D3(
        rn_reg[133]), .S0(n482), .S1(n489), .Y(n452) );
  MUX4XL U2237 ( .D0(rn_reg[26]), .D1(rn_reg[18]), .D2(rn_reg[10]), .D3(
        rn_reg[2]), .S0(n479), .S1(n486), .Y(n417) );
  MUX4XL U2238 ( .D0(rn_reg[154]), .D1(rn_reg[146]), .D2(rn_reg[138]), .D3(
        rn_reg[130]), .S0(n479), .S1(n486), .Y(n422) );
  MUX4XL U2239 ( .D0(rn_reg[24]), .D1(rn_reg[16]), .D2(rn_reg[8]), .D3(
        rn_reg[0]), .S0(N352), .S1(n484), .Y(n397) );
  NAND21X1 U2240 ( .B(n1319), .A(mempsrd), .Y(n1321) );
  NAND21X1 U2241 ( .B(stop_r), .A(n2124), .Y(n1320) );
  OA2222XL U2242 ( .A(n2117), .B(n2163), .C(n1318), .D(n2323), .E(n292), .F(
        n2118), .G(n2119), .H(n2120), .Y(n1319) );
  MUX2X1 U2243 ( .D0(n1187), .D1(n1186), .S(N345), .Y(n1204) );
  AO2222XL U2244 ( .A(n1786), .B(temp[1]), .C(n1816), .D(temp[0]), .E(n1769), 
        .F(temp[2]), .G(n2071), .H(temp[3]), .Y(n1187) );
  AO2222XL U2245 ( .A(n1786), .B(temp[5]), .C(n1816), .D(temp[4]), .E(n1769), 
        .F(temp[6]), .G(n2071), .H(temp[7]), .Y(n1186) );
  NAND21X1 U2246 ( .B(n548), .A(n2457), .Y(n2319) );
  AO2222XL U2247 ( .A(n656), .B(n1763), .C(n1945), .D(n657), .E(temp[5]), .F(
        n659), .G(n658), .H(ramsfraddr[5]), .Y(n640) );
  OAI22XL U2248 ( .A(n2060), .B(n1167), .C(n1569), .D(n1898), .Y(n1054) );
  AO21XL U2249 ( .B(ramdatao[3]), .C(n1142), .A(n1046), .Y(n1055) );
  OAI22XL U2250 ( .A(n1167), .B(n1921), .C(n1569), .D(n1225), .Y(n1123) );
  AO21XL U2251 ( .B(ramdatao[2]), .C(n1142), .A(n1115), .Y(n1124) );
  OAI22XL U2252 ( .A(n1167), .B(n1777), .C(n1569), .D(n1226), .Y(n934) );
  AO21XL U2253 ( .B(ramdatao[1]), .C(n1142), .A(n919), .Y(n935) );
  NAND21X1 U2254 ( .B(n155), .A(dec_accop[3]), .Y(n762) );
  XOR2XL U2255 ( .A(n1036), .B(acc[7]), .Y(n998) );
  NAND32XL U2256 ( .B(ramsfraddr[2]), .C(n2209), .A(n2211), .Y(n2214) );
  NAND21X1 U2257 ( .B(n495), .A(interrupt), .Y(n2371) );
  OAI221X1 U2258 ( .A(n837), .B(n496), .C(n2121), .D(n957), .E(n836), .Y(n1505) );
  AOI221XL U2259 ( .A(n1410), .B(n825), .C(instr[3]), .D(n783), .E(n782), .Y(
        n837) );
  AOI222XL U2260 ( .A(n127), .B(n835), .C(phase[3]), .D(n834), .E(phase[2]), 
        .F(n833), .Y(n836) );
  INVX1 U2261 ( .A(n734), .Y(n1170) );
  NAND21X1 U2262 ( .B(n1190), .A(dec_accop[14]), .Y(n734) );
  MUX2X1 U2263 ( .D0(n1964), .D1(temp[1]), .S(n1978), .Y(N12825) );
  MUX2XL U2264 ( .D0(n1962), .D1(temp[3]), .S(n1978), .Y(N12827) );
  MUX2XL U2265 ( .D0(n1174), .D1(n1171), .S(acc[7]), .Y(n983) );
  OAI221XL U2266 ( .A(n2456), .B(n822), .C(instr[7]), .D(n2320), .E(n1328), 
        .Y(n1308) );
  OA21XL U2267 ( .B(n821), .C(n1361), .A(n1366), .Y(n822) );
  INVX1 U2268 ( .A(n820), .Y(n821) );
  GEN2XL U2269 ( .D(n1093), .E(n1094), .C(n832), .B(n831), .A(n1313), .Y(n833)
         );
  INVX1 U2270 ( .A(n1312), .Y(n832) );
  MUX2XL U2271 ( .D0(n823), .D1(n1308), .S(instr[6]), .Y(n831) );
  AND2X1 U2272 ( .A(interrupt), .B(n2314), .Y(n823) );
  NAND21X1 U2273 ( .B(n1190), .A(dec_accop[4]), .Y(n763) );
  INVXL U2274 ( .A(n2452), .Y(n708) );
  MUX2BXL U2275 ( .D0(n1168), .D1(n278), .S(acc[1]), .Y(n919) );
  AOI21X1 U2276 ( .B(n1140), .C(n1480), .A(n1139), .Y(n278) );
  MUX2BXL U2277 ( .D0(n1168), .D1(n279), .S(acc[5]), .Y(n1141) );
  AOI21X1 U2278 ( .B(n1140), .C(n1789), .A(n1139), .Y(n279) );
  MUX2XL U2279 ( .D0(n1168), .D1(n1128), .S(acc[4]), .Y(n1129) );
  NAND21X1 U2280 ( .B(n1127), .A(n1126), .Y(n1128) );
  INVX1 U2281 ( .A(n1139), .Y(n1126) );
  MUX2XL U2282 ( .D0(n1140), .D1(n1125), .S(temp2_comb[4]), .Y(n1127) );
  MUX2BXL U2283 ( .D0(n1168), .D1(n280), .S(acc[3]), .Y(n1046) );
  AOI21X1 U2284 ( .B(n1140), .C(n1555), .A(n1139), .Y(n280) );
  MUX2BXL U2285 ( .D0(n1168), .D1(n281), .S(acc[2]), .Y(n1115) );
  AOI21X1 U2286 ( .B(n1140), .C(n1904), .A(n1139), .Y(n281) );
  MUX2BXL U2287 ( .D0(n1168), .D1(n282), .S(acc[6]), .Y(n1022) );
  AOI21X1 U2288 ( .B(n1140), .C(n2007), .A(n1139), .Y(n282) );
  MUX2XL U2289 ( .D0(n1174), .D1(n1171), .S(n2458), .Y(n930) );
  INVX1 U2290 ( .A(n605), .Y(n655) );
  NAND5XL U2291 ( .A(n604), .B(n603), .C(n602), .D(n2206), .E(n601), .Y(n605)
         );
  XOR2XL U2292 ( .A(n549), .B(ramsfraddr[0]), .Y(n604) );
  XOR2XL U2293 ( .A(n1807), .B(ramsfraddr[2]), .Y(n603) );
  AND4XL U2294 ( .A(ramwe), .B(n600), .C(n599), .D(n598), .Y(n601) );
  XOR2XL U2295 ( .A(n1596), .B(ramsfraddr[4]), .Y(n600) );
  XOR2XL U2296 ( .A(n1588), .B(ramsfraddr[3]), .Y(n599) );
  AOI211X1 U2297 ( .C(n1199), .D(n1198), .A(n1205), .B(n1197), .Y(n1200) );
  INVX1 U2298 ( .A(n1202), .Y(n1197) );
  OAI211XL U2299 ( .C(c), .D(n1196), .A(dec_cop[5]), .B(n1195), .Y(n1198) );
  INVXL U2300 ( .A(ramsfraddr[4]), .Y(n2218) );
  INVXL U2301 ( .A(acc[7]), .Y(n2060) );
  MUX2BXL U2302 ( .D0(sp[2]), .D1(n2333), .S(n235), .Y(n284) );
  MUX2BXL U2303 ( .D0(sp[3]), .D1(n1948), .S(n235), .Y(n285) );
  MUX2BXL U2304 ( .D0(sp[4]), .D1(n2336), .S(n235), .Y(n286) );
  INVXL U2305 ( .A(ramsfraddr[5]), .Y(n2207) );
  INVX1 U2306 ( .A(n728), .Y(n751) );
  NAND21XL U2307 ( .B(n154), .A(dec_accop[5]), .Y(n728) );
  INVX1 U2308 ( .A(n729), .Y(n750) );
  NAND21XL U2309 ( .B(n1190), .A(dec_accop[6]), .Y(n729) );
  AO21XL U2310 ( .B(n1050), .C(n1173), .A(n1555), .Y(n1051) );
  XOR3XL U2311 ( .A(n1049), .B(n274), .C(n1048), .Y(n1052) );
  MUX2XL U2312 ( .D0(n1174), .D1(n1171), .S(acc[3]), .Y(n1050) );
  AO21XL U2313 ( .B(n1119), .C(n1173), .A(n1904), .Y(n1120) );
  XOR3XL U2314 ( .A(n1118), .B(n271), .C(n1117), .Y(n1121) );
  MUX2XL U2315 ( .D0(n1174), .D1(n1171), .S(acc[2]), .Y(n1119) );
  NAND21X1 U2316 ( .B(n154), .A(dec_accop[1]), .Y(n730) );
  MUX4XL U2317 ( .D0(dpl_reg[4]), .D1(dpl_reg[12]), .D2(dpl_reg[20]), .D3(
        dpl_reg[28]), .S0(n392), .S1(n396), .Y(n383) );
  MUX4XL U2318 ( .D0(dpl_reg[5]), .D1(dpl_reg[13]), .D2(dpl_reg[21]), .D3(
        dpl_reg[29]), .S0(n392), .S1(n396), .Y(n385) );
  INVX1 U2319 ( .A(n725), .Y(n746) );
  NAND21XL U2320 ( .B(n154), .A(dec_accop[12]), .Y(n725) );
  INVX1 U2321 ( .A(n727), .Y(n748) );
  NAND21XL U2322 ( .B(n155), .A(dec_accop[11]), .Y(n727) );
  INVX1 U2323 ( .A(n2323), .Y(n497) );
  INVX1 U2324 ( .A(phase[0]), .Y(n2323) );
  INVX1 U2325 ( .A(n2163), .Y(n494) );
  INVX1 U2326 ( .A(phase[1]), .Y(n2163) );
  INVX1 U2327 ( .A(N344), .Y(n900) );
  INVXL U2328 ( .A(rs[0]), .Y(n1587) );
  NAND21XL U2329 ( .B(n1371), .A(n2453), .Y(n2318) );
  NAND43X1 U2330 ( .B(dec_accop[18]), .C(n1165), .D(n758), .A(dec_accop[17]), 
        .Y(n1979) );
  NAND21XL U2331 ( .B(n2453), .A(n1333), .Y(n1363) );
  MUX4X1 U2332 ( .D0(rn_reg[94]), .D1(rn_reg[86]), .D2(rn_reg[78]), .D3(
        rn_reg[70]), .S0(n482), .S1(n489), .Y(n459) );
  MUX4XL U2333 ( .D0(rn_reg[222]), .D1(rn_reg[214]), .D2(rn_reg[206]), .D3(
        rn_reg[198]), .S0(instr[0]), .S1(N353), .Y(n464) );
  MUX4X1 U2334 ( .D0(rn_reg[62]), .D1(rn_reg[54]), .D2(rn_reg[46]), .D3(
        rn_reg[38]), .S0(n482), .S1(n489), .Y(n458) );
  MUX4X1 U2335 ( .D0(rn_reg[190]), .D1(rn_reg[182]), .D2(rn_reg[174]), .D3(
        rn_reg[166]), .S0(n482), .S1(n489), .Y(n463) );
  MUX4X1 U2336 ( .D0(rn_reg[126]), .D1(rn_reg[118]), .D2(rn_reg[110]), .D3(
        rn_reg[102]), .S0(n482), .S1(n489), .Y(n460) );
  MUX4XL U2337 ( .D0(rn_reg[254]), .D1(rn_reg[246]), .D2(rn_reg[238]), .D3(
        rn_reg[230]), .S0(instr[0]), .S1(N353), .Y(n465) );
  MUX4XL U2338 ( .D0(dpl_reg[38]), .D1(dpl_reg[46]), .D2(dpl_reg[54]), .D3(
        dpl_reg[62]), .S0(n392), .S1(n396), .Y(n386) );
  MUX4X1 U2339 ( .D0(rn_reg[30]), .D1(rn_reg[22]), .D2(rn_reg[14]), .D3(
        rn_reg[6]), .S0(n482), .S1(n489), .Y(n457) );
  MUX4X1 U2340 ( .D0(rn_reg[158]), .D1(rn_reg[150]), .D2(rn_reg[142]), .D3(
        rn_reg[134]), .S0(n482), .S1(n489), .Y(n462) );
  NAND21XL U2341 ( .B(n1361), .A(n2452), .Y(n776) );
  NAND21XL U2342 ( .B(n2453), .A(n2452), .Y(n1327) );
  NAND21XL U2343 ( .B(n1167), .A(acc[4]), .Y(n1970) );
  NAND5XL U2344 ( .A(n797), .B(n1358), .C(n846), .D(n1107), .E(n674), .Y(n675)
         );
  NAND21XL U2345 ( .B(n154), .A(dec_accop[2]), .Y(n760) );
  MUX2XL U2346 ( .D0(n918), .D1(n287), .S(n2459), .Y(n1973) );
  AOI21XL U2347 ( .B(n1140), .C(n1872), .A(n1139), .Y(n287) );
  AO21XL U2348 ( .B(n752), .C(n1173), .A(n1872), .Y(n1971) );
  MUX2XL U2349 ( .D0(n1174), .D1(n1171), .S(n2459), .Y(n752) );
  AO21XL U2350 ( .B(temp2_comb[7]), .C(n997), .A(n992), .Y(n1156) );
  MUX4XL U2351 ( .D0(dpl_reg[6]), .D1(dpl_reg[14]), .D2(dpl_reg[22]), .D3(
        dpl_reg[30]), .S0(n392), .S1(n396), .Y(n387) );
  NAND21XL U2352 ( .B(n2305), .A(acc[2]), .Y(n1969) );
  XOR2XL U2353 ( .A(n1806), .B(ramsfraddr[1]), .Y(n602) );
  AOI21XL U2354 ( .B(dec_accop[18]), .C(accactv), .A(n1565), .Y(n288) );
  NOR5XL U2355 ( .A(dec_cop[5]), .B(n1192), .C(n1205), .D(n1191), .E(n154), 
        .Y(n1203) );
  MUX2XL U2356 ( .D0(n1189), .D1(n1188), .S(c), .Y(n1191) );
  NAND21X1 U2357 ( .B(dec_cop[6]), .A(dec_cop[7]), .Y(n1189) );
  INVX1 U2358 ( .A(ramdatao[2]), .Y(n2333) );
  INVX1 U2359 ( .A(ramdatao[1]), .Y(n2176) );
  INVX1 U2360 ( .A(ramdatao[4]), .Y(n2336) );
  MUX2BXL U2361 ( .D0(sp[6]), .D1(n2342), .S(n235), .Y(n289) );
  MUX2BXL U2362 ( .D0(sp[5]), .D1(n2339), .S(n235), .Y(n290) );
  INVX1 U2363 ( .A(n784), .Y(n1441) );
  AO2222XL U2364 ( .A(temp[6]), .B(n659), .C(n658), .D(ramsfraddr[6]), .E(
        n1944), .F(n657), .G(n656), .H(n2005), .Y(n644) );
  INVXL U2365 ( .A(ramsfraddr[2]), .Y(n2212) );
  INVX1 U2366 ( .A(n733), .Y(n754) );
  NAND21XL U2367 ( .B(n1190), .A(dec_accop[15]), .Y(n733) );
  INVX1 U2368 ( .A(N351), .Y(n547) );
  INVX1 U2369 ( .A(rs[1]), .Y(n1593) );
  GEN2XL U2370 ( .D(n860), .E(n859), .C(n1277), .B(n858), .A(n1908), .Y(n1798)
         );
  NAND32X1 U2371 ( .B(n493), .C(n477), .A(n1305), .Y(n860) );
  NAND21XL U2372 ( .B(n2315), .A(n2454), .Y(n1267) );
  NAND21XL U2373 ( .B(n2451), .A(n1100), .Y(n1415) );
  NAND21XL U2374 ( .B(n2452), .A(n1253), .Y(n1835) );
  NAND21XL U2375 ( .B(n2451), .A(n2452), .Y(n1365) );
  MUX2AXL U2376 ( .D0(sp[7]), .D1(n2344), .S(n235), .Y(n651) );
  NAND32XL U2377 ( .B(instr[5]), .C(n1835), .A(n2168), .Y(n973) );
  MUX2X1 U2378 ( .D0(n346), .D1(n345), .S(n349), .Y(dpc[1]) );
  MUX4X1 U2379 ( .D0(dpc_tab[1]), .D1(dpc_tab[7]), .D2(dpc_tab[13]), .D3(
        dpc_tab[19]), .S0(n357), .S1(n353), .Y(n346) );
  MUX4X1 U2380 ( .D0(dpc_tab[25]), .D1(dpc_tab[31]), .D2(dpc_tab[37]), .D3(
        dpc_tab[43]), .S0(n357), .S1(n353), .Y(n345) );
  AND2XL U2381 ( .A(b[1]), .B(n2459), .Y(N14337) );
  NAND21XL U2382 ( .B(instr[5]), .A(n2451), .Y(n709) );
  AO21XL U2383 ( .B(n1193), .C(n1164), .A(n155), .Y(n1195) );
  INVX1 U2384 ( .A(dec_cop[4]), .Y(n1164) );
  NAND21XL U2385 ( .B(n1190), .A(dec_cop[1]), .Y(n1202) );
  NAND21XL U2386 ( .B(n2453), .A(n794), .Y(n883) );
  NAND21X1 U2387 ( .B(n971), .A(phase[1]), .Y(n889) );
  MUX2BXL U2388 ( .D0(n16), .D1(n677), .S(n2457), .Y(n678) );
  NAND21X1 U2389 ( .B(n676), .A(n2313), .Y(n677) );
  INVX1 U2390 ( .A(n1163), .Y(n1205) );
  NAND21XL U2391 ( .B(n154), .A(dec_cop[2]), .Y(n1163) );
  NOR21XL U2392 ( .B(n1096), .A(n1095), .Y(n1108) );
  NOR43XL U2393 ( .B(interrupt), .C(n1094), .D(n1093), .A(n1092), .Y(n1095) );
  OAI22X1 U2394 ( .A(n1110), .B(n496), .C(n1109), .D(n493), .Y(n2310) );
  AOI221XL U2395 ( .A(n1372), .B(n1100), .C(n1370), .D(instr[6]), .E(n1099), 
        .Y(n1110) );
  AOI211X1 U2396 ( .C(n1362), .D(n1105), .A(n1104), .B(n1103), .Y(n1106) );
  AO21X1 U2397 ( .B(phase[1]), .C(n851), .A(n295), .Y(n857) );
  NAND43X1 U2398 ( .B(n1234), .C(n1288), .D(n1282), .A(n971), .Y(n851) );
  INVX1 U2399 ( .A(n788), .Y(n2121) );
  AOI32XL U2400 ( .A(n847), .B(n1493), .C(n786), .D(n1334), .E(instr[7]), .Y(
        n787) );
  AND2XL U2401 ( .A(b[0]), .B(n2459), .Y(N14336) );
  NAND21XL U2402 ( .B(n237), .A(acc[1]), .Y(n1965) );
  OAI31XL U2403 ( .A(n1097), .B(n1379), .C(n2319), .D(n1108), .Y(n1098) );
  INVX1 U2404 ( .A(n588), .Y(n606) );
  GEN2XL U2405 ( .D(n1493), .E(n1304), .C(n1362), .B(phase[0]), .A(n587), .Y(
        n588) );
  AND3X1 U2406 ( .A(n1841), .B(phase[1]), .C(n1294), .Y(n587) );
  INVXL U2407 ( .A(c), .Y(n1194) );
  XNOR2XL U2408 ( .A(n1036), .B(acc[6]), .Y(n291) );
  INVXL U2409 ( .A(N349), .Y(n543) );
  INVX1 U2410 ( .A(n717), .Y(n1093) );
  NOR2X1 U2411 ( .A(n1313), .B(n293), .Y(n292) );
  INVX1 U2412 ( .A(dec_cop[3]), .Y(n1193) );
  INVX1 U2413 ( .A(n1297), .Y(n2117) );
  OAI221XL U2414 ( .A(instr[5]), .B(n1435), .C(n1500), .D(n1371), .E(n1296), 
        .Y(n1297) );
  AOI211X1 U2415 ( .C(n1295), .D(n1304), .A(n1294), .B(n1298), .Y(n1296) );
  NAND21XL U2416 ( .B(n298), .A(ramsfraddr[7]), .Y(n1767) );
  NAND21XL U2417 ( .B(n2453), .A(n2157), .Y(n1434) );
  MUX2X1 U2418 ( .D0(n344), .D1(n343), .S(n349), .Y(dpc[2]) );
  MUX4X1 U2419 ( .D0(dpc_tab[2]), .D1(dpc_tab[8]), .D2(dpc_tab[14]), .D3(
        dpc_tab[20]), .S0(n357), .S1(n353), .Y(n344) );
  MUX4X1 U2420 ( .D0(dpc_tab[26]), .D1(dpc_tab[32]), .D2(dpc_tab[38]), .D3(
        dpc_tab[44]), .S0(n357), .S1(n353), .Y(n343) );
  NAND21XL U2421 ( .B(instr[4]), .A(n2453), .Y(n1268) );
  AOI32X1 U2422 ( .A(n30), .B(phase[1]), .C(n1252), .D(n1359), .E(n239), .Y(
        n1254) );
  INVX1 U2423 ( .A(n1251), .Y(n1252) );
  NAND21XL U2424 ( .B(n155), .A(dec_accop[16]), .Y(n1506) );
  AO21XL U2425 ( .B(n2452), .C(n1333), .A(n1493), .Y(n801) );
  AO21X1 U2426 ( .B(waitcnt[2]), .C(n2183), .A(n577), .Y(n2235) );
  OA21X1 U2427 ( .B(waitcnt[2]), .C(n2183), .A(n576), .Y(n577) );
  AO21X1 U2428 ( .B(waitcnt[1]), .C(n2184), .A(n575), .Y(n576) );
  OA22X1 U2429 ( .A(waitcnt[1]), .B(n2184), .C(waitcnt[0]), .D(n2187), .Y(n575) );
  INVX1 U2430 ( .A(n756), .Y(n1498) );
  NAND21XL U2431 ( .B(n154), .A(dec_accop[17]), .Y(n756) );
  MUX2X1 U2432 ( .D0(n348), .D1(n347), .S(n349), .Y(dpc[0]) );
  MUX4X1 U2433 ( .D0(dpc_tab[0]), .D1(dpc_tab[6]), .D2(dpc_tab[12]), .D3(
        dpc_tab[18]), .S0(n357), .S1(n353), .Y(n348) );
  MUX4X1 U2434 ( .D0(dpc_tab[24]), .D1(dpc_tab[30]), .D2(dpc_tab[36]), .D3(
        dpc_tab[42]), .S0(n357), .S1(n353), .Y(n347) );
  GEN2XL U2435 ( .D(n1406), .E(n30), .C(n781), .B(n780), .A(n779), .Y(n782) );
  OAI222XL U2436 ( .A(interrupt), .B(n2313), .C(N352), .D(n776), .E(instr[7]), 
        .F(n847), .Y(n780) );
  MUX2X1 U2437 ( .D0(n778), .D1(n240), .S(n777), .Y(n779) );
  OAI33XL U2438 ( .A(n2156), .B(n2315), .C(n1361), .D(n2457), .E(n1360), .F(
        n776), .Y(n781) );
  AND2XL U2439 ( .A(b[0]), .B(n2458), .Y(N14344) );
  MUX2X1 U2440 ( .D0(n334), .D1(n333), .S(n349), .Y(dph[1]) );
  MUX4X1 U2441 ( .D0(dph_reg[1]), .D1(dph_reg[9]), .D2(dph_reg[17]), .D3(
        dph_reg[25]), .S0(n356), .S1(n352), .Y(n334) );
  MUX4X1 U2442 ( .D0(dph_reg[33]), .D1(dph_reg[41]), .D2(dph_reg[49]), .D3(
        dph_reg[57]), .S0(n356), .S1(n352), .Y(n333) );
  MUX2X1 U2443 ( .D0(n332), .D1(n331), .S(n349), .Y(dph[2]) );
  MUX4X1 U2444 ( .D0(dph_reg[2]), .D1(dph_reg[10]), .D2(dph_reg[18]), .D3(
        dph_reg[26]), .S0(n356), .S1(n352), .Y(n332) );
  MUX4X1 U2445 ( .D0(dph_reg[34]), .D1(dph_reg[42]), .D2(dph_reg[50]), .D3(
        dph_reg[58]), .S0(n356), .S1(n352), .Y(n331) );
  MUX2BXL U2446 ( .D0(N352), .D1(n294), .S(n2451), .Y(n827) );
  OAI22XL U2447 ( .A(n1278), .B(n1092), .C(n2456), .D(n849), .Y(n294) );
  MUX2X1 U2448 ( .D0(n318), .D1(n317), .S(N351), .Y(dpl[1]) );
  MUX4X1 U2449 ( .D0(dpl_reg[1]), .D1(dpl_reg[9]), .D2(dpl_reg[17]), .D3(
        dpl_reg[25]), .S0(n354), .S1(n350), .Y(n318) );
  MUX4X1 U2450 ( .D0(dpl_reg[33]), .D1(dpl_reg[41]), .D2(dpl_reg[49]), .D3(
        dpl_reg[57]), .S0(n354), .S1(n350), .Y(n317) );
  MUX2X1 U2451 ( .D0(n316), .D1(n315), .S(N351), .Y(dpl[2]) );
  MUX4X1 U2452 ( .D0(dpl_reg[2]), .D1(dpl_reg[10]), .D2(dpl_reg[18]), .D3(
        dpl_reg[26]), .S0(n354), .S1(n350), .Y(n316) );
  MUX4X1 U2453 ( .D0(dpl_reg[34]), .D1(dpl_reg[42]), .D2(dpl_reg[50]), .D3(
        dpl_reg[58]), .S0(n354), .S1(n350), .Y(n315) );
  OA22X1 U2454 ( .A(waitcnt[1]), .B(n2177), .C(waitcnt[0]), .D(n2179), .Y(n573) );
  OAI22X1 U2455 ( .A(n492), .B(n2361), .C(n2162), .D(n496), .Y(n2326) );
  AND4X1 U2456 ( .A(n2161), .B(n2160), .C(n2159), .D(n2158), .Y(n2162) );
  OA22XL U2457 ( .A(n2151), .B(n2150), .C(instr[5]), .D(n2149), .Y(n2159) );
  OA2222XL U2458 ( .A(n2157), .B(n2156), .C(n2319), .D(n2155), .E(n2154), .F(
        n2153), .G(n16), .H(n2152), .Y(n2158) );
  AND2X1 U2459 ( .A(n1285), .B(phase[2]), .Y(n295) );
  INVX1 U2460 ( .A(n665), .Y(n2169) );
  AOI21AX1 U2461 ( .B(waitcnt[2]), .C(n2175), .A(n297), .Y(n296) );
  OAI21X1 U2462 ( .B(waitcnt[2]), .C(n2175), .A(n574), .Y(n297) );
  AND4X1 U2463 ( .A(n1160), .B(n1159), .C(n1158), .D(n1157), .Y(n1161) );
  INVX1 U2464 ( .A(dec_accop[1]), .Y(n1160) );
  INVX1 U2465 ( .A(dec_cop[6]), .Y(n1159) );
  INVX1 U2466 ( .A(dec_accop[4]), .Y(n1158) );
  INVX1 U2467 ( .A(ramdatao[7]), .Y(n2344) );
  INVX1 U2468 ( .A(ramdatao[6]), .Y(n2342) );
  INVX1 U2469 ( .A(ramdatao[5]), .Y(n2339) );
  INVX1 U2470 ( .A(phase[2]), .Y(n2118) );
  OAI31XL U2471 ( .A(n830), .B(n829), .C(n1327), .D(n828), .Y(n1313) );
  AO21XL U2472 ( .B(instr[7]), .C(n1101), .A(n824), .Y(n830) );
  AO21X1 U2473 ( .B(n2320), .C(n827), .A(n826), .Y(n828) );
  AOI32XL U2474 ( .A(n2148), .B(instr[6]), .C(n477), .D(n2147), .E(n2146), .Y(
        n2151) );
  INVX1 U2475 ( .A(temp2_comb[5]), .Y(n1789) );
  INVX1 U2476 ( .A(n664), .Y(n825) );
  NAND21XL U2477 ( .B(n2453), .A(n708), .Y(n664) );
  INVX1 U2478 ( .A(n841), .Y(n872) );
  OAI31XL U2479 ( .A(n840), .B(n839), .C(n1060), .D(phase[1]), .Y(n841) );
  INVX1 U2480 ( .A(n2160), .Y(n840) );
  INVX1 U2481 ( .A(n2362), .Y(n839) );
  INVX1 U2482 ( .A(dec_accop[17]), .Y(n1157) );
  INVX1 U2483 ( .A(ckcon[0]), .Y(n2179) );
  INVX1 U2484 ( .A(dec_cop[7]), .Y(n1162) );
  INVX1 U2485 ( .A(ckcon[4]), .Y(n2187) );
  NAND2XL U2486 ( .A(n299), .B(n1258), .Y(n1259) );
  GEN2XL U2487 ( .D(n723), .E(n722), .C(n2118), .B(n721), .A(n1142), .Y(n769)
         );
  AOI31XL U2488 ( .A(n1094), .B(instr[2]), .C(n1846), .D(n716), .Y(n722) );
  AOI32X1 U2489 ( .A(phase[3]), .B(n1339), .C(n1093), .D(phase[1]), .E(n720), 
        .Y(n721) );
  NAND21XL U2490 ( .B(n2451), .A(n800), .Y(n1385) );
  AO21X1 U2491 ( .B(N345), .C(n1780), .A(n1778), .Y(n1912) );
  NAND32XL U2492 ( .B(instr[4]), .C(n1255), .A(n1278), .Y(n2173) );
  OR2XL U2493 ( .A(instr[5]), .B(n1247), .Y(n1009) );
  NAND21XL U2494 ( .B(n2452), .A(n1339), .Y(n2153) );
  OAI211XL U2495 ( .C(n819), .D(n818), .A(n1100), .B(n1101), .Y(n1312) );
  XOR2XL U2496 ( .A(n2316), .B(n2451), .Y(n819) );
  XOR2XL U2497 ( .A(instr[7]), .B(n548), .Y(n818) );
  INVX1 U2498 ( .A(n1221), .Y(n1237) );
  OAI31XL U2499 ( .A(instr[7]), .B(n1367), .C(n1279), .D(n1408), .Y(n1221) );
  MUX2X1 U2500 ( .D0(n336), .D1(n335), .S(n349), .Y(dph[0]) );
  MUX4X1 U2501 ( .D0(dph_reg[0]), .D1(dph_reg[8]), .D2(dph_reg[16]), .D3(
        dph_reg[24]), .S0(n356), .S1(n352), .Y(n336) );
  MUX4X1 U2502 ( .D0(dph_reg[32]), .D1(dph_reg[40]), .D2(dph_reg[48]), .D3(
        dph_reg[56]), .S0(n356), .S1(n352), .Y(n335) );
  OA22XL U2503 ( .A(instr[7]), .B(n1279), .C(n1278), .D(n1277), .Y(n1281) );
  NAND21XL U2504 ( .B(n757), .A(ramdatao[0]), .Y(n1967) );
  INVX1 U2505 ( .A(n873), .Y(n2082) );
  OAI22XL U2506 ( .A(ramsfraddr[7]), .B(n874), .C(n872), .D(n871), .Y(n873) );
  INVXL U2507 ( .A(temp2_comb[2]), .Y(n1904) );
  INVXL U2508 ( .A(temp2_comb[1]), .Y(n1480) );
  INVX1 U2509 ( .A(temp2_comb[7]), .Y(n2096) );
  INVXL U2510 ( .A(temp2_comb[3]), .Y(n1555) );
  INVX1 U2511 ( .A(temp2_comb[6]), .Y(n2007) );
  INVX1 U2512 ( .A(n815), .Y(n965) );
  NOR2XL U2513 ( .A(dec_accop[9]), .B(dec_accop[10]), .Y(n300) );
  INVX1 U2514 ( .A(ckcon[1]), .Y(n2177) );
  INVX1 U2515 ( .A(ckcon[6]), .Y(n2183) );
  INVX1 U2516 ( .A(ckcon[5]), .Y(n2184) );
  INVX1 U2517 ( .A(ckcon[2]), .Y(n2175) );
  NAND21XL U2518 ( .B(instr[7]), .A(instr[5]), .Y(n1337) );
  NAND21XL U2519 ( .B(instr[4]), .A(n1100), .Y(n1251) );
  INVX1 U2520 ( .A(n1061), .Y(n869) );
  OR2X1 U2521 ( .A(memrd), .B(memwr), .Y(n2236) );
  OR2X1 U2522 ( .A(mempswr), .B(mempsrd), .Y(n2238) );
  INVX1 U2523 ( .A(n939), .Y(n949) );
  MUX2XL U2524 ( .D0(n2094), .D1(n2086), .S(pc_o[1]), .Y(n938) );
  OA22X1 U2525 ( .A(n2093), .B(n1475), .C(n2085), .D(n48), .Y(n937) );
  MUX2X1 U2526 ( .D0(n1230), .D1(n1229), .S(N345), .Y(n1231) );
  OA2222XL U2527 ( .A(n1228), .B(n1227), .C(n1898), .D(n1929), .E(n1868), .F(
        n1226), .G(n1225), .H(n2399), .Y(n1230) );
  OA2222XL U2528 ( .A(n2060), .B(n1228), .C(n1929), .D(n1921), .E(n1810), .F(
        n1868), .G(n2399), .H(n1777), .Y(n1229) );
  NAND21XL U2529 ( .B(n1003), .A(n2459), .Y(n1004) );
  INVXL U2530 ( .A(n2459), .Y(n1226) );
  INVXL U2531 ( .A(n2458), .Y(n1225) );
  INVXL U2532 ( .A(acc[4]), .Y(n1810) );
  INVXL U2533 ( .A(acc[3]), .Y(n1227) );
  INVXL U2534 ( .A(ramsfraddr[3]), .Y(n2220) );
  AND3X1 U2535 ( .A(n842), .B(n703), .C(n1363), .Y(n707) );
  OAI221X1 U2536 ( .A(n1092), .B(n1337), .C(n709), .D(n1302), .E(n705), .Y(
        n706) );
  INVXL U2537 ( .A(temp2_comb[4]), .Y(n1819) );
  AOI31XL U2538 ( .A(instr[6]), .B(n2456), .C(n1267), .D(n1334), .Y(n705) );
  NAND21XL U2539 ( .B(n876), .A(pc_o[0]), .Y(n1869) );
  NAND21X1 U2540 ( .B(n1307), .A(n1306), .Y(n1310) );
  AO21X1 U2541 ( .B(N352), .C(n1305), .A(n1304), .Y(n1306) );
  INVX1 U2542 ( .A(temp[0]), .Y(n1458) );
  INVX1 U2543 ( .A(temp[1]), .Y(n1481) );
  INVX1 U2544 ( .A(temp[3]), .Y(n1554) );
  INVX1 U2545 ( .A(temp[4]), .Y(n1809) );
  MUX2XL U2546 ( .D0(pc_o[11]), .D1(n2419), .S(n550), .Y(memaddr_comb[11]) );
  AO2222XL U2547 ( .A(n210), .B(ramdatao[3]), .C(n1534), .D(n2198), .E(
        memaddr[11]), .F(n2197), .G(p2[3]), .H(n211), .Y(n2419) );
  AO2222XL U2548 ( .A(pc_i[11]), .B(n2196), .C(n2195), .D(temp[3]), .E(n1983), 
        .F(n203), .G(alu_out[11]), .H(n114), .Y(n1534) );
  INVX1 U2549 ( .A(phase[3]), .Y(n2120) );
  INVX1 U2550 ( .A(n956), .Y(n1357) );
  INVX1 U2551 ( .A(temp[2]), .Y(n1897) );
  INVX1 U2552 ( .A(phase[4]), .Y(n957) );
  MUX2XL U2553 ( .D0(ramsfraddr[0]), .D1(n2348), .S(n551), .Y(
        ramsfraddr_comb[0]) );
  MUX2XL U2554 ( .D0(ramsfraddr[1]), .D1(n72), .S(n2450), .Y(
        ramsfraddr_comb[1]) );
  MUX2XL U2555 ( .D0(pc_o[13]), .D1(n2421), .S(n550), .Y(memaddr_comb[13]) );
  MUX2XL U2556 ( .D0(pc_o[7]), .D1(n2414), .S(n82), .Y(memaddr_comb[7]) );
  MUX2XL U2557 ( .D0(pc_o[12]), .D1(n2420), .S(n550), .Y(memaddr_comb[12]) );
  MUX2XL U2558 ( .D0(pc_o[14]), .D1(n2422), .S(n550), .Y(memaddr_comb[14]) );
  OR2X1 U2559 ( .A(state[2]), .B(state[1]), .Y(n2364) );
  NAND21X1 U2560 ( .B(state[0]), .A(n1086), .Y(n2109) );
  AO2222XL U2561 ( .A(n210), .B(ramdatao[4]), .C(n1537), .D(n2198), .E(
        pc_o[12]), .F(n2197), .G(p2[4]), .H(n211), .Y(n2420) );
  AO2222XL U2562 ( .A(pc_i[12]), .B(n2196), .C(n2195), .D(temp[4]), .E(n1982), 
        .F(n203), .G(alu_out[12]), .H(n114), .Y(n1537) );
  AO2222XL U2563 ( .A(n210), .B(ramdatao[6]), .C(n2026), .D(n2198), .E(
        pc_o[14]), .F(n2197), .G(p2[6]), .H(n211), .Y(n2422) );
  AO2222XL U2564 ( .A(pc_i[14]), .B(n2196), .C(n2195), .D(temp[6]), .E(n2025), 
        .F(n203), .G(alu_out[14]), .H(n114), .Y(n2026) );
  AO2222XL U2565 ( .A(n210), .B(ramdatao[5]), .C(n1953), .D(n2198), .E(
        pc_o[13]), .F(n2197), .G(p2[5]), .H(n211), .Y(n2421) );
  AO2222XL U2566 ( .A(pc_i[13]), .B(n2196), .C(n2195), .D(temp[5]), .E(n1981), 
        .F(n203), .G(alu_out[13]), .H(n114), .Y(n1953) );
  MUX2XL U2567 ( .D0(mempsrd), .D1(n2375), .S(n550), .Y(mempsrd_comb) );
  MUX2XL U2568 ( .D0(memaddr[8]), .D1(n2415), .S(n82), .Y(memaddr_comb[8]) );
  MUX2XL U2569 ( .D0(pc_o[9]), .D1(n2416), .S(n90), .Y(memaddr_comb[9]) );
  MUX2X1 U2570 ( .D0(pc_o[7]), .D1(n2049), .S(n1993), .Y(N12848) );
  AO21XL U2571 ( .B(n1974), .C(n2073), .A(n2439), .Y(N12831) );
  MUX2X1 U2572 ( .D0(memaddr[8]), .D1(n1986), .S(n1993), .Y(N12849) );
  MUX2X1 U2573 ( .D0(memaddr[9]), .D1(n1985), .S(n1993), .Y(N12850) );
  MUX2X1 U2574 ( .D0(memaddr[10]), .D1(n1984), .S(n109), .Y(N12851) );
  MUX2X1 U2575 ( .D0(pc_o[11]), .D1(n1983), .S(n109), .Y(N12852) );
  MUX2X1 U2576 ( .D0(memaddr[12]), .D1(n1982), .S(n109), .Y(N12853) );
  MUX2X1 U2577 ( .D0(memaddr[13]), .D1(n1981), .S(n109), .Y(N12854) );
  MUX2X1 U2578 ( .D0(memaddr[14]), .D1(n2025), .S(n109), .Y(N12855) );
  MUX2XL U2579 ( .D0(ramsfraddr[2]), .D1(n2350), .S(waitstaten), .Y(
        ramsfraddr_comb[2]) );
  MUX2X1 U2580 ( .D0(pc_o[15]), .D1(n2423), .S(waitstaten), .Y(
        memaddr_comb[15]) );
  AO2222XL U2581 ( .A(ramdatao[7]), .B(n210), .C(n2199), .D(n2198), .E(
        pc_o[15]), .F(n2197), .G(p2[7]), .H(n211), .Y(n2423) );
  AO2222XL U2582 ( .A(pc_i[15]), .B(n2196), .C(n2195), .D(temp[7]), .E(n2194), 
        .F(n203), .G(alu_out[15]), .H(n114), .Y(n2199) );
  INVX1 U2583 ( .A(idle), .Y(n2136) );
  MUX2XL U2584 ( .D0(pc_o[10]), .D1(n2418), .S(n90), .Y(memaddr_comb[10]) );
  NAND21X1 U2585 ( .B(n1471), .A(n1470), .Y(n2416) );
  OA2222XL U2586 ( .A(n48), .B(n1894), .C(n1481), .D(n1893), .E(n2176), .F(
        n1892), .G(n1891), .H(n1469), .Y(n1470) );
  AO2222XL U2587 ( .A(alu_out[9]), .B(n114), .C(n1889), .D(pc_i[9]), .E(n1985), 
        .F(n2193), .G(n1888), .H(instr[6]), .Y(n1471) );
  NAND21X1 U2588 ( .B(n1896), .A(n1895), .Y(n2418) );
  OA2222XL U2589 ( .A(n1894), .B(n1901), .C(n1897), .D(n1893), .E(n2333), .F(
        n1892), .G(n1891), .H(n1890), .Y(n1895) );
  AO2222XL U2590 ( .A(alu_out[10]), .B(n114), .C(pc_i[10]), .D(n1889), .E(
        n1984), .F(n203), .G(n1888), .H(instr[7]), .Y(n1896) );
  NAND21X1 U2591 ( .B(n1455), .A(n1454), .Y(n2415) );
  OA2222XL U2592 ( .A(n1894), .B(n40), .C(n1458), .D(n1893), .E(n2178), .F(
        n1892), .G(n1891), .H(n1453), .Y(n1454) );
  AO2222XL U2593 ( .A(alu_out[8]), .B(n114), .C(pc_i[8]), .D(n1889), .E(n1986), 
        .F(n2193), .G(n1888), .H(instr[5]), .Y(n1455) );
  INVXL U2594 ( .A(pc_o[0]), .Y(n1854) );
  INVX1 U2595 ( .A(pc_i[0]), .Y(n1871) );
  INVX1 U2596 ( .A(idle_r), .Y(n2137) );
  NAND21X1 U2597 ( .B(n1089), .A(n1088), .Y(n2133) );
  MUX2X1 U2598 ( .D0(cs_run), .D1(n2125), .S(codefetch_s), .Y(n1089) );
  NOR42XL U2599 ( .C(n2365), .D(n2125), .A(interrupt), .B(pdmode), .Y(n2126)
         );
  INVXL U2600 ( .A(pc_o[1]), .Y(n1479) );
  AO222X1 U2601 ( .A(n1684), .B(temp[1]), .C(dptr_inc[9]), .D(n147), .E(n1682), 
        .F(n18), .Y(n1985) );
  AO222X1 U2602 ( .A(n1684), .B(temp[0]), .C(dptr_inc[8]), .D(n147), .E(n1682), 
        .F(n19), .Y(n1986) );
  AO222X1 U2603 ( .A(n1666), .B(temp[7]), .C(dptr_inc[7]), .D(n1683), .E(n1665), .F(n17), .Y(n2049) );
  AO222X1 U2604 ( .A(n1684), .B(temp[2]), .C(dptr_inc[10]), .D(n147), .E(n1682), .F(n20), .Y(n1984) );
  AO222X1 U2605 ( .A(n1684), .B(temp[3]), .C(dptr_inc[11]), .D(n147), .E(n1682), .F(n21), .Y(n1983) );
  AO222X1 U2606 ( .A(n1684), .B(temp[4]), .C(dptr_inc[12]), .D(n147), .E(n1682), .F(n22), .Y(n1982) );
  MUX4XL U2607 ( .D0(dpl_reg[39]), .D1(dpl_reg[47]), .D2(dpl_reg[55]), .D3(
        dpl_reg[63]), .S0(n392), .S1(n396), .Y(n388) );
  MUX2XL U2608 ( .D0(ramdatao[0]), .D1(n2329), .S(n551), .Y(ramdatao_comb[0])
         );
  MUX2XL U2609 ( .D0(ramdatao[3]), .D1(n2335), .S(n551), .Y(ramdatao_comb[3])
         );
  MUX2X1 U2610 ( .D0(n1081), .D1(n2279), .S(n2331), .Y(n2335) );
  NAND32X1 U2611 ( .B(n1078), .C(n1077), .A(n1076), .Y(n1081) );
  AO2222XL U2612 ( .A(pc_i[11]), .B(n1058), .C(pc_o[11]), .D(n1057), .E(n2246), 
        .F(pc_o[3]), .G(temp2_comb[3]), .H(n1056), .Y(n1077) );
  MUX2X1 U2613 ( .D0(n308), .D1(n307), .S(N351), .Y(dpl[6]) );
  MUX4X1 U2614 ( .D0(dpl_reg[6]), .D1(dpl_reg[14]), .D2(dpl_reg[22]), .D3(
        dpl_reg[30]), .S0(N349), .S1(N350), .Y(n308) );
  MUX2X1 U2615 ( .D0(n326), .D1(n325), .S(dps[2]), .Y(dph[5]) );
  MUX4X1 U2616 ( .D0(dph_reg[5]), .D1(dph_reg[13]), .D2(dph_reg[21]), .D3(
        dph_reg[29]), .S0(n355), .S1(n351), .Y(n326) );
  MUX4X1 U2617 ( .D0(dph_reg[37]), .D1(dph_reg[45]), .D2(dph_reg[53]), .D3(
        dph_reg[61]), .S0(n355), .S1(n351), .Y(n325) );
  MUX2X1 U2618 ( .D0(n328), .D1(n327), .S(N351), .Y(dph[4]) );
  MUX4X1 U2619 ( .D0(dph_reg[4]), .D1(dph_reg[12]), .D2(dph_reg[20]), .D3(
        dph_reg[28]), .S0(n355), .S1(n351), .Y(n328) );
  MUX4X1 U2620 ( .D0(dph_reg[36]), .D1(dph_reg[44]), .D2(dph_reg[52]), .D3(
        dph_reg[60]), .S0(n355), .S1(n351), .Y(n327) );
  MUX4XL U2621 ( .D0(dpl_reg[7]), .D1(dpl_reg[15]), .D2(dpl_reg[23]), .D3(
        dpl_reg[31]), .S0(n392), .S1(n396), .Y(n389) );
  MUX2X1 U2622 ( .D0(n312), .D1(n311), .S(N351), .Y(dpl[4]) );
  MUX4X1 U2623 ( .D0(dpl_reg[4]), .D1(dpl_reg[12]), .D2(dpl_reg[20]), .D3(
        dpl_reg[28]), .S0(n354), .S1(n350), .Y(n312) );
  MUX4X1 U2624 ( .D0(dpl_reg[36]), .D1(dpl_reg[44]), .D2(dpl_reg[52]), .D3(
        dpl_reg[60]), .S0(n354), .S1(n350), .Y(n311) );
  AO222X1 U2625 ( .A(n1684), .B(temp[7]), .C(dptr_inc[15]), .D(n147), .E(n1682), .F(dph_current_7_), .Y(n2194) );
  INVX1 U2626 ( .A(n1667), .Y(dph_current_7_) );
  MUX2AXL U2627 ( .D0(N11845), .D1(n2344), .S(n1679), .Y(n1667) );
  AO222X1 U2628 ( .A(n1684), .B(temp[6]), .C(dptr_inc[14]), .D(n147), .E(n1682), .F(n24), .Y(n2025) );
  AO222X1 U2629 ( .A(n1684), .B(temp[5]), .C(dptr_inc[13]), .D(n147), .E(n1682), .F(n23), .Y(n1981) );
  MUX4X1 U2630 ( .D0(dph_reg[32]), .D1(dph_reg[40]), .D2(dph_reg[48]), .D3(
        dph_reg[56]), .S0(n541), .S1(n539), .Y(n358) );
  MUX2XL U2631 ( .D0(ramdatao[1]), .D1(n2330), .S(n551), .Y(ramdatao_comb[1])
         );
  MUX2X1 U2632 ( .D0(n322), .D1(n321), .S(N351), .Y(dph[7]) );
  MUX2X1 U2633 ( .D0(n306), .D1(n305), .S(dps[2]), .Y(dpl[7]) );
  AO222XL U2634 ( .A(n28), .B(memaddr[2]), .C(n27), .D(n2409), .E(pc_ini[2]), 
        .F(n556), .Y(N482) );
  AO222XL U2635 ( .A(n29), .B(pc_o[6]), .C(n2057), .D(n2413), .E(pc_ini[6]), 
        .F(n556), .Y(N486) );
  AO222XL U2636 ( .A(n28), .B(pc_o[5]), .C(n27), .D(n2412), .E(pc_ini[5]), .F(
        n556), .Y(N485) );
  AO222XL U2637 ( .A(n29), .B(memaddr[4]), .C(n2057), .D(n2411), .E(pc_ini[4]), 
        .F(n555), .Y(N484) );
  AO222XL U2638 ( .A(n28), .B(pc_o[3]), .C(n27), .D(n2410), .E(pc_ini[3]), .F(
        n556), .Y(N483) );
  AO222X1 U2639 ( .A(n29), .B(pc_o[8]), .C(n2057), .D(n2415), .E(pc_ini[8]), 
        .F(n555), .Y(N488) );
  AO222X1 U2640 ( .A(n28), .B(memaddr[7]), .C(n27), .D(n2414), .E(pc_ini[7]), 
        .F(n556), .Y(N487) );
  AO222X1 U2641 ( .A(n29), .B(pc_o[10]), .C(n2057), .D(n2418), .E(pc_ini[10]), 
        .F(n556), .Y(N490) );
  AO222X1 U2642 ( .A(n28), .B(pc_o[9]), .C(n27), .D(n2416), .E(pc_ini[9]), .F(
        n555), .Y(N489) );
  AO222XL U2643 ( .A(n29), .B(pc_o[1]), .C(n2057), .D(n2408), .E(pc_ini[1]), 
        .F(n555), .Y(N481) );
  AO222XL U2644 ( .A(n28), .B(pc_o[0]), .C(n27), .D(n2407), .E(pc_ini[0]), .F(
        n556), .Y(N480) );
  MUX2X1 U2645 ( .D0(n324), .D1(n323), .S(dps[2]), .Y(dph[6]) );
  MUX4X1 U2646 ( .D0(dph_reg[6]), .D1(dph_reg[14]), .D2(dph_reg[22]), .D3(
        dph_reg[30]), .S0(n355), .S1(n351), .Y(n324) );
  MUX4X1 U2647 ( .D0(dph_reg[38]), .D1(dph_reg[46]), .D2(dph_reg[54]), .D3(
        dph_reg[62]), .S0(n355), .S1(n351), .Y(n323) );
  MUX2X1 U2648 ( .D0(pc_o[15]), .D1(n2194), .S(n109), .Y(N12856) );
  AO21X1 U2649 ( .B(n2369), .C(n2368), .A(n2367), .Y(n1878) );
  INVX1 U2650 ( .A(n2363), .Y(n2369) );
  GEN2XL U2651 ( .D(n2366), .E(n2365), .C(n2364), .B(newinstrlock), .A(n561), 
        .Y(n2367) );
  AO22X1 U2652 ( .A(n502), .B(n2422), .C(pc_ini[14]), .D(n557), .Y(N494) );
  AO22X1 U2653 ( .A(n502), .B(n2421), .C(pc_ini[13]), .D(n557), .Y(N493) );
  AO22X1 U2654 ( .A(n507), .B(n2420), .C(pc_ini[12]), .D(n556), .Y(N492) );
  AO22X1 U2655 ( .A(n508), .B(n2419), .C(pc_ini[11]), .D(n556), .Y(N491) );
  AO22X1 U2656 ( .A(n502), .B(n2423), .C(pc_ini[15]), .D(n557), .Y(N495) );
  AND2XL U2657 ( .A(sfroe_r), .B(n551), .Y(sfroe) );
  MUX4X1 U2658 ( .D0(dph_reg[0]), .D1(dph_reg[8]), .D2(dph_reg[16]), .D3(
        dph_reg[24]), .S0(n42), .S1(N347), .Y(n359) );
  MUX2X1 U2659 ( .D0(n310), .D1(n309), .S(N351), .Y(dpl[5]) );
  MUX4X1 U2660 ( .D0(dpl_reg[5]), .D1(dpl_reg[13]), .D2(dpl_reg[21]), .D3(
        dpl_reg[29]), .S0(n354), .S1(n350), .Y(n310) );
  MUX4X1 U2661 ( .D0(dpl_reg[37]), .D1(dpl_reg[45]), .D2(dpl_reg[53]), .D3(
        dpl_reg[61]), .S0(n354), .S1(n350), .Y(n309) );
  MUX4X1 U2662 ( .D0(dph_reg[33]), .D1(dph_reg[41]), .D2(dph_reg[49]), .D3(
        dph_reg[57]), .S0(n390), .S1(n394), .Y(n360) );
  MUX4X1 U2663 ( .D0(dph_reg[34]), .D1(dph_reg[42]), .D2(dph_reg[50]), .D3(
        dph_reg[58]), .S0(n390), .S1(n394), .Y(n362) );
  NAND21X1 U2664 ( .B(pdmode), .A(n2368), .Y(n2108) );
  MUX2AXL U2665 ( .D0(n2116), .D1(pdmode), .S(n2115), .Y(n2446) );
  GEN2XL U2666 ( .D(n2111), .E(n2110), .C(n2109), .B(n2389), .A(n561), .Y(
        n2116) );
  AO21X1 U2667 ( .B(n2113), .C(n2137), .A(n2112), .Y(n2114) );
  MUX4X1 U2668 ( .D0(dph_reg[1]), .D1(dph_reg[9]), .D2(dph_reg[17]), .D3(
        dph_reg[25]), .S0(n390), .S1(n394), .Y(n361) );
  MUX4X1 U2669 ( .D0(dph_reg[2]), .D1(dph_reg[10]), .D2(dph_reg[18]), .D3(
        dph_reg[26]), .S0(n390), .S1(n394), .Y(n363) );
  MUX4X1 U2670 ( .D0(dph_reg[35]), .D1(dph_reg[43]), .D2(dph_reg[51]), .D3(
        dph_reg[59]), .S0(n390), .S1(n394), .Y(n364) );
  MUX2XL U2671 ( .D0(ramsfraddr[6]), .D1(n2354), .S(waitstaten), .Y(
        ramsfraddr_comb[6]) );
  MUX2X1 U2672 ( .D0(n342), .D1(n341), .S(n349), .Y(dpc[3]) );
  MUX4X1 U2673 ( .D0(dpc_tab[3]), .D1(dpc_tab[9]), .D2(dpc_tab[15]), .D3(
        dpc_tab[21]), .S0(n357), .S1(n353), .Y(n342) );
  MUX4X1 U2674 ( .D0(dpc_tab[27]), .D1(dpc_tab[33]), .D2(dpc_tab[39]), .D3(
        dpc_tab[45]), .S0(n357), .S1(n353), .Y(n341) );
  AO21X1 U2675 ( .B(waitstaten), .C(n1083), .A(n557), .Y(N520) );
  MUX2X1 U2676 ( .D0(p2sel), .D1(n2335), .S(n1082), .Y(n1083) );
  MUX4X1 U2677 ( .D0(dph_reg[3]), .D1(dph_reg[11]), .D2(dph_reg[19]), .D3(
        dph_reg[27]), .S0(n390), .S1(n394), .Y(n365) );
  MUX4X1 U2678 ( .D0(dph_reg[36]), .D1(dph_reg[44]), .D2(dph_reg[52]), .D3(
        dph_reg[60]), .S0(n390), .S1(n394), .Y(n366) );
  MUX4X1 U2679 ( .D0(dph_reg[37]), .D1(dph_reg[45]), .D2(dph_reg[53]), .D3(
        dph_reg[61]), .S0(n390), .S1(n394), .Y(n368) );
  MUX2X1 U2680 ( .D0(n314), .D1(n313), .S(N351), .Y(dpl[3]) );
  MUX4X1 U2681 ( .D0(dpl_reg[3]), .D1(dpl_reg[11]), .D2(dpl_reg[19]), .D3(
        dpl_reg[27]), .S0(n354), .S1(n350), .Y(n314) );
  MUX4X1 U2682 ( .D0(dpl_reg[35]), .D1(dpl_reg[43]), .D2(dpl_reg[51]), .D3(
        dpl_reg[59]), .S0(n354), .S1(n350), .Y(n313) );
  MUX2X1 U2683 ( .D0(n330), .D1(n329), .S(n349), .Y(dph[3]) );
  MUX4X1 U2684 ( .D0(dph_reg[3]), .D1(dph_reg[11]), .D2(dph_reg[19]), .D3(
        dph_reg[27]), .S0(n356), .S1(n352), .Y(n330) );
  MUX4X1 U2685 ( .D0(dph_reg[35]), .D1(dph_reg[43]), .D2(dph_reg[51]), .D3(
        dph_reg[59]), .S0(n356), .S1(n352), .Y(n329) );
  MUX4X1 U2686 ( .D0(dph_reg[4]), .D1(dph_reg[12]), .D2(dph_reg[20]), .D3(
        dph_reg[28]), .S0(n390), .S1(n394), .Y(n367) );
  MUX4X1 U2687 ( .D0(dph_reg[5]), .D1(dph_reg[13]), .D2(dph_reg[21]), .D3(
        dph_reg[29]), .S0(n390), .S1(n394), .Y(n369) );
  MUX4XL U2688 ( .D0(dph_reg[38]), .D1(dph_reg[46]), .D2(dph_reg[54]), .D3(
        dph_reg[62]), .S0(n391), .S1(n395), .Y(n370) );
  MUX2XL U2689 ( .D0(ramsfraddr[7]), .D1(n66), .S(n2450), .Y(
        ramsfraddr_comb[7]) );
  MUX2XL U2690 ( .D0(ramsfraddr[4]), .D1(n2352), .S(waitstaten), .Y(
        ramsfraddr_comb[4]) );
  MUX2X1 U2691 ( .D0(n373), .D1(n372), .S(n153), .Y(N11845) );
  MUX4XL U2692 ( .D0(dph_reg[7]), .D1(dph_reg[15]), .D2(dph_reg[23]), .D3(
        dph_reg[31]), .S0(n391), .S1(n395), .Y(n373) );
  MUX4XL U2693 ( .D0(dph_reg[39]), .D1(dph_reg[47]), .D2(dph_reg[55]), .D3(
        dph_reg[63]), .S0(n391), .S1(n395), .Y(n372) );
  MUX2XL U2694 ( .D0(ramsfraddr[3]), .D1(n2351), .S(n2450), .Y(
        ramsfraddr_comb[3]) );
  NOR3XL U2695 ( .A(n1451), .B(n2001), .C(p2sel), .Y(n301) );
  MUX4XL U2696 ( .D0(dph_reg[6]), .D1(dph_reg[14]), .D2(dph_reg[22]), .D3(
        dph_reg[30]), .S0(n391), .S1(n395), .Y(n371) );
  NAND21XL U2697 ( .B(ramsfraddr[2]), .A(n1441), .Y(n2248) );
  NAND5XL U2698 ( .A(n509), .B(ramwe), .C(n2207), .D(n2206), .E(n2205), .Y(
        n2219) );
  MUX2XL U2699 ( .D0(ramsfraddr[5]), .D1(n74), .S(n2450), .Y(
        ramsfraddr_comb[5]) );
  AO2222XL U2700 ( .A(multemp2[7]), .B(n1519), .C(n215), .D(b[5]), .E(n1520), 
        .F(n2430), .G(n1521), .H(n1514), .Y(N12482) );
  AO2222XL U2701 ( .A(n215), .B(b[3]), .C(n1521), .D(n1516), .E(n1520), .F(
        n532), .G(multemp2[5]), .H(n1519), .Y(N12480) );
  AO2222XL U2702 ( .A(n215), .B(b[1]), .C(n1521), .D(n1518), .E(n512), .F(
        n1520), .G(multemp2[3]), .H(n1519), .Y(N12478) );
  AO2222XL U2703 ( .A(n215), .B(b[6]), .C(n1521), .D(n1529), .E(n1520), .F(
        n2434), .G(multemp2[8]), .H(n1519), .Y(N12483) );
  AO2222XL U2704 ( .A(n215), .B(b[4]), .C(n1521), .D(n1515), .E(n1520), .F(
        n2436), .G(multemp2[6]), .H(n1519), .Y(N12481) );
  AO2222XL U2705 ( .A(n215), .B(b[2]), .C(n1521), .D(n1517), .E(n1520), .F(
        n516), .G(multemp2[4]), .H(n1519), .Y(N12479) );
  AO2222XL U2706 ( .A(n215), .B(b[0]), .C(n1521), .D(n303), .E(n535), .F(n1520), .G(multemp2[2]), .H(n1519), .Y(N12477) );
  MUX2X1 U2707 ( .D0(gf0), .D1(n516), .S(n302), .Y(n1881) );
  MUX2X1 U2708 ( .D0(n2430), .D1(f0), .S(n2273), .Y(n1882) );
  MUX2X1 U2709 ( .D0(n512), .D1(f1), .S(n2273), .Y(n1883) );
  NAND32X1 U2710 ( .B(finishdiv), .C(n506), .A(n1498), .Y(n2201) );
  NAND21X1 U2711 ( .B(n1019), .A(n1018), .Y(N12721) );
  NAND21X1 U2712 ( .B(n554), .A(n1017), .Y(n1018) );
  NOR21XL U2713 ( .B(sfrdatai[7]), .A(n2020), .Y(n1019) );
  AO2222XL U2714 ( .A(n1016), .B(ramdatai[7]), .C(n2073), .D(n1015), .E(n1014), 
        .F(n75), .G(pc_o[15]), .H(n1013), .Y(n1017) );
  OAI221X1 U2715 ( .A(n1536), .B(n2190), .C(n2189), .D(n1535), .E(n569), .Y(
        N12489) );
  INVX1 U2716 ( .A(p2[4]), .Y(n1536) );
  OAI221X1 U2717 ( .A(n1952), .B(n2190), .C(n2189), .D(n1951), .E(n568), .Y(
        N12490) );
  INVX1 U2718 ( .A(p2[5]), .Y(n1952) );
  OAI221X1 U2719 ( .A(n1531), .B(n2190), .C(n2189), .D(n1582), .E(n569), .Y(
        N12488) );
  INVX1 U2720 ( .A(p2[3]), .Y(n1531) );
  OAI221X1 U2721 ( .A(n2024), .B(n2190), .C(n2189), .D(n2023), .E(n568), .Y(
        N12491) );
  INVX1 U2722 ( .A(p2[6]), .Y(n2024) );
  OAI221X1 U2723 ( .A(n2191), .B(n2190), .C(n2189), .D(n2188), .E(n568), .Y(
        N12492) );
  INVX1 U2724 ( .A(p2[7]), .Y(n2191) );
  OAI22XL U2725 ( .A(n1572), .B(n2285), .C(n2271), .D(n2023), .Y(N12706) );
  AOI22XL U2726 ( .A(n236), .B(n1571), .C(ac), .D(n1570), .Y(n1572) );
  NAND6XL U2727 ( .A(n1569), .B(n1568), .C(n1567), .D(n2301), .E(n1566), .F(
        n1565), .Y(n1570) );
  MUX2XL U2728 ( .D0(n300), .D1(dec_accop[10]), .S(n1563), .Y(n1571) );
  OAI22X1 U2729 ( .A(n1528), .B(n1527), .C(n2188), .D(n1526), .Y(N12484) );
  OA21X1 U2730 ( .B(n1525), .C(n2286), .A(n1524), .Y(n1528) );
  AOI33X1 U2731 ( .A(finishdiv), .B(n2294), .C(n1523), .D(multemp2[9]), .E(
        finishmul), .F(n1522), .Y(n1524) );
  MUX2XL U2732 ( .D0(N13352), .D1(n276), .S(N13353), .Y(n1523) );
  OAI31XL U2733 ( .A(dps[0]), .B(n545), .C(n2256), .D(n562), .Y(N12679) );
  AND2XL U2734 ( .A(phase0_ff), .B(n551), .Y(newinstr) );
  OA21X1 U2735 ( .B(n2037), .C(n2036), .A(n507), .Y(N12730) );
  AO2222XL U2736 ( .A(n2029), .B(n75), .C(n2028), .D(n2047), .E(intvect[4]), 
        .F(n2246), .G(n2027), .H(ramdatai[7]), .Y(n2037) );
  OAI221X1 U2737 ( .A(n2090), .B(n2035), .C(n2039), .D(n2034), .E(n2033), .Y(
        n2036) );
  OA222X1 U2738 ( .A(n2096), .B(n2032), .C(n50), .D(n2031), .E(n2059), .F(
        n2030), .Y(n2033) );
  OA21X1 U2739 ( .B(n1766), .C(n1765), .A(n507), .Y(N12728) );
  OAI221X1 U2740 ( .A(n1787), .B(n2035), .C(n1954), .D(n2034), .E(n1764), .Y(
        n1765) );
  AO2222XL U2741 ( .A(n2029), .B(memdatai[5]), .C(n2028), .D(n1763), .E(
        intvect[2]), .F(n2246), .G(n2027), .H(ramdatai[5]), .Y(n1766) );
  OA222X1 U2742 ( .A(n1789), .B(n2032), .C(n44), .D(n2031), .E(n1776), .F(
        n2030), .Y(n1764) );
  OA21X1 U2743 ( .B(n1545), .C(n1544), .A(n507), .Y(N12727) );
  OAI221X1 U2744 ( .A(n1817), .B(n2035), .C(n1824), .D(n2034), .E(n1543), .Y(
        n1544) );
  AO2222XL U2745 ( .A(n2029), .B(memdatai[4]), .C(n2028), .D(n1542), .E(
        intvect[1]), .F(n2246), .G(n2027), .H(ramdatai[4]), .Y(n1545) );
  OA222X1 U2746 ( .A(n1819), .B(n2032), .C(n34), .D(n2031), .E(n1809), .F(
        n2030), .Y(n1543) );
  OA21X1 U2747 ( .B(n1559), .C(n1558), .A(n507), .Y(N12726) );
  OAI221X1 U2748 ( .A(n1677), .B(n2035), .C(n1557), .D(n2034), .E(n1556), .Y(
        n1558) );
  AO2222XL U2749 ( .A(n2029), .B(n58), .C(n2028), .D(n1553), .E(intvect[0]), 
        .F(n2246), .G(n2027), .H(ramdatai[3]), .Y(n1559) );
  OA222X1 U2750 ( .A(n1555), .B(n2032), .C(n54), .D(n2031), .E(n1554), .F(
        n2030), .Y(n1556) );
  OA21X1 U2751 ( .B(n2011), .C(n2010), .A(n507), .Y(N12729) );
  OAI221X1 U2752 ( .A(n2009), .B(n2035), .C(n2013), .D(n2034), .E(n2008), .Y(
        n2010) );
  AO2222XL U2753 ( .A(n2029), .B(n59), .C(n2028), .D(n2005), .E(intvect[3]), 
        .F(n2246), .G(n2027), .H(ramdatai[6]), .Y(n2011) );
  OA222X1 U2754 ( .A(n2007), .B(n2032), .C(n36), .D(n2031), .E(n2006), .F(
        n2030), .Y(n2008) );
  NOR32XL U2755 ( .B(n509), .C(n497), .A(newinstrlock), .Y(N689) );
  AND2X1 U2756 ( .A(n2134), .B(n127), .Y(N681) );
  AND2X1 U2757 ( .A(state[1]), .B(n501), .Y(N589) );
  AND2X1 U2758 ( .A(n2134), .B(phase[2]), .Y(N682) );
  AND2X1 U2759 ( .A(n2134), .B(phase[3]), .Y(N683) );
  AND2X1 U2760 ( .A(n2134), .B(phase[4]), .Y(N684) );
  AND2X1 U2761 ( .A(state[2]), .B(n501), .Y(N590) );
  INVX1 U2762 ( .A(temp[7]), .Y(n2059) );
  MUX4X1 U2763 ( .D0(dph_reg[7]), .D1(dph_reg[15]), .D2(dph_reg[23]), .D3(
        dph_reg[31]), .S0(n355), .S1(n351), .Y(n322) );
  MUX4X1 U2764 ( .D0(dpl_reg[7]), .D1(dpl_reg[15]), .D2(dpl_reg[23]), .D3(
        dpl_reg[31]), .S0(dps[0]), .S1(N350), .Y(n306) );
  MUX4X1 U2765 ( .D0(dph_reg[39]), .D1(dph_reg[47]), .D2(dph_reg[55]), .D3(
        dph_reg[63]), .S0(n355), .S1(n351), .Y(n321) );
  MUX4X1 U2766 ( .D0(dpl_reg[38]), .D1(dpl_reg[46]), .D2(dpl_reg[54]), .D3(
        dpl_reg[62]), .S0(N349), .S1(N350), .Y(n307) );
  MUX4X1 U2767 ( .D0(dpl_reg[39]), .D1(dpl_reg[47]), .D2(dpl_reg[55]), .D3(
        dpl_reg[63]), .S0(dps[0]), .S1(dps[1]), .Y(n305) );
  MUX2X1 U2768 ( .D0(n338), .D1(n337), .S(n349), .Y(dpc[5]) );
  MUX4X1 U2769 ( .D0(dpc_tab[5]), .D1(dpc_tab[11]), .D2(dpc_tab[17]), .D3(
        dpc_tab[23]), .S0(n356), .S1(n352), .Y(n338) );
  MUX4X1 U2770 ( .D0(dpc_tab[29]), .D1(dpc_tab[35]), .D2(dpc_tab[41]), .D3(
        dpc_tab[47]), .S0(n356), .S1(n352), .Y(n337) );
  MUX2X1 U2771 ( .D0(n340), .D1(n339), .S(n349), .Y(dpc[4]) );
  MUX4X1 U2772 ( .D0(dpc_tab[4]), .D1(dpc_tab[10]), .D2(dpc_tab[16]), .D3(
        dpc_tab[22]), .S0(n357), .S1(n353), .Y(n340) );
  MUX4X1 U2773 ( .D0(dpc_tab[28]), .D1(dpc_tab[34]), .D2(dpc_tab[40]), .D3(
        dpc_tab[46]), .S0(n357), .S1(n353), .Y(n339) );
  NOR2X1 U2774 ( .A(n1025), .B(n1024), .Y(N12975) );
  XNOR2XL U2775 ( .A(waitcnt[1]), .B(waitcnt[0]), .Y(n1025) );
  NOR2X1 U2776 ( .A(waitcnt[0]), .B(n1024), .Y(N12974) );
  NOR2X1 U2777 ( .A(n1023), .B(n1024), .Y(N12976) );
  AOI21X1 U2778 ( .B(waitcnt[0]), .C(waitcnt[1]), .A(waitcnt[2]), .Y(n1023) );
  NAND5XL U2779 ( .A(n1439), .B(n2233), .C(n2205), .D(ramsfraddr[5]), .E(n1438), .Y(n2189) );
  AOI32XL U2780 ( .A(n236), .B(n2302), .C(n2301), .D(ov), .E(n2300), .Y(n2303)
         );
  NAND43X1 U2781 ( .B(n2299), .C(n2298), .D(n2297), .A(n2296), .Y(n2300) );
  XOR2XL U2782 ( .A(n261), .B(n231), .Y(n2302) );
  INVX1 U2783 ( .A(n2301), .Y(n2298) );
  MUX2BXL U2784 ( .D0(N13345), .D1(n1921), .S(N13353), .Y(n303) );
  INVX1 U2785 ( .A(stop), .Y(n1849) );
  AOI21BX1 U2786 ( .C(cpu_hold), .B(d_hold), .A(cpu_resume_fff), .Y(n726) );
  INVX1 U2787 ( .A(n1705), .Y(n1759) );
  OAI211X1 U2788 ( .C(n1873), .D(n108), .A(n1703), .B(n1702), .Y(n1705) );
  OA22X1 U2789 ( .A(add_5280_3_carry_9_), .B(n1701), .C(add_5280_4_carry[9]), 
        .D(n1700), .Y(n1702) );
  MUX2X1 U2790 ( .D0(n1699), .D1(n1698), .S(memaddr[8]), .Y(n1703) );
  INVX1 U2791 ( .A(memaddr[10]), .Y(n1901) );
  INVX1 U2792 ( .A(n1636), .Y(n1729) );
  OAI211X1 U2793 ( .C(n1818), .D(n108), .A(n1635), .B(n1634), .Y(n1636) );
  OA222X1 U2794 ( .A(n1828), .B(n1656), .C(n1633), .D(n34), .E(n1632), .F(
        n1700), .Y(n1634) );
  AOI221XL U2795 ( .A(n1697), .B(n1631), .C(n1693), .D(pc_o[3]), .E(n1637), 
        .Y(n1633) );
  INVX1 U2796 ( .A(n1618), .Y(n1725) );
  OAI211X1 U2797 ( .C(n1940), .D(n108), .A(n1617), .B(n1616), .Y(n1618) );
  OA222X1 U2798 ( .A(n1941), .B(n1656), .C(n1615), .D(n36), .E(n1614), .F(
        n1700), .Y(n1616) );
  AOI221XL U2799 ( .A(n1697), .B(n1613), .C(n1693), .D(memaddr[5]), .E(n1620), 
        .Y(n1615) );
  AOI221XL U2800 ( .A(n104), .B(n1696), .C(n1695), .D(n2200), .E(n1694), .Y(
        n1698) );
  AO21X1 U2801 ( .B(n1693), .C(memaddr[7]), .A(n1692), .Y(n1694) );
  INVX1 U2802 ( .A(p2[1]), .Y(n1469) );
  INVX1 U2803 ( .A(p2[0]), .Y(n1453) );
  INVX1 U2804 ( .A(p2[2]), .Y(n1890) );
  AND2XL U2805 ( .A(b[7]), .B(acc[1]), .Y(N14351) );
  AND2XL U2806 ( .A(b[2]), .B(acc[1]), .Y(N14346) );
  AND2XL U2807 ( .A(b[4]), .B(acc[0]), .Y(N14340) );
  AND2XL U2808 ( .A(b[3]), .B(acc[1]), .Y(N14347) );
  AND2XL U2809 ( .A(b[5]), .B(acc[0]), .Y(N14341) );
  AND2XL U2810 ( .A(b[4]), .B(acc[1]), .Y(N14348) );
  AND2XL U2811 ( .A(b[6]), .B(acc[0]), .Y(N14342) );
  AND2XL U2812 ( .A(b[5]), .B(acc[1]), .Y(N14349) );
  AND2XL U2813 ( .A(b[6]), .B(acc[1]), .Y(N14350) );
  AND2XL U2814 ( .A(b[1]), .B(acc[1]), .Y(N14345) );
  AND2XL U2815 ( .A(b[2]), .B(acc[0]), .Y(N14338) );
  AND2XL U2816 ( .A(b[3]), .B(acc[0]), .Y(N14339) );
  AND2XL U2817 ( .A(b[7]), .B(acc[0]), .Y(N14343) );
  AO21XL U2818 ( .B(n1693), .C(pc_o[0]), .A(n1661), .Y(n1657) );
  AOI21BX1 U2819 ( .C(n108), .B(pc_i[1]), .A(n1659), .Y(n304) );
  INVX1 U2820 ( .A(n1648), .Y(n1731) );
  OAI211X1 U2821 ( .C(n1647), .D(n108), .A(n1646), .B(n1645), .Y(n1648) );
  AOI22X1 U2822 ( .A(n104), .B(n1644), .C(n1695), .D(n1643), .Y(n1645) );
  INVX1 U2823 ( .A(n1629), .Y(n1727) );
  OAI211X1 U2824 ( .C(n1788), .D(n108), .A(n1628), .B(n1627), .Y(n1629) );
  AOI22X1 U2825 ( .A(n104), .B(n1626), .C(n101), .D(n1625), .Y(n1627) );
  MUX2X1 U2826 ( .D0(n1635), .D1(n1621), .S(memaddr[5]), .Y(n1628) );
  INVX1 U2827 ( .A(n1610), .Y(n1724) );
  OAI211X1 U2828 ( .C(n2092), .D(n108), .A(n1609), .B(n1608), .Y(n1610) );
  AOI22X1 U2829 ( .A(n104), .B(n1607), .C(n101), .D(n1606), .Y(n1608) );
  MUX2X1 U2830 ( .D0(n1617), .D1(n1601), .S(pc_o[7]), .Y(n1609) );
  INVX1 U2831 ( .A(n1688), .Y(n1750) );
  OAI221X1 U2832 ( .A(n1687), .B(n48), .C(n1686), .D(n1704), .E(n1685), .Y(
        n1688) );
  AOI222XL U2833 ( .A(N11787), .B(n1695), .C(N11804), .D(n1693), .E(N11821), 
        .F(n1697), .Y(n1685) );
  INVX1 U2834 ( .A(n1681), .Y(n1748) );
  OAI221X1 U2835 ( .A(n1687), .B(n1901), .C(n1916), .D(n1704), .E(n1680), .Y(
        n1681) );
  AOI222XL U2836 ( .A(N11788), .B(n1695), .C(N11805), .D(n1693), .E(N11822), 
        .F(n1697), .Y(n1680) );
  INVX1 U2837 ( .A(n1678), .Y(n1746) );
  OAI221X1 U2838 ( .A(n1687), .B(n52), .C(n1677), .D(n1704), .E(n1676), .Y(
        n1678) );
  AOI222XL U2839 ( .A(N11789), .B(n1695), .C(N11806), .D(n1693), .E(N11823), 
        .F(n1697), .Y(n1676) );
  INVX1 U2840 ( .A(n1675), .Y(n1744) );
  OAI221X1 U2841 ( .A(n1687), .B(n1827), .C(n1817), .D(n1704), .E(n1674), .Y(
        n1675) );
  AOI222XL U2842 ( .A(N11790), .B(n1695), .C(N11807), .D(n135), .E(N11824), 
        .F(n1697), .Y(n1674) );
  INVX1 U2843 ( .A(n1673), .Y(n1742) );
  OAI221X1 U2844 ( .A(n1687), .B(n1955), .C(n1787), .D(n1704), .E(n1672), .Y(
        n1673) );
  AOI222XL U2845 ( .A(N11791), .B(n1695), .C(N11808), .D(n135), .E(N11825), 
        .F(n1697), .Y(n1672) );
  INVX1 U2846 ( .A(n1671), .Y(n1740) );
  OAI221X1 U2847 ( .A(n1687), .B(n2015), .C(n2009), .D(n1704), .E(n1670), .Y(
        n1671) );
  AOI222XL U2848 ( .A(N11792), .B(n1695), .C(N11809), .D(n135), .E(N11826), 
        .F(n1697), .Y(n1670) );
  INVX1 U2849 ( .A(n1669), .Y(n1738) );
  OAI221X1 U2850 ( .A(n1687), .B(n38), .C(n2090), .D(n1704), .E(n1668), .Y(
        n1669) );
  AOI222XL U2851 ( .A(N11793), .B(n1695), .C(N11810), .D(n135), .E(N11827), 
        .F(n1697), .Y(n1668) );
  MUX2IXL U2852 ( .D0(n1664), .D1(n1663), .S(pc_o[0]), .Y(n1736) );
  NAND21X1 U2853 ( .B(n135), .A(n1704), .Y(n1664) );
  NAND21X1 U2854 ( .B(n1662), .A(n1687), .Y(n1663) );
  NAND21X1 U2855 ( .B(memaddr[4]), .A(n1640), .Y(n1632) );
  NAND21X1 U2856 ( .B(memaddr[6]), .A(n1622), .Y(n1614) );
  OR2X1 U2857 ( .A(memaddr[7]), .B(n1614), .Y(n1696) );
  XOR2XL U2858 ( .A(n32), .B(pc_o[1]), .Y(n1903) );
  NAND21XL U2859 ( .B(pc_o[1]), .A(n32), .Y(n1641) );
  OR2X1 U2860 ( .A(pc_o[5]), .B(n1632), .Y(n1613) );
  NAND21XL U2861 ( .B(pc_o[0]), .A(n1602), .Y(n1650) );
  NAND32X1 U2862 ( .B(pc_o[7]), .C(n1689), .A(n40), .Y(add_5280_3_carry_9_) );
  NAND32X1 U2863 ( .B(memaddr[5]), .C(n1619), .A(n36), .Y(n1689) );
  NAND21X1 U2864 ( .B(pc_o[8]), .A(n1690), .Y(add_5280_4_carry[9]) );
  INVX1 U2865 ( .A(n1084), .Y(cs_run) );
  NAND21X1 U2866 ( .B(n2364), .A(state[0]), .Y(n1084) );
  INVX1 U2867 ( .A(temp[5]), .Y(n1776) );
  INVX1 U2868 ( .A(N345), .Y(n1779) );
  INVX1 U2869 ( .A(stop_r), .Y(n2113) );
  NAND21XL U2870 ( .B(n32), .A(pc_o[1]), .Y(n1649) );
  AO21X1 U2871 ( .B(n127), .C(n1012), .A(n1011), .Y(n2245) );
  XOR2X1 U2872 ( .A(n1605), .B(pc_o[7]), .Y(n2095) );
  NAND21X1 U2873 ( .B(n36), .A(n1691), .Y(n1605) );
  OAI31XL U2874 ( .A(n1345), .B(n1344), .C(n1343), .D(phase[0]), .Y(n2034) );
  GEN2XL U2875 ( .D(instr[2]), .E(n1342), .C(n2314), .B(n1341), .A(n1340), .Y(
        n1343) );
  XOR2X1 U2876 ( .A(n1612), .B(memaddr[6]), .Y(n1941) );
  XOR2X1 U2877 ( .A(n1630), .B(pc_o[4]), .Y(n1828) );
  XOR2X1 U2878 ( .A(n1624), .B(pc_o[5]), .Y(n1790) );
  NAND21X1 U2879 ( .B(n34), .A(n1623), .Y(n1624) );
  AOI32XL U2880 ( .A(n1329), .B(instr[2]), .C(n103), .D(n1432), .E(n30), .Y(
        n1330) );
  INVX1 U2881 ( .A(temp[6]), .Y(n2006) );
  NOR21XL U2882 ( .B(n2322), .A(n981), .Y(n2019) );
  NOR43XL U2883 ( .B(n2017), .C(n127), .D(n1012), .A(ramsfraddr[7]), .Y(n981)
         );
  NAND5XL U2884 ( .A(ramsfraddr[7]), .B(n127), .C(n564), .D(n980), .E(n1012), 
        .Y(n2020) );
  INVX1 U2885 ( .A(n1011), .Y(n980) );
  INVX1 U2886 ( .A(memaddr[13]), .Y(n1955) );
  INVX1 U2887 ( .A(memaddr[12]), .Y(n1827) );
  INVX1 U2888 ( .A(memaddr[14]), .Y(n2015) );
  INVX1 U2889 ( .A(n2170), .Y(n2180) );
  OAI211X1 U2890 ( .C(n2169), .D(n2168), .A(n2167), .B(n2166), .Y(n2170) );
  AO21X1 U2891 ( .B(n1347), .C(n127), .A(n1346), .Y(n1350) );
  AO21X1 U2892 ( .B(pc_o[7]), .C(n1614), .A(n1690), .Y(n1607) );
  GEN2XL U2893 ( .D(n2147), .E(n111), .C(n979), .B(n978), .A(n1838), .Y(n1012)
         );
  AND2XL U2894 ( .A(n30), .B(instr[5]), .Y(n979) );
  NAND21XL U2895 ( .B(dec_accop[10]), .A(dec_accop[9]), .Y(n2301) );
  AO21X1 U2896 ( .B(pc_o[5]), .C(n1632), .A(n1622), .Y(n1626) );
  OAI22XL U2897 ( .A(n2186), .B(n1949), .C(n1948), .D(n2185), .Y(N12968) );
  INVX1 U2898 ( .A(ckcon[3]), .Y(n1949) );
  OAI22X1 U2899 ( .A(n2186), .B(n1950), .C(n2344), .D(n2185), .Y(N12972) );
  INVX1 U2900 ( .A(ckcon[7]), .Y(n1950) );
  NAND43X1 U2901 ( .B(ramsfraddr[4]), .C(n1946), .D(n2249), .A(ramsfraddr[3]), 
        .Y(n1947) );
  AND2X1 U2902 ( .A(cpu_resume_ff1), .B(n563), .Y(N13380) );
  INVXL U2903 ( .A(b[4]), .Y(n2288) );
  INVXL U2904 ( .A(b[2]), .Y(n2287) );
  INVXL U2905 ( .A(b[7]), .Y(n2286) );
  INVXL U2906 ( .A(b[1]), .Y(n2290) );
  INVXL U2907 ( .A(b[6]), .Y(n2291) );
  INVXL U2908 ( .A(b[5]), .Y(n2293) );
  INVXL U2909 ( .A(b[3]), .Y(n2292) );
  INVX1 U2910 ( .A(finishmul), .Y(n2204) );
  INVX1 U2911 ( .A(finishdiv), .Y(n2202) );
  INVX1 U2912 ( .A(n2213), .Y(n2229) );
  NAND32XL U2913 ( .B(ramsfraddr[0]), .C(n2212), .A(n2211), .Y(n2213) );
  NAND21XL U2914 ( .B(n89), .A(n912), .Y(n2104) );
  NAND21X1 U2915 ( .B(n903), .A(n1773), .Y(n905) );
  OAI211X1 U2916 ( .C(n1485), .D(n2038), .A(n941), .B(n940), .Y(n2274) );
  OAI32X1 U2917 ( .A(n85), .B(n1868), .C(n905), .D(n904), .E(n905), .Y(n908)
         );
  OAI211XL U2918 ( .C(n1868), .D(n1914), .A(n56), .B(n64), .Y(n1870) );
  OAI22XL U2919 ( .A(n554), .B(n1457), .C(n98), .D(n2020), .Y(N12714) );
  NAND21XL U2920 ( .B(n93), .A(n911), .Y(n912) );
  MAJ3XL U2921 ( .A(n2077), .B(n1064), .C(n1063), .Y(n1902) );
  NOR21X1 U2922 ( .B(n2384), .A(n2385), .Y(n2403) );
  NAND42X4 U2923 ( .C(n866), .D(idle_r), .A(n865), .B(n864), .Y(n867) );
  MAJ3X1 U2924 ( .A(n1034), .B(n1033), .C(n1032), .Y(n1035) );
  MAJ3X1 U2925 ( .A(n2077), .B(n1902), .C(n249), .Y(n1794) );
  GEN2X1 U2926 ( .D(n1845), .E(n1222), .C(n1217), .B(n1216), .A(n1215), .Y(
        n1243) );
  MAJ3X1 U2927 ( .A(n2077), .B(n1795), .C(n1794), .Y(n1823) );
  MAJ3X1 U2928 ( .A(n2077), .B(n1796), .C(n1823), .Y(n1936) );
  MAJ3X1 U2929 ( .A(n2077), .B(n1937), .C(n1936), .Y(n2076) );
  MAJ3X1 U2930 ( .A(n2077), .B(n2076), .C(n250), .Y(n2083) );
  XNOR2XL U2931 ( .A(pc_o[15]), .B(add_5280_3_carry_15_), .Y(N11810) );
  OR2X1 U2932 ( .A(add_5280_3_carry_14_), .B(pc_o[14]), .Y(
        add_5280_3_carry_15_) );
  XNOR2XL U2933 ( .A(add_5280_3_carry_14_), .B(pc_o[14]), .Y(N11809) );
  OR2X1 U2934 ( .A(add_5280_3_carry_13_), .B(pc_o[13]), .Y(
        add_5280_3_carry_14_) );
  XNOR2XL U2935 ( .A(add_5280_3_carry_13_), .B(pc_o[13]), .Y(N11808) );
  OR2X1 U2936 ( .A(add_5280_3_carry_12_), .B(pc_o[12]), .Y(
        add_5280_3_carry_13_) );
  XNOR2XL U2937 ( .A(add_5280_3_carry_12_), .B(pc_o[12]), .Y(N11807) );
  OR2X1 U2938 ( .A(add_5280_3_carry_11_), .B(pc_o[11]), .Y(
        add_5280_3_carry_12_) );
  XNOR2XL U2939 ( .A(add_5280_3_carry_11_), .B(pc_o[11]), .Y(N11806) );
  OR2X1 U2940 ( .A(add_5280_3_carry_10_), .B(pc_o[10]), .Y(
        add_5280_3_carry_11_) );
  XNOR2XL U2941 ( .A(add_5280_3_carry_10_), .B(pc_o[10]), .Y(N11805) );
  OR2X1 U2942 ( .A(add_5280_3_carry_9_), .B(memaddr[9]), .Y(
        add_5280_3_carry_10_) );
  XNOR2XL U2943 ( .A(add_5280_3_carry_9_), .B(memaddr[9]), .Y(N11804) );
  XNOR2XL U2944 ( .A(pc_o[15]), .B(add_5280_4_carry[15]), .Y(N11827) );
  OR2X1 U2945 ( .A(add_5280_4_carry[14]), .B(pc_o[14]), .Y(
        add_5280_4_carry[15]) );
  XNOR2XL U2946 ( .A(add_5280_4_carry[14]), .B(pc_o[14]), .Y(N11826) );
  OR2X1 U2947 ( .A(add_5280_4_carry[13]), .B(pc_o[13]), .Y(
        add_5280_4_carry[14]) );
  XNOR2XL U2948 ( .A(add_5280_4_carry[13]), .B(pc_o[13]), .Y(N11825) );
  OR2X1 U2949 ( .A(add_5280_4_carry[12]), .B(pc_o[12]), .Y(
        add_5280_4_carry[13]) );
  XNOR2XL U2950 ( .A(add_5280_4_carry[12]), .B(pc_o[12]), .Y(N11824) );
  OR2X1 U2951 ( .A(add_5280_4_carry[11]), .B(memaddr[11]), .Y(
        add_5280_4_carry[12]) );
  XNOR2XL U2952 ( .A(add_5280_4_carry[11]), .B(memaddr[11]), .Y(N11823) );
  OR2X1 U2953 ( .A(add_5280_4_carry[10]), .B(pc_o[10]), .Y(
        add_5280_4_carry[11]) );
  XNOR2XL U2954 ( .A(add_5280_4_carry[10]), .B(pc_o[10]), .Y(N11822) );
  OR2X1 U2955 ( .A(add_5280_4_carry[9]), .B(pc_o[9]), .Y(add_5280_4_carry[10])
         );
  XNOR2XL U2956 ( .A(add_5280_4_carry[9]), .B(pc_o[9]), .Y(N11821) );
  XOR2X1 U2957 ( .A(pc_o[15]), .B(add_5280_2_carry[15]), .Y(N11793) );
  AND2X1 U2958 ( .A(pc_o[14]), .B(add_5280_2_carry[14]), .Y(
        add_5280_2_carry[15]) );
  XOR2X1 U2959 ( .A(add_5280_2_carry[14]), .B(pc_o[14]), .Y(N11792) );
  AND2X1 U2960 ( .A(pc_o[13]), .B(add_5280_2_carry[13]), .Y(
        add_5280_2_carry[14]) );
  XOR2X1 U2961 ( .A(add_5280_2_carry[13]), .B(pc_o[13]), .Y(N11791) );
  AND2X1 U2962 ( .A(pc_o[12]), .B(add_5280_2_carry[12]), .Y(
        add_5280_2_carry[13]) );
  XOR2X1 U2963 ( .A(add_5280_2_carry[12]), .B(pc_o[12]), .Y(N11790) );
  AND2X1 U2964 ( .A(pc_o[11]), .B(add_5280_2_carry[11]), .Y(
        add_5280_2_carry[12]) );
  XOR2X1 U2965 ( .A(add_5280_2_carry[11]), .B(pc_o[11]), .Y(N11789) );
  AND2X1 U2966 ( .A(pc_o[10]), .B(add_5280_2_carry[10]), .Y(
        add_5280_2_carry[11]) );
  XOR2X1 U2967 ( .A(add_5280_2_carry[10]), .B(pc_o[10]), .Y(N11788) );
  AND2X1 U2968 ( .A(pc_o[9]), .B(n257), .Y(add_5280_2_carry[10]) );
  XOR2X1 U2969 ( .A(n257), .B(pc_o[9]), .Y(N11787) );
endmodule


module mcu51_cpu_a0_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n15, n16, n17, n18, n19,
         n23, n24, n25, n26, n27, n28, n29, n30, n63;

  FAD1X1 U3 ( .A(n24), .B(A[6]), .CI(n6), .CO(n5), .SO(DIFF[6]) );
  FAD1X1 U4 ( .A(n25), .B(A[5]), .CI(n7), .CO(n6), .SO(DIFF[5]) );
  FAD1X1 U5 ( .A(n26), .B(A[4]), .CI(n8), .CO(n7), .SO(DIFF[4]) );
  OAI21X1 U7 ( .B(n11), .C(n9), .A(n10), .Y(n8) );
  NOR2X1 U10 ( .A(n27), .B(A[3]), .Y(n9) );
  XOR2X1 U20 ( .A(n3), .B(n19), .Y(DIFF[1]) );
  OAI21X1 U21 ( .B(n17), .C(n19), .A(n18), .Y(n16) );
  NOR2X1 U24 ( .A(n29), .B(A[1]), .Y(n17) );
  INVX1 U39 ( .A(B[4]), .Y(n26) );
  INVX1 U40 ( .A(B[3]), .Y(n27) );
  INVX1 U41 ( .A(B[5]), .Y(n25) );
  XNOR2XL U42 ( .A(n2), .B(n16), .Y(DIFF[2]) );
  XNOR2XL U43 ( .A(A[0]), .B(n30), .Y(DIFF[0]) );
  OR2X1 U44 ( .A(n28), .B(A[2]), .Y(n63) );
  XOR2XL U45 ( .A(n11), .B(n1), .Y(DIFF[3]) );
  NOR2X2 U46 ( .A(n30), .B(A[0]), .Y(n19) );
  INVX1 U47 ( .A(B[6]), .Y(n24) );
  INVX2 U48 ( .A(n4), .Y(DIFF[8]) );
  NAND2X1 U49 ( .A(n29), .B(A[1]), .Y(n18) );
  NAND2XL U50 ( .A(n28), .B(A[2]), .Y(n15) );
  AOI21AX1 U51 ( .B(n16), .C(n63), .A(n15), .Y(n11) );
  NAND2X1 U52 ( .A(n63), .B(n15), .Y(n2) );
  NAND21XL U53 ( .B(n17), .A(n18), .Y(n3) );
  NAND21XL U54 ( .B(n9), .A(n10), .Y(n1) );
  MAJ3X1 U55 ( .A(n23), .B(A[7]), .C(n5), .Y(n4) );
  INVX1 U56 ( .A(B[7]), .Y(n23) );
  INVX3 U57 ( .A(B[1]), .Y(n29) );
  INVX3 U58 ( .A(B[2]), .Y(n28) );
  INVX3 U59 ( .A(B[0]), .Y(n30) );
  NAND2XL U60 ( .A(n27), .B(A[3]), .Y(n10) );
endmodule


module mcu51_cpu_a0_DW01_add_10 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n24, n25, n26, n27, n28, n29, n81;

  XOR2X1 U2 ( .A(A[8]), .B(B[15]), .Y(n1) );
  FAD1X1 U3 ( .A(B[14]), .B(A[8]), .CI(n7), .CO(n6), .SO(SUM[14]) );
  FAD1X1 U4 ( .A(B[13]), .B(A[8]), .CI(n8), .CO(n7), .SO(SUM[13]) );
  FAD1X1 U5 ( .A(B[12]), .B(A[8]), .CI(n9), .CO(n8), .SO(SUM[12]) );
  FAD1X1 U6 ( .A(B[11]), .B(A[8]), .CI(n10), .CO(n9), .SO(SUM[11]) );
  FAD1X1 U7 ( .A(B[10]), .B(A[8]), .CI(n11), .CO(n10), .SO(SUM[10]) );
  FAD1X1 U8 ( .A(B[9]), .B(A[8]), .CI(n12), .CO(n11), .SO(SUM[9]) );
  FAD1X1 U9 ( .A(B[8]), .B(A[8]), .CI(n13), .CO(n12), .SO(SUM[8]) );
  FAD1X1 U10 ( .A(B[7]), .B(A[7]), .CI(n14), .CO(n13), .SO(SUM[7]) );
  FAD1X1 U11 ( .A(B[6]), .B(A[6]), .CI(n15), .CO(n14), .SO(SUM[6]) );
  FAD1X1 U12 ( .A(B[5]), .B(A[5]), .CI(n16), .CO(n15), .SO(SUM[5]) );
  FAD1X1 U13 ( .A(B[4]), .B(A[4]), .CI(n17), .CO(n16), .SO(SUM[4]) );
  XOR2X1 U14 ( .A(n20), .B(n2), .Y(SUM[3]) );
  OAI21X1 U15 ( .B(n20), .C(n18), .A(n19), .Y(n17) );
  NOR2X1 U18 ( .A(B[3]), .B(A[3]), .Y(n18) );
  XOR2X1 U28 ( .A(n29), .B(n4), .Y(SUM[1]) );
  OAI21X1 U29 ( .B(n29), .C(n26), .A(n27), .Y(n25) );
  NOR2X1 U32 ( .A(A[1]), .B(B[1]), .Y(n26) );
  NOR2X1 U37 ( .A(A[0]), .B(B[0]), .Y(n28) );
  NAND2XL U42 ( .A(n81), .B(n24), .Y(n3) );
  NAND21XL U43 ( .B(n26), .A(n27), .Y(n4) );
  NAND21XL U44 ( .B(n28), .A(n29), .Y(n5) );
  NAND2XL U45 ( .A(B[3]), .B(A[3]), .Y(n19) );
  AOI21AX1 U46 ( .B(n25), .C(n81), .A(n24), .Y(n20) );
  XNOR2XL U47 ( .A(n3), .B(n25), .Y(SUM[2]) );
  NAND21XL U48 ( .B(n18), .A(n19), .Y(n2) );
  NAND2X1 U49 ( .A(A[0]), .B(B[0]), .Y(n29) );
  NAND2X1 U50 ( .A(B[2]), .B(A[2]), .Y(n24) );
  OR2X1 U51 ( .A(B[2]), .B(A[2]), .Y(n81) );
  NAND2X1 U52 ( .A(A[1]), .B(B[1]), .Y(n27) );
  INVX1 U53 ( .A(n5), .Y(SUM[0]) );
  XOR2X1 U54 ( .A(n6), .B(n1), .Y(SUM[15]) );
endmodule


module mcu51_cpu_a0_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n15, n16, n17, n18, n19,
         n23, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n74, n75;

  FAD1X1 U2 ( .A(A[7]), .B(n33), .CI(n7), .CO(n6), .SO(DIFF[7]) );
  FAD1X1 U3 ( .A(A[6]), .B(n34), .CI(n8), .CO(n7), .SO(DIFF[6]) );
  OAI21X1 U5 ( .B(n11), .C(n9), .A(n10), .Y(n8) );
  NOR2X1 U8 ( .A(A[5]), .B(n35), .Y(n9) );
  OAI21X1 U19 ( .B(n19), .C(n17), .A(n18), .Y(n16) );
  NOR2X1 U22 ( .A(A[3]), .B(n37), .Y(n17) );
  XOR2X1 U32 ( .A(n5), .B(n27), .Y(DIFF[1]) );
  OAI21X1 U33 ( .B(n25), .C(n27), .A(n26), .Y(n24) );
  NOR2X1 U39 ( .A(n40), .B(A[0]), .Y(n27) );
  OR2X1 U51 ( .A(A[4]), .B(n36), .Y(n75) );
  XNOR2XL U52 ( .A(A[0]), .B(n40), .Y(DIFF[0]) );
  XOR2XL U53 ( .A(n19), .B(n3), .Y(DIFF[3]) );
  XOR2XL U54 ( .A(n11), .B(n1), .Y(DIFF[5]) );
  NAND2XL U55 ( .A(A[1]), .B(n39), .Y(n26) );
  NOR2XL U56 ( .A(A[1]), .B(n39), .Y(n25) );
  NAND2XL U57 ( .A(A[3]), .B(n37), .Y(n18) );
  NAND2XL U58 ( .A(A[5]), .B(n35), .Y(n10) );
  NAND2XL U59 ( .A(A[4]), .B(n36), .Y(n15) );
  INVXL U60 ( .A(n17), .Y(n30) );
  NAND2XL U61 ( .A(n30), .B(n18), .Y(n3) );
  INVXL U62 ( .A(n9), .Y(n28) );
  NAND2XL U63 ( .A(n28), .B(n10), .Y(n1) );
  AOI21AX1 U64 ( .B(n16), .C(n75), .A(n15), .Y(n11) );
  AOI21AX1 U65 ( .B(n24), .C(n74), .A(n23), .Y(n19) );
  INVX2 U66 ( .A(n6), .Y(DIFF[8]) );
  OR2X1 U67 ( .A(A[2]), .B(n38), .Y(n74) );
  NAND2X1 U68 ( .A(A[2]), .B(n38), .Y(n23) );
  NAND2X1 U69 ( .A(n32), .B(n26), .Y(n5) );
  INVX1 U70 ( .A(n25), .Y(n32) );
  XNOR2XL U71 ( .A(n2), .B(n16), .Y(DIFF[4]) );
  NAND2XL U72 ( .A(n75), .B(n15), .Y(n2) );
  XNOR2XL U73 ( .A(n4), .B(n24), .Y(DIFF[2]) );
  NAND2XL U74 ( .A(n74), .B(n23), .Y(n4) );
  INVX1 U75 ( .A(B[7]), .Y(n33) );
  INVX1 U76 ( .A(B[6]), .Y(n34) );
  INVXL U77 ( .A(B[1]), .Y(n39) );
  INVXL U78 ( .A(B[2]), .Y(n38) );
  INVXL U79 ( .A(B[0]), .Y(n40) );
  INVXL U80 ( .A(B[4]), .Y(n36) );
  INVXL U81 ( .A(B[3]), .Y(n37) );
  INVXL U82 ( .A(B[5]), .Y(n35) );
endmodule


module mcu51_cpu_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  NOR21XL U2 ( .B(A[0]), .A(n1), .Y(carry[1]) );
  INVX1 U3 ( .A(B[0]), .Y(n1) );
endmodule


module mcu51_cpu_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  NOR21XL U1 ( .B(A[0]), .A(n1), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n1) );
  XOR2X1 U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  HAD1XL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mpb_a0 ( i_rd, i_wr, wdat0, wdat1, addr0, addr1, r_i2c_attr, esfrm_oe, 
        esfrm_we, sfrack, esfrm_wdat, esfrm_adr, mcu_esfr_rdat, delay_rdat, 
        delay_rrdy, esfrm_rrdy, esfrm_rdat, channel_sel, r_pg0_sel, dma_w, 
        dma_r, dma_addr, dma_wdat, dma_ack, memaddr, memaddr_c, memwr, memrd, 
        memrd_c, cpurst, memdatao, memack, hit_xd, hit_xr, hit_ps, hit_ps_c, 
        idat_r, idat_w, idat_adr, idat_wdat, iram_ce, xram_ce, regx_re, 
        iram_we, xram_we, regx_we, iram_a, xram_a, iram_d, xram_d, iram_rdat, 
        xram_rdat, regx_rdat, bist_en, bist_wr, bist_adr, bist_wdat, bist_xram, 
        mclk, srstz );
  input [1:0] i_rd;
  input [1:0] i_wr;
  input [7:0] wdat0;
  input [7:0] wdat1;
  input [7:0] addr0;
  input [7:0] addr1;
  output [7:0] esfrm_wdat;
  output [6:0] esfrm_adr;
  input [7:0] mcu_esfr_rdat;
  input [7:0] delay_rdat;
  output [7:0] esfrm_rdat;
  input [3:0] r_pg0_sel;
  input [10:0] dma_addr;
  input [7:0] dma_wdat;
  input [15:0] memaddr;
  input [15:0] memaddr_c;
  input [7:0] memdatao;
  input [7:0] idat_adr;
  input [7:0] idat_wdat;
  output [10:0] iram_a;
  output [10:0] xram_a;
  output [7:0] iram_d;
  output [7:0] xram_d;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  input [7:0] regx_rdat;
  input [10:0] bist_adr;
  input [7:0] bist_wdat;
  input r_i2c_attr, delay_rrdy, channel_sel, dma_w, dma_r, memwr, memrd,
         memrd_c, cpurst, idat_r, idat_w, bist_en, bist_wr, bist_xram, mclk,
         srstz;
  output esfrm_oe, esfrm_we, sfrack, esfrm_rrdy, dma_ack, memack, hit_xd,
         hit_xr, hit_ps, hit_ps_c, iram_ce, xram_ce, regx_re, iram_we, xram_we,
         regx_we;
  wire   dma_hit_x, pg0_rdwait, pg0_wrwait, N44, N45, r_pg0_rdrdy, N46,
         net128106, net153111, net153117, net153118, net153134, net153137,
         net153139, net153149, net153150, net153155, net153160, net153170,
         net153175, net153178, net153180, net153181, net153187, net153188,
         net153189, net153191, net153192, net153194, net153195, net153205,
         net153231, net153232, net153258, net153273, net153274, net153276,
         net153277, net153278, net153279, net153288, net153289, net153293,
         net153306, net153307, net153308, net166703, net166897, net166998,
         net169106, net169799, net169798, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238;
  wire   [1:0] xram_rdsel;

  DFFRQX1 r_pg0_rdrdy_reg ( .D(N46), .C(mclk), .XR(srstz), .Q(r_pg0_rdrdy) );
  DFFRQX1 xram_rdsel_reg_0_ ( .D(n203), .C(mclk), .XR(srstz), .Q(xram_rdsel[0]) );
  DFFRQX1 xram_rdsel_reg_1_ ( .D(net128106), .C(mclk), .XR(srstz), .Q(
        xram_rdsel[1]) );
  DFFRQX1 pg0_rdwait_reg ( .D(N45), .C(mclk), .XR(srstz), .Q(pg0_rdwait) );
  DFFRQX1 pg0_wrwait_reg ( .D(N44), .C(mclk), .XR(srstz), .Q(pg0_wrwait) );
  AO21X4 U3 ( .B(memaddr_c[0]), .C(net153188), .A(n130), .Y(xram_a[0]) );
  INVX1 U4 ( .A(n43), .Y(n12) );
  INVX1 U5 ( .A(i_wr[0]), .Y(n15) );
  INVX1 U6 ( .A(net153293), .Y(net153289) );
  NAND42X1 U7 ( .C(n2), .D(net153188), .A(n33), .B(n31), .Y(n18) );
  NAND21X1 U8 ( .B(n2), .A(n33), .Y(n28) );
  MUX2IX2 U9 ( .D0(n29), .D1(n30), .S(net153205), .Y(esfrm_adr[6]) );
  INVX1 U10 ( .A(addr1[6]), .Y(n29) );
  INVX1 U11 ( .A(addr0[6]), .Y(n30) );
  INVX1 U12 ( .A(addr0[3]), .Y(n46) );
  INVX1 U13 ( .A(addr1[3]), .Y(n45) );
  INVX1 U14 ( .A(net153180), .Y(net153187) );
  NAND31X1 U15 ( .C(net153139), .A(n9), .B(net153232), .Y(net153181) );
  INVX1 U16 ( .A(net153231), .Y(n9) );
  INVX3 U17 ( .A(net153181), .Y(net153188) );
  NAND21X2 U18 ( .B(net153117), .A(n11), .Y(net153277) );
  NAND21X1 U19 ( .B(n24), .A(n41), .Y(n11) );
  NAND21X1 U20 ( .B(n12), .A(n40), .Y(n41) );
  NAND21X1 U21 ( .B(n43), .A(n6), .Y(net153180) );
  NAND21X1 U22 ( .B(n21), .A(net153194), .Y(n27) );
  INVX1 U23 ( .A(dma_addr[6]), .Y(n21) );
  NOR21XL U24 ( .B(n27), .A(n32), .Y(n31) );
  INVX1 U25 ( .A(n26), .Y(n32) );
  NAND21X1 U26 ( .B(net153180), .A(esfrm_adr[6]), .Y(n33) );
  NAND21X1 U27 ( .B(n20), .A(net153195), .Y(n26) );
  INVX1 U28 ( .A(memaddr[6]), .Y(n20) );
  INVX1 U29 ( .A(n180), .Y(n195) );
  INVX1 U30 ( .A(memrd_c), .Y(n90) );
  NAND21X1 U31 ( .B(n23), .A(n39), .Y(n40) );
  NAND21X1 U32 ( .B(net153150), .A(n38), .Y(n39) );
  NAND21X1 U33 ( .B(xram_rdsel[1]), .A(xram_rdsel[0]), .Y(n38) );
  NAND21X1 U34 ( .B(net153306), .A(addr1[7]), .Y(n59) );
  NAND21X1 U35 ( .B(net153192), .A(net153195), .Y(n34) );
  INVX1 U36 ( .A(bist_adr[6]), .Y(n22) );
  INVX1 U37 ( .A(net153175), .Y(net153194) );
  NAND21X1 U38 ( .B(pg0_wrwait), .A(n76), .Y(n79) );
  NAND32X1 U39 ( .B(n81), .C(n110), .A(n177), .Y(net153117) );
  NAND31X1 U40 ( .C(xram_rdsel[0]), .A(net153289), .B(n12), .Y(net153288) );
  NOR21XL U41 ( .B(n7), .A(n8), .Y(net153189) );
  NAND21X1 U42 ( .B(n25), .A(n34), .Y(n8) );
  NAND21X1 U43 ( .B(net153191), .A(net153188), .Y(n7) );
  NOR21XL U44 ( .B(dma_addr[8]), .A(net153175), .Y(n25) );
  NAND21X1 U45 ( .B(n16), .A(n17), .Y(iram_a[6]) );
  NAND21X1 U46 ( .B(net153134), .A(esfrm_adr[6]), .Y(n17) );
  OAI22X1 U47 ( .A(net153137), .B(net153160), .C(n6), .D(n22), .Y(n16) );
  AOI221X1 U48 ( .A(net153187), .B(esfrm_adr[5]), .C(memaddr[5]), .D(net153195), .E(n144), .Y(n145) );
  INVX1 U49 ( .A(esfrm_adr[3]), .Y(n167) );
  OA222X1 U50 ( .A(n205), .B(net153178), .C(n157), .D(net153180), .E(n207), 
        .F(net153181), .Y(n158) );
  NAND21X1 U51 ( .B(net153139), .A(n42), .Y(net153175) );
  NAND31X1 U52 ( .C(net153118), .A(n43), .B(n35), .Y(n14) );
  INVX1 U53 ( .A(net169799), .Y(n35) );
  NAND21X1 U54 ( .B(xram_rdsel[0]), .A(xram_rdsel[1]), .Y(n13) );
  OAI211X1 U55 ( .C(n95), .D(n108), .A(n114), .B(n94), .Y(xram_d[1]) );
  NAND2X1 U56 ( .A(n13), .B(n14), .Y(dma_ack) );
  NAND21X2 U57 ( .B(net153306), .A(addr1[7]), .Y(n60) );
  INVX1 U58 ( .A(net169798), .Y(n10) );
  INVX3 U59 ( .A(n37), .Y(net153205) );
  AND2X1 U60 ( .A(n57), .B(n58), .Y(n1) );
  AND2X1 U61 ( .A(bist_adr[6]), .B(bist_en), .Y(n2) );
  OA33X1 U62 ( .A(n182), .B(net153134), .C(n181), .D(n180), .E(bist_en), .F(
        n179), .Y(n3) );
  INVX1 U63 ( .A(n42), .Y(net153232) );
  NAND31X1 U64 ( .C(n4), .A(net153274), .B(n42), .Y(net153273) );
  INVX1 U65 ( .A(bist_en), .Y(net166703) );
  INVXL U66 ( .A(net166703), .Y(n4) );
  INVXL U67 ( .A(n4), .Y(n5) );
  INVXL U68 ( .A(n4), .Y(n6) );
  OAI211X1 U69 ( .C(n101), .D(n108), .A(n120), .B(n100), .Y(xram_d[4]) );
  NAND21X1 U70 ( .B(net153117), .A(n86), .Y(n87) );
  INVX4 U71 ( .A(net153178), .Y(net153195) );
  NAND31X2 U72 ( .C(net153139), .A(net153231), .B(n10), .Y(net153178) );
  NAND21X1 U73 ( .B(net153307), .A(i_wr[1]), .Y(n61) );
  NAND21X2 U74 ( .B(i_wr[1]), .A(n15), .Y(net153111) );
  INVX3 U75 ( .A(i_rd[1]), .Y(net153306) );
  INVX1 U76 ( .A(i_rd[1]), .Y(n36) );
  INVX1 U77 ( .A(net153279), .Y(n24) );
  INVX1 U78 ( .A(net153278), .Y(n23) );
  NOR42X2 U79 ( .C(n26), .D(n27), .A(memaddr_c[6]), .B(n28), .Y(n19) );
  BUFXL U80 ( .A(net153149), .Y(n43) );
  INVX1 U81 ( .A(n10), .Y(n42) );
  NOR21X2 U82 ( .B(n18), .A(n19), .Y(xram_a[6]) );
  NAND31X2 U83 ( .C(i_wr[1]), .A(net153306), .B(addr0[7]), .Y(net153308) );
  NAND21X2 U84 ( .B(i_wr[1]), .A(n36), .Y(n37) );
  AND2X2 U85 ( .A(memaddr_c[4]), .B(net153188), .Y(n142) );
  MUX2IX2 U86 ( .D0(addr1[5]), .D1(addr0[5]), .S(net153205), .Y(n170) );
  AOI21X1 U87 ( .B(net153277), .C(net153118), .A(n203), .Y(net169798) );
  BUFXL U88 ( .A(net153117), .Y(net169799) );
  INVX2 U89 ( .A(idat_w), .Y(n183) );
  INVXL U90 ( .A(esfrm_we), .Y(n202) );
  NAND31X1 U91 ( .C(n48), .A(n200), .B(net153111), .Y(n76) );
  AO21XL U92 ( .B(n197), .C(n196), .A(pg0_rdwait), .Y(net153293) );
  MUX2IX2 U93 ( .D0(n46), .D1(n45), .S(n37), .Y(esfrm_adr[3]) );
  OR3X4 U94 ( .A(n142), .B(n143), .C(n47), .Y(xram_a[4]) );
  OAI21AXL U95 ( .B(net153178), .C(n141), .A(n140), .Y(n47) );
  BUFXL U96 ( .A(i_wr[1]), .Y(net169106) );
  AOI21XL U97 ( .B(xram_rdsel[0]), .C(xram_rdsel[1]), .A(n195), .Y(n62) );
  INVX2 U98 ( .A(n170), .Y(esfrm_adr[5]) );
  BUFXL U99 ( .A(n199), .Y(n48) );
  AND2XL U100 ( .A(n74), .B(n110), .Y(N45) );
  INVXL U101 ( .A(n110), .Y(n111) );
  OAI211X1 U102 ( .C(n129), .D(net153180), .A(n160), .B(n128), .Y(n130) );
  AOI21BBX1 U103 ( .B(n89), .C(n88), .A(n87), .Y(n203) );
  AND2X2 U104 ( .A(n199), .B(n196), .Y(esfrm_oe) );
  NAND3X2 U105 ( .A(n59), .B(net153308), .C(n61), .Y(n67) );
  INVX1 U106 ( .A(n129), .Y(esfrm_adr[0]) );
  MUX2IX1 U107 ( .D0(addr1[0]), .D1(addr0[0]), .S(net153205), .Y(n129) );
  MUX2XL U108 ( .D0(wdat0[3]), .D1(wdat1[3]), .S(net169106), .Y(esfrm_wdat[3])
         );
  MUX2XL U109 ( .D0(wdat0[7]), .D1(wdat1[7]), .S(net169106), .Y(esfrm_wdat[7])
         );
  MUX2XL U110 ( .D0(wdat0[1]), .D1(wdat1[1]), .S(net169106), .Y(esfrm_wdat[1])
         );
  MUX2XL U111 ( .D0(wdat0[5]), .D1(wdat1[5]), .S(net169106), .Y(esfrm_wdat[5])
         );
  MUX2XL U112 ( .D0(wdat0[2]), .D1(wdat1[2]), .S(net169106), .Y(esfrm_wdat[2])
         );
  MUX2XL U113 ( .D0(wdat0[6]), .D1(wdat1[6]), .S(net169106), .Y(esfrm_wdat[6])
         );
  MUX2XL U114 ( .D0(addr1[2]), .D1(addr0[2]), .S(net153205), .Y(esfrm_adr[2])
         );
  OAI21BBX1 U115 ( .A(memaddr_c[3]), .B(net153188), .C(n137), .Y(xram_a[3]) );
  AND2X2 U116 ( .A(n51), .B(n67), .Y(esfrm_we) );
  OA21X1 U117 ( .B(n201), .C(n200), .A(net153111), .Y(n51) );
  BUFXL U118 ( .A(esfrm_oe), .Y(n52) );
  INVXL U119 ( .A(n52), .Y(n53) );
  AOI221X1 U120 ( .A(net153187), .B(esfrm_adr[2]), .C(memaddr[2]), .D(
        net153195), .E(n133), .Y(n134) );
  OAI21BBX1 U121 ( .A(memaddr_c[1]), .B(net153188), .C(n132), .Y(xram_a[1]) );
  NAND3X2 U122 ( .A(n60), .B(net153308), .C(n61), .Y(n199) );
  AOI221X1 U123 ( .A(net153187), .B(esfrm_adr[1]), .C(memaddr[1]), .D(
        net153195), .E(n131), .Y(n132) );
  MUX2X1 U124 ( .D0(addr1[1]), .D1(addr0[1]), .S(net153205), .Y(esfrm_adr[1])
         );
  NAND21XL U125 ( .B(i_rd[0]), .A(n36), .Y(n196) );
  OAI21BBX1 U126 ( .A(memaddr_c[5]), .B(net153188), .C(n145), .Y(xram_a[5]) );
  INVX1 U127 ( .A(n72), .Y(n54) );
  AO21X1 U128 ( .B(net153289), .C(n182), .A(n83), .Y(net153149) );
  NAND21X2 U129 ( .B(net153289), .A(n83), .Y(n177) );
  NAND21X2 U130 ( .B(n182), .A(n83), .Y(n185) );
  NAND2X1 U131 ( .A(r_pg0_sel[2]), .B(n71), .Y(n66) );
  INVX1 U132 ( .A(n66), .Y(n55) );
  INVX1 U133 ( .A(n66), .Y(n56) );
  INVX1 U134 ( .A(net153134), .Y(net166998) );
  INVX1 U135 ( .A(net153137), .Y(net166897) );
  NAND21XL U136 ( .B(bist_en), .A(n110), .Y(net153137) );
  NAND2X1 U137 ( .A(addr1[4]), .B(n37), .Y(n57) );
  NAND2XL U138 ( .A(addr0[4]), .B(net153205), .Y(n58) );
  OAI221XL U139 ( .A(n1), .B(net153134), .C(n219), .D(net153137), .E(n168), 
        .Y(iram_a[4]) );
  INVX1 U140 ( .A(n1), .Y(esfrm_adr[4]) );
  OAI21BBX1 U141 ( .A(memaddr_c[2]), .B(net153188), .C(n134), .Y(xram_a[2]) );
  AND2XL U142 ( .A(n202), .B(n53), .Y(sfrack) );
  INVXL U143 ( .A(addr1[7]), .Y(net153307) );
  INVXL U144 ( .A(n67), .Y(n197) );
  OAI221XL U145 ( .A(n210), .B(net153180), .C(n211), .D(n6), .E(net153189), 
        .Y(xram_a[8]) );
  AND2X1 U146 ( .A(xram_rdsel[0]), .B(n82), .Y(n80) );
  NAND21XL U147 ( .B(bist_en), .A(net153276), .Y(n108) );
  NAND21X2 U148 ( .B(idat_r), .A(n183), .Y(n110) );
  NAND31X1 U149 ( .C(net166998), .A(n211), .B(net153137), .Y(iram_a[8]) );
  OAI21BBX1 U150 ( .A(dma_addr[1]), .B(net153194), .C(n162), .Y(n131) );
  AOI221X1 U151 ( .A(net153187), .B(esfrm_adr[3]), .C(memaddr[3]), .D(
        net153195), .E(n136), .Y(n137) );
  OAI21BBX1 U152 ( .A(dma_addr[2]), .B(net153194), .C(n164), .Y(n133) );
  OAI21BBX1 U153 ( .A(dma_addr[5]), .B(net153194), .C(n169), .Y(n144) );
  AOI21XL U154 ( .B(net153150), .C(n90), .A(xram_rdsel[1]), .Y(n65) );
  NAND31XL U155 ( .C(dma_w), .A(n65), .B(xram_rdsel[0]), .Y(net153279) );
  NAND6X1 U156 ( .A(memwr), .B(n185), .C(n177), .D(net153149), .E(net153150), 
        .F(net153118), .Y(n180) );
  NOR2XL U157 ( .A(n62), .B(n68), .Y(memack) );
  NAND21X1 U158 ( .B(n85), .A(n84), .Y(n86) );
  NAND21X1 U159 ( .B(xram_rdsel[1]), .A(net153288), .Y(n84) );
  NAND21XL U160 ( .B(n5), .A(bist_adr[1]), .Y(n162) );
  OAI211XL U161 ( .C(n172), .D(net153180), .A(n171), .B(n151), .Y(xram_a[7])
         );
  NAND21XL U162 ( .B(n5), .A(bist_adr[0]), .Y(n160) );
  INVX1 U163 ( .A(n69), .Y(n68) );
  INVX1 U164 ( .A(net153137), .Y(net153170) );
  INVX1 U165 ( .A(net153134), .Y(net153155) );
  INVX1 U166 ( .A(n185), .Y(n81) );
  INVX1 U167 ( .A(n91), .Y(n106) );
  NAND32XL U168 ( .B(bist_en), .C(net153276), .A(net153232), .Y(n91) );
  INVX1 U169 ( .A(net153274), .Y(net153276) );
  NAND21XL U170 ( .B(bist_en), .A(n43), .Y(net153139) );
  INVX1 U171 ( .A(cpurst), .Y(n69) );
  NAND21X1 U172 ( .B(net166703), .A(bist_wdat[0]), .Y(n112) );
  NAND21X1 U173 ( .B(n6), .A(bist_wdat[4]), .Y(n120) );
  NAND21X1 U174 ( .B(bist_en), .A(n111), .Y(net153134) );
  AO21X1 U175 ( .B(n111), .C(n74), .A(n189), .Y(N46) );
  NAND21X1 U176 ( .B(n6), .A(bist_wdat[1]), .Y(n114) );
  NAND21X1 U177 ( .B(n5), .A(bist_wdat[5]), .Y(n122) );
  NAND21X1 U178 ( .B(n6), .A(bist_wdat[2]), .Y(n116) );
  NAND21X1 U179 ( .B(net166703), .A(bist_wdat[3]), .Y(n118) );
  NAND21X1 U180 ( .B(n5), .A(bist_wr), .Y(n184) );
  INVX1 U181 ( .A(n208), .Y(n148) );
  INVX1 U182 ( .A(net153273), .Y(net153258) );
  NOR21XL U183 ( .B(net153187), .A(n1), .Y(n143) );
  NAND21XL U184 ( .B(n83), .A(n79), .Y(net153274) );
  AO21X1 U185 ( .B(n195), .C(hit_xr), .A(n187), .Y(regx_we) );
  INVX1 U186 ( .A(n72), .Y(n83) );
  NAND21X1 U187 ( .B(n55), .A(n181), .Y(n72) );
  INVX1 U188 ( .A(n157), .Y(n71) );
  INVX1 U189 ( .A(n178), .Y(n187) );
  NAND21XL U190 ( .B(n182), .A(n56), .Y(n178) );
  INVX1 U191 ( .A(n93), .Y(esfrm_wdat[0]) );
  INVX1 U192 ( .A(n101), .Y(esfrm_wdat[4]) );
  INVX1 U193 ( .A(idat_adr[6]), .Y(net153160) );
  OAI211X1 U194 ( .C(net128106), .D(n3), .A(n193), .B(n192), .Y(xram_ce) );
  MUX3IX1 U195 ( .D0(n191), .D1(n190), .D2(bist_xram), .S0(n203), .S1(bist_en), 
        .Y(n192) );
  AND2X1 U196 ( .A(net128106), .B(dma_hit_x), .Y(n191) );
  OAI31XL U197 ( .A(memaddr_c[15]), .B(memaddr_c[14]), .C(n206), .D(net128106), 
        .Y(n190) );
  OAI221X1 U198 ( .A(n167), .B(net153134), .C(n220), .D(net153137), .E(n166), 
        .Y(iram_a[3]) );
  OAI221X1 U199 ( .A(n170), .B(net153134), .C(n218), .D(net153137), .E(n169), 
        .Y(iram_a[5]) );
  OAI211X1 U200 ( .C(n176), .D(net153137), .A(net153134), .B(n175), .Y(
        iram_a[10]) );
  OAI211X1 U201 ( .C(net153175), .D(n159), .A(n175), .B(n158), .Y(xram_a[10])
         );
  NOR32XL U202 ( .B(n174), .C(n173), .A(n221), .Y(n176) );
  NAND21X1 U203 ( .B(n125), .A(n124), .Y(iram_d[6]) );
  AO22X1 U204 ( .A(idat_wdat[6]), .B(net153170), .C(esfrm_wdat[6]), .D(
        net153155), .Y(n125) );
  NAND21X1 U205 ( .B(n127), .A(n126), .Y(iram_d[7]) );
  AO22X1 U206 ( .A(idat_wdat[7]), .B(net153170), .C(esfrm_wdat[7]), .D(
        net153155), .Y(n127) );
  NAND21X1 U207 ( .B(n121), .A(n120), .Y(iram_d[4]) );
  AO22X1 U208 ( .A(idat_wdat[4]), .B(net153170), .C(net153155), .D(
        esfrm_wdat[4]), .Y(n121) );
  NAND21X1 U209 ( .B(n123), .A(n122), .Y(iram_d[5]) );
  AO22X1 U210 ( .A(idat_wdat[5]), .B(net153170), .C(esfrm_wdat[5]), .D(
        net153155), .Y(n123) );
  NAND21X1 U211 ( .B(n119), .A(n118), .Y(iram_d[3]) );
  AO22X1 U212 ( .A(idat_wdat[3]), .B(net153170), .C(esfrm_wdat[3]), .D(
        net153155), .Y(n119) );
  NAND21X1 U213 ( .B(n117), .A(n116), .Y(iram_d[2]) );
  AO22X1 U214 ( .A(idat_wdat[2]), .B(net153170), .C(esfrm_wdat[2]), .D(
        net153155), .Y(n117) );
  NAND21X1 U215 ( .B(n113), .A(n112), .Y(iram_d[0]) );
  AO22X1 U216 ( .A(idat_wdat[0]), .B(net153170), .C(net153155), .D(
        esfrm_wdat[0]), .Y(n113) );
  NAND21X1 U217 ( .B(n189), .A(n188), .Y(regx_re) );
  NAND43X1 U218 ( .B(n216), .C(n187), .D(n207), .A(n186), .Y(n188) );
  AND4XL U219 ( .A(memaddr_c[9]), .B(memaddr_c[8]), .C(n203), .D(net128106), 
        .Y(n186) );
  NAND21X1 U220 ( .B(n115), .A(n114), .Y(iram_d[1]) );
  AO22X1 U221 ( .A(idat_wdat[1]), .B(net153170), .C(esfrm_wdat[1]), .D(
        net166998), .Y(n115) );
  INVX1 U222 ( .A(hit_xd), .Y(n179) );
  MUX2XL U223 ( .D0(net169799), .D1(n194), .S(bist_en), .Y(iram_ce) );
  NAND21XL U224 ( .B(n198), .A(n53), .Y(esfrm_rrdy) );
  OAI211X1 U225 ( .C(n184), .D(n194), .A(n3), .B(n193), .Y(xram_we) );
  INVX1 U226 ( .A(n198), .Y(n204) );
  OAI222XL U227 ( .A(net153134), .B(n185), .C(bist_xram), .D(n184), .E(
        net153137), .F(n183), .Y(iram_we) );
  NOR21XL U228 ( .B(n110), .A(n78), .Y(N44) );
  NOR21XL U229 ( .B(n185), .A(n77), .Y(n78) );
  NOR21XL U230 ( .B(n79), .A(n181), .Y(n77) );
  NAND21X1 U231 ( .B(net166703), .A(bist_wdat[6]), .Y(n124) );
  OAI21BBXL U232 ( .A(n75), .B(net153293), .C(n177), .Y(n74) );
  INVX1 U233 ( .A(n73), .Y(n189) );
  NAND21XL U234 ( .B(net153289), .A(n56), .Y(n73) );
  INVX1 U235 ( .A(iram_a[9]), .Y(n152) );
  INVX1 U236 ( .A(n181), .Y(n75) );
  NAND43X1 U237 ( .B(net169799), .C(net153139), .D(net153118), .A(dma_hit_x), 
        .Y(n193) );
  INVX1 U238 ( .A(n213), .Y(n173) );
  AOI22X1 U239 ( .A(memaddr[0]), .B(net153195), .C(dma_addr[0]), .D(net153194), 
        .Y(n128) );
  AO21X1 U240 ( .B(dma_addr[3]), .C(net153194), .A(n135), .Y(n136) );
  INVX1 U241 ( .A(n166), .Y(n135) );
  NAND21XL U242 ( .B(dma_w), .A(memrd_c), .Y(net153278) );
  NOR21XL U243 ( .B(net153293), .A(n80), .Y(n88) );
  NOR2XL U244 ( .A(net153278), .B(dma_r), .Y(n89) );
  OAI211X1 U245 ( .C(n93), .D(n108), .A(n112), .B(n92), .Y(xram_d[0]) );
  AOI22X1 U246 ( .A(memdatao[0]), .B(n106), .C(dma_wdat[0]), .D(net153258), 
        .Y(n92) );
  AOI22XL U247 ( .A(memdatao[4]), .B(n106), .C(dma_wdat[4]), .D(net153258), 
        .Y(n100) );
  NAND21X1 U248 ( .B(net153276), .A(xram_rdsel[1]), .Y(n82) );
  INVXL U249 ( .A(n82), .Y(n85) );
  INVX1 U250 ( .A(memaddr[12]), .Y(n224) );
  AO21XL U251 ( .B(r_pg0_sel[1]), .C(n71), .A(n55), .Y(n181) );
  OAI211XL U252 ( .C(r_pg0_sel[1]), .D(r_pg0_sel[0]), .A(r_pg0_sel[2]), .B(
        r_pg0_sel[3]), .Y(n201) );
  NAND2XL U253 ( .A(n201), .B(r_pg0_sel[3]), .Y(n157) );
  NAND6XL U254 ( .A(memaddr[14]), .B(memaddr[15]), .C(memaddr[13]), .D(
        memaddr[11]), .E(memaddr[12]), .F(n70), .Y(n215) );
  AND4X1 U255 ( .A(memaddr[9]), .B(memaddr[10]), .C(memaddr[7]), .D(memaddr[8]), .Y(n70) );
  INVX1 U256 ( .A(memaddr[10]), .Y(n205) );
  INVX1 U257 ( .A(r_i2c_attr), .Y(n200) );
  MUX2IXL U258 ( .D0(wdat0[0]), .D1(wdat1[0]), .S(net169106), .Y(n93) );
  MUX2IXL U259 ( .D0(wdat0[4]), .D1(wdat1[4]), .S(net169106), .Y(n101) );
  NAND21X1 U260 ( .B(net166703), .A(bist_adr[2]), .Y(n164) );
  NAND21X1 U261 ( .B(n6), .A(bist_adr[5]), .Y(n169) );
  NAND21X1 U262 ( .B(n5), .A(bist_adr[3]), .Y(n166) );
  NAND21X1 U263 ( .B(n161), .A(n160), .Y(iram_a[0]) );
  AO22XL U264 ( .A(idat_adr[0]), .B(net153170), .C(net153155), .D(esfrm_adr[0]), .Y(n161) );
  NAND21X1 U265 ( .B(n163), .A(n162), .Y(iram_a[1]) );
  AO22XL U266 ( .A(idat_adr[1]), .B(net153170), .C(net153155), .D(esfrm_adr[1]), .Y(n163) );
  INVX1 U267 ( .A(esfrm_wdat[1]), .Y(n95) );
  AOI22XL U268 ( .A(memdatao[1]), .B(n106), .C(dma_wdat[1]), .D(net153258), 
        .Y(n94) );
  NAND21X1 U269 ( .B(n5), .A(bist_adr[4]), .Y(n168) );
  NAND21X1 U270 ( .B(n139), .A(n138), .Y(n140) );
  NAND21X1 U271 ( .B(net153175), .A(dma_addr[4]), .Y(n138) );
  INVX1 U272 ( .A(n168), .Y(n139) );
  OAI211X1 U273 ( .C(n109), .D(n108), .A(n126), .B(n107), .Y(xram_d[7]) );
  INVX1 U274 ( .A(esfrm_wdat[7]), .Y(n109) );
  AOI22XL U275 ( .A(memdatao[7]), .B(n106), .C(dma_wdat[7]), .D(net153258), 
        .Y(n107) );
  OAI211X1 U276 ( .C(n103), .D(n108), .A(n122), .B(n102), .Y(xram_d[5]) );
  INVX1 U277 ( .A(esfrm_wdat[5]), .Y(n103) );
  AOI22XL U278 ( .A(memdatao[5]), .B(n106), .C(dma_wdat[5]), .D(net153258), 
        .Y(n102) );
  OAI211X1 U279 ( .C(n97), .D(n108), .A(n116), .B(n96), .Y(xram_d[2]) );
  INVX1 U280 ( .A(esfrm_wdat[2]), .Y(n97) );
  AOI22XL U281 ( .A(memdatao[2]), .B(n106), .C(dma_wdat[2]), .D(net153258), 
        .Y(n96) );
  OAI211X1 U282 ( .C(n99), .D(n108), .A(n118), .B(n98), .Y(xram_d[3]) );
  INVX1 U283 ( .A(esfrm_wdat[3]), .Y(n99) );
  AOI22XL U284 ( .A(memdatao[3]), .B(n106), .C(dma_wdat[3]), .D(net153258), 
        .Y(n98) );
  OAI211X1 U285 ( .C(n105), .D(n108), .A(n124), .B(n104), .Y(xram_d[6]) );
  INVX1 U286 ( .A(esfrm_wdat[6]), .Y(n105) );
  AOI22XL U287 ( .A(memdatao[6]), .B(n106), .C(dma_wdat[6]), .D(net153258), 
        .Y(n104) );
  OAI221X1 U288 ( .A(net153134), .B(n172), .C(net153137), .D(n174), .E(n171), 
        .Y(iram_a[7]) );
  INVXL U289 ( .A(r_pg0_sel[0]), .Y(n172) );
  NAND21X1 U290 ( .B(n165), .A(n164), .Y(iram_a[2]) );
  AO22XL U291 ( .A(idat_adr[2]), .B(net166897), .C(net153155), .D(esfrm_adr[2]), .Y(n165) );
  OAI211XL U292 ( .C(n156), .D(net153178), .A(n155), .B(n154), .Y(xram_a[9])
         );
  INVX1 U293 ( .A(memaddr[9]), .Y(n156) );
  OA21X1 U294 ( .B(net153175), .C(n153), .A(n152), .Y(n154) );
  OR2X1 U295 ( .A(memrd), .B(memwr), .Y(net153231) );
  INVX1 U296 ( .A(memaddr[4]), .Y(n141) );
  AOI222XL U297 ( .A(dma_addr[7]), .B(net153194), .C(net153195), .D(n150), .E(
        net153188), .F(n149), .Y(n151) );
  OAI31XL U298 ( .A(n213), .B(memaddr[10]), .C(n147), .D(n146), .Y(n150) );
  OAI31XL U299 ( .A(n213), .B(n148), .C(memaddr_c[10]), .D(n212), .Y(n149) );
  INVX1 U300 ( .A(n214), .Y(n147) );
  INVX1 U301 ( .A(memaddr[8]), .Y(net153192) );
  INVX1 U302 ( .A(memaddr_c[8]), .Y(net153191) );
  AOI32XL U303 ( .A(net153187), .B(r_pg0_sel[2]), .C(n201), .D(net153188), .E(
        memaddr_c[9]), .Y(n155) );
  OR2X1 U304 ( .A(delay_rrdy), .B(r_pg0_rdrdy), .Y(n198) );
  AO222XL U305 ( .A(xram_rdat[7]), .B(n75), .C(iram_rdat[7]), .D(n83), .E(
        regx_rdat[7]), .F(n56), .Y(n231) );
  AO222XL U306 ( .A(xram_rdat[1]), .B(n75), .C(iram_rdat[1]), .D(n83), .E(
        regx_rdat[1]), .F(n56), .Y(n237) );
  AO222XL U307 ( .A(xram_rdat[2]), .B(n75), .C(iram_rdat[2]), .D(n83), .E(
        regx_rdat[2]), .F(n56), .Y(n236) );
  AO222XL U308 ( .A(xram_rdat[0]), .B(n75), .C(iram_rdat[0]), .D(n54), .E(
        regx_rdat[0]), .F(n56), .Y(n238) );
  INVX1 U309 ( .A(idat_adr[7]), .Y(n174) );
  AO222XL U310 ( .A(xram_rdat[4]), .B(n75), .C(iram_rdat[4]), .D(n83), .E(
        regx_rdat[4]), .F(n56), .Y(n234) );
  AO222XL U311 ( .A(xram_rdat[5]), .B(n75), .C(iram_rdat[5]), .D(n83), .E(
        regx_rdat[5]), .F(n56), .Y(n233) );
  AO222XL U312 ( .A(xram_rdat[3]), .B(n75), .C(iram_rdat[3]), .D(n54), .E(
        regx_rdat[3]), .F(n56), .Y(n235) );
  AO222XL U313 ( .A(xram_rdat[6]), .B(n75), .C(iram_rdat[6]), .D(n83), .E(
        regx_rdat[6]), .F(n56), .Y(n232) );
  NAND21X1 U314 ( .B(n5), .A(bist_wdat[7]), .Y(n126) );
  NAND21X1 U315 ( .B(net166703), .A(bist_adr[7]), .Y(n171) );
  NAND21X1 U316 ( .B(net166703), .A(bist_adr[10]), .Y(n175) );
  INVX1 U317 ( .A(memaddr[7]), .Y(n146) );
  INVX1 U318 ( .A(dma_w), .Y(net153118) );
  INVX1 U319 ( .A(dma_r), .Y(net153150) );
  INVX1 U320 ( .A(bist_xram), .Y(n194) );
  INVX1 U321 ( .A(dma_addr[10]), .Y(n159) );
  INVX1 U322 ( .A(dma_addr[9]), .Y(n153) );
  INVXL U323 ( .A(net153277), .Y(net128106) );
  AO222XL U324 ( .A(delay_rdat[2]), .B(n230), .C(r_pg0_rdrdy), .D(n236), .E(
        mcu_esfr_rdat[2]), .F(n204), .Y(esfrm_rdat[2]) );
  INVX3 U325 ( .A(n79), .Y(n182) );
  AO222XL U326 ( .A(delay_rdat[1]), .B(n230), .C(r_pg0_rdrdy), .D(n237), .E(
        mcu_esfr_rdat[1]), .F(n204), .Y(esfrm_rdat[1]) );
  AO222XL U327 ( .A(delay_rdat[0]), .B(n230), .C(r_pg0_rdrdy), .D(n238), .E(
        mcu_esfr_rdat[0]), .F(n204), .Y(esfrm_rdat[0]) );
  OAI21X1 U328 ( .B(dma_addr[9]), .C(dma_addr[8]), .A(dma_addr[10]), .Y(
        dma_hit_x) );
  OAI21X1 U329 ( .B(n207), .C(n208), .A(n209), .Y(n206) );
  INVX1 U330 ( .A(r_pg0_sel[1]), .Y(n210) );
  NAND4X1 U331 ( .A(memaddr_c[14]), .B(memaddr_c[13]), .C(memaddr_c[15]), .D(
        n217), .Y(n216) );
  NOR32XL U332 ( .B(memaddr_c[12]), .C(memaddr_c[11]), .A(n212), .Y(n217) );
  NOR21XL U333 ( .B(bist_adr[9]), .A(n5), .Y(iram_a[9]) );
  INVX1 U334 ( .A(bist_adr[8]), .Y(n211) );
  INVX1 U335 ( .A(channel_sel), .Y(n213) );
  MUX2IX1 U336 ( .D0(n222), .D1(n223), .S(idat_adr[6]), .Y(n221) );
  NAND2X1 U337 ( .A(idat_adr[4]), .B(idat_adr[5]), .Y(n223) );
  AOI21X1 U338 ( .B(n220), .C(n219), .A(n218), .Y(n222) );
  INVX1 U339 ( .A(idat_adr[5]), .Y(n218) );
  INVX1 U340 ( .A(idat_adr[4]), .Y(n219) );
  INVX1 U341 ( .A(idat_adr[3]), .Y(n220) );
  INVX1 U342 ( .A(n215), .Y(hit_xr) );
  NOR4XL U343 ( .A(memaddr[14]), .B(memaddr[15]), .C(memaddr[13]), .D(n225), 
        .Y(hit_xd) );
  OAI211X1 U344 ( .C(n205), .D(n214), .A(n224), .B(n226), .Y(n225) );
  AOI211X1 U345 ( .C(memaddr_c[14]), .D(n227), .A(memaddr_c[15]), .B(n68), .Y(
        hit_ps_c) );
  NAND4X1 U346 ( .A(n208), .B(n209), .C(n207), .D(n212), .Y(n227) );
  INVX1 U347 ( .A(memaddr_c[7]), .Y(n212) );
  INVX1 U348 ( .A(memaddr_c[10]), .Y(n207) );
  NOR3XL U349 ( .A(memaddr_c[12]), .B(memaddr_c[13]), .C(memaddr_c[11]), .Y(
        n209) );
  NOR2X1 U350 ( .A(memaddr_c[8]), .B(memaddr_c[9]), .Y(n208) );
  AOI211X1 U351 ( .C(memaddr[14]), .D(n228), .A(memaddr[15]), .B(n68), .Y(
        hit_ps) );
  NAND4X1 U352 ( .A(n205), .B(n226), .C(n214), .D(n229), .Y(n228) );
  NOR3XL U353 ( .A(memaddr[12]), .B(memaddr[7]), .C(memaddr[13]), .Y(n229) );
  NOR2X1 U354 ( .A(memaddr[8]), .B(memaddr[9]), .Y(n214) );
  INVX1 U355 ( .A(memaddr[11]), .Y(n226) );
  AO222X1 U356 ( .A(delay_rdat[7]), .B(n230), .C(r_pg0_rdrdy), .D(n231), .E(
        mcu_esfr_rdat[7]), .F(n204), .Y(esfrm_rdat[7]) );
  AO222X1 U357 ( .A(delay_rdat[6]), .B(n230), .C(r_pg0_rdrdy), .D(n232), .E(
        mcu_esfr_rdat[6]), .F(n204), .Y(esfrm_rdat[6]) );
  AO222X1 U358 ( .A(delay_rdat[5]), .B(n230), .C(r_pg0_rdrdy), .D(n233), .E(
        mcu_esfr_rdat[5]), .F(n204), .Y(esfrm_rdat[5]) );
  AO222X1 U359 ( .A(delay_rdat[4]), .B(n230), .C(r_pg0_rdrdy), .D(n234), .E(
        mcu_esfr_rdat[4]), .F(n204), .Y(esfrm_rdat[4]) );
  AO222X1 U360 ( .A(delay_rdat[3]), .B(n230), .C(r_pg0_rdrdy), .D(n235), .E(
        mcu_esfr_rdat[3]), .F(n204), .Y(esfrm_rdat[3]) );
  NOR21XL U361 ( .B(delay_rrdy), .A(r_pg0_rdrdy), .Y(n230) );
endmodule

