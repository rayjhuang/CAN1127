//
// Copyright 2021 MACRONIX INTERNATIONAL Co., Ltd.  All Rights Reserved.
//
// CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF MACRONIX INTERNATIONAL Co., Ltd
//      Process:                MXIC 0.18um CMOS 1P6M LOGIC (1.8V/5V)
//      Design Rule Doc.:       3105-L18B     V17
//      Spice model Doc.:       3126-L18B     V13
//      XRC cmd file    :       3213-L18B     V18
//      Date            :       2021/04/15
//      Author          :       izzieduan
//      VERSION         :       V2.0
//



// type: AND2 
`timescale 1ns/10ps
`celldefine
module AND2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0746912:0.195864:1.3566;
		specparam tpd_A_Y_f = 0.087472:0.238957:1.65799;
		specparam tpd_B_Y_r = 0.0818553:0.196286:1.33563;
		specparam tpd_B_Y_f = 0.098421:0.256274:1.70569;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND2 
`timescale 1ns/10ps
`celldefine
module AND2X12 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.236753:0.358363:1.4943;
		specparam tpd_A_Y_f = 0.223373:0.346777:1.16478;
		specparam tpd_B_Y_r = 0.24415:0.358203:1.46702;
		specparam tpd_B_Y_f = 0.235625:0.363947:1.21873;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND2 
`timescale 1ns/10ps
`celldefine
module AND2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0858498:0.217238:1.3806;
		specparam tpd_A_Y_f = 0.0954939:0.235953:1.30943;
		specparam tpd_B_Y_r = 0.092697:0.213967:1.34676;
		specparam tpd_B_Y_f = 0.106133:0.251154:1.35731;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND2 
`timescale 1ns/10ps
`celldefine
module AND2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.108843:0.253745:1.45939;
		specparam tpd_A_Y_f = 0.126471:0.281405:1.44256;
		specparam tpd_B_Y_r = 0.115667:0.24723:1.40735;
		specparam tpd_B_Y_f = 0.14033:0.299447:1.50547;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND2 
`timescale 1ns/10ps
`celldefine
module AND2X6 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.140729:0.299052:1.57254;
		specparam tpd_A_Y_f = 0.164244:0.329305:1.56942;
		specparam tpd_B_Y_r = 0.148145:0.293688:1.53041;
		specparam tpd_B_Y_f = 0.174917:0.343519:1.60503;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND2 
`timescale 1ns/10ps
`celldefine
module AND2X8 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.167051:0.329728:1.61333;
		specparam tpd_A_Y_f = 0.197017:0.367197:1.61534;
		specparam tpd_B_Y_r = 0.174459:0.324761:1.56439;
		specparam tpd_B_Y_f = 0.207628:0.379746:1.64863;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND2 
`timescale 1ns/10ps
`celldefine
module AND2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.108266:0.235876:1.39847;
		specparam tpd_A_Y_f = 0.113174:0.257795:1.45875;
		specparam tpd_B_Y_r = 0.116167:0.232615:1.36406;
		specparam tpd_B_Y_f = 0.127155:0.276874:1.51734;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND3 
`timescale 1ns/10ps
`celldefine
module AND3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.100812:0.23625:1.45403;
		specparam tpd_A_Y_f = 0.0975328:0.255213:1.66191;
		specparam tpd_B_Y_r = 0.114744:0.241418:1.43821;
		specparam tpd_B_Y_f = 0.110345:0.273121:1.7128;
		specparam tpd_C_Y_r = 0.122159:0.24118:1.39862;
		specparam tpd_C_Y_f = 0.119122:0.28631:1.75507;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND3 
`timescale 1ns/10ps
`celldefine
module AND3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.10847:0.250958:1.4591;
		specparam tpd_A_Y_f = 0.109137:0.273772:1.66567;
		specparam tpd_B_Y_r = 0.122094:0.253802:1.43556;
		specparam tpd_B_Y_f = 0.122114:0.290866:1.71737;
		specparam tpd_C_Y_r = 0.12911:0.25105:1.38363;
		specparam tpd_C_Y_f = 0.131768:0.303829:1.76035;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND3 
`timescale 1ns/10ps
`celldefine
module AND3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.14559:0.301277:1.57302;
		specparam tpd_A_Y_f = 0.137113:0.296445:1.47066;
		specparam tpd_B_Y_r = 0.159178:0.303157:1.54111;
		specparam tpd_B_Y_f = 0.149781:0.311718:1.51845;
		specparam tpd_C_Y_r = 0.166187:0.299152:1.48203;
		specparam tpd_C_Y_f = 0.159729:0.323701:1.55698;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND3 
`timescale 1ns/10ps
`celldefine
module AND3X8 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.210882:0.375539:1.66746;
		specparam tpd_A_Y_f = 0.197596:0.364723:1.55776;
		specparam tpd_B_Y_r = 0.224383:0.377848:1.62172;
		specparam tpd_B_Y_f = 0.215166:0.385453:1.61186;
		specparam tpd_C_Y_r = 0.231404:0.373067:1.54648;
		specparam tpd_C_Y_f = 0.224235:0.395509:1.64338;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND3 
`timescale 1ns/10ps
`celldefine
module AND3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.11594:0.249346:1.45429;
		specparam tpd_A_Y_f = 0.107693:0.25296:1.46803;
		specparam tpd_B_Y_r = 0.12994:0.254745:1.43921;
		specparam tpd_B_Y_f = 0.120986:0.271307:1.5218;
		specparam tpd_C_Y_r = 0.13694:0.253484:1.39739;
		specparam tpd_C_Y_f = 0.132432:0.286742:1.56791;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND4 
`timescale 1ns/10ps
`celldefine
module AND4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	and (Y, A, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.115641:0.256782:1.46611;
		specparam tpd_A_Y_f = 0.112433:0.27805:1.71907;
		specparam tpd_B_Y_r = 0.135309:0.267844:1.46164;
		specparam tpd_B_Y_f = 0.12827:0.298319:1.77473;
		specparam tpd_C_Y_r = 0.148692:0.273673:1.4315;
		specparam tpd_C_Y_f = 0.141121:0.314486:1.81975;
		specparam tpd_D_Y_r = 0.156531:0.278647:1.39802;
		specparam tpd_D_Y_f = 0.151021:0.327367:1.85764;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND4 
`timescale 1ns/10ps
`celldefine
module AND4X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	and (Y, A, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.126245:0.277891:1.5175;
		specparam tpd_A_Y_f = 0.125909:0.300877:1.76713;
		specparam tpd_B_Y_r = 0.145775:0.287332:1.50797;
		specparam tpd_B_Y_f = 0.14197:0.320736:1.82155;
		specparam tpd_C_Y_r = 0.158332:0.291219:1.47113;
		specparam tpd_C_Y_f = 0.154725:0.335356:1.86494;
		specparam tpd_D_Y_r = 0.166432:0.295187:1.42695;
		specparam tpd_D_Y_f = 0.16608:0.350277:1.90795;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND4 
`timescale 1ns/10ps
`celldefine
module AND4X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	and (Y, A, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.176208:0.336319:1.60395;
		specparam tpd_A_Y_f = 0.163971:0.328744:1.54731;
		specparam tpd_B_Y_r = 0.1956:0.345353:1.58374;
		specparam tpd_B_Y_f = 0.17974:0.348381:1.59461;
		specparam tpd_C_Y_r = 0.208104:0.348169:1.53684;
		specparam tpd_C_Y_f = 0.192728:0.362969:1.63371;
		specparam tpd_D_Y_r = 0.215798:0.350835:1.48347;
		specparam tpd_D_Y_f = 0.204495:0.376203:1.67178;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AND4 
`timescale 1ns/10ps
`celldefine
module AND4XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	and (Y, A, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.130519:0.265508:1.44948;
		specparam tpd_A_Y_f = 0.125093:0.274199:1.48031;
		specparam tpd_B_Y_r = 0.148942:0.276324:1.44087;
		specparam tpd_B_Y_f = 0.147078:0.301079:1.55278;
		specparam tpd_C_Y_r = 0.163729:0.283956:1.41412;
		specparam tpd_C_Y_f = 0.165278:0.322355:1.61028;
		specparam tpd_D_Y_r = 0.170451:0.286588:1.37967;
		specparam tpd_D_Y_f = 0.174446:0.332203:1.64418;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: ANT 
`timescale 1ns/10ps
`celldefine
module ANT (A);
	input A;
	// Timing
	specify

	endspecify
endmodule
`endcelldefine

// type: AO21 
`timescale 1ns/10ps
`celldefine
module AO21X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, B, C);
	or (Y, A, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0825084:0.22058:1.36411;
		specparam tpd_A_Y_f = 0.187488:0.379442:2.03748;
		specparam tpd_B_Y_r = 0.135366:0.286271:1.54006;
		specparam tpd_B_Y_f = 0.208316:0.38265:1.91653;
		specparam tpd_C_Y_r = 0.142804:0.279484:1.48461;
		specparam tpd_C_Y_f = 0.230349:0.409501:1.97507;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO21 
`timescale 1ns/10ps
`celldefine
module AO21X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, B, C);
	or (Y, A, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.100974:0.252785:1.43223;
		specparam tpd_A_Y_f = 0.25924:0.448626:1.9358;
		specparam tpd_B_Y_r = 0.167768:0.32876:1.61856;
		specparam tpd_B_Y_f = 0.281377:0.455353:1.79763;
		specparam tpd_C_Y_r = 0.174981:0.321843:1.5541;
		specparam tpd_C_Y_f = 0.298659:0.476051:1.83929;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO21 
`timescale 1ns/10ps
`celldefine
module AO21XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, B, C);
	or (Y, A, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.109075:0.236477:1.31917;
		specparam tpd_A_Y_f = 0.206834:0.384578:1.88287;
		specparam tpd_B_Y_r = 0.181025:0.323472:1.54881;
		specparam tpd_B_Y_f = 0.240061:0.402311:1.74141;
		specparam tpd_C_Y_r = 0.190116:0.313506:1.46304;
		specparam tpd_C_Y_f = 0.26455:0.432157:1.80926;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO2222 
`timescale 1ns/10ps
`celldefine
module AO2222X1 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	and (int_fwire_0, G, H);
	and (int_fwire_1, E, F);
	and (int_fwire_2, C, D);
	and (int_fwire_3, A, B);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.128796:0.269162:1.47932;
		specparam tpd_A_Y_f = 0.157839:0.31664:1.63735;
		specparam tpd_B_Y_r = 0.137705:0.267671:1.45457;
		specparam tpd_B_Y_f = 0.1741:0.334961:1.67764;
		specparam tpd_C_Y_r = 0.184413:0.328091:1.63439;
		specparam tpd_C_Y_f = 0.210413:0.357423:1.58829;
		specparam tpd_D_Y_r = 0.192487:0.325603:1.59063;
		specparam tpd_D_Y_f = 0.225993:0.37689:1.62899;
		specparam tpd_E_Y_r = 0.141425:0.278133:1.48775;
		specparam tpd_E_Y_f = 0.163195:0.316413:1.63025;
		specparam tpd_F_Y_r = 0.14999:0.276075:1.46036;
		specparam tpd_F_Y_f = 0.178705:0.33387:1.67155;
		specparam tpd_G_Y_r = 0.197484:0.338513:1.64331;
		specparam tpd_G_Y_f = 0.215216:0.356583:1.5749;
		specparam tpd_H_Y_r = 0.2056:0.335408:1.59979;
		specparam tpd_H_Y_f = 0.230495:0.375697:1.61626;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO2222 
`timescale 1ns/10ps
`celldefine
module AO2222X4 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	and (int_fwire_0, G, H);
	and (int_fwire_1, E, F);
	and (int_fwire_2, C, D);
	and (int_fwire_3, A, B);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.180885:0.337077:1.63306;
		specparam tpd_A_Y_f = 0.232609:0.40124:1.7641;
		specparam tpd_B_Y_r = 0.189566:0.334432:1.59596;
		specparam tpd_B_Y_f = 0.247927:0.418316:1.79975;
		specparam tpd_C_Y_r = 0.238989:0.394206:1.77107;
		specparam tpd_C_Y_f = 0.284447:0.442444:1.68855;
		specparam tpd_D_Y_r = 0.24711:0.391968:1.7167;
		specparam tpd_D_Y_f = 0.299821:0.461634:1.72599;
		specparam tpd_E_Y_r = 0.188934:0.338082:1.61358;
		specparam tpd_E_Y_f = 0.240823:0.405383:1.77889;
		specparam tpd_F_Y_r = 0.196987:0.332488:1.56365;
		specparam tpd_F_Y_f = 0.256461:0.42284:1.82261;
		specparam tpd_G_Y_r = 0.252611:0.401726:1.77058;
		specparam tpd_G_Y_f = 0.293415:0.446708:1.69121;
		specparam tpd_H_Y_r = 0.26054:0.399658:1.71738;
		specparam tpd_H_Y_f = 0.308477:0.465451:1.72788;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO2222 
`timescale 1ns/10ps
`celldefine
module AO2222XL (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	and (int_fwire_0, G, H);
	and (int_fwire_1, E, F);
	and (int_fwire_2, C, D);
	and (int_fwire_3, A, B);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.168323:0.301809:1.44041;
		specparam tpd_A_Y_f = 0.218331:0.386147:1.84741;
		specparam tpd_B_Y_r = 0.177383:0.295567:1.3908;
		specparam tpd_B_Y_f = 0.237482:0.407889:1.89732;
		specparam tpd_C_Y_r = 0.237205:0.373023:1.60973;
		specparam tpd_C_Y_f = 0.294177:0.454928:1.79524;
		specparam tpd_D_Y_r = 0.246419:0.367186:1.54362;
		specparam tpd_D_Y_f = 0.313087:0.477758:1.83605;
		specparam tpd_E_Y_r = 0.199269:0.333524:1.50761;
		specparam tpd_E_Y_f = 0.226531:0.387147:1.82773;
		specparam tpd_F_Y_r = 0.21679:0.338941:1.4913;
		specparam tpd_F_Y_f = 0.249914:0.41175:1.86834;
		specparam tpd_G_Y_r = 0.252265:0.389056:1.63533;
		specparam tpd_G_Y_f = 0.315956:0.471316:1.80889;
		specparam tpd_H_Y_r = 0.267463:0.385255:1.56893;
		specparam tpd_H_Y_f = 0.327358:0.485471:1.83244;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO222 
`timescale 1ns/10ps
`celldefine
module AO222X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	and (int_fwire_0, E, F);
	and (int_fwire_1, C, D);
	and (int_fwire_2, A, B);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.123713:0.278604:1.48252;
		specparam tpd_A_Y_f = 0.221827:0.423806:2.04748;
		specparam tpd_B_Y_r = 0.132633:0.276832:1.45816;
		specparam tpd_B_Y_f = 0.246779:0.450945:2.09768;
		specparam tpd_C_Y_r = 0.181523:0.338405:1.62647;
		specparam tpd_C_Y_f = 0.336175:0.525276:2.05609;
		specparam tpd_D_Y_r = 0.189541:0.335758:1.58712;
		specparam tpd_D_Y_f = 0.35884:0.551807:2.09504;
		specparam tpd_E_Y_r = 0.215908:0.375695:1.74684;
		specparam tpd_E_Y_f = 0.380837:0.56977:1.98675;
		specparam tpd_F_Y_r = 0.223142:0.370288:1.67072;
		specparam tpd_F_Y_f = 0.402317:0.595152:2.02697;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO222 
`timescale 1ns/10ps
`celldefine
module AO222X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	and (int_fwire_0, E, F);
	and (int_fwire_1, C, D);
	and (int_fwire_2, A, B);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.198289:0.371778:1.67805;
		specparam tpd_A_Y_f = 0.394748:0.594558:2.06473;
		specparam tpd_B_Y_r = 0.206715:0.369916:1.6394;
		specparam tpd_B_Y_f = 0.416561:0.619702:2.10249;
		specparam tpd_C_Y_r = 0.242113:0.412916:1.76604;
		specparam tpd_C_Y_f = 0.495601:0.686077:2.03396;
		specparam tpd_D_Y_r = 0.249823:0.409584:1.70135;
		specparam tpd_D_Y_f = 0.516491:0.711308:2.0722;
		specparam tpd_E_Y_r = 0.290425:0.463756:1.89234;
		specparam tpd_E_Y_f = 0.54446:0.737347:1.94953;
		specparam tpd_F_Y_r = 0.29808:0.458987:1.79894;
		specparam tpd_F_Y_f = 0.565423:0.762655:1.99023;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO222 
`timescale 1ns/10ps
`celldefine
module AO222XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	and (int_fwire_0, E, F);
	and (int_fwire_1, C, D);
	and (int_fwire_2, A, B);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.183657:0.334868:1.50877;
		specparam tpd_A_Y_f = 0.308626:0.504192:2.05599;
		specparam tpd_B_Y_r = 0.193501:0.330229:1.46992;
		specparam tpd_B_Y_f = 0.329346:0.528633:2.09307;
		specparam tpd_C_Y_r = 0.260503:0.411097:1.67021;
		specparam tpd_C_Y_f = 0.48171:0.667047:2.07213;
		specparam tpd_D_Y_r = 0.271602:0.409876:1.61889;
		specparam tpd_D_Y_f = 0.503173:0.693998:2.10165;
		specparam tpd_E_Y_r = 0.290147:0.443135:1.77505;
		specparam tpd_E_Y_f = 0.525486:0.710284:1.9889;
		specparam tpd_F_Y_r = 0.29937:0.435032:1.66532;
		specparam tpd_F_Y_f = 0.562108:0.754228:2.05926;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22A 
`timescale 1ns/10ps
`celldefine
module AO22AX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	and (int_fwire_0, C, D__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.105892:0.261167:1.49688;
		specparam tpd_A_Y_f = 0.17109:0.358588:1.99736;
		specparam tpd_B_Y_r = 0.113027:0.256211:1.45152;
		specparam tpd_B_Y_f = 0.18597:0.375918:2.04012;
		specparam tpd_C_Y_r = 0.166005:0.319383:1.64571;
		specparam tpd_C_Y_f = 0.199835:0.373105:1.8943;
		specparam tpd_D_Y_r = 0.235805:0.381512:1.6092;
		specparam tpd_D_Y_f = 0.286332:0.458109:1.86775;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22A 
`timescale 1ns/10ps
`celldefine
module AO22AX4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	and (int_fwire_0, C, D__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.173231:0.348684:1.68435;
		specparam tpd_A_Y_f = 0.267886:0.446772:1.77946;
		specparam tpd_B_Y_r = 0.180363:0.342917:1.62493;
		specparam tpd_B_Y_f = 0.280646:0.461922:1.81379;
		specparam tpd_C_Y_r = 0.240951:0.410904:1.82677;
		specparam tpd_C_Y_f = 0.297331:0.46513:1.65244;
		specparam tpd_D_Y_r = 0.310894:0.473724:1.72024;
		specparam tpd_D_Y_f = 0.380753:0.54581:1.56615;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22A 
`timescale 1ns/10ps
`celldefine
module AO22AXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	and (int_fwire_0, C, D__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.157141:0.312443:1.51678;
		specparam tpd_A_Y_f = 0.247427:0.429392:1.9498;
		specparam tpd_B_Y_r = 0.166469:0.305791:1.45643;
		specparam tpd_B_Y_f = 0.267941:0.453177:1.99988;
		specparam tpd_C_Y_r = 0.222422:0.370131:1.65891;
		specparam tpd_C_Y_f = 0.277043:0.447155:1.80126;
		specparam tpd_D_Y_r = 0.314232:0.476612:1.8278;
		specparam tpd_D_Y_f = 0.387846:0.54349:1.59773;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22B 
`timescale 1ns/10ps
`celldefine
module AO22BX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire B__bar, D__bar, int_fwire_0;
	wire int_fwire_1;

	not (D__bar, D);
	and (int_fwire_0, C, D__bar);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.108925:0.253438:1.45457;
		specparam tpd_A_Y_f = 0.15971:0.343603:1.9354;
		specparam tpd_B_Y_r = 0.163666:0.308883:1.55391;
		specparam tpd_B_Y_f = 0.220189:0.383834:1.7206;
		specparam tpd_C_Y_r = 0.157552:0.306652:1.59128;
		specparam tpd_C_Y_f = 0.207885:0.379529:1.88255;
		specparam tpd_D_Y_r = 0.213143:0.357781:1.60654;
		specparam tpd_D_Y_f = 0.270423:0.435044:1.7582;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22B 
`timescale 1ns/10ps
`celldefine
module AO22BX4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire B__bar, D__bar, int_fwire_0;
	wire int_fwire_1;

	not (D__bar, D);
	and (int_fwire_0, C, D__bar);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.173348:0.339077:1.63955;
		specparam tpd_A_Y_f = 0.253722:0.431197:1.74424;
		specparam tpd_B_Y_r = 0.228723:0.389756:1.64926;
		specparam tpd_B_Y_f = 0.31344:0.470896:1.45284;
		specparam tpd_C_Y_r = 0.223721:0.38819:1.75689;
		specparam tpd_C_Y_f = 0.301991:0.468547:1.65927;
		specparam tpd_D_Y_r = 0.279244:0.439301:1.6991;
		specparam tpd_D_Y_f = 0.363025:0.522156:1.48995;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22B 
`timescale 1ns/10ps
`celldefine
module AO22BXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire B__bar, D__bar, int_fwire_0;
	wire int_fwire_1;

	not (D__bar, D);
	and (int_fwire_0, C, D__bar);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.155919:0.298996:1.47872;
		specparam tpd_A_Y_f = 0.216061:0.396593:1.90027;
		specparam tpd_B_Y_r = 0.225505:0.386255:1.75165;
		specparam tpd_B_Y_f = 0.285233:0.435702:1.48966;
		specparam tpd_C_Y_r = 0.225841:0.371033:1.64927;
		specparam tpd_C_Y_f = 0.289971:0.462305:1.84068;
		specparam tpd_D_Y_r = 0.294802:0.456083:1.81662;
		specparam tpd_D_Y_f = 0.358504:0.511425:1.56493;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22 
`timescale 1ns/10ps
`celldefine
module AO22X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, C, D);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.113153:0.260871:1.48268;
		specparam tpd_A_Y_f = 0.159138:0.34473:1.93396;
		specparam tpd_B_Y_r = 0.12004:0.254026:1.43668;
		specparam tpd_B_Y_f = 0.170958:0.35811:1.96918;
		specparam tpd_C_Y_r = 0.167824:0.319324:1.63455;
		specparam tpd_C_Y_f = 0.209013:0.384018:1.88698;
		specparam tpd_D_Y_r = 0.175203:0.313119:1.56986;
		specparam tpd_D_Y_f = 0.223221:0.40099:1.92787;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22 
`timescale 1ns/10ps
`celldefine
module AO22X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, C, D);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.179618:0.346925:1.65516;
		specparam tpd_A_Y_f = 0.253556:0.430797:1.73478;
		specparam tpd_B_Y_r = 0.186599:0.339491:1.59117;
		specparam tpd_B_Y_f = 0.262435:0.441077:1.75805;
		specparam tpd_C_Y_r = 0.236995:0.403452:1.78334;
		specparam tpd_C_Y_f = 0.301626:0.469701:1.6493;
		specparam tpd_D_Y_r = 0.244325:0.397608:1.70395;
		specparam tpd_D_Y_f = 0.31446:0.485408:1.68489;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO22 
`timescale 1ns/10ps
`celldefine
module AO22XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, C, D);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.15934:0.304988:1.49598;
		specparam tpd_A_Y_f = 0.222602:0.404429:1.91434;
		specparam tpd_B_Y_r = 0.167795:0.294616:1.41908;
		specparam tpd_B_Y_f = 0.246286:0.432889:1.98459;
		specparam tpd_C_Y_r = 0.227419:0.374827:1.66132;
		specparam tpd_C_Y_f = 0.300378:0.475751:1.85862;
		specparam tpd_D_Y_r = 0.236337:0.365402:1.56553;
		specparam tpd_D_Y_f = 0.323617:0.504348:1.91843;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO33 
`timescale 1ns/10ps
`celldefine
module AO33X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, D, E, F);
	and (int_fwire_1, A, B, C);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.116306:0.241762:1.42184;
		specparam tpd_A_Y_f = 0.109912:0.251158:1.52116;
		specparam tpd_B_Y_r = 0.129135:0.246993:1.40897;
		specparam tpd_B_Y_f = 0.122588:0.269064:1.57178;
		specparam tpd_C_Y_r = 0.136243:0.246663:1.37326;
		specparam tpd_C_Y_f = 0.132356:0.282978:1.61379;
		specparam tpd_D_Y_r = 0.128279:0.252133:1.42998;
		specparam tpd_D_Y_f = 0.116096:0.255242:1.51638;
		specparam tpd_E_Y_r = 0.140889:0.256853:1.41426;
		specparam tpd_E_Y_f = 0.128453:0.27266:1.57059;
		specparam tpd_F_Y_r = 0.148602:0.257207:1.37873;
		specparam tpd_F_Y_f = 0.138771:0.287268:1.61428;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO33 
`timescale 1ns/10ps
`celldefine
module AO33X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, D, E, F);
	and (int_fwire_1, A, B, C);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.153587:0.299877:1.53656;
		specparam tpd_A_Y_f = 0.151018:0.310254:1.61204;
		specparam tpd_B_Y_r = 0.167105:0.302976:1.5119;
		specparam tpd_B_Y_f = 0.165253:0.327414:1.65955;
		specparam tpd_C_Y_r = 0.174886:0.301848:1.46803;
		specparam tpd_C_Y_f = 0.177226:0.340732:1.69584;
		specparam tpd_D_Y_r = 0.169563:0.311061:1.54682;
		specparam tpd_D_Y_f = 0.159389:0.316255:1.61358;
		specparam tpd_E_Y_r = 0.183089:0.313963:1.52242;
		specparam tpd_E_Y_f = 0.173374:0.332734:1.66267;
		specparam tpd_F_Y_r = 0.190711:0.312685:1.47721;
		specparam tpd_F_Y_f = 0.185142:0.345649:1.69926;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO33 
`timescale 1ns/10ps
`celldefine
module AO33XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, D, E, F);
	and (int_fwire_1, A, B, C);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.130585:0.258256:1.44589;
		specparam tpd_A_Y_f = 0.116954:0.252423:1.40239;
		specparam tpd_B_Y_r = 0.143866:0.26358:1.43249;
		specparam tpd_B_Y_f = 0.130599:0.271041:1.45502;
		specparam tpd_C_Y_r = 0.151174:0.263056:1.39767;
		specparam tpd_C_Y_f = 0.138552:0.281979:1.48779;
		specparam tpd_D_Y_r = 0.141737:0.266556:1.44954;
		specparam tpd_D_Y_f = 0.120327:0.252293:1.38825;
		specparam tpd_E_Y_r = 0.155969:0.272537:1.43469;
		specparam tpd_E_Y_f = 0.13355:0.270721:1.44598;
		specparam tpd_F_Y_r = 0.162675:0.270962:1.39184;
		specparam tpd_F_Y_f = 0.145367:0.286335:1.4948;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO44 
`timescale 1ns/10ps
`celldefine
module AO44X1 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, E, F, G, H);
	and (int_fwire_1, A, B, C, D);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.131775:0.263878:1.46151;
		specparam tpd_A_Y_f = 0.117846:0.263663:1.54401;
		specparam tpd_B_Y_r = 0.15357:0.277222:1.46202;
		specparam tpd_B_Y_f = 0.135018:0.285954:1.6047;
		specparam tpd_C_Y_r = 0.165799:0.282554:1.43378;
		specparam tpd_C_Y_f = 0.146435:0.300623:1.6472;
		specparam tpd_D_Y_r = 0.17265:0.28589:1.40034;
		specparam tpd_D_Y_f = 0.155282:0.312384:1.68225;
		specparam tpd_E_Y_r = 0.147996:0.277354:1.47589;
		specparam tpd_E_Y_f = 0.124785:0.268222:1.54106;
		specparam tpd_F_Y_r = 0.16586:0.286935:1.47058;
		specparam tpd_F_Y_f = 0.138942:0.286869:1.59575;
		specparam tpd_G_Y_r = 0.177741:0.290597:1.43842;
		specparam tpd_G_Y_f = 0.150345:0.301303:1.64175;
		specparam tpd_H_Y_r = 0.186244:0.296183:1.40377;
		specparam tpd_H_Y_f = 0.16068:0.314646:1.68434;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO44 
`timescale 1ns/10ps
`celldefine
module AO44X4 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, E, F, G, H);
	and (int_fwire_1, A, B, C, D);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.189668:0.342905:1.62767;
		specparam tpd_A_Y_f = 0.16364:0.326934:1.6462;
		specparam tpd_B_Y_r = 0.207971:0.351563:1.61183;
		specparam tpd_B_Y_f = 0.1781:0.343278:1.69087;
		specparam tpd_C_Y_r = 0.220312:0.353996:1.56741;
		specparam tpd_C_Y_f = 0.190314:0.357387:1.72995;
		specparam tpd_D_Y_r = 0.229184:0.360716:1.5324;
		specparam tpd_D_Y_f = 0.202306:0.370695:1.7621;
		specparam tpd_E_Y_r = 0.202766:0.349388:1.6222;
		specparam tpd_E_Y_f = 0.17197:0.33214:1.65125;
		specparam tpd_F_Y_r = 0.220343:0.356943:1.60469;
		specparam tpd_F_Y_f = 0.186151:0.348223:1.69762;
		specparam tpd_G_Y_r = 0.232706:0.359279:1.55904;
		specparam tpd_G_Y_f = 0.198931:0.362111:1.73941;
		specparam tpd_H_Y_r = 0.240981:0.364749:1.5273;
		specparam tpd_H_Y_f = 0.210127:0.374073:1.76739;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AO44 
`timescale 1ns/10ps
`celldefine
module AO44XL (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, E, F, G, H);
	and (int_fwire_1, A, B, C, D);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.159047:0.283203:1.42685;
		specparam tpd_A_Y_f = 0.13956:0.271079:1.34357;
		specparam tpd_B_Y_r = 0.17807:0.295327:1.42424;
		specparam tpd_B_Y_f = 0.159552:0.295164:1.40685;
		specparam tpd_C_Y_r = 0.191658:0.302004:1.40063;
		specparam tpd_C_Y_f = 0.175166:0.313178:1.45675;
		specparam tpd_D_Y_r = 0.198739:0.30595:1.37516;
		specparam tpd_D_Y_f = 0.180991:0.319822:1.47674;
		specparam tpd_E_Y_r = 0.177864:0.300878:1.44882;
		specparam tpd_E_Y_f = 0.143723:0.272212:1.32869;
		specparam tpd_F_Y_r = 0.197577:0.313027:1.44068;
		specparam tpd_F_Y_f = 0.166726:0.299764:1.40726;
		specparam tpd_G_Y_r = 0.211942:0.320538:1.41496;
		specparam tpd_G_Y_f = 0.184598:0.319692:1.46423;
		specparam tpd_H_Y_r = 0.219398:0.324349:1.38366;
		specparam tpd_H_Y_f = 0.195015:0.33179:1.49997;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI211 
`timescale 1ns/10ps
`celldefine
module AOI211X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, D__bar);
	not (C__bar, C);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0889251:0.219095:1.70049;
		specparam tpd_A_Y_f = 0.0364747:0.103021:0.770934;
		specparam tpd_B_Y_r = 0.143724:0.256634:1.61853;
		specparam tpd_B_Y_f = 0.0473057:0.121747:0.77715;
		specparam tpd_C_Y_r = 0.161084:0.276353:1.48517;
		specparam tpd_C_Y_f = 0.0860295:0.184386:1.09611;
		specparam tpd_D_Y_r = 0.178263:0.293062:1.49053;
		specparam tpd_D_Y_f = 0.0931192:0.17563:0.973825;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI211 
`timescale 1ns/10ps
`celldefine
module AOI211X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, D__bar);
	not (C__bar, C);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.277439:0.42477:1.91069;
		specparam tpd_A_Y_f = 0.173942:0.289821:0.893675;
		specparam tpd_B_Y_r = 0.332989:0.463809:1.88908;
		specparam tpd_B_Y_f = 0.185668:0.304762:0.934975;
		specparam tpd_C_Y_r = 0.348525:0.481081:1.75484;
		specparam tpd_C_Y_f = 0.25767:0.376391:1.13311;
		specparam tpd_D_Y_r = 0.367653:0.501066:1.79441;
		specparam tpd_D_Y_f = 0.264852:0.368683:1.06389;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI211 
`timescale 1ns/10ps
`celldefine
module AOI211XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, D__bar);
	not (C__bar, C);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0934256:0.224309:1.71908;
		specparam tpd_A_Y_f = 0.0561208:0.134764:0.976037;
		specparam tpd_B_Y_r = 0.149509:0.264414:1.63367;
		specparam tpd_B_Y_f = 0.0821938:0.166142:1.01486;
		specparam tpd_C_Y_r = 0.171935:0.290443:1.49992;
		specparam tpd_C_Y_f = 0.18355:0.29285:1.57879;
		specparam tpd_D_Y_r = 0.188819:0.307357:1.50745;
		specparam tpd_D_Y_f = 0.197911:0.289972:1.4145;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21A 
`timescale 1ns/10ps
`celldefine
module AOI21AX1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire B__bar, C__bar, int_fwire_0;
	wire int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, A, C__bar);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.115201:0.234451:1.38558;
		specparam tpd_A_Y_f = 0.0788401:0.163705:0.760029;
		specparam tpd_B_Y_r = 0.0938968:0.217002:1.62842;
		specparam tpd_B_Y_f = 0.0736083:0.185843:1.39592;
		specparam tpd_C_Y_r = 0.106776:0.230977:1.64449;
		specparam tpd_C_Y_f = 0.0811231:0.17796:1.26496;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21A 
`timescale 1ns/10ps
`celldefine
module AOI21AX4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire B__bar, C__bar, int_fwire_0;
	wire int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, A, C__bar);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.263216:0.389251:1.60622;
		specparam tpd_A_Y_f = 0.217691:0.330209:1.04041;
		specparam tpd_B_Y_r = 0.243662:0.37761:1.69686;
		specparam tpd_B_Y_f = 0.235646:0.351876:1.08791;
		specparam tpd_C_Y_r = 0.258548:0.394669:1.74776;
		specparam tpd_C_Y_f = 0.243258:0.344578:1.02374;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21A 
`timescale 1ns/10ps
`celldefine
module AOI21AXL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire B__bar, C__bar, int_fwire_0;
	wire int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, A, C__bar);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.156194:0.263665:1.3116;
		specparam tpd_A_Y_f = 0.104001:0.195822:0.84352;
		specparam tpd_B_Y_r = 0.143004:0.270861:1.70453;
		specparam tpd_B_Y_f = 0.0959801:0.188076:1.17294;
		specparam tpd_C_Y_r = 0.16337:0.293499:1.74547;
		specparam tpd_C_Y_f = 0.105134:0.177172:1.00821;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21BB 
`timescale 1ns/10ps
`celldefine
module AOI21BBX1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, int_fwire_0, int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, C);
	and (int_fwire_1, A__bar, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0706427:0.18956:1.61601;
		specparam tpd_A_Y_f = 0.0439126:0.140575:1.15452;
		specparam tpd_B_Y_r = 0.0983801:0.217231:1.30354;
		specparam tpd_B_Y_f = 0.126755:0.23929:1.06023;
		specparam tpd_C_Y_r = 0.110606:0.236846:1.36037;
		specparam tpd_C_Y_f = 0.150093:0.247607:1.02755;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21BB 
`timescale 1ns/10ps
`celldefine
module AOI21BBX4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, int_fwire_0, int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, C);
	and (int_fwire_1, A__bar, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0738122:0.191443:1.59896;
		specparam tpd_A_Y_f = 0.042036:0.140535:1.1532;
		specparam tpd_B_Y_r = 0.142717:0.281186:1.44551;
		specparam tpd_B_Y_f = 0.227349:0.354602:1.26843;
		specparam tpd_C_Y_r = 0.158158:0.298892:1.50309;
		specparam tpd_C_Y_f = 0.250621:0.362036:1.18472;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21BB 
`timescale 1ns/10ps
`celldefine
module AOI21BBXL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, int_fwire_0, int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, C);
	and (int_fwire_1, A__bar, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0775706:0.199452:1.64277;
		specparam tpd_A_Y_f = 0.0651734:0.167425:1.32234;
		specparam tpd_B_Y_r = 0.12605:0.239172:1.28318;
		specparam tpd_B_Y_f = 0.171018:0.30793:1.47591;
		specparam tpd_C_Y_r = 0.141427:0.258671:1.33811;
		specparam tpd_C_Y_f = 0.197549:0.319075:1.42824;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21B 
`timescale 1ns/10ps
`celldefine
module AOI21BX1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, C);
	not (B__bar, B);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.085859:0.224358:1.79242;
		specparam tpd_A_Y_f = 0.027119:0.0825378:0.696871;
		specparam tpd_B_Y_r = 0.103525:0.223267:1.60257;
		specparam tpd_B_Y_f = 0.0495574:0.133996:0.959736;
		specparam tpd_C_Y_r = 0.179042:0.296134:1.37417;
		specparam tpd_C_Y_f = 0.109115:0.196853:0.785727;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21B 
`timescale 1ns/10ps
`celldefine
module AOI21BX4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, C);
	not (B__bar, B);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.20128:0.350305:1.77083;
		specparam tpd_A_Y_f = 0.171789:0.283965:0.905704;
		specparam tpd_B_Y_r = 0.226226:0.360512:1.6527;
		specparam tpd_B_Y_f = 0.250669:0.365198:1.11725;
		specparam tpd_C_Y_r = 0.286948:0.417494:1.64686;
		specparam tpd_C_Y_f = 0.302269:0.409038:1.0775;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21B 
`timescale 1ns/10ps
`celldefine
module AOI21BXL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, C);
	not (B__bar, B);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.106076:0.244455:1.82617;
		specparam tpd_A_Y_f = 0.0448383:0.109208:0.789891;
		specparam tpd_B_Y_r = 0.141254:0.26585:1.64408;
		specparam tpd_B_Y_f = 0.0942015:0.184203:1.12693;
		specparam tpd_C_Y_r = 0.213448:0.320683:1.30608;
		specparam tpd_C_Y_f = 0.163163:0.268227:1.08335;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21 
`timescale 1ns/10ps
`celldefine
module AOI21X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1;

	not (C__bar, C);
	not (A__bar, A);
	and (int_fwire_0, A__bar, C__bar);
	not (B__bar, B);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0928044:0.224569:1.73295;
		specparam tpd_A_Y_f = 0.0365734:0.108375:0.862466;
		specparam tpd_B_Y_r = 0.11865:0.240201:1.61778;
		specparam tpd_B_Y_f = 0.0740015:0.169916:1.13845;
		specparam tpd_C_Y_r = 0.138154:0.263142:1.67333;
		specparam tpd_C_Y_f = 0.0812192:0.162794:1.01805;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21 
`timescale 1ns/10ps
`celldefine
module AOI21X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1;

	not (C__bar, C);
	not (A__bar, A);
	and (int_fwire_0, A__bar, C__bar);
	not (B__bar, B);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.238256:0.39028:1.87775;
		specparam tpd_A_Y_f = 0.16508:0.275525:0.852526;
		specparam tpd_B_Y_r = 0.259853:0.395646:1.74212;
		specparam tpd_B_Y_f = 0.224624:0.340539:1.03305;
		specparam tpd_C_Y_r = 0.278155:0.415801:1.79515;
		specparam tpd_C_Y_f = 0.231912:0.333528:0.975246;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI21 
`timescale 1ns/10ps
`celldefine
module AOI21XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1;

	not (C__bar, C);
	not (A__bar, A);
	and (int_fwire_0, A__bar, C__bar);
	not (B__bar, B);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0724576:0.209931:1.76297;
		specparam tpd_A_Y_f = 0.0397968:0.121368:1.0252;
		specparam tpd_B_Y_r = 0.103096:0.22507:1.56895;
		specparam tpd_B_Y_f = 0.0922732:0.201495:1.40349;
		specparam tpd_C_Y_r = 0.118902:0.243764:1.61818;
		specparam tpd_C_Y_f = 0.100677:0.193055:1.25576;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI221 
`timescale 1ns/10ps
`celldefine
module AOI221X1 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	not (E__bar, E);
	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar, E__bar);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar, E__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar, E__bar);
	and (int_fwire_3, A__bar, C__bar, E__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0882046:0.217653:1.67671;
		specparam tpd_A_Y_f = 0.0587355:0.14224:0.991477;
		specparam tpd_B_Y_r = 0.10756:0.236579:1.69802;
		specparam tpd_B_Y_f = 0.0669815:0.14029:0.911464;
		specparam tpd_C_Y_r = 0.19378:0.310145:1.62929;
		specparam tpd_C_Y_f = 0.111129:0.200451:1.05193;
		specparam tpd_D_Y_r = 0.214712:0.332254:1.65326;
		specparam tpd_D_Y_f = 0.11913:0.195521:0.950563;
		specparam tpd_E_Y_r = 0.251484:0.366048:1.54023;
		specparam tpd_E_Y_f = 0.0836923:0.176036:0.884312;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI221 
`timescale 1ns/10ps
`celldefine
module AOI221X4 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	not (E__bar, E);
	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar, E__bar);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar, E__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar, E__bar);
	and (int_fwire_3, A__bar, C__bar, E__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.26768:0.41902:1.91742;
		specparam tpd_A_Y_f = 0.228983:0.351314:1.11779;
		specparam tpd_B_Y_r = 0.289824:0.44107:1.96112;
		specparam tpd_B_Y_f = 0.237472:0.348587:1.08625;
		specparam tpd_C_Y_r = 0.377784:0.514872:1.90722;
		specparam tpd_C_Y_f = 0.28723:0.40999:1.26369;
		specparam tpd_D_Y_r = 0.399746:0.539006:1.95044;
		specparam tpd_D_Y_f = 0.295048:0.405866:1.20693;
		specparam tpd_E_Y_r = 0.436931:0.573093:1.87074;
		specparam tpd_E_Y_f = 0.243198:0.375111:1.25029;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI221 
`timescale 1ns/10ps
`celldefine
module AOI221XL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	not (E__bar, E);
	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar, E__bar);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar, E__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar, E__bar);
	and (int_fwire_3, A__bar, C__bar, E__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.150263:0.277273:1.73571;
		specparam tpd_A_Y_f = 0.0774174:0.146052:0.742234;
		specparam tpd_B_Y_r = 0.180519:0.307452:1.78684;
		specparam tpd_B_Y_f = 0.0859209:0.135567:0.612256;
		specparam tpd_C_Y_r = 0.308952:0.424809:1.71878;
		specparam tpd_C_Y_f = 0.139512:0.21124:0.836415;
		specparam tpd_D_Y_r = 0.34361:0.462387:1.77194;
		specparam tpd_D_Y_f = 0.14917:0.202605:0.701327;
		specparam tpd_E_Y_r = 0.393128:0.509765:1.67673;
		specparam tpd_E_Y_f = 0.11685:0.19108:0.736004;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI222 
`timescale 1ns/10ps
`celldefine
module AOI222X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7;

	not (F__bar, F);
	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar, F__bar);
	not (E__bar, E);
	and (int_fwire_1, B__bar, D__bar, E__bar);
	not (C__bar, C);
	and (int_fwire_2, B__bar, C__bar, F__bar);
	and (int_fwire_3, B__bar, C__bar, E__bar);
	not (A__bar, A);
	and (int_fwire_4, A__bar, D__bar, F__bar);
	and (int_fwire_5, A__bar, D__bar, E__bar);
	and (int_fwire_6, A__bar, C__bar, F__bar);
	and (int_fwire_7, A__bar, C__bar, E__bar);
	or (Y, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.375303:0.521755:2.14173;
		specparam tpd_A_Y_f = 0.172285:0.277395:0.869512;
		specparam tpd_B_Y_r = 0.414367:0.562256:2.19522;
		specparam tpd_B_Y_f = 0.180387:0.277534:0.865461;
		specparam tpd_C_Y_r = 0.476151:0.607401:2.10384;
		specparam tpd_C_Y_f = 0.192004:0.301428:0.941688;
		specparam tpd_D_Y_r = 0.514585:0.649464:2.16074;
		specparam tpd_D_Y_f = 0.199221:0.29697:0.911714;
		specparam tpd_E_Y_r = 0.525299:0.658496:2.01274;
		specparam tpd_E_Y_f = 0.212431:0.326322:1.04458;
		specparam tpd_F_Y_r = 0.563348:0.700824:2.07433;
		specparam tpd_F_Y_f = 0.219609:0.318776:0.983488;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI222 
`timescale 1ns/10ps
`celldefine
module AOI222X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7;

	not (F__bar, F);
	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar, F__bar);
	not (E__bar, E);
	and (int_fwire_1, B__bar, D__bar, E__bar);
	not (C__bar, C);
	and (int_fwire_2, B__bar, C__bar, F__bar);
	and (int_fwire_3, B__bar, C__bar, E__bar);
	not (A__bar, A);
	and (int_fwire_4, A__bar, D__bar, F__bar);
	and (int_fwire_5, A__bar, D__bar, E__bar);
	and (int_fwire_6, A__bar, C__bar, F__bar);
	and (int_fwire_7, A__bar, C__bar, E__bar);
	or (Y, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.337248:0.488151:2.05077;
		specparam tpd_A_Y_f = 0.246856:0.366393:1.0677;
		specparam tpd_B_Y_r = 0.36133:0.512689:2.09104;
		specparam tpd_B_Y_f = 0.255286:0.36384:1.03853;
		specparam tpd_C_Y_r = 0.438124:0.576308:2.02593;
		specparam tpd_C_Y_f = 0.29072:0.410232:1.17861;
		specparam tpd_D_Y_r = 0.461532:0.602115:2.06862;
		specparam tpd_D_Y_f = 0.298451:0.405826:1.12287;
		specparam tpd_E_Y_r = 0.487159:0.627709:1.94989;
		specparam tpd_E_Y_f = 0.335578:0.455279:1.31168;
		specparam tpd_F_Y_r = 0.510432:0.653246:1.99377;
		specparam tpd_F_Y_f = 0.343278:0.44977:1.22439;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI222 
`timescale 1ns/10ps
`celldefine
module AOI222XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7;

	not (F__bar, F);
	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar, F__bar);
	not (E__bar, E);
	and (int_fwire_1, B__bar, D__bar, E__bar);
	not (C__bar, C);
	and (int_fwire_2, B__bar, C__bar, F__bar);
	and (int_fwire_3, B__bar, C__bar, E__bar);
	not (A__bar, A);
	and (int_fwire_4, A__bar, D__bar, F__bar);
	and (int_fwire_5, A__bar, D__bar, E__bar);
	and (int_fwire_6, A__bar, C__bar, F__bar);
	and (int_fwire_7, A__bar, C__bar, E__bar);
	or (Y, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.164703:0.288464:1.71989;
		specparam tpd_A_Y_f = 0.0709735:0.148027:0.848277;
		specparam tpd_B_Y_r = 0.189899:0.314106:1.74294;
		specparam tpd_B_Y_f = 0.0796121:0.14585:0.776942;
		specparam tpd_C_Y_r = 0.274052:0.386686:1.67093;
		specparam tpd_C_Y_f = 0.115176:0.196012:0.897982;
		specparam tpd_D_Y_r = 0.299029:0.413393:1.69833;
		specparam tpd_D_Y_f = 0.123306:0.191021:0.803904;
		specparam tpd_E_Y_r = 0.326394:0.441839:1.58172;
		specparam tpd_E_Y_f = 0.149266:0.233132:1.00781;
		specparam tpd_F_Y_r = 0.351143:0.468405:1.61228;
		specparam tpd_F_Y_f = 0.157151:0.226907:0.882501;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22A 
`timescale 1ns/10ps
`celldefine
module AOI22AX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (B__bar, B);
	and (int_fwire_0, B__bar, D);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0808486:0.214745:1.71378;
		specparam tpd_A_Y_f = 0.0506754:0.151765:1.30283;
		specparam tpd_B_Y_r = 0.0940241:0.227654:1.73086;
		specparam tpd_B_Y_f = 0.057694:0.146088:1.18731;
		specparam tpd_C_Y_r = 0.111012:0.229476:1.51992;
		specparam tpd_C_Y_f = 0.108915:0.220098:1.45622;
		specparam tpd_D_Y_r = 0.192676:0.307862:1.35402;
		specparam tpd_D_Y_f = 0.180144:0.28521:1.16366;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22A 
`timescale 1ns/10ps
`celldefine
module AOI22AX4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (B__bar, B);
	and (int_fwire_0, B__bar, D);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.273532:0.425849:1.93009;
		specparam tpd_A_Y_f = 0.235658:0.352456:1.06877;
		specparam tpd_B_Y_r = 0.290539:0.443387:1.97715;
		specparam tpd_B_Y_f = 0.243228:0.346389:1.01098;
		specparam tpd_C_Y_r = 0.295496:0.436707:1.78381;
		specparam tpd_C_Y_f = 0.293463:0.411649:1.22705;
		specparam tpd_D_Y_r = 0.39125:0.522899:1.75052;
		specparam tpd_D_Y_f = 0.364412:0.475545:1.18202;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22A 
`timescale 1ns/10ps
`celldefine
module AOI22AXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (B__bar, B);
	and (int_fwire_0, B__bar, D);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.131229:0.266644:1.80468;
		specparam tpd_A_Y_f = 0.0618295:0.142935:1.03485;
		specparam tpd_B_Y_r = 0.151517:0.286902:1.82847;
		specparam tpd_B_Y_f = 0.0709742:0.136041:0.904265;
		specparam tpd_C_Y_r = 0.165337:0.290173:1.61452;
		specparam tpd_C_Y_f = 0.124375:0.213721:1.17002;
		specparam tpd_D_Y_r = 0.271698:0.377045:1.33012;
		specparam tpd_D_Y_f = 0.21606:0.31966:1.12623;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22B 
`timescale 1ns/10ps
`celldefine
module AOI22BX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, C__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	and (int_fwire_0, B, D);
	not (C__bar, C);
	and (int_fwire_1, B, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0739717:0.208587:1.73125;
		specparam tpd_A_Y_f = 0.0498246:0.145268:1.21889;
		specparam tpd_B_Y_r = 0.132561:0.242515:1.29272;
		specparam tpd_B_Y_f = 0.103265:0.199556:0.979752;
		specparam tpd_C_Y_r = 0.121928:0.242662:1.58463;
		specparam tpd_C_Y_f = 0.0950118:0.197451:1.28593;
		specparam tpd_D_Y_r = 0.183216:0.294656:1.33296;
		specparam tpd_D_Y_f = 0.150581:0.24787:1.03104;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22B 
`timescale 1ns/10ps
`celldefine
module AOI22BX4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, C__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	and (int_fwire_0, B, D);
	not (C__bar, C);
	and (int_fwire_1, B, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.259467:0.409712:1.87742;
		specparam tpd_A_Y_f = 0.228552:0.342611:1.01365;
		specparam tpd_B_Y_r = 0.319371:0.444547:1.63136;
		specparam tpd_B_Y_f = 0.279906:0.390076:1.09599;
		specparam tpd_C_Y_r = 0.311233:0.450057:1.79895;
		specparam tpd_C_Y_f = 0.279899:0.395408:1.1564;
		specparam tpd_D_Y_r = 0.373391:0.499559:1.67408;
		specparam tpd_D_Y_f = 0.332149:0.441884:1.14845;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22B 
`timescale 1ns/10ps
`celldefine
module AOI22BXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, C__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	and (int_fwire_0, B, D);
	not (C__bar, C);
	and (int_fwire_1, B, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0999417:0.238841:1.85144;
		specparam tpd_A_Y_f = 0.0634629:0.149545:1.09718;
		specparam tpd_B_Y_r = 0.167321:0.273956:1.30144;
		specparam tpd_B_Y_f = 0.13136:0.236677:1.07768;
		specparam tpd_C_Y_r = 0.173207:0.305244:1.73937;
		specparam tpd_C_Y_f = 0.126127:0.216734:1.20533;
		specparam tpd_D_Y_r = 0.241396:0.351126:1.38238;
		specparam tpd_D_Y_f = 0.195071:0.301376:1.15218;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22C 
`timescale 1ns/10ps
`celldefine
module AOI22CX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire C__bar, D__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	not (D__bar, D);
	and (int_fwire_0, B, D__bar);
	not (C__bar, C);
	and (int_fwire_1, B, C__bar);
	and (int_fwire_2, A, D__bar);
	and (int_fwire_3, A, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.12747:0.238504:1.20807;
		specparam tpd_A_Y_f = 0.151969:0.257046:0.964858;
		specparam tpd_B_Y_r = 0.143658:0.266914:1.32458;
		specparam tpd_B_Y_f = 0.17695:0.262618:0.869198;
		specparam tpd_C_Y_r = 0.095417:0.218979:1.66235;
		specparam tpd_C_Y_f = 0.0436529:0.126435:0.953455;
		specparam tpd_D_Y_r = 0.119401:0.242516:1.66925;
		specparam tpd_D_Y_f = 0.0525115:0.126608:0.879973;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22C 
`timescale 1ns/10ps
`celldefine
module AOI22CX4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire C__bar, D__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	not (D__bar, D);
	and (int_fwire_0, B, D__bar);
	not (C__bar, C);
	and (int_fwire_1, B, C__bar);
	and (int_fwire_2, A, D__bar);
	and (int_fwire_3, A, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.287036:0.410103:1.49029;
		specparam tpd_A_Y_f = 0.291734:0.423513:1.38591;
		specparam tpd_B_Y_r = 0.304375:0.439749:1.61118;
		specparam tpd_B_Y_f = 0.31654:0.429087:1.27694;
		specparam tpd_C_Y_r = 0.249075:0.382323:1.77944;
		specparam tpd_C_Y_f = 0.182668:0.291341:0.893545;
		specparam tpd_D_Y_r = 0.277184:0.412102:1.82811;
		specparam tpd_D_Y_f = 0.191596:0.293447:0.882017;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22C 
`timescale 1ns/10ps
`celldefine
module AOI22CXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire C__bar, D__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	not (D__bar, D);
	and (int_fwire_0, B, D__bar);
	not (C__bar, C);
	and (int_fwire_1, B, C__bar);
	and (int_fwire_2, A, D__bar);
	and (int_fwire_3, A, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.133128:0.235978:1.14147;
		specparam tpd_A_Y_f = 0.206601:0.328967:1.28004;
		specparam tpd_B_Y_r = 0.154876:0.268297:1.26607;
		specparam tpd_B_Y_f = 0.238314:0.342354:1.16749;
		specparam tpd_C_Y_r = 0.09976:0.227694:1.68257;
		specparam tpd_C_Y_f = 0.0653969:0.166405:1.22393;
		specparam tpd_D_Y_r = 0.117961:0.24578:1.68485;
		specparam tpd_D_Y_f = 0.0755491:0.164703:1.12722;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22 
`timescale 1ns/10ps
`celldefine
module AOI22X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2, int_fwire_3;

	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0820397:0.215811:1.73534;
		specparam tpd_A_Y_f = 0.0468169:0.133826:1.08735;
		specparam tpd_B_Y_r = 0.0977378:0.231445:1.7475;
		specparam tpd_B_Y_f = 0.0533042:0.127399:0.969269;
		specparam tpd_C_Y_r = 0.1325:0.25351:1.58766;
		specparam tpd_C_Y_f = 0.0842717:0.180931:1.14681;
		specparam tpd_D_Y_r = 0.14901:0.271071:1.60815;
		specparam tpd_D_Y_f = 0.091315:0.173124:1.02422;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22 
`timescale 1ns/10ps
`celldefine
module AOI22X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2, int_fwire_3;

	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.242663:0.395315:1.87557;
		specparam tpd_A_Y_f = 0.226055:0.341265:1.03043;
		specparam tpd_B_Y_r = 0.258975:0.412372:1.91689;
		specparam tpd_B_Y_f = 0.234113:0.337307:0.992201;
		specparam tpd_C_Y_r = 0.298566:0.441341:1.8091;
		specparam tpd_C_Y_f = 0.285643:0.402291:1.18994;
		specparam tpd_D_Y_r = 0.314406:0.458771:1.84454;
		specparam tpd_D_Y_f = 0.293865:0.399173:1.13803;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI22 
`timescale 1ns/10ps
`celldefine
module AOI22XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2, int_fwire_3;

	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.115915:0.249013:1.76993;
		specparam tpd_A_Y_f = 0.0723768:0.155374:1.03336;
		specparam tpd_B_Y_r = 0.137695:0.272568:1.8184;
		specparam tpd_B_Y_f = 0.0807842:0.144569:0.878029;
		specparam tpd_C_Y_r = 0.193212:0.319554:1.65988;
		specparam tpd_C_Y_f = 0.134676:0.220791:1.13193;
		specparam tpd_D_Y_r = 0.214952:0.343867:1.70546;
		specparam tpd_D_Y_f = 0.143601:0.210672:0.966684;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI31 
`timescale 1ns/10ps
`celldefine
module AOI31X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_1, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.102141:0.223311:1.59516;
		specparam tpd_A_Y_f = 0.0564063:0.145344:1.03989;
		specparam tpd_B_Y_r = 0.127739:0.249275:1.62436;
		specparam tpd_B_Y_f = 0.0695419:0.148683:0.979247;
		specparam tpd_C_Y_r = 0.149878:0.27408:1.65301;
		specparam tpd_C_Y_f = 0.0777035:0.148552:0.878364;
		specparam tpd_D_Y_r = 0.103781:0.242916:1.81052;
		specparam tpd_D_Y_f = 0.0254866:0.079406:0.694264;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI31 
`timescale 1ns/10ps
`celldefine
module AOI31X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_1, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.246373:0.381169:1.74895;
		specparam tpd_A_Y_f = 0.211027:0.32526:1.05982;
		specparam tpd_B_Y_r = 0.274489:0.410623:1.80665;
		specparam tpd_B_Y_f = 0.224004:0.329915:1.04349;
		specparam tpd_C_Y_r = 0.300248:0.438256:1.85403;
		specparam tpd_C_Y_f = 0.232124:0.330111:1.00134;
		specparam tpd_D_Y_r = 0.25479:0.407774:1.93597;
		specparam tpd_D_Y_f = 0.153744:0.265786:0.918767;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI31 
`timescale 1ns/10ps
`celldefine
module AOI31XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_1, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.114304:0.242392:1.68271;
		specparam tpd_A_Y_f = 0.0635408:0.156311:1.09293;
		specparam tpd_B_Y_r = 0.140674:0.268448:1.71094;
		specparam tpd_B_Y_f = 0.0773628:0.160121:1.02956;
		specparam tpd_C_Y_r = 0.157987:0.286447:1.69699;
		specparam tpd_C_Y_f = 0.0853321:0.159309:0.926565;
		specparam tpd_D_Y_r = 0.0856457:0.227923:1.84991;
		specparam tpd_D_Y_f = 0.0280366:0.0871345:0.748982;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI32 
`timescale 1ns/10ps
`celldefine
module AOI32X1 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;
	wire int_fwire_4, int_fwire_5;

	not (E__bar, E);
	not (C__bar, C);
	and (int_fwire_0, C__bar, E__bar);
	not (D__bar, D);
	and (int_fwire_1, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_2, B__bar, E__bar);
	and (int_fwire_3, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_4, A__bar, E__bar);
	and (int_fwire_5, A__bar, D__bar);
	or (Y, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.106697:0.237334:1.73616;
		specparam tpd_A_Y_f = 0.0548275:0.134501:0.975399;
		specparam tpd_B_Y_r = 0.134339:0.2647:1.76542;
		specparam tpd_B_Y_f = 0.0692507:0.140486:0.923705;
		specparam tpd_C_Y_r = 0.157023:0.287904:1.78854;
		specparam tpd_C_Y_f = 0.077328:0.141078:0.830807;
		specparam tpd_D_Y_r = 0.194513:0.315339:1.63029;
		specparam tpd_D_Y_f = 0.0895281:0.174519:0.950554;
		specparam tpd_E_Y_r = 0.215894:0.337657:1.65322;
		specparam tpd_E_Y_f = 0.0967355:0.170968:0.872885;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI32 
`timescale 1ns/10ps
`celldefine
module AOI32X4 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;
	wire int_fwire_4, int_fwire_5;

	not (E__bar, E);
	not (C__bar, C);
	and (int_fwire_0, C__bar, E__bar);
	not (D__bar, D);
	and (int_fwire_1, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_2, B__bar, E__bar);
	and (int_fwire_3, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_4, A__bar, E__bar);
	and (int_fwire_5, A__bar, D__bar);
	or (Y, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.265597:0.416612:1.93141;
		specparam tpd_A_Y_f = 0.214922:0.321249:0.905313;
		specparam tpd_B_Y_r = 0.295922:0.446541:1.9913;
		specparam tpd_B_Y_f = 0.229361:0.327704:0.896402;
		specparam tpd_C_Y_r = 0.32116:0.472083:2.03588;
		specparam tpd_C_Y_f = 0.237453:0.328496:0.865486;
		specparam tpd_D_Y_r = 0.35726:0.496993:1.90621;
		specparam tpd_D_Y_f = 0.241368:0.356866:1.03145;
		specparam tpd_E_Y_r = 0.380389:0.522177:1.94388;
		specparam tpd_E_Y_f = 0.248607:0.353283:0.996964;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI32 
`timescale 1ns/10ps
`celldefine
module AOI32XL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;
	wire int_fwire_4, int_fwire_5;

	not (E__bar, E);
	not (C__bar, C);
	and (int_fwire_0, C__bar, E__bar);
	not (D__bar, D);
	and (int_fwire_1, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_2, B__bar, E__bar);
	and (int_fwire_3, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_4, A__bar, E__bar);
	and (int_fwire_5, A__bar, D__bar);
	or (Y, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0821782:0.221565:1.81152;
		specparam tpd_A_Y_f = 0.0599524:0.147423:1.08763;
		specparam tpd_B_Y_r = 0.112199:0.250091:1.84069;
		specparam tpd_B_Y_f = 0.0774139:0.155443:1.03007;
		specparam tpd_C_Y_r = 0.129537:0.267499:1.84723;
		specparam tpd_C_Y_f = 0.0846287:0.15366:0.924515;
		specparam tpd_D_Y_r = 0.212361:0.344016:1.7452;
		specparam tpd_D_Y_f = 0.116822:0.207809:1.1139;
		specparam tpd_E_Y_r = 0.226147:0.356919:1.72442;
		specparam tpd_E_Y_f = 0.125016:0.205674:1.02386;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI33 
`timescale 1ns/10ps
`celldefine
module AOI33X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;

	not (F__bar, F);
	not (C__bar, C);
	and (int_fwire_0, C__bar, F__bar);
	not (E__bar, E);
	and (int_fwire_1, C__bar, E__bar);
	not (D__bar, D);
	and (int_fwire_2, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_3, B__bar, F__bar);
	and (int_fwire_4, B__bar, E__bar);
	and (int_fwire_5, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_6, A__bar, F__bar);
	and (int_fwire_7, A__bar, E__bar);
	and (int_fwire_8, A__bar, D__bar);
	or (Y, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.208976:0.330655:1.63579;
		specparam tpd_A_Y_f = 0.12365:0.212266:1.11741;
		specparam tpd_B_Y_r = 0.232534:0.354901:1.66333;
		specparam tpd_B_Y_f = 0.135752:0.214048:1.03409;
		specparam tpd_C_Y_r = 0.254737:0.378613:1.68997;
		specparam tpd_C_Y_f = 0.143317:0.209918:0.908621;
		specparam tpd_D_Y_r = 0.138084:0.26855:1.75873;
		specparam tpd_D_Y_f = 0.0614139:0.14517:1.0299;
		specparam tpd_E_Y_r = 0.165687:0.2945:1.79164;
		specparam tpd_E_Y_f = 0.0756509:0.147522:0.949415;
		specparam tpd_F_Y_r = 0.188193:0.319163:1.81657;
		specparam tpd_F_Y_f = 0.0833433:0.145232:0.830759;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI33 
`timescale 1ns/10ps
`celldefine
module AOI33X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;

	not (F__bar, F);
	not (C__bar, C);
	and (int_fwire_0, C__bar, F__bar);
	not (E__bar, E);
	and (int_fwire_1, C__bar, E__bar);
	not (D__bar, D);
	and (int_fwire_2, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_3, B__bar, F__bar);
	and (int_fwire_4, B__bar, E__bar);
	and (int_fwire_5, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_6, A__bar, F__bar);
	and (int_fwire_7, A__bar, E__bar);
	and (int_fwire_8, A__bar, D__bar);
	or (Y, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.37523:0.517041:1.92498;
		specparam tpd_A_Y_f = 0.293534:0.406061:1.13558;
		specparam tpd_B_Y_r = 0.400473:0.543803:1.97406;
		specparam tpd_B_Y_f = 0.305587:0.407402:1.09171;
		specparam tpd_C_Y_r = 0.424513:0.569439:2.01845;
		specparam tpd_C_Y_f = 0.313135:0.403515:1.01319;
		specparam tpd_D_Y_r = 0.304165:0.455607:1.99457;
		specparam tpd_D_Y_f = 0.235955:0.347151:0.988998;
		specparam tpd_E_Y_r = 0.333844:0.485579:2.05962;
		specparam tpd_E_Y_f = 0.250143:0.350362:0.953468;
		specparam tpd_F_Y_r = 0.358537:0.51049:2.11031;
		specparam tpd_F_Y_f = 0.257842:0.347758:0.893708;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: AOI33 
`timescale 1ns/10ps
`celldefine
module AOI33XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;

	not (F__bar, F);
	not (C__bar, C);
	and (int_fwire_0, C__bar, F__bar);
	not (E__bar, E);
	and (int_fwire_1, C__bar, E__bar);
	not (D__bar, D);
	and (int_fwire_2, C__bar, D__bar);
	not (B__bar, B);
	and (int_fwire_3, B__bar, F__bar);
	and (int_fwire_4, B__bar, E__bar);
	and (int_fwire_5, B__bar, D__bar);
	not (A__bar, A);
	and (int_fwire_6, A__bar, F__bar);
	and (int_fwire_7, A__bar, E__bar);
	and (int_fwire_8, A__bar, D__bar);
	or (Y, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.274327:0.392678:1.63717;
		specparam tpd_A_Y_f = 0.121576:0.200189:0.902956;
		specparam tpd_B_Y_r = 0.312171:0.432685:1.70226;
		specparam tpd_B_Y_f = 0.134076:0.201877:0.83049;
		specparam tpd_C_Y_r = 0.347643:0.470705:1.74926;
		specparam tpd_C_Y_f = 0.142434:0.199059:0.713217;
		specparam tpd_D_Y_r = 0.192818:0.318594:1.76867;
		specparam tpd_D_Y_f = 0.0654736:0.137247:0.811463;
		specparam tpd_E_Y_r = 0.234414:0.360533:1.82821;
		specparam tpd_E_Y_f = 0.0803489:0.14092:0.744326;
		specparam tpd_F_Y_r = 0.265773:0.392306:1.86533;
		specparam tpd_F_Y_f = 0.0879229:0.138968:0.635341;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BKEEP 
`timescale 1ns/10ps
`celldefine
module BKEEP (Y);
	inout Y;
	//Function
	wire io_wire;
	buf(weak0,weak1) I0(Y, io_wire);
	buf              I1(io_wire, Y);
	// Timing
	specify

	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX1 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0717461:0.192509:1.33359;
		specparam tpd_A_Y_f = 0.0804106:0.197769:1.07408;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX12 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0873623:0.224895:1.4169;
		specparam tpd_A_Y_f = 0.0943118:0.219778:1.04193;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX16 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0915989:0.233201:1.44065;
		specparam tpd_A_Y_f = 0.10836:0.242622:1.13018;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX2 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0627298:0.176239:1.26226;
		specparam tpd_A_Y_f = 0.0817201:0.201476:1.07523;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX20 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0929329:0.235338:1.44169;
		specparam tpd_A_Y_f = 0.113758:0.253274:1.20121;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX24 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.091824:0.231192:1.41656;
		specparam tpd_A_Y_f = 0.106918:0.238774:1.09652;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX3 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0646799:0.186413:1.30902;
		specparam tpd_A_Y_f = 0.0881781:0.215296:1.11469;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX30 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.101776:0.247737:1.46576;
		specparam tpd_A_Y_f = 0.122784:0.261747:1.17638;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX36 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.112497:0.262414:1.49208;
		specparam tpd_A_Y_f = 0.138746:0.281999:1.22689;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX4 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0751946:0.205456:1.35104;
		specparam tpd_A_Y_f = 0.107612:0.243353:1.18205;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX6 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0794808:0.211863:1.41168;
		specparam tpd_A_Y_f = 0.082333:0.203914:1.04713;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFX8 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.073856:0.203175:1.34339;
		specparam tpd_A_Y_f = 0.0993963:0.229456:1.11141;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: BUF 
`timescale 1ns/10ps
`celldefine
module BUFXL (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0925589:0.207856:1.28375;
		specparam tpd_A_Y_f = 0.117787:0.260989:1.37088;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKAND2 
`timescale 1ns/10ps
`celldefine
module CKAND2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0943631:0.225447:1.41534;
		specparam tpd_A_Y_f = 0.0979449:0.246797:1.51513;
		specparam tpd_B_Y_r = 0.101874:0.221516:1.37612;
		specparam tpd_B_Y_f = 0.109807:0.264336:1.5738;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKAND2 
`timescale 1ns/10ps
`celldefine
module CKAND2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.109648:0.252161:1.45611;
		specparam tpd_A_Y_f = 0.119526:0.281851:1.59417;
		specparam tpd_B_Y_r = 0.117299:0.246498:1.40584;
		specparam tpd_B_Y_f = 0.133009:0.299639:1.65094;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKAND2 
`timescale 1ns/10ps
`celldefine
module CKAND2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.139928:0.297144:1.55957;
		specparam tpd_A_Y_f = 0.156052:0.326559:1.64905;
		specparam tpd_B_Y_r = 0.147418:0.289591:1.50057;
		specparam tpd_B_Y_f = 0.171026:0.346533:1.7068;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKAND2 
`timescale 1ns/10ps
`celldefine
module CKAND2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.107373:0.238554:1.37223;
		specparam tpd_A_Y_f = 0.13672:0.311666:1.85198;
		specparam tpd_B_Y_r = 0.115529:0.233975:1.32657;
		specparam tpd_B_Y_f = 0.154973:0.333979:1.91986;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKAND3 
`timescale 1ns/10ps
`celldefine
module CKAND3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0996915:0.231011:1.42166;
		specparam tpd_A_Y_f = 0.100683:0.249341:1.51452;
		specparam tpd_B_Y_r = 0.114127:0.237502:1.40442;
		specparam tpd_B_Y_f = 0.115841:0.270197:1.57278;
		specparam tpd_C_Y_r = 0.121135:0.237403:1.36918;
		specparam tpd_C_Y_f = 0.125917:0.284402:1.61493;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKAND3 
`timescale 1ns/10ps
`celldefine
module CKAND3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.10407:0.241136:1.41921;
		specparam tpd_A_Y_f = 0.111026:0.267728:1.53594;
		specparam tpd_B_Y_r = 0.117805:0.246006:1.39982;
		specparam tpd_B_Y_f = 0.126102:0.286985:1.59082;
		specparam tpd_C_Y_r = 0.124893:0.244142:1.35426;
		specparam tpd_C_Y_f = 0.137392:0.301268:1.63669;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKAND3 
`timescale 1ns/10ps
`celldefine
module CKAND3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.124959:0.274664:1.49037;
		specparam tpd_A_Y_f = 0.135761:0.30013:1.57176;
		specparam tpd_B_Y_r = 0.138829:0.27636:1.45526;
		specparam tpd_B_Y_f = 0.151241:0.319418:1.62797;
		specparam tpd_C_Y_r = 0.14558:0.272838:1.40003;
		specparam tpd_C_Y_f = 0.162685:0.330867:1.67038;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKAND3 
`timescale 1ns/10ps
`celldefine
module CKAND3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.132908:0.274387:1.48187;
		specparam tpd_A_Y_f = 0.133106:0.30482:1.79704;
		specparam tpd_B_Y_r = 0.147492:0.278507:1.45474;
		specparam tpd_B_Y_f = 0.152247:0.329227:1.86391;
		specparam tpd_C_Y_r = 0.15536:0.276296:1.4021;
		specparam tpd_C_Y_f = 0.166521:0.345438:1.91551;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX1 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0717543:0.191244:1.34963;
		specparam tpd_A_Y_f = 0.0728464:0.181832:1.03353;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX12 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0817996:0.219841:1.4381;
		specparam tpd_A_Y_f = 0.0893235:0.232234:1.37326;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX16 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0941527:0.241599:1.50027;
		specparam tpd_A_Y_f = 0.101267:0.250929:1.40921;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX2 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0872703:0.224361:1.49615;
		specparam tpd_A_Y_f = 0.0767152:0.203664:1.25554;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX20 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.092842:0.240339:1.49883;
		specparam tpd_A_Y_f = 0.102634:0.254522:1.43246;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX24 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0908246:0.237125:1.49084;
		specparam tpd_A_Y_f = 0.102948:0.255184:1.44802;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX3 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0740797:0.204606:1.37776;
		specparam tpd_A_Y_f = 0.0899133:0.22807:1.3183;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX30 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.102283:0.253209:1.51601;
		specparam tpd_A_Y_f = 0.116295:0.272087:1.45387;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX36 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.113214:0.268297:1.5379;
		specparam tpd_A_Y_f = 0.129711:0.288972:1.48094;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX4 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.070809:0.199207:1.34107;
		specparam tpd_A_Y_f = 0.105056:0.245192:1.26772;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX6 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0836768:0.221094:1.43487;
		specparam tpd_A_Y_f = 0.0912495:0.234453:1.38618;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFX8 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0800476:0.217616:1.43634;
		specparam tpd_A_Y_f = 0.0884087:0.231305:1.38284;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKBUF 
`timescale 1ns/10ps
`celldefine
module CKBUFXL (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0897882:0.217644:1.43879;
		specparam tpd_A_Y_f = 0.0921425:0.244911:1.71938;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX1 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0291324:0.170319:1.78355;
		specparam tpd_A_Y_f = 0.0290559:0.156066:1.6515;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX12 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.203818:0.363839:1.76928;
		specparam tpd_A_Y_f = 0.196614:0.336085:1.34252;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX16 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.219473:0.383495:1.81241;
		specparam tpd_A_Y_f = 0.212306:0.360901:1.46374;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX2 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0268728:0.167532:1.78176;
		specparam tpd_A_Y_f = 0.0262293:0.152046:1.62902;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX20 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.24068:0.404656:1.85517;
		specparam tpd_A_Y_f = 0.231317:0.37932:1.45948;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX24 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.258427:0.424058:1.86801;
		specparam tpd_A_Y_f = 0.251139:0.405374:1.57627;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX3 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0263758:0.167445:1.78259;
		specparam tpd_A_Y_f = 0.0253771:0.147185:1.58466;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX30 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.272838:0.441614:1.904;
		specparam tpd_A_Y_f = 0.271761:0.429662:1.60385;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX36 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.289906:0.460447:1.91175;
		specparam tpd_A_Y_f = 0.292166:0.452467:1.6177;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX4 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0254963:0.165262:1.77186;
		specparam tpd_A_Y_f = 0.024213:0.144218:1.56108;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX6 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.169288:0.323663:1.67894;
		specparam tpd_A_Y_f = 0.165969:0.30294:1.37463;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVX8 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.170226:0.325398:1.70097;
		specparam tpd_A_Y_f = 0.169799:0.30896:1.39087;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKINV 
`timescale 1ns/10ps
`celldefine
module CKINVXL (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0304831:0.171036:1.7717;
		specparam tpd_A_Y_f = 0.0340005:0.170179:1.79973;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKMUX2 
`timescale 1ns/10ps
`celldefine
module CKMUX2X1 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire int_fwire_0, int_fwire_1, S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.147496:0.296386:1.55909;
		specparam tpd_D0_Y_f = 0.154923:0.316071:1.50529;
		specparam tpd_D1_Y_r = 0.148503:0.29891:1.5623;
		specparam tpd_D1_Y_f = 0.158917:0.320922:1.51786;
		specparam tpd_S_Y_posedge_r = 0.10881:0.249189:1.45256;
		specparam tpd_S_Y_posedge_f = 0.126836:0.281192:1.47751;
		specparam tpd_S_Y_negedge_r = 0.141578:0.298986:1.61443;
		specparam tpd_S_Y_negedge_f = 0.140527:0.290322:1.25729;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: CKMUX2 
`timescale 1ns/10ps
`celldefine
module CKMUX2X2 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire int_fwire_0, int_fwire_1, S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.156873:0.315111:1.61347;
		specparam tpd_D0_Y_f = 0.169729:0.340053:1.54575;
		specparam tpd_D1_Y_r = 0.159879:0.320145:1.62366;
		specparam tpd_D1_Y_f = 0.174742:0.346167:1.5596;
		specparam tpd_S_Y_posedge_r = 0.121825:0.274988:1.52528;
		specparam tpd_S_Y_posedge_f = 0.145536:0.310896:1.52927;
		specparam tpd_S_Y_negedge_r = 0.151165:0.318183:1.65953;
		specparam tpd_S_Y_negedge_f = 0.153499:0.313986:1.28333;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: CKMUX2 
`timescale 1ns/10ps
`celldefine
module CKMUX2X4 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire int_fwire_0, int_fwire_1, S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.194455:0.362086:1.68674;
		specparam tpd_D0_Y_f = 0.220096:0.40228:1.65762;
		specparam tpd_D1_Y_r = 0.196389:0.36595:1.69323;
		specparam tpd_D1_Y_f = 0.22369:0.406252:1.66867;
		specparam tpd_S_Y_posedge_r = 0.160357:0.323756:1.61538;
		specparam tpd_S_Y_posedge_f = 0.197037:0.372716:1.63784;
		specparam tpd_S_Y_negedge_r = 0.184461:0.36062:1.68901;
		specparam tpd_S_Y_negedge_f = 0.198748:0.370421:1.36858;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: CKMUX2 
`timescale 1ns/10ps
`celldefine
module CKMUX2XL (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire int_fwire_0, int_fwire_1, S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.165487:0.310976:1.55107;
		specparam tpd_D0_Y_f = 0.164545:0.331196:1.60297;
		specparam tpd_D1_Y_r = 0.165566:0.31194:1.55918;
		specparam tpd_D1_Y_f = 0.165696:0.331551:1.59542;
		specparam tpd_S_Y_posedge_r = 0.123723:0.264105:1.4559;
		specparam tpd_S_Y_posedge_f = 0.139583:0.300399:1.58146;
		specparam tpd_S_Y_negedge_r = 0.157988:0.322178:1.68299;
		specparam tpd_S_Y_negedge_f = 0.144691:0.2955:1.27139;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: CKMUX3 
`timescale 1ns/10ps
`celldefine
module CKMUX3X1 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	and (int_fwire_0, D2, S1);
	not (S1__bar, S1);
	and (int_fwire_1, D1, S0, S1__bar);
	not (S0__bar, S0);
	and (int_fwire_2, D0, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.242607:0.400475:1.69618;
		specparam tpd_D0_Y_f = 0.273072:0.461152:1.7201;
		specparam tpd_D1_Y_r = 0.252986:0.416375:1.7683;
		specparam tpd_D1_Y_f = 0.258113:0.434445:1.60557;
		specparam tpd_D2_Y_r = 0.137053:0.280388:1.55011;
		specparam tpd_D2_Y_f = 0.14004:0.284203:1.34854;
		specparam tpd_S0_Y_posedge_r = 0.22289:0.383536:1.69188;
		specparam tpd_S0_Y_posedge_f = 0.26344:0.451156:1.76816;
		specparam tpd_S0_Y_negedge_r = 0.257198:0.437284:1.8685;
		specparam tpd_S0_Y_negedge_f = 0.248685:0.42407:1.35533;
		specparam tpd_S1_Y_posedge_r = 0.109054:0.247177:1.37746;
		specparam tpd_S1_Y_posedge_f = 0.150802:0.329258:1.63201;
		specparam tpd_S1_Y_negedge_r = 0.169734:0.346529:1.75374;
		specparam tpd_S1_Y_negedge_f = 0.137715:0.282021:1.14749;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: CKMUX3 
`timescale 1ns/10ps
`celldefine
module CKMUX3X2 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	and (int_fwire_0, D2, S1);
	not (S1__bar, S1);
	and (int_fwire_1, D1, S0, S1__bar);
	not (S0__bar, S0);
	and (int_fwire_2, D0, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.265424:0.433366:1.75727;
		specparam tpd_D0_Y_f = 0.304209:0.499504:1.73317;
		specparam tpd_D1_Y_r = 0.277237:0.450752:1.83083;
		specparam tpd_D1_Y_f = 0.287558:0.470908:1.61464;
		specparam tpd_D2_Y_r = 0.150847:0.304612:1.5992;
		specparam tpd_D2_Y_f = 0.158116:0.311631:1.35028;
		specparam tpd_S0_Y_posedge_r = 0.247582:0.418551:1.76408;
		specparam tpd_S0_Y_posedge_f = 0.295626:0.490784:1.78272;
		specparam tpd_S0_Y_negedge_r = 0.27937:0.469441:1.91489;
		specparam tpd_S0_Y_negedge_f = 0.277269:0.459934:1.35904;
		specparam tpd_S1_Y_posedge_r = 0.125559:0.278147:1.46439;
		specparam tpd_S1_Y_posedge_f = 0.184013:0.373336:1.65832;
		specparam tpd_S1_Y_negedge_r = 0.189012:0.378052:1.80447;
		specparam tpd_S1_Y_negedge_f = 0.152659:0.308212:1.13302;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: CKMUX3 
`timescale 1ns/10ps
`celldefine
module CKMUX3X4 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	and (int_fwire_0, D2, S1);
	not (S1__bar, S1);
	and (int_fwire_1, D1, S0, S1__bar);
	not (S0__bar, S0);
	and (int_fwire_2, D0, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.329728:0.504448:1.83853;
		specparam tpd_D0_Y_f = 0.390144:0.587706:1.80642;
		specparam tpd_D1_Y_r = 0.34498:0.525185:1.91433;
		specparam tpd_D1_Y_f = 0.369618:0.555315:1.68146;
		specparam tpd_D2_Y_r = 0.196513:0.35925:1.66323;
		specparam tpd_D2_Y_f = 0.210674:0.371524:1.38822;
		specparam tpd_S0_Y_posedge_r = 0.315802:0.493089:1.86412;
		specparam tpd_S0_Y_posedge_f = 0.38268:0.580222:1.85457;
		specparam tpd_S0_Y_negedge_r = 0.342483:0.539157:1.97074;
		specparam tpd_S0_Y_negedge_f = 0.358245:0.542942:1.41782;
		specparam tpd_S1_Y_posedge_r = 0.174133:0.336496:1.58105;
		specparam tpd_S1_Y_posedge_f = 0.277467:0.472011:1.74362;
		specparam tpd_S1_Y_negedge_r = 0.251597:0.448138:1.86915;
		specparam tpd_S1_Y_negedge_f = 0.202052:0.364308:1.16077;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND2 
`timescale 1ns/10ps
`celldefine
module CKNAND2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0390359:0.180113:1.7745;
		specparam tpd_A_Y_f = 0.039952:0.162432:1.62956;
		specparam tpd_B_Y_r = 0.0485842:0.192805:1.8029;
		specparam tpd_B_Y_f = 0.048035:0.15761:1.51451;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND2 
`timescale 1ns/10ps
`celldefine
module CKNAND2X12 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.191932:0.35276:1.77263;
		specparam tpd_A_Y_f = 0.191324:0.333129:1.48673;
		specparam tpd_B_Y_r = 0.205853:0.368456:1.83019;
		specparam tpd_B_Y_f = 0.19798:0.326479:1.43242;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND2 
`timescale 1ns/10ps
`celldefine
module CKNAND2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0371177:0.179243:1.78483;
		specparam tpd_A_Y_f = 0.0418465:0.175581:1.77549;
		specparam tpd_B_Y_r = 0.0445969:0.188433:1.79429;
		specparam tpd_B_Y_f = 0.0492201:0.170034:1.6667;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND2 
`timescale 1ns/10ps
`celldefine
module CKNAND2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0343618:0.175297:1.77462;
		specparam tpd_A_Y_f = 0.0334824:0.151615:1.5675;
		specparam tpd_B_Y_r = 0.0433792:0.186637:1.78579;
		specparam tpd_B_Y_f = 0.0410603:0.147032:1.45547;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND2 
`timescale 1ns/10ps
`celldefine
module CKNAND2X6 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.192348:0.349556:1.71467;
		specparam tpd_A_Y_f = 0.203035:0.360188:1.7657;
		specparam tpd_B_Y_r = 0.20741:0.366241:1.77047;
		specparam tpd_B_Y_f = 0.210482:0.353485:1.70793;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND2 
`timescale 1ns/10ps
`celldefine
module CKNAND2X8 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.171902:0.328312:1.71799;
		specparam tpd_A_Y_f = 0.177344:0.315884:1.46329;
		specparam tpd_B_Y_r = 0.182186:0.341707:1.76673;
		specparam tpd_B_Y_f = 0.184193:0.310696:1.41914;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND2 
`timescale 1ns/10ps
`celldefine
module CKNAND2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0434059:0.189024:1.8265;
		specparam tpd_A_Y_f = 0.0461742:0.171425:1.69368;
		specparam tpd_B_Y_r = 0.0523847:0.19941:1.83741;
		specparam tpd_B_Y_f = 0.0547571:0.165067:1.56401;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND3 
`timescale 1ns/10ps
`celldefine
module CKNAND3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0469567:0.18922:1.78741;
		specparam tpd_A_Y_f = 0.0450553:0.162928:1.57603;
		specparam tpd_B_Y_r = 0.0606402:0.204286:1.80384;
		specparam tpd_B_Y_f = 0.0594444:0.166075:1.49224;
		specparam tpd_C_Y_r = 0.0699165:0.215301:1.81639;
		specparam tpd_C_Y_f = 0.0670532:0.164815:1.38239;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND3 
`timescale 1ns/10ps
`celldefine
module CKNAND3X12 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.235878:0.399485:1.881;
		specparam tpd_A_Y_f = 0.218681:0.354519:1.45412;
		specparam tpd_B_Y_r = 0.252327:0.417492:1.93215;
		specparam tpd_B_Y_f = 0.232033:0.356671:1.41979;
		specparam tpd_C_Y_r = 0.265714:0.431316:1.9725;
		specparam tpd_C_Y_f = 0.23894:0.352543:1.35655;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND3 
`timescale 1ns/10ps
`celldefine
module CKNAND3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0442016:0.186334:1.77932;
		specparam tpd_A_Y_f = 0.0407098:0.153311:1.50836;
		specparam tpd_B_Y_r = 0.0573544:0.200936:1.79299;
		specparam tpd_B_Y_f = 0.0543523:0.157789:1.44221;
		specparam tpd_C_Y_r = 0.0666801:0.211805:1.80617;
		specparam tpd_C_Y_f = 0.0617624:0.156219:1.33366;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND3 
`timescale 1ns/10ps
`celldefine
module CKNAND3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.159482:0.309313:1.68198;
		specparam tpd_A_Y_f = 0.187757:0.296552:1.00991;
		specparam tpd_B_Y_r = 0.174894:0.32854:1.74317;
		specparam tpd_B_Y_f = 0.200843:0.300963:0.988068;
		specparam tpd_C_Y_r = 0.187991:0.343877:1.79274;
		specparam tpd_C_Y_f = 0.208596:0.30037:0.940847;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND3 
`timescale 1ns/10ps
`celldefine
module CKNAND3X8 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.20341:0.364338:1.82378;
		specparam tpd_A_Y_f = 0.19854:0.331982:1.41364;
		specparam tpd_B_Y_r = 0.21965:0.382682:1.87923;
		specparam tpd_B_Y_f = 0.212124:0.334949:1.38337;
		specparam tpd_C_Y_r = 0.232729:0.396291:1.91953;
		specparam tpd_C_Y_f = 0.219324:0.332255:1.32947;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNAND3 
`timescale 1ns/10ps
`celldefine
module CKNAND3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0615725:0.204812:1.8021;
		specparam tpd_A_Y_f = 0.0601018:0.175104:1.55268;
		specparam tpd_B_Y_r = 0.0785668:0.223098:1.84042;
		specparam tpd_B_Y_f = 0.0769944:0.180044:1.4645;
		specparam tpd_C_Y_r = 0.0854254:0.228856:1.81383;
		specparam tpd_C_Y_f = 0.0847021:0.177862:1.34783;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR2 
`timescale 1ns/10ps
`celldefine
module CKNOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0413049:0.171852:1.69114;
		specparam tpd_A_Y_f = 0.0478632:0.170477:1.6209;
		specparam tpd_B_Y_r = 0.0630866:0.176423:1.52041;
		specparam tpd_B_Y_f = 0.0754587:0.201907:1.65501;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR2 
`timescale 1ns/10ps
`celldefine
module CKNOR2X12 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.195115:0.341407:1.67023;
		specparam tpd_A_Y_f = 0.196399:0.33936:1.46366;
		specparam tpd_B_Y_r = 0.217447:0.348689:1.59215;
		specparam tpd_B_Y_f = 0.234082:0.381437:1.5931;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR2 
`timescale 1ns/10ps
`celldefine
module CKNOR2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.036202:0.165838:1.68399;
		specparam tpd_A_Y_f = 0.0371376:0.153798:1.49529;
		specparam tpd_B_Y_r = 0.0584387:0.171199:1.50807;
		specparam tpd_B_Y_f = 0.0584426:0.182086:1.52548;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR2 
`timescale 1ns/10ps
`celldefine
module CKNOR2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.182321:0.324893:1.64542;
		specparam tpd_A_Y_f = 0.198007:0.318452:1.17403;
		specparam tpd_B_Y_r = 0.203772:0.332881:1.58396;
		specparam tpd_B_Y_f = 0.233227:0.358511:1.28798;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR2 
`timescale 1ns/10ps
`celldefine
module CKNOR2X6 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.205884:0.356413:1.73599;
		specparam tpd_A_Y_f = 0.214225:0.359594:1.58183;
		specparam tpd_B_Y_r = 0.228058:0.362885:1.67188;
		specparam tpd_B_Y_f = 0.239713:0.388169:1.663;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR2 
`timescale 1ns/10ps
`celldefine
module CKNOR2X8 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.173537:0.314639:1.59582;
		specparam tpd_A_Y_f = 0.174738:0.319113:1.51257;
		specparam tpd_B_Y_r = 0.196122:0.324045:1.52635;
		specparam tpd_B_Y_f = 0.211314:0.363043:1.64925;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR2 
`timescale 1ns/10ps
`celldefine
module CKNOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0470974:0.181329:1.72779;
		specparam tpd_A_Y_f = 0.0489352:0.157641:1.46299;
		specparam tpd_B_Y_r = 0.0707864:0.187836:1.56019;
		specparam tpd_B_Y_f = 0.0754667:0.18902:1.49879;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR3 
`timescale 1ns/10ps
`celldefine
module CKNOR3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.045382:0.169825:1.62616;
		specparam tpd_A_Y_f = 0.0553433:0.171476:1.46945;
		specparam tpd_B_Y_r = 0.0936315:0.207238:1.53702;
		specparam tpd_B_Y_f = 0.0921218:0.206733:1.47885;
		specparam tpd_C_Y_r = 0.113875:0.223515:1.39306;
		specparam tpd_C_Y_f = 0.114647:0.236145:1.5581;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR3 
`timescale 1ns/10ps
`celldefine
module CKNOR3X12 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.268845:0.418833:1.8038;
		specparam tpd_A_Y_f = 0.235153:0.378758:1.54665;
		specparam tpd_B_Y_r = 0.320456:0.458668:1.78388;
		specparam tpd_B_Y_f = 0.2778:0.420026:1.64543;
		specparam tpd_C_Y_r = 0.341314:0.475102:1.68909;
		specparam tpd_C_Y_f = 0.325704:0.469075:1.77481;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR3 
`timescale 1ns/10ps
`celldefine
module CKNOR3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0512258:0.17908:1.65193;
		specparam tpd_A_Y_f = 0.0480445:0.1447:1.1939;
		specparam tpd_B_Y_r = 0.105249:0.221233:1.5773;
		specparam tpd_B_Y_f = 0.0780113:0.181046:1.24536;
		specparam tpd_C_Y_r = 0.127059:0.239806:1.43825;
		specparam tpd_C_Y_f = 0.0927718:0.207254:1.35392;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR3 
`timescale 1ns/10ps
`celldefine
module CKNOR3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.191065:0.329272:1.6295;
		specparam tpd_A_Y_f = 0.19812:0.315825:1.03227;
		specparam tpd_B_Y_r = 0.24791:0.378265:1.6455;
		specparam tpd_B_Y_f = 0.243689:0.362353:1.14619;
		specparam tpd_C_Y_r = 0.269837:0.397902:1.58238;
		specparam tpd_C_Y_f = 0.273398:0.393644:1.24311;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR3 
`timescale 1ns/10ps
`celldefine
module CKNOR3X8 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.299908:0.429676:1.61055;
		specparam tpd_A_Y_f = 0.291444:0.432669:1.69666;
		specparam tpd_B_Y_r = 0.279771:0.414219:1.69398;
		specparam tpd_B_Y_f = 0.253347:0.393521:1.58382;
		specparam tpd_C_Y_r = 0.229956:0.375966:1.70901;
		specparam tpd_C_Y_f = 0.210625:0.351305:1.47935;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKNOR3 
`timescale 1ns/10ps
`celldefine
module CKNOR3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.063784:0.192005:1.6616;
		specparam tpd_A_Y_f = 0.0701247:0.17408:1.36699;
		specparam tpd_B_Y_r = 0.113894:0.227078:1.56937;
		specparam tpd_B_Y_f = 0.101307:0.200718:1.32203;
		specparam tpd_C_Y_r = 0.135363:0.245479:1.43834;
		specparam tpd_C_Y_f = 0.126873:0.232411:1.41399;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKOR2 
`timescale 1ns/10ps
`celldefine
module CKOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0990305:0.232111:1.46191;
		specparam tpd_A_Y_f = 0.108082:0.254387:1.50855;
		specparam tpd_B_Y_r = 0.12089:0.260371:1.53405;
		specparam tpd_B_Y_f = 0.130167:0.264423:1.48147;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKOR2 
`timescale 1ns/10ps
`celldefine
module CKOR2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.123814:0.270721:1.57681;
		specparam tpd_A_Y_f = 0.130489:0.288684:1.5462;
		specparam tpd_B_Y_r = 0.146393:0.296143:1.63951;
		specparam tpd_B_Y_f = 0.152318:0.295922:1.50571;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKOR2 
`timescale 1ns/10ps
`celldefine
module CKOR2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.156238:0.313884:1.64837;
		specparam tpd_A_Y_f = 0.172513:0.338506:1.60519;
		specparam tpd_B_Y_r = 0.175514:0.33322:1.69241;
		specparam tpd_B_Y_f = 0.194478:0.346792:1.5468;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKOR2 
`timescale 1ns/10ps
`celldefine
module CKOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.125708:0.259479:1.49393;
		specparam tpd_A_Y_f = 0.134163:0.2997:1.79257;
		specparam tpd_B_Y_r = 0.168106:0.310187:1.6294;
		specparam tpd_B_Y_f = 0.158263:0.310646:1.72821;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKOR3 
`timescale 1ns/10ps
`celldefine
module CKOR3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.105681:0.245229:1.51442;
		specparam tpd_A_Y_f = 0.105921:0.252619:1.42949;
		specparam tpd_B_Y_r = 0.14678:0.291846:1.62408;
		specparam tpd_B_Y_f = 0.156256:0.295051:1.45379;
		specparam tpd_C_Y_r = 0.170829:0.322186:1.72559;
		specparam tpd_C_Y_f = 0.176613:0.313135:1.39814;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKOR3 
`timescale 1ns/10ps
`celldefine
module CKOR3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.113724:0.261369:1.55557;
		specparam tpd_A_Y_f = 0.11792:0.273886:1.46188;
		specparam tpd_B_Y_r = 0.153712:0.304428:1.65627;
		specparam tpd_B_Y_f = 0.169097:0.315019:1.47733;
		specparam tpd_C_Y_r = 0.177215:0.333193:1.75115;
		specparam tpd_C_Y_f = 0.189675:0.332583:1.41687;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKOR3 
`timescale 1ns/10ps
`celldefine
module CKOR3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.137322:0.294211:1.62644;
		specparam tpd_A_Y_f = 0.153169:0.318757:1.52594;
		specparam tpd_B_Y_r = 0.176315:0.334314:1.71585;
		specparam tpd_B_Y_f = 0.204623:0.358622:1.52831;
		specparam tpd_C_Y_r = 0.201245:0.363782:1.80185;
		specparam tpd_C_Y_f = 0.225312:0.37521:1.45726;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CKOR3 
`timescale 1ns/10ps
`celldefine
module CKOR3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.132172:0.266674:1.46862;
		specparam tpd_A_Y_f = 0.151475:0.304285:1.4571;
		specparam tpd_B_Y_r = 0.165495:0.302412:1.55179;
		specparam tpd_B_Y_f = 0.20448:0.342205:1.45106;
		specparam tpd_C_Y_r = 0.187428:0.328128:1.63905;
		specparam tpd_C_Y_f = 0.226379:0.360106:1.37172;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: CLKDLN 
`timescale 1ns/10ps
`celldefine
module CLKDLNX1 (ECK, E, SE, CKN);
	output ECK;
	input E, SE, CKN;
	reg notifier;
	wire delayed_E, delayed_SE, delayed_CKN;

	// Function
	wire int_fwire_clk, int_fwire_INTERNAL6, int_fwire_INTERNAL6__bar;
	wire int_fwire_test;

	buf (int_fwire_clk, delayed_CKN);
	or (int_fwire_test, delayed_E, delayed_SE);
	altos_latch (int_fwire_INTERNAL6, notifier, int_fwire_clk, int_fwire_test);
	not (int_fwire_INTERNAL6__bar, int_fwire_INTERNAL6);
	or (ECK, delayed_CKN, int_fwire_INTERNAL6__bar);

	// Timing
	specify
		specparam tpd_CKN_ECK_r = 0.28216:0.387556:1.32424;
		specparam tpd_CKN_ECK_f = 0.31173:0.464819:1.60573;
		specparam tsetup_E_CKN_NTB_SE_posedge_NTB_SE_negedge = 0.0893992:0.0376004:-0.506993;
		specparam thold_E_CKN_NTB_SE_posedge_NTB_SE_negedge = 0.0564178:0.0968976:0.590061;
		specparam tsetup_E_CKN_NTB_SE_negedge_NTB_SE_negedge = 0.0893992:0.0376004:-0.506993;
		specparam thold_E_CKN_NTB_SE_negedge_NTB_SE_negedge = 0.0564178:0.0968976:0.590061;
		specparam tsetup_SE_CKN_NTB_E_posedge_NTB_E_negedge = 0.0760352:0.0257694:-0.55584;
		specparam thold_SE_CKN_NTB_E_posedge_NTB_E_negedge = 0.0587:0.103636:0.630439;
		specparam tsetup_SE_CKN_NTB_E_negedge_NTB_E_negedge = 0.0760352:0.0257694:-0.55584;
		specparam thold_SE_CKN_NTB_E_negedge_NTB_E_negedge = 0.0587:0.103636:0.630439;
		specparam tpw_CKN_posedge = 0.29668:0.330811:2.72095;
		specparam tpw_CKN_negedge = 0.29668:0.330811:2.72095;

		(CKN => ECK) = ( tpd_CKN_ECK_r , tpd_CKN_ECK_f );
		$setuphold (negedge CKN &&& ~SE, posedge E &&& ~SE, 
			 tsetup_E_CKN_NTB_SE_posedge_NTB_SE_negedge, 
			 thold_E_CKN_NTB_SE_posedge_NTB_SE_negedge, notifier,,, delayed_CKN, delayed_E);
		$setuphold (negedge CKN &&& ~SE, negedge E &&& ~SE, 
			 tsetup_E_CKN_NTB_SE_negedge_NTB_SE_negedge, 
			 thold_E_CKN_NTB_SE_negedge_NTB_SE_negedge, notifier,,, delayed_CKN, delayed_E);
		$setuphold (negedge CKN &&& ~E, posedge SE &&& ~E, 
			 tsetup_SE_CKN_NTB_E_posedge_NTB_E_negedge, 
			 thold_SE_CKN_NTB_E_posedge_NTB_E_negedge, notifier,,, delayed_CKN, delayed_SE);
		$setuphold (negedge CKN &&& ~E, negedge SE &&& ~E, 
			 tsetup_SE_CKN_NTB_E_negedge_NTB_E_negedge, 
			 thold_SE_CKN_NTB_E_negedge_NTB_E_negedge, notifier,,, delayed_CKN, delayed_SE);
		$width (posedge CKN, tpw_CKN_posedge, 0, notifier);
		$width (negedge CKN, tpw_CKN_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: CLKDLN 
`timescale 1ns/10ps
`celldefine
module CLKDLNX2 (ECK, E, SE, CKN);
	output ECK;
	input E, SE, CKN;
	reg notifier;
	wire delayed_E, delayed_SE, delayed_CKN;

	// Function
	wire int_fwire_clk, int_fwire_INTERNAL6, int_fwire_INTERNAL6__bar;
	wire int_fwire_test;

	buf (int_fwire_clk, delayed_CKN);
	or (int_fwire_test, delayed_E, delayed_SE);
	altos_latch (int_fwire_INTERNAL6, notifier, int_fwire_clk, int_fwire_test);
	not (int_fwire_INTERNAL6__bar, int_fwire_INTERNAL6);
	or (ECK, delayed_CKN, int_fwire_INTERNAL6__bar);

	// Timing
	specify
		specparam tpd_CKN_ECK_r = 0.293711:0.402027:1.34036;
		specparam tpd_CKN_ECK_f = 0.339881:0.501295:1.6344;
		specparam tsetup_E_CKN_NTB_SE_posedge_NTB_SE_negedge = 0.0831675:0.0327551:-0.510394;
		specparam thold_E_CKN_NTB_SE_posedge_NTB_SE_negedge = 0.0546101:0.0947078:0.588252;
		specparam tsetup_E_CKN_NTB_SE_negedge_NTB_SE_negedge = 0.0831675:0.0327551:-0.510394;
		specparam thold_E_CKN_NTB_SE_negedge_NTB_SE_negedge = 0.0546101:0.0947078:0.588252;
		specparam tsetup_SE_CKN_NTB_E_posedge_NTB_E_negedge = 0.0745416:0.0202171:-0.556879;
		specparam thold_SE_CKN_NTB_E_posedge_NTB_E_negedge = 0.0587:0.103636:0.630439;
		specparam tsetup_SE_CKN_NTB_E_negedge_NTB_E_negedge = 0.0745416:0.0202171:-0.556879;
		specparam thold_SE_CKN_NTB_E_negedge_NTB_E_negedge = 0.0587:0.103636:0.630439;
		specparam tpw_CKN_posedge = 0.294079:0.330811:2.72095;
		specparam tpw_CKN_negedge = 0.294079:0.330811:2.72095;

		(CKN => ECK) = ( tpd_CKN_ECK_r , tpd_CKN_ECK_f );
		$setuphold (negedge CKN &&& ~SE, posedge E &&& ~SE, 
			 tsetup_E_CKN_NTB_SE_posedge_NTB_SE_negedge, 
			 thold_E_CKN_NTB_SE_posedge_NTB_SE_negedge, notifier,,, delayed_CKN, delayed_E);
		$setuphold (negedge CKN &&& ~SE, negedge E &&& ~SE, 
			 tsetup_E_CKN_NTB_SE_negedge_NTB_SE_negedge, 
			 thold_E_CKN_NTB_SE_negedge_NTB_SE_negedge, notifier,,, delayed_CKN, delayed_E);
		$setuphold (negedge CKN &&& ~E, posedge SE &&& ~E, 
			 tsetup_SE_CKN_NTB_E_posedge_NTB_E_negedge, 
			 thold_SE_CKN_NTB_E_posedge_NTB_E_negedge, notifier,,, delayed_CKN, delayed_SE);
		$setuphold (negedge CKN &&& ~E, negedge SE &&& ~E, 
			 tsetup_SE_CKN_NTB_E_negedge_NTB_E_negedge, 
			 thold_SE_CKN_NTB_E_negedge_NTB_E_negedge, notifier,,, delayed_CKN, delayed_SE);
		$width (posedge CKN, tpw_CKN_posedge, 0, notifier);
		$width (negedge CKN, tpw_CKN_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: CLKDLN 
`timescale 1ns/10ps
`celldefine
module CLKDLNX4 (ECK, E, SE, CKN);
	output ECK;
	input E, SE, CKN;
	reg notifier;
	wire delayed_E, delayed_SE, delayed_CKN;

	// Function
	wire int_fwire_clk, int_fwire_INTERNAL6, int_fwire_INTERNAL6__bar;
	wire int_fwire_test;

	buf (int_fwire_clk, delayed_CKN);
	or (int_fwire_test, delayed_E, delayed_SE);
	altos_latch (int_fwire_INTERNAL6, notifier, int_fwire_clk, int_fwire_test);
	not (int_fwire_INTERNAL6__bar, int_fwire_INTERNAL6);
	or (ECK, delayed_CKN, int_fwire_INTERNAL6__bar);

	// Timing
	specify
		specparam tpd_CKN_ECK_r = 0.322479:0.434033:1.3679;
		specparam tpd_CKN_ECK_f = 0.407895:0.578016:1.71128;
		specparam tsetup_E_CKN_NTB_SE_posedge_NTB_SE_negedge = 0.0734748:0.0230679:-0.517225;
		specparam thold_E_CKN_NTB_SE_posedge_NTB_SE_negedge = 0.0546101:0.0947078:0.588252;
		specparam tsetup_E_CKN_NTB_SE_negedge_NTB_SE_negedge = 0.0734748:0.0230679:-0.517225;
		specparam thold_E_CKN_NTB_SE_negedge_NTB_SE_negedge = 0.0546101:0.0947078:0.588252;
		specparam tsetup_SE_CKN_NTB_E_posedge_NTB_E_negedge = 0.0629735:0.01256:-0.563398;
		specparam thold_SE_CKN_NTB_E_posedge_NTB_E_negedge = 0.0587:0.103636:0.630439;
		specparam tsetup_SE_CKN_NTB_E_negedge_NTB_E_negedge = 0.0629735:0.01256:-0.563398;
		specparam thold_SE_CKN_NTB_E_negedge_NTB_E_negedge = 0.0587:0.103636:0.630439;
		specparam tpw_CKN_posedge = 0.28397:0.330811:2.72095;
		specparam tpw_CKN_negedge = 0.28397:0.330811:2.72095;

		(CKN => ECK) = ( tpd_CKN_ECK_r , tpd_CKN_ECK_f );
		$setuphold (negedge CKN &&& ~SE, posedge E &&& ~SE, 
			 tsetup_E_CKN_NTB_SE_posedge_NTB_SE_negedge, 
			 thold_E_CKN_NTB_SE_posedge_NTB_SE_negedge, notifier,,, delayed_CKN, delayed_E);
		$setuphold (negedge CKN &&& ~SE, negedge E &&& ~SE, 
			 tsetup_E_CKN_NTB_SE_negedge_NTB_SE_negedge, 
			 thold_E_CKN_NTB_SE_negedge_NTB_SE_negedge, notifier,,, delayed_CKN, delayed_E);
		$setuphold (negedge CKN &&& ~E, posedge SE &&& ~E, 
			 tsetup_SE_CKN_NTB_E_posedge_NTB_E_negedge, 
			 thold_SE_CKN_NTB_E_posedge_NTB_E_negedge, notifier,,, delayed_CKN, delayed_SE);
		$setuphold (negedge CKN &&& ~E, negedge SE &&& ~E, 
			 tsetup_SE_CKN_NTB_E_negedge_NTB_E_negedge, 
			 thold_SE_CKN_NTB_E_negedge_NTB_E_negedge, notifier,,, delayed_CKN, delayed_SE);
		$width (posedge CKN, tpw_CKN_posedge, 0, notifier);
		$width (negedge CKN, tpw_CKN_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: CLKDLN 
`timescale 1ns/10ps
`celldefine
module CLKDLNXL (ECK, E, SE, CKN);
	output ECK;
	input E, SE, CKN;
	reg notifier;
	wire delayed_E, delayed_SE, delayed_CKN;

	// Function
	wire int_fwire_clk, int_fwire_INTERNAL6, int_fwire_INTERNAL6__bar;
	wire int_fwire_test;

	buf (int_fwire_clk, delayed_CKN);
	or (int_fwire_test, delayed_E, delayed_SE);
	altos_latch (int_fwire_INTERNAL6, notifier, int_fwire_clk, int_fwire_test);
	not (int_fwire_INTERNAL6__bar, int_fwire_INTERNAL6);
	or (ECK, delayed_CKN, int_fwire_INTERNAL6__bar);

	// Timing
	specify
		specparam tpd_CKN_ECK_r = 0.28131:0.385827:1.32763;
		specparam tpd_CKN_ECK_f = 0.301605:0.449132:1.59287;
		specparam tsetup_E_CKN_NTB_SE_posedge_NTB_SE_negedge = 0.0900044:0.0397081:-0.505803;
		specparam thold_E_CKN_NTB_SE_posedge_NTB_SE_negedge = 0.0546101:0.0947078:0.588252;
		specparam tsetup_E_CKN_NTB_SE_negedge_NTB_SE_negedge = 0.0900044:0.0397081:-0.505803;
		specparam thold_E_CKN_NTB_SE_negedge_NTB_SE_negedge = 0.0546101:0.0947078:0.588252;
		specparam tsetup_SE_CKN_NTB_E_posedge_NTB_E_negedge = 0.0756151:0.0257694:-0.555578;
		specparam thold_SE_CKN_NTB_E_posedge_NTB_E_negedge = 0.0587:0.103636:0.630439;
		specparam tsetup_SE_CKN_NTB_E_negedge_NTB_E_negedge = 0.0756151:0.0257694:-0.555578;
		specparam thold_SE_CKN_NTB_E_negedge_NTB_E_negedge = 0.0587:0.103636:0.630439;
		specparam tpw_CKN_posedge = 0.296984:0.330811:2.72095;
		specparam tpw_CKN_negedge = 0.296984:0.330811:2.72095;

		(CKN => ECK) = ( tpd_CKN_ECK_r , tpd_CKN_ECK_f );
		$setuphold (negedge CKN &&& ~SE, posedge E &&& ~SE, 
			 tsetup_E_CKN_NTB_SE_posedge_NTB_SE_negedge, 
			 thold_E_CKN_NTB_SE_posedge_NTB_SE_negedge, notifier,,, delayed_CKN, delayed_E);
		$setuphold (negedge CKN &&& ~SE, negedge E &&& ~SE, 
			 tsetup_E_CKN_NTB_SE_negedge_NTB_SE_negedge, 
			 thold_E_CKN_NTB_SE_negedge_NTB_SE_negedge, notifier,,, delayed_CKN, delayed_E);
		$setuphold (negedge CKN &&& ~E, posedge SE &&& ~E, 
			 tsetup_SE_CKN_NTB_E_posedge_NTB_E_negedge, 
			 thold_SE_CKN_NTB_E_posedge_NTB_E_negedge, notifier,,, delayed_CKN, delayed_SE);
		$setuphold (negedge CKN &&& ~E, negedge SE &&& ~E, 
			 tsetup_SE_CKN_NTB_E_negedge_NTB_E_negedge, 
			 thold_SE_CKN_NTB_E_negedge_NTB_E_negedge, notifier,,, delayed_CKN, delayed_SE);
		$width (posedge CKN, tpw_CKN_posedge, 0, notifier);
		$width (negedge CKN, tpw_CKN_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: CLKDL 
`timescale 1ns/10ps
`celldefine
module CLKDLX1 (ECK, E, SE, CK);
	output ECK;
	input E, SE, CK;
	reg notifier;
	wire delayed_E, delayed_SE, delayed_CK;

	// Function
	wire int_fwire_clk, int_fwire_INTERNAL6, int_fwire_test;

	not (int_fwire_clk, delayed_CK);
	or (int_fwire_test, delayed_E, delayed_SE);
	altos_latch (int_fwire_INTERNAL6, notifier, int_fwire_clk, int_fwire_test);
	and (ECK, delayed_CK, int_fwire_INTERNAL6);

	// Timing
	specify
		specparam tpd_CK_ECK_r = 0.252335:0.382065:1.50617;
		specparam tpd_CK_ECK_f = 0.253227:0.387023:1.38244;
		specparam tsetup_E_CK_NTB_SE_posedge_NTB_SE_posedge = 0.129226:0.154501:0.32349;
		specparam thold_E_CK_NTB_SE_posedge_NTB_SE_posedge = -0.0961486:-0.127126:-0.290561;
		specparam tsetup_E_CK_NTB_SE_negedge_NTB_SE_posedge = 0.129226:0.154501:0.32349;
		specparam thold_E_CK_NTB_SE_negedge_NTB_SE_posedge = -0.0961486:-0.127126:-0.290561;
		specparam tsetup_SE_CK_NTB_E_posedge_NTB_E_posedge = 0.105482:0.128767:0.235965;
		specparam thold_SE_CK_NTB_E_posedge_NTB_E_posedge = -0.0812875:-0.107701:-0.198359;
		specparam tsetup_SE_CK_NTB_E_negedge_NTB_E_posedge = 0.105482:0.128767:0.235965;
		specparam thold_SE_CK_NTB_E_negedge_NTB_E_posedge = -0.0812875:-0.107701:-0.198359;
		specparam tpw_CK_posedge = 0.13546:0.330811:2.72095;
		specparam tpw_CK_negedge = 0.13546:0.330811:2.72095;

		(CK => ECK) = ( tpd_CK_ECK_r , tpd_CK_ECK_f );
		$setuphold (posedge CK &&& ~SE, posedge E &&& ~SE, 
			 tsetup_E_CK_NTB_SE_posedge_NTB_SE_posedge, 
			 thold_E_CK_NTB_SE_posedge_NTB_SE_posedge, notifier,,, delayed_CK, delayed_E);
		$setuphold (posedge CK &&& ~SE, negedge E &&& ~SE, 
			 tsetup_E_CK_NTB_SE_negedge_NTB_SE_posedge, 
			 thold_E_CK_NTB_SE_negedge_NTB_SE_posedge, notifier,,, delayed_CK, delayed_E);
		$setuphold (posedge CK &&& ~E, posedge SE &&& ~E, 
			 tsetup_SE_CK_NTB_E_posedge_NTB_E_posedge, 
			 thold_SE_CK_NTB_E_posedge_NTB_E_posedge, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK &&& ~E, negedge SE &&& ~E, 
			 tsetup_SE_CK_NTB_E_negedge_NTB_E_posedge, 
			 thold_SE_CK_NTB_E_negedge_NTB_E_posedge, notifier,,, delayed_CK, delayed_SE);
		$width (posedge CK, tpw_CK_posedge, 0, notifier);
		$width (negedge CK, tpw_CK_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: CLKDL 
`timescale 1ns/10ps
`celldefine
module CLKDLX2 (ECK, E, SE, CK);
	output ECK;
	input E, SE, CK;
	reg notifier;
	wire delayed_E, delayed_SE, delayed_CK;

	// Function
	wire int_fwire_clk, int_fwire_INTERNAL6, int_fwire_test;

	not (int_fwire_clk, delayed_CK);
	or (int_fwire_test, delayed_E, delayed_SE);
	altos_latch (int_fwire_INTERNAL6, notifier, int_fwire_clk, int_fwire_test);
	and (ECK, delayed_CK, int_fwire_INTERNAL6);

	// Timing
	specify
		specparam tpd_CK_ECK_r = 0.266746:0.399356:1.49899;
		specparam tpd_CK_ECK_f = 0.269307:0.407167:1.36266;
		specparam tsetup_E_CK_NTB_SE_posedge_NTB_SE_posedge = 0.129226:0.154501:0.324327;
		specparam thold_E_CK_NTB_SE_posedge_NTB_SE_posedge = -0.0961486:-0.127126:-0.286564;
		specparam tsetup_E_CK_NTB_SE_negedge_NTB_SE_posedge = 0.129226:0.154501:0.324327;
		specparam thold_E_CK_NTB_SE_negedge_NTB_SE_posedge = -0.0961486:-0.127126:-0.286564;
		specparam tsetup_SE_CK_NTB_E_posedge_NTB_E_posedge = 0.10664:0.126767:0.236036;
		specparam thold_SE_CK_NTB_E_posedge_NTB_E_posedge = -0.0790145:-0.103888:-0.195339;
		specparam tsetup_SE_CK_NTB_E_negedge_NTB_E_posedge = 0.10664:0.126767:0.236036;
		specparam thold_SE_CK_NTB_E_negedge_NTB_E_posedge = -0.0790145:-0.103888:-0.195339;
		specparam tpw_CK_posedge = 0.145683:0.330811:2.72095;
		specparam tpw_CK_negedge = 0.145683:0.330811:2.72095;

		(CK => ECK) = ( tpd_CK_ECK_r , tpd_CK_ECK_f );
		$setuphold (posedge CK &&& ~SE, posedge E &&& ~SE, 
			 tsetup_E_CK_NTB_SE_posedge_NTB_SE_posedge, 
			 thold_E_CK_NTB_SE_posedge_NTB_SE_posedge, notifier,,, delayed_CK, delayed_E);
		$setuphold (posedge CK &&& ~SE, negedge E &&& ~SE, 
			 tsetup_E_CK_NTB_SE_negedge_NTB_SE_posedge, 
			 thold_E_CK_NTB_SE_negedge_NTB_SE_posedge, notifier,,, delayed_CK, delayed_E);
		$setuphold (posedge CK &&& ~E, posedge SE &&& ~E, 
			 tsetup_SE_CK_NTB_E_posedge_NTB_E_posedge, 
			 thold_SE_CK_NTB_E_posedge_NTB_E_posedge, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK &&& ~E, negedge SE &&& ~E, 
			 tsetup_SE_CK_NTB_E_negedge_NTB_E_posedge, 
			 thold_SE_CK_NTB_E_negedge_NTB_E_posedge, notifier,,, delayed_CK, delayed_SE);
		$width (posedge CK, tpw_CK_posedge, 0, notifier);
		$width (negedge CK, tpw_CK_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: CLKDL 
`timescale 1ns/10ps
`celldefine
module CLKDLX4 (ECK, E, SE, CK);
	output ECK;
	input E, SE, CK;
	reg notifier;
	wire delayed_E, delayed_SE, delayed_CK;

	// Function
	wire int_fwire_clk, int_fwire_INTERNAL6, int_fwire_test;

	not (int_fwire_clk, delayed_CK);
	or (int_fwire_test, delayed_E, delayed_SE);
	altos_latch (int_fwire_INTERNAL6, notifier, int_fwire_clk, int_fwire_test);
	and (ECK, delayed_CK, int_fwire_INTERNAL6);

	// Timing
	specify
		specparam tpd_CK_ECK_r = 0.304171:0.443956:1.55683;
		specparam tpd_CK_ECK_f = 0.3098:0.455997:1.40075;
		specparam tsetup_E_CK_NTB_SE_posedge_NTB_SE_posedge = 0.129226:0.154501:0.322751;
		specparam thold_E_CK_NTB_SE_posedge_NTB_SE_posedge = -0.0962354:-0.131037:-0.290648;
		specparam tsetup_E_CK_NTB_SE_negedge_NTB_SE_posedge = 0.129226:0.154501:0.322751;
		specparam thold_E_CK_NTB_SE_negedge_NTB_SE_posedge = -0.0962354:-0.131037:-0.290648;
		specparam tsetup_SE_CK_NTB_E_posedge_NTB_E_posedge = 0.105402:0.128481:0.237598;
		specparam thold_SE_CK_NTB_E_posedge_NTB_E_posedge = -0.0814852:-0.105485:-0.196964;
		specparam tsetup_SE_CK_NTB_E_negedge_NTB_E_posedge = 0.105402:0.128481:0.237598;
		specparam thold_SE_CK_NTB_E_negedge_NTB_E_posedge = -0.0814852:-0.105485:-0.196964;
		specparam tpw_CK_posedge = 0.171413:0.330811:2.72095;
		specparam tpw_CK_negedge = 0.171413:0.330811:2.72095;

		(CK => ECK) = ( tpd_CK_ECK_r , tpd_CK_ECK_f );
		$setuphold (posedge CK &&& ~SE, posedge E &&& ~SE, 
			 tsetup_E_CK_NTB_SE_posedge_NTB_SE_posedge, 
			 thold_E_CK_NTB_SE_posedge_NTB_SE_posedge, notifier,,, delayed_CK, delayed_E);
		$setuphold (posedge CK &&& ~SE, negedge E &&& ~SE, 
			 tsetup_E_CK_NTB_SE_negedge_NTB_SE_posedge, 
			 thold_E_CK_NTB_SE_negedge_NTB_SE_posedge, notifier,,, delayed_CK, delayed_E);
		$setuphold (posedge CK &&& ~E, posedge SE &&& ~E, 
			 tsetup_SE_CK_NTB_E_posedge_NTB_E_posedge, 
			 thold_SE_CK_NTB_E_posedge_NTB_E_posedge, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK &&& ~E, negedge SE &&& ~E, 
			 tsetup_SE_CK_NTB_E_negedge_NTB_E_posedge, 
			 thold_SE_CK_NTB_E_negedge_NTB_E_posedge, notifier,,, delayed_CK, delayed_SE);
		$width (posedge CK, tpw_CK_posedge, 0, notifier);
		$width (negedge CK, tpw_CK_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: CLKDL 
`timescale 1ns/10ps
`celldefine
module CLKDLXL (ECK, E, SE, CK);
	output ECK;
	input E, SE, CK;
	reg notifier;
	wire delayed_E, delayed_SE, delayed_CK;

	// Function
	wire int_fwire_clk, int_fwire_INTERNAL6, int_fwire_test;

	not (int_fwire_clk, delayed_CK);
	or (int_fwire_test, delayed_E, delayed_SE);
	altos_latch (int_fwire_INTERNAL6, notifier, int_fwire_clk, int_fwire_test);
	and (ECK, delayed_CK, int_fwire_INTERNAL6);

	// Timing
	specify
		specparam tpd_CK_ECK_r = 0.253082:0.379253:1.48233;
		specparam tpd_CK_ECK_f = 0.248957:0.377365:1.35825;
		specparam tsetup_E_CK_NTB_SE_posedge_NTB_SE_posedge = 0.129226:0.154501:0.323687;
		specparam thold_E_CK_NTB_SE_posedge_NTB_SE_posedge = -0.0961486:-0.127126:-0.290561;
		specparam tsetup_E_CK_NTB_SE_negedge_NTB_SE_posedge = 0.129226:0.154501:0.323687;
		specparam thold_E_CK_NTB_SE_negedge_NTB_SE_posedge = -0.0961486:-0.127126:-0.290561;
		specparam tsetup_SE_CK_NTB_E_posedge_NTB_E_posedge = 0.107054:0.128767:0.235965;
		specparam thold_SE_CK_NTB_E_posedge_NTB_E_posedge = -0.0799933:-0.105485:-0.196964;
		specparam tsetup_SE_CK_NTB_E_negedge_NTB_E_posedge = 0.107054:0.128767:0.235965;
		specparam thold_SE_CK_NTB_E_negedge_NTB_E_posedge = -0.0799933:-0.105485:-0.196964;
		specparam tpw_CK_posedge = 0.132486:0.330811:2.72095;
		specparam tpw_CK_negedge = 0.132486:0.330811:2.72095;

		(CK => ECK) = ( tpd_CK_ECK_r , tpd_CK_ECK_f );
		$setuphold (posedge CK &&& ~SE, posedge E &&& ~SE, 
			 tsetup_E_CK_NTB_SE_posedge_NTB_SE_posedge, 
			 thold_E_CK_NTB_SE_posedge_NTB_SE_posedge, notifier,,, delayed_CK, delayed_E);
		$setuphold (posedge CK &&& ~SE, negedge E &&& ~SE, 
			 tsetup_E_CK_NTB_SE_negedge_NTB_SE_posedge, 
			 thold_E_CK_NTB_SE_negedge_NTB_SE_posedge, notifier,,, delayed_CK, delayed_E);
		$setuphold (posedge CK &&& ~E, posedge SE &&& ~E, 
			 tsetup_SE_CK_NTB_E_posedge_NTB_E_posedge, 
			 thold_SE_CK_NTB_E_posedge_NTB_E_posedge, notifier,,, delayed_CK, delayed_SE);
		$setuphold (posedge CK &&& ~E, negedge SE &&& ~E, 
			 tsetup_SE_CK_NTB_E_negedge_NTB_E_posedge, 
			 thold_SE_CK_NTB_E_negedge_NTB_E_posedge, notifier,,, delayed_CK, delayed_SE);
		$width (posedge CK, tpw_CK_posedge, 0, notifier);
		$width (negedge CK, tpw_CK_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNQ 
`timescale 1ns/10ps
`celldefine
module DFFNQX1 (Q, D, XC);
	output Q;
	input D, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, xcr_0;

	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, delayed_D);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XC_Q_negedge_r = 0.361954:0.525104:1.96469;
		specparam tpd_XC_Q_negedge_f = 0.329871:0.487575:1.64448;
		specparam tsetup_D_XC_posedge_negedge = 0.0897988:0.0457279:-0.314214;
		specparam thold_D_XC_posedge_negedge = 0.0606207:0.105071:0.519914;
		specparam tsetup_D_XC_negedge_negedge = 0.0897988:0.0457279:-0.314214;
		specparam thold_D_XC_negedge_negedge = 0.0606207:0.105071:0.519914;
		specparam tpw_XC_posedge = 0.275026:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.275026:0.330811:2.72095;

		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC, posedge D, 
			 tsetup_D_XC_posedge_negedge, 
			 thold_D_XC_posedge_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC, negedge D, 
			 tsetup_D_XC_negedge_negedge, 
			 thold_D_XC_negedge_negedge, notifier,,, delayed_XC, delayed_D);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNQ 
`timescale 1ns/10ps
`celldefine
module DFFNQX2 (Q, D, XC);
	output Q;
	input D, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, xcr_0;

	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, delayed_D);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XC_Q_negedge_r = 0.35664:0.521862:1.94079;
		specparam tpd_XC_Q_negedge_f = 0.322517:0.481937:1.62697;
		specparam tsetup_D_XC_posedge_negedge = 0.048816:0.00807721:-0.334243;
		specparam thold_D_XC_posedge_negedge = 0.061882:0.111727:0.5127;
		specparam tsetup_D_XC_negedge_negedge = 0.048816:0.00807721:-0.334243;
		specparam thold_D_XC_negedge_negedge = 0.061882:0.111727:0.5127;
		specparam tpw_XC_posedge = 0.23878:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.23878:0.330811:2.72095;

		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC, posedge D, 
			 tsetup_D_XC_posedge_negedge, 
			 thold_D_XC_posedge_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC, negedge D, 
			 tsetup_D_XC_negedge_negedge, 
			 thold_D_XC_negedge_negedge, notifier,,, delayed_XC, delayed_D);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNQ 
`timescale 1ns/10ps
`celldefine
module DFFNQX4 (Q, D, XC);
	output Q;
	input D, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, xcr_0;

	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, delayed_D);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XC_Q_negedge_r = 0.40881:0.573786:2.0077;
		specparam tpd_XC_Q_negedge_f = 0.350906:0.491089:1.36926;
		specparam tsetup_D_XC_posedge_negedge = 0.0344184:-0.0118349:-0.36479;
		specparam thold_D_XC_posedge_negedge = 0.0715268:0.126002:0.541069;
		specparam tsetup_D_XC_negedge_negedge = 0.0344184:-0.0118349:-0.36479;
		specparam thold_D_XC_negedge_negedge = 0.0715268:0.126002:0.541069;
		specparam tpw_XC_posedge = 0.212948:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.212948:0.330811:2.72095;

		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC, posedge D, 
			 tsetup_D_XC_posedge_negedge, 
			 thold_D_XC_posedge_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC, negedge D, 
			 tsetup_D_XC_negedge_negedge, 
			 thold_D_XC_negedge_negedge, notifier,,, delayed_XC, delayed_D);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNQ 
`timescale 1ns/10ps
`celldefine
module DFFNQXL (Q, D, XC);
	output Q;
	input D, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, xcr_0;

	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, delayed_D);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XC_Q_negedge_r = 0.393793:0.5593:2.05776;
		specparam tpd_XC_Q_negedge_f = 0.357512:0.521912:1.84185;
		specparam tsetup_D_XC_posedge_negedge = 0.0596308:0.00962617:-0.408687;
		specparam thold_D_XC_posedge_negedge = 0.0876961:0.14193:0.620217;
		specparam tsetup_D_XC_negedge_negedge = 0.0596308:0.00962617:-0.408687;
		specparam thold_D_XC_negedge_negedge = 0.0876961:0.14193:0.620217;
		specparam tpw_XC_posedge = 0.275026:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.275026:0.330811:2.72095;

		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC, posedge D, 
			 tsetup_D_XC_posedge_negedge, 
			 thold_D_XC_posedge_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC, negedge D, 
			 tsetup_D_XC_negedge_negedge, 
			 thold_D_XC_negedge_negedge, notifier,,, delayed_XC, delayed_D);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNQX 
`timescale 1ns/10ps
`celldefine
module DFFNQXX1 (Q, XQ, D, XC);
	output Q, XQ;
	input D, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, delayed_D);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XC_Q_negedge_r = 0.361689:0.522735:1.94329;
		specparam tpd_XC_Q_negedge_f = 0.326723:0.483623:1.61128;
		specparam tpd_XC_XQ_negedge_r = 0.404124:0.555437:1.97723;
		specparam tpd_XC_XQ_negedge_f = 0.471602:0.619308:1.75278;
		specparam tsetup_D_XC_posedge_negedge = 0.0913555:0.0453576:-0.307883;
		specparam thold_D_XC_posedge_negedge = 0.0605643:0.11:0.525024;
		specparam tsetup_D_XC_negedge_negedge = 0.0913555:0.0453576:-0.307883;
		specparam thold_D_XC_negedge_negedge = 0.0605643:0.11:0.525024;
		specparam tpw_XC_posedge = 0.269808:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.269808:0.330811:2.72095;

		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC, posedge D, 
			 tsetup_D_XC_posedge_negedge, 
			 thold_D_XC_posedge_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC, negedge D, 
			 tsetup_D_XC_negedge_negedge, 
			 thold_D_XC_negedge_negedge, notifier,,, delayed_XC, delayed_D);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNQX 
`timescale 1ns/10ps
`celldefine
module DFFNQXX2 (Q, XQ, D, XC);
	output Q, XQ;
	input D, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, delayed_D);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XC_Q_negedge_r = 0.35414:0.515364:1.90806;
		specparam tpd_XC_Q_negedge_f = 0.314858:0.467257:1.51803;
		specparam tpd_XC_XQ_negedge_r = 0.40389:0.552692:1.93476;
		specparam tpd_XC_XQ_negedge_f = 0.4612:0.601995:1.64715;
		specparam tsetup_D_XC_posedge_negedge = 0.0545913:0.0105639:-0.3139;
		specparam thold_D_XC_posedge_negedge = 0.0620273:0.109174:0.499564;
		specparam tsetup_D_XC_negedge_negedge = 0.0545913:0.0105639:-0.3139;
		specparam thold_D_XC_negedge_negedge = 0.0620273:0.109174:0.499564;
		specparam tpw_XC_posedge = 0.236454:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.236454:0.330811:2.72095;

		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC, posedge D, 
			 tsetup_D_XC_posedge_negedge, 
			 thold_D_XC_posedge_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC, negedge D, 
			 tsetup_D_XC_negedge_negedge, 
			 thold_D_XC_negedge_negedge, notifier,,, delayed_XC, delayed_D);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNQX 
`timescale 1ns/10ps
`celldefine
module DFFNQXX4 (Q, XQ, D, XC);
	output Q, XQ;
	input D, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, delayed_D);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XC_Q_negedge_r = 0.408319:0.570713:1.96684;
		specparam tpd_XC_Q_negedge_f = 0.34366:0.482727:1.34113;
		specparam tpd_XC_XQ_negedge_r = 0.441524:0.587562:1.98234;
		specparam tpd_XC_XQ_negedge_f = 0.499628:0.622012:1.4712;
		specparam tsetup_D_XC_posedge_negedge = 0.0381904:-0.001:-0.331206;
		specparam thold_D_XC_posedge_negedge = 0.0695783:0.119171:0.514237;
		specparam tsetup_D_XC_negedge_negedge = 0.0381904:-0.001:-0.331206;
		specparam thold_D_XC_negedge_negedge = 0.0695783:0.119171:0.514237;
		specparam tpw_XC_posedge = 0.212948:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.212948:0.330811:2.72095;

		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC, posedge D, 
			 tsetup_D_XC_posedge_negedge, 
			 thold_D_XC_posedge_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC, negedge D, 
			 tsetup_D_XC_negedge_negedge, 
			 thold_D_XC_negedge_negedge, notifier,,, delayed_XC, delayed_D);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNQX 
`timescale 1ns/10ps
`celldefine
module DFFNQXXL (Q, XQ, D, XC);
	output Q, XQ;
	input D, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, delayed_D);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XC_Q_negedge_r = 0.397053:0.55979:2.02483;
		specparam tpd_XC_Q_negedge_f = 0.352674:0.504464:1.60978;
		specparam tpd_XC_XQ_negedge_r = 0.427539:0.581011:2.049;
		specparam tpd_XC_XQ_negedge_f = 0.494965:0.639547:1.76122;
		specparam tsetup_D_XC_posedge_negedge = 0.0618491:0.0128323:-0.391495;
		specparam thold_D_XC_posedge_negedge = 0.0832981:0.137091:0.60438;
		specparam tsetup_D_XC_negedge_negedge = 0.0618491:0.0128323:-0.391495;
		specparam thold_D_XC_negedge_negedge = 0.0832981:0.137091:0.60438;
		specparam tpw_XC_posedge = 0.272717:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.272717:0.330811:2.72095;

		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC, posedge D, 
			 tsetup_D_XC_posedge_negedge, 
			 thold_D_XC_posedge_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC, negedge D, 
			 tsetup_D_XC_negedge_negedge, 
			 thold_D_XC_negedge_negedge, notifier,,, delayed_XC, delayed_D);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNRQ 
`timescale 1ns/10ps
`celldefine
module DFFNRQX1 (Q, D, XR, XC);
	output Q;
	input D, XR, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.119116:0.259614:1.23346;
		specparam tpd_XR_Q_negedge_f = 0.119116:0.259614:1.23346;
		specparam tpd_XC_Q_negedge_r = 0.411103:0.580177:2.03325;
		specparam tpd_XC_Q_negedge_f = 0.325031:0.465557:1.42986;
		specparam tsetup_D_XC_XR_posedge_XR_negedge = 0.048994:-0.000901656:-0.390933;
		specparam thold_D_XC_XR_posedge_XR_negedge = 0.0798552:0.133048:0.580951;
		specparam tsetup_D_XC_XR_negedge_XR_negedge = 0.048994:-0.000901656:-0.390933;
		specparam thold_D_XC_XR_negedge_XR_negedge = 0.0798552:0.133048:0.580951;
		specparam trecovery_XR_XC_D_posedge_D_negedge = -0.280772:-0.34714:-0.514649;
		specparam tremoval_XR_XC_D_posedge_D_negedge = 0.363912:0.482092:1.18277;
		specparam tpw_XR_negedge = 0.299603:0.393753:2.72095;
		specparam tpw_XC_posedge = 0.301119:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.301119:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& XR, posedge D &&& XR, 
			 tsetup_D_XC_XR_posedge_XR_negedge, 
			 thold_D_XC_XR_posedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XR, negedge D &&& XR, 
			 tsetup_D_XC_XR_negedge_XR_negedge, 
			 thold_D_XC_XR_negedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XR &&& D, negedge XC &&& D, 
			 trecovery_XR_XC_D_posedge_D_negedge, notifier);
		$hold (negedge XC &&& D, posedge XR &&& D, 
			 tremoval_XR_XC_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNRQ 
`timescale 1ns/10ps
`celldefine
module DFFNRQX2 (Q, D, XR, XC);
	output Q;
	input D, XR, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.135635:0.282112:1.23015;
		specparam tpd_XR_Q_negedge_f = 0.135635:0.282112:1.23015;
		specparam tpd_XC_Q_negedge_r = 0.406195:0.578323:1.99066;
		specparam tpd_XC_Q_negedge_f = 0.319575:0.461222:1.31664;
		specparam tsetup_D_XC_XR_posedge_XR_negedge = 0.0571988:0.015:-0.316325;
		specparam thold_D_XC_XR_posedge_XR_negedge = 0.0639626:0.111421:0.506869;
		specparam tsetup_D_XC_XR_negedge_XR_negedge = 0.0571988:0.015:-0.316325;
		specparam thold_D_XC_XR_negedge_XR_negedge = 0.0639626:0.111421:0.506869;
		specparam trecovery_XR_XC_D_posedge_D_negedge = -0.248618:-0.310484:-0.333944;
		specparam tremoval_XR_XC_D_posedge_D_negedge = 0.341391:0.453372:1.10718;
		specparam tpw_XR_negedge = 0.304423:0.398998:2.72095;
		specparam tpw_XC_posedge = 0.249513:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.249513:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& XR, posedge D &&& XR, 
			 tsetup_D_XC_XR_posedge_XR_negedge, 
			 thold_D_XC_XR_posedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XR, negedge D &&& XR, 
			 tsetup_D_XC_XR_negedge_XR_negedge, 
			 thold_D_XC_XR_negedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XR &&& D, negedge XC &&& D, 
			 trecovery_XR_XC_D_posedge_D_negedge, notifier);
		$hold (negedge XC &&& D, posedge XR &&& D, 
			 tremoval_XR_XC_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNRQ 
`timescale 1ns/10ps
`celldefine
module DFFNRQX4 (Q, D, XR, XC);
	output Q;
	input D, XR, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.135714:0.28473:1.26379;
		specparam tpd_XR_Q_negedge_f = 0.135714:0.28473:1.26379;
		specparam tpd_XC_Q_negedge_r = 0.458925:0.633421:2.05363;
		specparam tpd_XC_Q_negedge_f = 0.36281:0.507681:1.39791;
		specparam tsetup_D_XC_XR_posedge_XR_negedge = 0.0468435:0.004:-0.332858;
		specparam thold_D_XC_XR_posedge_XR_negedge = 0.069446:0.120584:0.51357;
		specparam tsetup_D_XC_XR_negedge_XR_negedge = 0.0468435:0.004:-0.332858;
		specparam thold_D_XC_XR_negedge_XR_negedge = 0.069446:0.120584:0.51357;
		specparam trecovery_XR_XC_D_posedge_D_negedge = -0.264293:-0.345281:-0.436509;
		specparam tremoval_XR_XC_D_posedge_D_negedge = 0.332275:0.448551:1.10018;
		specparam tpw_XR_negedge = 0.319351:0.412111:2.72095;
		specparam tpw_XC_posedge = 0.223395:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.223395:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& XR, posedge D &&& XR, 
			 tsetup_D_XC_XR_posedge_XR_negedge, 
			 thold_D_XC_XR_posedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XR, negedge D &&& XR, 
			 tsetup_D_XC_XR_negedge_XR_negedge, 
			 thold_D_XC_XR_negedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XR &&& D, negedge XC &&& D, 
			 trecovery_XR_XC_D_posedge_D_negedge, notifier);
		$hold (negedge XC &&& D, posedge XR &&& D, 
			 tremoval_XR_XC_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNRQ 
`timescale 1ns/10ps
`celldefine
module DFFNRQXL (Q, D, XR, XC);
	output Q;
	input D, XR, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.11628:0.25537:1.29239;
		specparam tpd_XR_Q_negedge_f = 0.11628:0.25537:1.29239;
		specparam tpd_XC_Q_negedge_r = 0.405471:0.571559:2.02993;
		specparam tpd_XC_Q_negedge_f = 0.32131:0.462157:1.50692;
		specparam tsetup_D_XC_XR_posedge_XR_negedge = 0.0481601:-0.000897984:-0.390572;
		specparam thold_D_XC_XR_posedge_XR_negedge = 0.0792763:0.131028:0.583632;
		specparam tsetup_D_XC_XR_negedge_XR_negedge = 0.0481601:-0.000897984:-0.390572;
		specparam thold_D_XC_XR_negedge_XR_negedge = 0.0792763:0.131028:0.583632;
		specparam trecovery_XR_XC_D_posedge_D_negedge = -0.28196:-0.343356:-0.532708;
		specparam tremoval_XR_XC_D_posedge_D_negedge = 0.363912:0.482092:1.18277;
		specparam tpw_XR_negedge = 0.299603:0.393753:2.72095;
		specparam tpw_XC_posedge = 0.301119:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.301119:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& XR, posedge D &&& XR, 
			 tsetup_D_XC_XR_posedge_XR_negedge, 
			 thold_D_XC_XR_posedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XR, negedge D &&& XR, 
			 tsetup_D_XC_XR_negedge_XR_negedge, 
			 thold_D_XC_XR_negedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XR &&& D, negedge XC &&& D, 
			 trecovery_XR_XC_D_posedge_D_negedge, notifier);
		$hold (negedge XC &&& D, posedge XR &&& D, 
			 tremoval_XR_XC_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNRQX 
`timescale 1ns/10ps
`celldefine
module DFFNRQXX1 (Q, XQ, D, XR, XC);
	output Q, XQ;
	input D, XR, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.116923:0.254417:1.20241;
		specparam tpd_XR_Q_negedge_f = 0.116923:0.254417:1.20241;
		specparam tpd_XC_Q_negedge_r = 0.374674:0.537119:1.94963;
		specparam tpd_XC_Q_negedge_f = 0.29003:0.424492:1.31526;
		specparam tpd_XR_XQ_negedge_r = 0.231137:0.39785:1.83629;
		specparam tpd_XR_XQ_negedge_f = 0.231137:0.39785:1.83629;
		specparam tpd_XC_XQ_negedge_r = 0.377994:0.528645:1.93413;
		specparam tpd_XC_XQ_negedge_f = 0.461013:0.590008:1.47556;
		specparam tsetup_D_XC_XR_posedge_XR_negedge = 0.0717744:0.029:-0.313265;
		specparam thold_D_XC_XR_posedge_XR_negedge = 0.0564074:0.102923:0.506274;
		specparam tsetup_D_XC_XR_negedge_XR_negedge = 0.0717744:0.029:-0.313265;
		specparam thold_D_XC_XR_negedge_XR_negedge = 0.0564074:0.102923:0.506274;
		specparam trecovery_XR_XC_D_posedge_D_negedge = -0.247264:-0.302884:-0.406232;
		specparam tremoval_XR_XC_D_posedge_D_negedge = 0.344531:0.455729:1.1122;
		specparam tpw_XR_negedge = 0.297904:0.39113:2.72095;
		specparam tpw_XC_posedge = 0.296211:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.296211:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& XR, posedge D &&& XR, 
			 tsetup_D_XC_XR_posedge_XR_negedge, 
			 thold_D_XC_XR_posedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XR, negedge D &&& XR, 
			 tsetup_D_XC_XR_negedge_XR_negedge, 
			 thold_D_XC_XR_negedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XR &&& D, negedge XC &&& D, 
			 trecovery_XR_XC_D_posedge_D_negedge, notifier);
		$hold (negedge XC &&& D, posedge XR &&& D, 
			 tremoval_XR_XC_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNRQX 
`timescale 1ns/10ps
`celldefine
module DFFNRQXX2 (Q, XQ, D, XR, XC);
	output Q, XQ;
	input D, XR, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.136191:0.283312:1.25644;
		specparam tpd_XR_Q_negedge_f = 0.136191:0.283312:1.25644;
		specparam tpd_XC_Q_negedge_r = 0.391009:0.560505:1.98077;
		specparam tpd_XC_Q_negedge_f = 0.308919:0.450328:1.33357;
		specparam tpd_XR_XQ_negedge_r = 0.284668:0.456369:1.94332;
		specparam tpd_XR_XQ_negedge_f = 0.284668:0.456369:1.94332;
		specparam tpd_XC_XQ_negedge_r = 0.429335:0.582586:1.99792;
		specparam tpd_XC_XQ_negedge_f = 0.51835:0.651582:1.55369;
		specparam tsetup_D_XC_XR_posedge_XR_negedge = 0.0626671:0.02:-0.314417;
		specparam thold_D_XC_XR_posedge_XR_negedge = 0.0568065:0.10399:0.497005;
		specparam tsetup_D_XC_XR_negedge_XR_negedge = 0.0626671:0.02:-0.314417;
		specparam thold_D_XC_XR_negedge_XR_negedge = 0.0568065:0.10399:0.497005;
		specparam trecovery_XR_XC_D_posedge_D_negedge = -0.239312:-0.29928:-0.332429;
		specparam tremoval_XR_XC_D_posedge_D_negedge = 0.337069:0.447981:1.10632;
		specparam tpw_XR_negedge = 0.303215:0.398998:2.72095;
		specparam tpw_XC_posedge = 0.238781:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.238781:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& XR, posedge D &&& XR, 
			 tsetup_D_XC_XR_posedge_XR_negedge, 
			 thold_D_XC_XR_posedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XR, negedge D &&& XR, 
			 tsetup_D_XC_XR_negedge_XR_negedge, 
			 thold_D_XC_XR_negedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XR &&& D, negedge XC &&& D, 
			 trecovery_XR_XC_D_posedge_D_negedge, notifier);
		$hold (negedge XC &&& D, posedge XR &&& D, 
			 tremoval_XR_XC_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNRQX 
`timescale 1ns/10ps
`celldefine
module DFFNRQXX4 (Q, XQ, D, XR, XC);
	output Q, XQ;
	input D, XR, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.135059:0.28228:1.25586;
		specparam tpd_XR_Q_negedge_f = 0.135059:0.28228:1.25586;
		specparam tpd_XC_Q_negedge_r = 0.461629:0.632571:2.04951;
		specparam tpd_XC_Q_negedge_f = 0.365774:0.508469:1.39986;
		specparam tpd_XR_XQ_negedge_r = 0.257782:0.420478:1.89871;
		specparam tpd_XR_XQ_negedge_f = 0.257782:0.420478:1.89871;
		specparam tpd_XC_XQ_negedge_r = 0.471375:0.619632:2.03989;
		specparam tpd_XC_XQ_negedge_f = 0.574504:0.698681:1.57528;
		specparam tsetup_D_XC_XR_posedge_XR_negedge = 0.0526127:0.0100777:-0.329428;
		specparam thold_D_XC_XR_posedge_XR_negedge = 0.0661056:0.114017:0.504253;
		specparam tsetup_D_XC_XR_negedge_XR_negedge = 0.0526127:0.0100777:-0.329428;
		specparam thold_D_XC_XR_negedge_XR_negedge = 0.0661056:0.114017:0.504253;
		specparam trecovery_XR_XC_D_posedge_D_negedge = -0.2577:-0.341884:-0.444391;
		specparam tremoval_XR_XC_D_posedge_D_negedge = 0.325073:0.438791:1.09877;
		specparam tpw_XR_negedge = 0.320483:0.412111:2.72095;
		specparam tpw_XC_posedge = 0.212948:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.212948:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& XR, posedge D &&& XR, 
			 tsetup_D_XC_XR_posedge_XR_negedge, 
			 thold_D_XC_XR_posedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XR, negedge D &&& XR, 
			 tsetup_D_XC_XR_negedge_XR_negedge, 
			 thold_D_XC_XR_negedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XR &&& D, negedge XC &&& D, 
			 trecovery_XR_XC_D_posedge_D_negedge, notifier);
		$hold (negedge XC &&& D, posedge XR &&& D, 
			 tremoval_XR_XC_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNRQX 
`timescale 1ns/10ps
`celldefine
module DFFNRQXXL (Q, XQ, D, XR, XC);
	output Q, XQ;
	input D, XR, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.115505:0.257292:1.31411;
		specparam tpd_XR_Q_negedge_f = 0.115505:0.257292:1.31411;
		specparam tpd_XC_Q_negedge_r = 0.395058:0.560291:2.01159;
		specparam tpd_XC_Q_negedge_f = 0.31719:0.460266:1.5193;
		specparam tpd_XR_XQ_negedge_r = 0.214605:0.381805:1.82308;
		specparam tpd_XR_XQ_negedge_f = 0.214605:0.381805:1.82308;
		specparam tpd_XC_XQ_negedge_r = 0.390927:0.545998:2.01238;
		specparam tpd_XC_XQ_negedge_f = 0.474374:0.61501:1.67623;
		specparam tsetup_D_XC_XR_posedge_XR_negedge = 0.0482801:-0.00161798:-0.393715;
		specparam thold_D_XC_XR_posedge_XR_negedge = 0.0783702:0.13195:0.585736;
		specparam tsetup_D_XC_XR_negedge_XR_negedge = 0.0482801:-0.00161798:-0.393715;
		specparam thold_D_XC_XR_negedge_XR_negedge = 0.0783702:0.13195:0.585736;
		specparam trecovery_XR_XC_D_posedge_D_negedge = -0.27714:-0.340126:-0.531822;
		specparam tremoval_XR_XC_D_posedge_D_negedge = 0.366186:0.485391:1.18391;
		specparam tpw_XR_negedge = 0.297904:0.39113:2.72095;
		specparam tpw_XC_posedge = 0.298509:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.298509:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& XR, posedge D &&& XR, 
			 tsetup_D_XC_XR_posedge_XR_negedge, 
			 thold_D_XC_XR_posedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XR, negedge D &&& XR, 
			 tsetup_D_XC_XR_negedge_XR_negedge, 
			 thold_D_XC_XR_negedge_XR_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XR &&& D, negedge XC &&& D, 
			 trecovery_XR_XC_D_posedge_D_negedge, notifier);
		$hold (negedge XC &&& D, posedge XR &&& D, 
			 tremoval_XR_XC_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSQ 
`timescale 1ns/10ps
`celldefine
module DFFNSQX1 (Q, D, XS, XC);
	output Q;
	input D, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_s;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.305805:0.466083:1.93578;
		specparam tpd_XS_Q_negedge_f = 0.305805:0.466083:1.93578;
		specparam tpd_XC_Q_negedge_r = 0.370201:0.533516:2.00539;
		specparam tpd_XC_Q_negedge_f = 0.330754:0.469762:1.4123;
		specparam tsetup_D_XC_XS_posedge_XS_negedge = 0.0467337:-0.00358131:-0.38468;
		specparam thold_D_XC_XS_posedge_XS_negedge = 0.06951:0.119035:0.555611;
		specparam tsetup_D_XC_XS_negedge_XS_negedge = 0.0467337:-0.00358131:-0.38468;
		specparam thold_D_XC_XS_negedge_XS_negedge = 0.06951:0.119035:0.555611;
		specparam trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge = -0.00311354:-0.0504841:-0.258485;
		specparam tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0778331:0.129147:0.450172;
		specparam tpw_XS_negedge = 0.180304:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.324279:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.324279:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& XS, posedge D &&& XS, 
			 tsetup_D_XC_XS_posedge_XS_negedge, 
			 thold_D_XC_XS_posedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XS, negedge D &&& XS, 
			 tsetup_D_XC_XS_negedge_XS_negedge, 
			 thold_D_XC_XS_negedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XS &&& ~D, negedge XC &&& ~D, 
			 trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge XC &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSQ 
`timescale 1ns/10ps
`celldefine
module DFFNSQX2 (Q, D, XS, XC);
	output Q;
	input D, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_s;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.324878:0.489849:1.95836;
		specparam tpd_XS_Q_negedge_f = 0.324878:0.489849:1.95836;
		specparam tpd_XC_Q_negedge_r = 0.358351:0.522918:1.94381;
		specparam tpd_XC_Q_negedge_f = 0.330707:0.474285:1.36155;
		specparam tsetup_D_XC_XS_posedge_XS_negedge = 0.0546817:0.0103515:-0.316687;
		specparam thold_D_XC_XS_posedge_XS_negedge = 0.0554475:0.100307:0.482781;
		specparam tsetup_D_XC_XS_negedge_XS_negedge = 0.0546817:0.0103515:-0.316687;
		specparam thold_D_XC_XS_negedge_XS_negedge = 0.0554475:0.100307:0.482781;
		specparam trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0123409:-0.0335759:-0.17484;
		specparam tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0625424:0.107112:0.385752;
		specparam tpw_XS_negedge = 0.188262:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.27212:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.27212:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& XS, posedge D &&& XS, 
			 tsetup_D_XC_XS_posedge_XS_negedge, 
			 thold_D_XC_XS_posedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XS, negedge D &&& XS, 
			 tsetup_D_XC_XS_negedge_XS_negedge, 
			 thold_D_XC_XS_negedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XS &&& ~D, negedge XC &&& ~D, 
			 trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge XC &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSQ 
`timescale 1ns/10ps
`celldefine
module DFFNSQX4 (Q, D, XS, XC);
	output Q;
	input D, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_s;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.352596:0.518103:2.00268;
		specparam tpd_XS_Q_negedge_f = 0.352596:0.518103:2.00268;
		specparam tpd_XC_Q_negedge_r = 0.388457:0.554731:1.98183;
		specparam tpd_XC_Q_negedge_f = 0.36204:0.508575:1.43854;
		specparam tsetup_D_XC_XS_posedge_XS_negedge = 0.0402943:-0.005:-0.334634;
		specparam thold_D_XC_XS_posedge_XS_negedge = 0.0632114:0.112317:0.494925;
		specparam tsetup_D_XC_XS_negedge_XS_negedge = 0.0402943:-0.005:-0.334634;
		specparam thold_D_XC_XS_negedge_XS_negedge = 0.0632114:0.112317:0.494925;
		specparam trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.00013008:-0.0394561:-0.18689;
		specparam tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0629623:0.110385:0.388329;
		specparam tpw_XS_negedge = 0.203815:0.349169:2.72095;
		specparam tpw_XC_posedge = 0.243715:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.243715:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& XS, posedge D &&& XS, 
			 tsetup_D_XC_XS_posedge_XS_negedge, 
			 thold_D_XC_XS_posedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XS, negedge D &&& XS, 
			 tsetup_D_XC_XS_negedge_XS_negedge, 
			 thold_D_XC_XS_negedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XS &&& ~D, negedge XC &&& ~D, 
			 trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge XC &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSQ 
`timescale 1ns/10ps
`celldefine
module DFFNSQXL (Q, D, XS, XC);
	output Q;
	input D, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_s;
	wire xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.299127:0.45701:1.92741;
		specparam tpd_XS_Q_negedge_f = 0.299127:0.45701:1.92741;
		specparam tpd_XC_Q_negedge_r = 0.365478:0.526738:2.00138;
		specparam tpd_XC_Q_negedge_f = 0.328054:0.469889:1.53701;
		specparam tsetup_D_XC_XS_posedge_XS_negedge = 0.0453076:-0.00424123:-0.385072;
		specparam thold_D_XC_XS_posedge_XS_negedge = 0.070214:0.12:0.55073;
		specparam tsetup_D_XC_XS_negedge_XS_negedge = 0.0453076:-0.00424123:-0.385072;
		specparam thold_D_XC_XS_negedge_XS_negedge = 0.070214:0.12:0.55073;
		specparam trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge = -0.00561974:-0.0510399:-0.264186;
		specparam tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.078318:0.129147:0.455949;
		specparam tpw_XS_negedge = 0.176886:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.323956:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.323956:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& XS, posedge D &&& XS, 
			 tsetup_D_XC_XS_posedge_XS_negedge, 
			 thold_D_XC_XS_posedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XS, negedge D &&& XS, 
			 tsetup_D_XC_XS_negedge_XS_negedge, 
			 thold_D_XC_XS_negedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XS &&& ~D, negedge XC &&& ~D, 
			 trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge XC &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSQX 
`timescale 1ns/10ps
`celldefine
module DFFNSQXX1 (Q, XQ, D, XS, XC);
	output Q, XQ;
	input D, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.324806:0.483595:1.96209;
		specparam tpd_XS_Q_negedge_f = 0.324806:0.483595:1.96209;
		specparam tpd_XC_Q_negedge_r = 0.372218:0.536263:2.02044;
		specparam tpd_XC_Q_negedge_f = 0.333714:0.475141:1.44412;
		specparam tpd_XS_XQ_negedge_r = 0.140055:0.28683:1.2561;
		specparam tpd_XS_XQ_negedge_f = 0.140055:0.28683:1.2561;
		specparam tpd_XC_XQ_negedge_r = 0.450708:0.610421:2.08212;
		specparam tpd_XC_XQ_negedge_f = 0.457854:0.591564:1.52239;
		specparam tsetup_D_XC_XS_posedge_XS_negedge = 0.0490722:0.000640091:-0.381925;
		specparam thold_D_XC_XS_posedge_XS_negedge = 0.0712583:0.118295:0.551595;
		specparam tsetup_D_XC_XS_negedge_XS_negedge = 0.0490722:0.000640091:-0.381925;
		specparam thold_D_XC_XS_negedge_XS_negedge = 0.0712583:0.118295:0.551595;
		specparam trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge = -0.000690663:-0.0471914:-0.256439;
		specparam tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0764637:0.127725:0.450334;
		specparam tpw_XS_negedge = 0.205948:0.341301:2.72095;
		specparam tpw_XC_posedge = 0.324279:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.324279:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& XS, posedge D &&& XS, 
			 tsetup_D_XC_XS_posedge_XS_negedge, 
			 thold_D_XC_XS_posedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XS, negedge D &&& XS, 
			 tsetup_D_XC_XS_negedge_XS_negedge, 
			 thold_D_XC_XS_negedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XS &&& ~D, negedge XC &&& ~D, 
			 trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge XC &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSQX 
`timescale 1ns/10ps
`celldefine
module DFFNSQXX2 (Q, XQ, D, XS, XC);
	output Q, XQ;
	input D, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.381165:0.543331:2.03919;
		specparam tpd_XS_Q_negedge_f = 0.381165:0.543331:2.03919;
		specparam tpd_XC_Q_negedge_r = 0.362102:0.526311:1.95398;
		specparam tpd_XC_Q_negedge_f = 0.3336:0.477024:1.36398;
		specparam tpd_XS_XQ_negedge_r = 0.158555:0.310574:1.29146;
		specparam tpd_XS_XQ_negedge_f = 0.158555:0.310574:1.29146;
		specparam tpd_XC_XQ_negedge_r = 0.487037:0.648314:2.07415;
		specparam tpd_XC_XQ_negedge_f = 0.479545:0.612237:1.47665;
		specparam tsetup_D_XC_XS_posedge_XS_negedge = 0.0549488:0.00982899:-0.31704;
		specparam thold_D_XC_XS_posedge_XS_negedge = 0.0585376:0.103485:0.482842;
		specparam tsetup_D_XC_XS_negedge_XS_negedge = 0.0549488:0.00982899:-0.31704;
		specparam thold_D_XC_XS_negedge_XS_negedge = 0.0585376:0.103485:0.482842;
		specparam trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0103548:-0.0306228:-0.177079;
		specparam tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0625424:0.107112:0.385752;
		specparam tpw_XS_negedge = 0.247865:0.385885:2.72095;
		specparam tpw_XC_posedge = 0.27212:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.27212:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& XS, posedge D &&& XS, 
			 tsetup_D_XC_XS_posedge_XS_negedge, 
			 thold_D_XC_XS_posedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XS, negedge D &&& XS, 
			 tsetup_D_XC_XS_negedge_XS_negedge, 
			 thold_D_XC_XS_negedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XS &&& ~D, negedge XC &&& ~D, 
			 trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge XC &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSQX 
`timescale 1ns/10ps
`celldefine
module DFFNSQXX4 (Q, XQ, D, XS, XC);
	output Q, XQ;
	input D, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.378205:0.539606:2.01983;
		specparam tpd_XS_Q_negedge_f = 0.378205:0.539606:2.01983;
		specparam tpd_XC_Q_negedge_r = 0.391151:0.55631:1.98788;
		specparam tpd_XC_Q_negedge_f = 0.363384:0.508429:1.42516;
		specparam tpd_XS_XQ_negedge_r = 0.147546:0.297019:1.28454;
		specparam tpd_XS_XQ_negedge_f = 0.147546:0.297019:1.28454;
		specparam tpd_XC_XQ_negedge_r = 0.500593:0.657678:2.07391;
		specparam tpd_XC_XQ_negedge_f = 0.501226:0.632559:1.52456;
		specparam tsetup_D_XC_XS_posedge_XS_negedge = 0.0401973:-0.005:-0.334694;
		specparam thold_D_XC_XS_posedge_XS_negedge = 0.0658254:0.111441:0.494058;
		specparam tsetup_D_XC_XS_negedge_XS_negedge = 0.0401973:-0.005:-0.334694;
		specparam thold_D_XC_XS_negedge_XS_negedge = 0.0658254:0.111441:0.494058;
		specparam trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.000469937:-0.0399001:-0.186219;
		specparam tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0629623:0.110385:0.388329;
		specparam tpw_XS_negedge = 0.242438:0.372772:2.72095;
		specparam tpw_XC_posedge = 0.241391:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.241391:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& XS, posedge D &&& XS, 
			 tsetup_D_XC_XS_posedge_XS_negedge, 
			 thold_D_XC_XS_posedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XS, negedge D &&& XS, 
			 tsetup_D_XC_XS_negedge_XS_negedge, 
			 thold_D_XC_XS_negedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XS &&& ~D, negedge XC &&& ~D, 
			 trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge XC &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSQX 
`timescale 1ns/10ps
`celldefine
module DFFNSQXXL (Q, XQ, D, XS, XC);
	output Q, XQ;
	input D, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.304439:0.463252:1.9401;
		specparam tpd_XS_Q_negedge_f = 0.304439:0.463252:1.9401;
		specparam tpd_XC_Q_negedge_r = 0.36704:0.528559:2.00819;
		specparam tpd_XC_Q_negedge_f = 0.328126:0.470363:1.53249;
		specparam tpd_XS_XQ_negedge_r = 0.13752:0.286095:1.33615;
		specparam tpd_XS_XQ_negedge_f = 0.13752:0.286095:1.33615;
		specparam tpd_XC_XQ_negedge_r = 0.427952:0.58668:2.06377;
		specparam tpd_XC_XQ_negedge_f = 0.438735:0.575582:1.60969;
		specparam tsetup_D_XC_XS_posedge_XS_negedge = 0.0499535:-0.00221248:-0.383551;
		specparam thold_D_XC_XS_posedge_XS_negedge = 0.0727257:0.12:0.553603;
		specparam tsetup_D_XC_XS_negedge_XS_negedge = 0.0499535:-0.00221248:-0.383551;
		specparam thold_D_XC_XS_negedge_XS_negedge = 0.0727257:0.12:0.553603;
		specparam trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge = -0.00136368:-0.0486447:-0.256704;
		specparam tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge = 0.0769737:0.124088:0.445976;
		specparam tpw_XS_negedge = 0.18568:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.324279:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.324279:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& XS, posedge D &&& XS, 
			 tsetup_D_XC_XS_posedge_XS_negedge, 
			 thold_D_XC_XS_posedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& XS, negedge D &&& XS, 
			 tsetup_D_XC_XS_negedge_XS_negedge, 
			 thold_D_XC_XS_negedge_XS_negedge, notifier,,, delayed_XC, delayed_D);
		$recovery (posedge XS &&& ~D, negedge XC &&& ~D, 
			 trecovery_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge XC &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XC_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSRQ 
`timescale 1ns/10ps
`celldefine
module DFFNSRQX1 (Q, D, XR, XS, XC);
	output Q;
	input D, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.125318:0.251128:1.43307;
		specparam tpd_XR_Q_negedge_f = 0.118481:0.255585:1.17831;
		specparam tpd_XS_Q_negedge_r = 0.338619:0.503932:1.97576;
		specparam tpd_XS_Q_negedge_f = 0.338619:0.503932:1.97576;
		specparam tpd_XC_Q_negedge_r = 0.400368:0.569222:2.02856;
		specparam tpd_XC_Q_negedge_f = 0.344352:0.482064:1.39287;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.0348314:-0.0137623:-0.405054;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = 0.0755102:0.125804:0.574726;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.0348314:-0.0137623:-0.405054;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = 0.0755102:0.125804:0.574726;
		specparam trecovery_XR_XC_adacond1_posedge_adacond1_negedge = -0.281472:-0.337:-0.485315;
		specparam tremoval_XR_XC_adacond1_posedge_adacond1_negedge = 0.410307:0.521259:1.21857;
		specparam tpw_XR_negedge = 0.337323:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0127215:0.00120794:0.0222495;
		specparam thold_XR_XS_posedge_posedge = 0.0468551:0.0581851:0.131098;
		specparam trecovery_XS_XC_adacond2_posedge_adacond2_negedge = 0.00208896:-0.0427328:-0.216796;
		specparam tremoval_XS_XC_adacond2_posedge_adacond2_negedge = 0.0843182:0.134582:0.430291;
		specparam tsetup_XS_XR_posedge_posedge = 0.0381898:0.0572803:0.180262;
		specparam thold_XS_XR_posedge_posedge = 0.0476258:0.0581153:0.0487559;
		specparam tpw_XS_negedge = 0.204446:0.338678:2.72095;
		specparam tpw_XC_posedge = 0.344478:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.344478:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge XC &&& adacond1, 
			 trecovery_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge XC &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge XC &&& adacond2, 
			 trecovery_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge XC &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSRQ 
`timescale 1ns/10ps
`celldefine
module DFFNSRQX2 (Q, D, XR, XS, XC);
	output Q;
	input D, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.140825:0.274422:1.46356;
		specparam tpd_XR_Q_negedge_f = 0.137247:0.283402:1.23785;
		specparam tpd_XS_Q_negedge_r = 0.359534:0.529839:1.99013;
		specparam tpd_XS_Q_negedge_f = 0.359534:0.529839:1.99013;
		specparam tpd_XC_Q_negedge_r = 0.390022:0.560025:1.95512;
		specparam tpd_XC_Q_negedge_f = 0.341976:0.483776:1.34033;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.046846:0.005:-0.325287;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = 0.0576643:0.104399:0.489618;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.046846:0.005:-0.325287;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = 0.0576643:0.104399:0.489618;
		specparam trecovery_XR_XC_adacond1_posedge_adacond1_negedge = -0.249375:-0.298877:-0.317216;
		specparam tremoval_XR_XC_adacond1_posedge_adacond1_negedge = 0.389283:0.495131:1.14882;
		specparam tpw_XR_negedge = 0.342486:0.435715:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0151904:0.00527768:0.0528624;
		specparam thold_XR_XS_posedge_posedge = 0.0317232:0.040574:0.111665;
		specparam trecovery_XS_XC_adacond2_posedge_adacond2_negedge = 0.0144528:-0.0264003:-0.127341;
		specparam tremoval_XS_XC_adacond2_posedge_adacond2_negedge = 0.0694549:0.112874:0.358727;
		specparam tsetup_XS_XR_posedge_posedge = 0.0300076:0.0466011:0.179852;
		specparam thold_XS_XR_posedge_posedge = 0.0506115:0.0585097:0.0844956;
		specparam tpw_XS_negedge = 0.212135:0.346546:2.72095;
		specparam tpw_XC_posedge = 0.293291:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.293291:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge XC &&& adacond1, 
			 trecovery_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge XC &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge XC &&& adacond2, 
			 trecovery_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge XC &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSRQ 
`timescale 1ns/10ps
`celldefine
module DFFNSRQX4 (Q, D, XR, XS, XC);
	output Q;
	input D, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.14274:0.275182:1.45718;
		specparam tpd_XR_Q_negedge_f = 0.136952:0.283423:1.23793;
		specparam tpd_XS_Q_negedge_r = 0.40274:0.573972:2.04474;
		specparam tpd_XS_Q_negedge_f = 0.40274:0.573972:2.04474;
		specparam tpd_XC_Q_negedge_r = 0.442042:0.613942:2.01101;
		specparam tpd_XC_Q_negedge_f = 0.392397:0.535765:1.40287;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.0275397:-0.014:-0.344434;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = 0.0659517:0.115792:0.503199;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.0275397:-0.014:-0.344434;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = 0.0659517:0.115792:0.503199;
		specparam trecovery_XR_XC_adacond1_posedge_adacond1_negedge = -0.273142:-0.34072:-0.408067;
		specparam tremoval_XR_XC_adacond1_posedge_adacond1_negedge = 0.383714:0.491133:1.1495;
		specparam tpw_XR_negedge = 0.36097:0.446205:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0160492:0.0200938:0.10914;
		specparam thold_XR_XS_posedge_posedge = 0.0376927:0.0521995:0.135159;
		specparam trecovery_XS_XC_adacond2_posedge_adacond2_negedge = -0.00159063:-0.041279:-0.140072;
		specparam tremoval_XS_XC_adacond2_posedge_adacond2_negedge = 0.071037:0.115673:0.358562;
		specparam tsetup_XS_XR_posedge_posedge = 0.0153897:0.0186358:0.169299;
		specparam thold_XS_XR_posedge_posedge = 0.0554021:0.0623464:0.138932;
		specparam tpw_XS_negedge = 0.237915:0.37015:2.72095;
		specparam tpw_XC_posedge = 0.259664:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.259664:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge XC &&& adacond1, 
			 trecovery_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge XC &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge XC &&& adacond2, 
			 trecovery_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge XC &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSRQ 
`timescale 1ns/10ps
`celldefine
module DFFNSRQXL (Q, D, XR, XS, XC);
	output Q;
	input D, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.123302:0.24493:1.41795;
		specparam tpd_XR_Q_negedge_f = 0.116984:0.254377:1.26016;
		specparam tpd_XS_Q_negedge_r = 0.332953:0.494898:1.9605;
		specparam tpd_XS_Q_negedge_f = 0.332953:0.494898:1.9605;
		specparam tpd_XC_Q_negedge_r = 0.39601:0.561612:2.01582;
		specparam tpd_XC_Q_negedge_f = 0.340822:0.480568:1.49566;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.0336667:-0.0135164:-0.408257;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = 0.075698:0.126486:0.576142;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.0336667:-0.0135164:-0.408257;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = 0.075698:0.126486:0.576142;
		specparam trecovery_XR_XC_adacond1_posedge_adacond1_negedge = -0.280745:-0.335531:-0.499644;
		specparam tremoval_XR_XC_adacond1_posedge_adacond1_negedge = 0.414304:0.521259:1.21857;
		specparam tpw_XR_negedge = 0.339738:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0119051:0.00333537:0.00604527;
		specparam thold_XR_XS_posedge_posedge = 0.0502978:0.0666707:0.138895;
		specparam trecovery_XS_XC_adacond2_posedge_adacond2_negedge = 0.000780342:-0.0456846:-0.217404;
		specparam tremoval_XS_XC_adacond2_posedge_adacond2_negedge = 0.0834175:0.133903:0.431198;
		specparam tsetup_XS_XR_posedge_posedge = 0.0386664:0.0624279:0.180063;
		specparam thold_XS_XR_posedge_posedge = 0.0486497:0.0584917:0.0499985;
		specparam tpw_XS_negedge = 0.201502:0.336056:2.72095;
		specparam tpw_XC_posedge = 0.344478:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.344478:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge XC &&& adacond1, 
			 trecovery_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge XC &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge XC &&& adacond2, 
			 trecovery_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge XC &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSRQX 
`timescale 1ns/10ps
`celldefine
module DFFNSRQXX1 (Q, XQ, D, XR, XS, XC);
	output Q, XQ;
	input D, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.12573:0.250009:1.40919;
		specparam tpd_XR_Q_negedge_f = 0.119096:0.254735:1.16747;
		specparam tpd_XS_Q_negedge_r = 0.34522:0.508925:1.96177;
		specparam tpd_XS_Q_negedge_f = 0.34522:0.508925:1.96177;
		specparam tpd_XC_Q_negedge_r = 0.405712:0.572077:2.01109;
		specparam tpd_XC_Q_negedge_f = 0.350702:0.48718:1.38931;
		specparam tpd_XR_XQ_negedge_r = 0.276965:0.454653:1.89292;
		specparam tpd_XR_XQ_negedge_f = 0.276965:0.454653:1.89292;
		specparam tpd_XS_XQ_negedge_r = 0.152247:0.302567:1.54904;
		specparam tpd_XS_XQ_negedge_f = 0.142634:0.289973:1.31135;
		specparam tpd_XC_XQ_negedge_r = 0.470625:0.628851:2.07375;
		specparam tpd_XC_XQ_negedge_f = 0.494512:0.628365:1.584;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.0352384:-0.013951:-0.404853;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = 0.0759414:0.126296:0.574872;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.0352384:-0.013951:-0.404853;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = 0.0759414:0.126296:0.574872;
		specparam trecovery_XR_XC_adacond1_posedge_adacond1_negedge = -0.283768:-0.341419:-0.492626;
		specparam tremoval_XR_XC_adacond1_posedge_adacond1_negedge = 0.410513:0.521259:1.21982;
		specparam tpw_XR_negedge = 0.341604:0.427847:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0121601:-2.70039e-05:-0.00874389;
		specparam thold_XR_XS_posedge_posedge = 0.0560964:0.0771004:0.155663;
		specparam trecovery_XS_XC_adacond2_posedge_adacond2_negedge = 0.00162942:-0.0432596:-0.215816;
		specparam tremoval_XS_XC_adacond2_posedge_adacond2_negedge = 0.0843182:0.134582:0.427324;
		specparam tsetup_XS_XR_posedge_posedge = 0.0576627:0.0896626:0.245299;
		specparam thold_XS_XR_posedge_posedge = 0.0112432:-2.70039e-05:-0.0965731;
		specparam tpw_XS_negedge = 0.217712:0.346546:2.72095;
		specparam tpw_XC_posedge = 0.344478:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.344478:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge XC &&& adacond1, 
			 trecovery_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge XC &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge XC &&& adacond2, 
			 trecovery_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge XC &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSRQX 
`timescale 1ns/10ps
`celldefine
module DFFNSRQXX2 (Q, XQ, D, XR, XS, XC);
	output Q, XQ;
	input D, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.143536:0.277411:1.46315;
		specparam tpd_XR_Q_negedge_f = 0.139554:0.285546:1.24199;
		specparam tpd_XS_Q_negedge_r = 0.412581:0.58041:2.05377;
		specparam tpd_XS_Q_negedge_f = 0.412581:0.58041:2.05377;
		specparam tpd_XC_Q_negedge_r = 0.399735:0.568802:1.9616;
		specparam tpd_XC_Q_negedge_f = 0.351541:0.493511:1.35277;
		specparam tpd_XR_XQ_negedge_r = 0.33584:0.519288:2.01002;
		specparam tpd_XR_XQ_negedge_f = 0.33584:0.519288:2.01002;
		specparam tpd_XS_XQ_negedge_r = 0.170181:0.327892:1.6131;
		specparam tpd_XS_XQ_negedge_f = 0.158786:0.311015:1.33023;
		specparam tpd_XC_XQ_negedge_r = 0.50708:0.667645:2.07237;
		specparam tpd_XC_XQ_negedge_f = 0.523452:0.654141:1.52616;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.0465245:0.001:-0.327431;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = 0.0597737:0.104757:0.490697;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.0465245:0.001:-0.327431;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = 0.0597737:0.104757:0.490697;
		specparam trecovery_XR_XC_adacond1_posedge_adacond1_negedge = -0.251662:-0.304823:-0.326564;
		specparam tremoval_XR_XC_adacond1_posedge_adacond1_negedge = 0.38553:0.492755:1.14527;
		specparam tpw_XR_negedge = 0.344728:0.435715:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0137748:0.00294929:0.00179658;
		specparam thold_XR_XS_posedge_posedge = 0.0595707:0.0772882:0.157577;
		specparam trecovery_XS_XC_adacond2_posedge_adacond2_negedge = 0.0139126:-0.0284322:-0.128852;
		specparam tremoval_XS_XC_adacond2_posedge_adacond2_negedge = 0.0672198:0.110502:0.359116;
		specparam tsetup_XS_XR_posedge_posedge = 0.0673878:0.100953:0.258484;
		specparam thold_XS_XR_posedge_posedge = 0.0157497:0.00294929:-0.0960501;
		specparam tpw_XS_negedge = 0.26099:0.393753:2.72095;
		specparam tpw_XC_posedge = 0.293291:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.293291:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge XC &&& adacond1, 
			 trecovery_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge XC &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge XC &&& adacond2, 
			 trecovery_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge XC &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSRQX 
`timescale 1ns/10ps
`celldefine
module DFFNSRQXX4 (Q, XQ, D, XR, XS, XC);
	output Q, XQ;
	input D, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.145125:0.279511:1.48168;
		specparam tpd_XR_Q_negedge_f = 0.138741:0.28583:1.25411;
		specparam tpd_XS_Q_negedge_r = 0.432135:0.602691:2.09388;
		specparam tpd_XS_Q_negedge_f = 0.432135:0.602691:2.09388;
		specparam tpd_XC_Q_negedge_r = 0.454048:0.626717:2.04866;
		specparam tpd_XC_Q_negedge_f = 0.40456:0.548904:1.43046;
		specparam tpd_XR_XQ_negedge_r = 0.304453:0.478842:1.97152;
		specparam tpd_XR_XQ_negedge_f = 0.304453:0.478842:1.97152;
		specparam tpd_XS_XQ_negedge_r = 0.141546:0.288194:1.52686;
		specparam tpd_XS_XQ_negedge_f = 0.144289:0.291328:1.26892;
		specparam tpd_XC_XQ_negedge_r = 0.548407:0.705732:2.12627;
		specparam tpd_XC_XQ_negedge_f = 0.569249:0.694891:1.5411;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.026855:-0.014:-0.345073;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = 0.066581:0.118197:0.503675;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.026855:-0.014:-0.345073;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = 0.066581:0.118197:0.503675;
		specparam trecovery_XR_XC_adacond1_posedge_adacond1_negedge = -0.277032:-0.35089:-0.412972;
		specparam tremoval_XR_XC_adacond1_posedge_adacond1_negedge = 0.379962:0.488738:1.14996;
		specparam tpw_XR_negedge = 0.364896:0.448828:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0156056:0.00124518:0.0507074;
		specparam thold_XR_XS_posedge_posedge = 0.0509401:0.0625699:0.141378;
		specparam trecovery_XS_XC_adacond2_posedge_adacond2_negedge = -0.00412171:-0.0436374:-0.140867;
		specparam tremoval_XS_XC_adacond2_posedge_adacond2_negedge = 0.071037:0.115673:0.3556;
		specparam tsetup_XS_XR_posedge_posedge = 0.0475644:0.0718983:0.206819;
		specparam thold_XS_XR_posedge_posedge = 0.014624:0.0012982:-0.0630279;
		specparam tpw_XS_negedge = 0.271157:0.388508:2.72095;
		specparam tpw_XC_posedge = 0.259371:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.259371:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge XC &&& adacond1, 
			 trecovery_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge XC &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge XC &&& adacond2, 
			 trecovery_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge XC &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFNSRQX 
`timescale 1ns/10ps
`celldefine
module DFFNSRQXXL (Q, XQ, D, XR, XS, XC);
	output Q, XQ;
	input D, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.123872:0.246131:1.42468;
		specparam tpd_XR_Q_negedge_f = 0.117316:0.254569:1.26582;
		specparam tpd_XS_Q_negedge_r = 0.340042:0.502437:1.97372;
		specparam tpd_XS_Q_negedge_f = 0.340042:0.502437:1.97372;
		specparam tpd_XC_Q_negedge_r = 0.401427:0.56668:2.02478;
		specparam tpd_XC_Q_negedge_f = 0.346921:0.486905:1.51203;
		specparam tpd_XR_XQ_negedge_r = 0.258783:0.435109:1.86992;
		specparam tpd_XR_XQ_negedge_f = 0.258783:0.435109:1.86992;
		specparam tpd_XS_XQ_negedge_r = 0.15052:0.299224:1.55533;
		specparam tpd_XS_XQ_negedge_f = 0.138808:0.285471:1.34911;
		specparam tpd_XC_XQ_negedge_r = 0.44974:0.607732:2.07022;
		specparam tpd_XC_XQ_negedge_f = 0.474872:0.610211:1.62833;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.0324728:-0.0131933:-0.405445;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = 0.0758393:0.126589:0.573554;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.0324728:-0.0131933:-0.405445;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = 0.0758393:0.126589:0.573554;
		specparam trecovery_XR_XC_adacond1_posedge_adacond1_negedge = -0.28347:-0.338343:-0.505211;
		specparam tremoval_XR_XC_adacond1_posedge_adacond1_negedge = 0.414304:0.521259:1.21982;
		specparam tpw_XR_negedge = 0.343448:0.427847:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0110957:-2.70039e-05:-0.0114676;
		specparam thold_XR_XS_posedge_posedge = 0.0537842:0.0747337:0.145756;
		specparam trecovery_XS_XC_adacond2_posedge_adacond2_negedge = -0.000643911:-0.0430113:-0.218823;
		specparam tremoval_XS_XC_adacond2_posedge_adacond2_negedge = 0.0821221:0.132054:0.429464;
		specparam tsetup_XS_XR_posedge_posedge = 0.0540697:0.0878454:0.22611;
		specparam thold_XS_XR_posedge_posedge = 0.0110957:-2.70039e-05:-0.0925756;
		specparam tpw_XS_negedge = 0.20314:0.341301:2.72095;
		specparam tpw_XC_posedge = 0.344478:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.344478:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:D)) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:D)) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge XC &&& adacond1, 
			 trecovery_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge XC &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XC_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge XC &&& adacond2, 
			 trecovery_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge XC &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XC_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFQ 
`timescale 1ns/10ps
`celldefine
module DFFQX1 (Q, D, C);
	output Q;
	input D, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, xcr_0;

	altos_dff_err (xcr_0, delayed_C, delayed_D);
	altos_dff (int_fwire_IQ, notifier, delayed_C, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_C_Q_posedge_r = 0.340521:0.481889:1.65266;
		specparam tpd_C_Q_posedge_f = 0.35686:0.486679:1.23992;
		specparam tsetup_D_C_posedge_posedge = 0.133727:0.117885:0.137624;
		specparam thold_D_C_posedge_posedge = -0.0498018:-0.0590555:-0.0827271;
		specparam tsetup_D_C_negedge_posedge = 0.133727:0.117885:0.137624;
		specparam thold_D_C_negedge_posedge = -0.0498018:-0.0590555:-0.0827271;
		specparam tpw_C_posedge = 0.192788:0.330811:2.72095;
		specparam tpw_C_negedge = 0.192788:0.330811:2.72095;

		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C, posedge D, 
			 tsetup_D_C_posedge_posedge, 
			 thold_D_C_posedge_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C, negedge D, 
			 tsetup_D_C_negedge_posedge, 
			 thold_D_C_negedge_posedge, notifier,,, delayed_C, delayed_D);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFQ 
`timescale 1ns/10ps
`celldefine
module DFFQX2 (Q, D, C);
	output Q;
	input D, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, xcr_0;

	altos_dff_err (xcr_0, delayed_C, delayed_D);
	altos_dff (int_fwire_IQ, notifier, delayed_C, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_C_Q_posedge_r = 0.326804:0.469366:1.6528;
		specparam tpd_C_Q_posedge_f = 0.334618:0.460657:1.17225;
		specparam tsetup_D_C_posedge_posedge = 0.109831:0.10614:0.145363;
		specparam thold_D_C_posedge_posedge = -0.0450546:-0.0582791:-0.0953827;
		specparam tsetup_D_C_negedge_posedge = 0.109831:0.10614:0.145363;
		specparam thold_D_C_negedge_posedge = -0.0450546:-0.0582791:-0.0953827;
		specparam tpw_C_posedge = 0.195087:0.330811:2.72095;
		specparam tpw_C_negedge = 0.195087:0.330811:2.72095;

		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C, posedge D, 
			 tsetup_D_C_posedge_posedge, 
			 thold_D_C_posedge_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C, negedge D, 
			 tsetup_D_C_negedge_posedge, 
			 thold_D_C_negedge_posedge, notifier,,, delayed_C, delayed_D);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFQ 
`timescale 1ns/10ps
`celldefine
module DFFQX4 (Q, D, C);
	output Q;
	input D, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, xcr_0;

	altos_dff_err (xcr_0, delayed_C, delayed_D);
	altos_dff (int_fwire_IQ, notifier, delayed_C, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_C_Q_posedge_r = 0.380111:0.521999:1.67508;
		specparam tpd_C_Q_posedge_f = 0.356062:0.475254:1.10958;
		specparam tsetup_D_C_posedge_posedge = 0.0880327:0.089487:0.130348;
		specparam thold_D_C_posedge_posedge = -0.0393427:-0.049409:-0.0864595;
		specparam tsetup_D_C_negedge_posedge = 0.0880327:0.089487:0.130348;
		specparam thold_D_C_negedge_posedge = -0.0393427:-0.049409:-0.0864595;
		specparam tpw_C_posedge = 0.247192:0.330811:2.72095;
		specparam tpw_C_negedge = 0.247192:0.330811:2.72095;

		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C, posedge D, 
			 tsetup_D_C_posedge_posedge, 
			 thold_D_C_posedge_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C, negedge D, 
			 tsetup_D_C_negedge_posedge, 
			 thold_D_C_negedge_posedge, notifier,,, delayed_C, delayed_D);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFQ 
`timescale 1ns/10ps
`celldefine
module DFFQXL (Q, D, C);
	output Q;
	input D, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, xcr_0;

	altos_dff_err (xcr_0, delayed_C, delayed_D);
	altos_dff (int_fwire_IQ, notifier, delayed_C, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_C_Q_posedge_r = 0.339308:0.479845:1.67047;
		specparam tpd_C_Q_posedge_f = 0.349686:0.474497:1.20993;
		specparam tsetup_D_C_posedge_posedge = 0.135542:0.117885:0.137496;
		specparam thold_D_C_posedge_posedge = -0.0490312:-0.0590375:-0.0823977;
		specparam tsetup_D_C_negedge_posedge = 0.135542:0.117885:0.137496;
		specparam thold_D_C_negedge_posedge = -0.0490312:-0.0590375:-0.0823977;
		specparam tpw_C_posedge = 0.190377:0.330811:2.72095;
		specparam tpw_C_negedge = 0.190377:0.330811:2.72095;

		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C, posedge D, 
			 tsetup_D_C_posedge_posedge, 
			 thold_D_C_posedge_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C, negedge D, 
			 tsetup_D_C_negedge_posedge, 
			 thold_D_C_negedge_posedge, notifier,,, delayed_C, delayed_D);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFQX 
`timescale 1ns/10ps
`celldefine
module DFFQXX1 (Q, XQ, D, C);
	output Q, XQ;
	input D, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, xcr_0;

	altos_dff_err (xcr_0, delayed_C, delayed_D);
	altos_dff (int_fwire_IQ, notifier, delayed_C, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_C_Q_posedge_r = 0.336453:0.477262:1.66788;
		specparam tpd_C_Q_posedge_f = 0.35462:0.483265:1.24111;
		specparam tpd_C_XQ_posedge_r = 0.436449:0.56917:1.73483;
		specparam tpd_C_XQ_posedge_f = 0.438:0.560632:1.35309;
		specparam tsetup_D_C_posedge_posedge = 0.141053:0.125665:0.148462;
		specparam thold_D_C_posedge_posedge = -0.0534608:-0.062618:-0.0931804;
		specparam tsetup_D_C_negedge_posedge = 0.141053:0.125665:0.148462;
		specparam thold_D_C_negedge_posedge = -0.0534608:-0.062618:-0.0931804;
		specparam tpw_C_posedge = 0.19899:0.330811:2.72095;
		specparam tpw_C_negedge = 0.19899:0.330811:2.72095;

		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C, posedge D, 
			 tsetup_D_C_posedge_posedge, 
			 thold_D_C_posedge_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C, negedge D, 
			 tsetup_D_C_negedge_posedge, 
			 thold_D_C_negedge_posedge, notifier,,, delayed_C, delayed_D);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFQX 
`timescale 1ns/10ps
`celldefine
module DFFQXX2 (Q, XQ, D, C);
	output Q, XQ;
	input D, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, xcr_0;

	altos_dff_err (xcr_0, delayed_C, delayed_D);
	altos_dff (int_fwire_IQ, notifier, delayed_C, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_C_Q_posedge_r = 0.327482:0.466531:1.63782;
		specparam tpd_C_Q_posedge_f = 0.33587:0.458908:1.16359;
		specparam tpd_C_XQ_posedge_r = 0.430292:0.561216:1.72572;
		specparam tpd_C_XQ_posedge_f = 0.425584:0.540688:1.25675;
		specparam tsetup_D_C_posedge_posedge = 0.111298:0.10614:0.14643;
		specparam thold_D_C_posedge_posedge = -0.0451315:-0.0585159:-0.0963364;
		specparam tsetup_D_C_negedge_posedge = 0.111298:0.10614:0.14643;
		specparam thold_D_C_negedge_posedge = -0.0451315:-0.0585159:-0.0963364;
		specparam tpw_C_posedge = 0.205376:0.330811:2.72095;
		specparam tpw_C_negedge = 0.205376:0.330811:2.72095;

		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C, posedge D, 
			 tsetup_D_C_posedge_posedge, 
			 thold_D_C_posedge_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C, negedge D, 
			 tsetup_D_C_negedge_posedge, 
			 thold_D_C_negedge_posedge, notifier,,, delayed_C, delayed_D);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFQX 
`timescale 1ns/10ps
`celldefine
module DFFQXX4 (Q, XQ, D, C);
	output Q, XQ;
	input D, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, xcr_0;

	altos_dff_err (xcr_0, delayed_C, delayed_D);
	altos_dff (int_fwire_IQ, notifier, delayed_C, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_C_Q_posedge_r = 0.392892:0.538453:1.73302;
		specparam tpd_C_Q_posedge_f = 0.369369:0.491995:1.14276;
		specparam tpd_C_XQ_posedge_r = 0.467156:0.596019:1.76921;
		specparam tpd_C_XQ_posedge_f = 0.484029:0.589065:1.22781;
		specparam tsetup_D_C_posedge_posedge = 0.084267:0.0836083:0.0980512;
		specparam thold_D_C_posedge_posedge = -0.0359078:-0.0470833:-0.0585818;
		specparam tsetup_D_C_negedge_posedge = 0.084267:0.0836083:0.0980512;
		specparam thold_D_C_negedge_posedge = -0.0359078:-0.0470833:-0.0585818;
		specparam tpw_C_posedge = 0.275936:0.330811:2.72095;
		specparam tpw_C_negedge = 0.275936:0.330811:2.72095;

		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C, posedge D, 
			 tsetup_D_C_posedge_posedge, 
			 thold_D_C_posedge_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C, negedge D, 
			 tsetup_D_C_negedge_posedge, 
			 thold_D_C_negedge_posedge, notifier,,, delayed_C, delayed_D);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFQX 
`timescale 1ns/10ps
`celldefine
module DFFQXXL (Q, XQ, D, C);
	output Q, XQ;
	input D, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, xcr_0;

	altos_dff_err (xcr_0, delayed_C, delayed_D);
	altos_dff (int_fwire_IQ, notifier, delayed_C, delayed_D, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_C_Q_posedge_r = 0.335805:0.473245:1.64684;
		specparam tpd_C_Q_posedge_f = 0.348235:0.470145:1.19185;
		specparam tpd_C_XQ_posedge_r = 0.424223:0.557304:1.72941;
		specparam tpd_C_XQ_posedge_f = 0.422255:0.542043:1.32972;
		specparam tsetup_D_C_posedge_posedge = 0.139786:0.125669:0.14828;
		specparam thold_D_C_posedge_posedge = -0.0497372:-0.0627406:-0.0918572;
		specparam tsetup_D_C_negedge_posedge = 0.139786:0.125669:0.14828;
		specparam thold_D_C_negedge_posedge = -0.0497372:-0.0627406:-0.0918572;
		specparam tpw_C_posedge = 0.192759:0.330811:2.72095;
		specparam tpw_C_negedge = 0.192759:0.330811:2.72095;

		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C, posedge D, 
			 tsetup_D_C_posedge_posedge, 
			 thold_D_C_posedge_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C, negedge D, 
			 tsetup_D_C_negedge_posedge, 
			 thold_D_C_negedge_posedge, notifier,,, delayed_C, delayed_D);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFRQ 
`timescale 1ns/10ps
`celldefine
module DFFRQX1 (Q, D, XR, C);
	output Q;
	input D, XR, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_r, xcr_0;

	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.119322:0.259519:1.23144;
		specparam tpd_XR_Q_negedge_f = 0.119322:0.259519:1.23144;
		specparam tpd_C_Q_posedge_r = 0.363879:0.510765:1.69829;
		specparam tpd_C_Q_posedge_f = 0.351691:0.472544:1.1681;
		specparam tsetup_D_C_XR_posedge_XR_posedge = 0.144194:0.131587:0.155098;
		specparam thold_D_C_XR_posedge_XR_posedge = -0.0617841:-0.0734618:-0.0966717;
		specparam tsetup_D_C_XR_negedge_XR_posedge = 0.144194:0.131587:0.155098;
		specparam thold_D_C_XR_negedge_XR_posedge = -0.0617841:-0.0734618:-0.0966717;
		specparam trecovery_XR_C_D_posedge_D_posedge = -0.196657:-0.256799:0.0177881;
		specparam tremoval_XR_C_D_posedge_D_posedge = 0.255857:0.354139:0.800991;
		specparam tpw_XR_negedge = 0.304423:0.398998:2.72095;
		specparam tpw_C_posedge = 0.211647:0.330811:2.72095;
		specparam tpw_C_negedge = 0.211647:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& XR, posedge D &&& XR, 
			 tsetup_D_C_XR_posedge_XR_posedge, 
			 thold_D_C_XR_posedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XR, negedge D &&& XR, 
			 tsetup_D_C_XR_negedge_XR_posedge, 
			 thold_D_C_XR_negedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XR &&& D, posedge C &&& D, 
			 trecovery_XR_C_D_posedge_D_posedge, notifier);
		$hold (posedge C &&& D, posedge XR &&& D, 
			 tremoval_XR_C_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFRQ 
`timescale 1ns/10ps
`celldefine
module DFFRQX2 (Q, D, XR, C);
	output Q;
	input D, XR, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_r, xcr_0;

	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.135603:0.282001:1.22936;
		specparam tpd_XR_Q_negedge_f = 0.135603:0.282001:1.22936;
		specparam tpd_C_Q_posedge_r = 0.373575:0.527097:1.72774;
		specparam tpd_C_Q_posedge_f = 0.338963:0.46292:1.10122;
		specparam tsetup_D_C_XR_posedge_XR_posedge = 0.122378:0.113047:0.133363;
		specparam thold_D_C_XR_posedge_XR_posedge = -0.052623:-0.0655302:-0.0842735;
		specparam tsetup_D_C_XR_negedge_XR_posedge = 0.122378:0.113047:0.133363;
		specparam thold_D_C_XR_negedge_XR_posedge = -0.052623:-0.0655302:-0.0842735;
		specparam trecovery_XR_C_D_posedge_D_posedge = -0.186878:-0.241203:0.0934334;
		specparam tremoval_XR_C_D_posedge_D_posedge = 0.25225:0.346674:0.809844;
		specparam tpw_XR_negedge = 0.309858:0.404243:2.72095;
		specparam tpw_C_posedge = 0.228933:0.330811:2.72095;
		specparam tpw_C_negedge = 0.228933:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& XR, posedge D &&& XR, 
			 tsetup_D_C_XR_posedge_XR_posedge, 
			 thold_D_C_XR_posedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XR, negedge D &&& XR, 
			 tsetup_D_C_XR_negedge_XR_posedge, 
			 thold_D_C_XR_negedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XR &&& D, posedge C &&& D, 
			 trecovery_XR_C_D_posedge_D_posedge, notifier);
		$hold (posedge C &&& D, posedge XR &&& D, 
			 tremoval_XR_C_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFRQ 
`timescale 1ns/10ps
`celldefine
module DFFRQX4 (Q, D, XR, C);
	output Q;
	input D, XR, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_r, xcr_0;

	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.135735:0.284561:1.26181;
		specparam tpd_XR_Q_negedge_f = 0.135735:0.284561:1.26181;
		specparam tpd_C_Q_posedge_r = 0.436395:0.59223:1.79229;
		specparam tpd_C_Q_posedge_f = 0.375582:0.502534:1.16641;
		specparam tsetup_D_C_XR_posedge_XR_posedge = 0.100795:0.0990951:0.126395;
		specparam thold_D_C_XR_posedge_XR_posedge = -0.0449106:-0.0563548:-0.078795;
		specparam tsetup_D_C_XR_negedge_XR_posedge = 0.100795:0.0990951:0.126395;
		specparam thold_D_C_XR_negedge_XR_posedge = -0.0449106:-0.0563548:-0.078795;
		specparam trecovery_XR_C_D_posedge_D_posedge = -0.185605:-0.26658:-0.0248395;
		specparam tremoval_XR_C_D_posedge_D_posedge = 0.239555:0.336971:0.799518;
		specparam tpw_XR_negedge = 0.324051:0.417356:2.72095;
		specparam tpw_C_posedge = 0.291615:0.330811:2.72095;
		specparam tpw_C_negedge = 0.291615:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& XR, posedge D &&& XR, 
			 tsetup_D_C_XR_posedge_XR_posedge, 
			 thold_D_C_XR_posedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XR, negedge D &&& XR, 
			 tsetup_D_C_XR_negedge_XR_posedge, 
			 thold_D_C_XR_negedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XR &&& D, posedge C &&& D, 
			 trecovery_XR_C_D_posedge_D_posedge, notifier);
		$hold (posedge C &&& D, posedge XR &&& D, 
			 tremoval_XR_C_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFRQ 
`timescale 1ns/10ps
`celldefine
module DFFRQXL (Q, D, XR, C);
	output Q;
	input D, XR, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_r, xcr_0;

	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.119103:0.255818:1.27363;
		specparam tpd_XR_Q_negedge_f = 0.119103:0.255818:1.27363;
		specparam tpd_C_Q_posedge_r = 0.362929:0.505589:1.69545;
		specparam tpd_C_Q_posedge_f = 0.350504:0.469573:1.2275;
		specparam tsetup_D_C_XR_posedge_XR_posedge = 0.143922:0.131606:0.157555;
		specparam thold_D_C_XR_posedge_XR_posedge = -0.0628089:-0.0740062:-0.0992781;
		specparam tsetup_D_C_XR_negedge_XR_posedge = 0.143922:0.131606:0.157555;
		specparam thold_D_C_XR_negedge_XR_posedge = -0.0628089:-0.0740062:-0.0992781;
		specparam trecovery_XR_C_D_posedge_D_posedge = -0.199649:-0.25729:-0.00176561;
		specparam tremoval_XR_C_D_posedge_D_posedge = 0.257384:0.35521:0.803457;
		specparam tpw_XR_negedge = 0.304423:0.398998:2.72095;
		specparam tpw_C_posedge = 0.206584:0.330811:2.72095;
		specparam tpw_C_negedge = 0.206584:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& XR, posedge D &&& XR, 
			 tsetup_D_C_XR_posedge_XR_posedge, 
			 thold_D_C_XR_posedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XR, negedge D &&& XR, 
			 tsetup_D_C_XR_negedge_XR_posedge, 
			 thold_D_C_XR_negedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XR &&& D, posedge C &&& D, 
			 trecovery_XR_C_D_posedge_D_posedge, notifier);
		$hold (posedge C &&& D, posedge XR &&& D, 
			 tremoval_XR_C_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFRQX 
`timescale 1ns/10ps
`celldefine
module DFFRQXX1 (Q, XQ, D, XR, C);
	output Q, XQ;
	input D, XR, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire xcr_0;

	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.116947:0.254219:1.20004;
		specparam tpd_XR_Q_negedge_f = 0.116947:0.254219:1.20004;
		specparam tpd_C_Q_posedge_r = 0.351291:0.495872:1.68179;
		specparam tpd_C_Q_posedge_f = 0.346609:0.464504:1.13268;
		specparam tpd_XR_XQ_negedge_r = 0.231244:0.398658:1.84679;
		specparam tpd_XR_XQ_negedge_f = 0.231244:0.398658:1.84679;
		specparam tpd_C_XQ_posedge_r = 0.434636:0.569581:1.76412;
		specparam tpd_C_XQ_posedge_f = 0.437378:0.549404:1.21778;
		specparam tsetup_D_C_XR_posedge_XR_posedge = 0.147136:0.133333:0.162359;
		specparam thold_D_C_XR_posedge_XR_posedge = -0.060874:-0.0716673:-0.0990706;
		specparam tsetup_D_C_XR_negedge_XR_posedge = 0.147136:0.133333:0.162359;
		specparam thold_D_C_XR_negedge_XR_posedge = -0.060874:-0.0716673:-0.0990706;
		specparam trecovery_XR_C_D_posedge_D_posedge = -0.195786:-0.249867:0.0284831;
		specparam tremoval_XR_C_D_posedge_D_posedge = 0.257488:0.356241:0.804677;
		specparam tpw_XR_negedge = 0.302705:0.396376:2.72095;
		specparam tpw_C_posedge = 0.209115:0.330811:2.72095;
		specparam tpw_C_negedge = 0.209115:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& XR, posedge D &&& XR, 
			 tsetup_D_C_XR_posedge_XR_posedge, 
			 thold_D_C_XR_posedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XR, negedge D &&& XR, 
			 tsetup_D_C_XR_negedge_XR_posedge, 
			 thold_D_C_XR_negedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XR &&& D, posedge C &&& D, 
			 trecovery_XR_C_D_posedge_D_posedge, notifier);
		$hold (posedge C &&& D, posedge XR &&& D, 
			 tremoval_XR_C_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFRQX 
`timescale 1ns/10ps
`celldefine
module DFFRQXX2 (Q, XQ, D, XR, C);
	output Q, XQ;
	input D, XR, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire xcr_0;

	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.134751:0.27977:1.22925;
		specparam tpd_XR_Q_negedge_f = 0.134751:0.27977:1.22925;
		specparam tpd_C_Q_posedge_r = 0.36241:0.513531:1.71618;
		specparam tpd_C_Q_posedge_f = 0.335201:0.45781:1.09796;
		specparam tpd_XR_XQ_negedge_r = 0.283646:0.454976:1.93391;
		specparam tpd_XR_XQ_negedge_f = 0.283646:0.454976:1.93391;
		specparam tpd_C_XQ_posedge_r = 0.455791:0.59164:1.78142;
		specparam tpd_C_XQ_posedge_f = 0.485933:0.599244:1.25585;
		specparam tsetup_D_C_XR_posedge_XR_posedge = 0.123888:0.118437:0.138263;
		specparam thold_D_C_XR_posedge_XR_posedge = -0.0512505:-0.0626565:-0.0849358;
		specparam tsetup_D_C_XR_negedge_XR_posedge = 0.123888:0.118437:0.138263;
		specparam thold_D_C_XR_negedge_XR_posedge = -0.0512505:-0.0626565:-0.0849358;
		specparam trecovery_XR_C_D_posedge_D_posedge = -0.184859:-0.237318:0.0983524;
		specparam tremoval_XR_C_D_posedge_D_posedge = 0.249893:0.348786:0.807733;
		specparam tpw_XR_negedge = 0.306142:0.401621:2.72095;
		specparam tpw_C_posedge = 0.239353:0.330811:2.72095;
		specparam tpw_C_negedge = 0.239353:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& XR, posedge D &&& XR, 
			 tsetup_D_C_XR_posedge_XR_posedge, 
			 thold_D_C_XR_posedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XR, negedge D &&& XR, 
			 tsetup_D_C_XR_negedge_XR_posedge, 
			 thold_D_C_XR_negedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XR &&& D, posedge C &&& D, 
			 trecovery_XR_C_D_posedge_D_posedge, notifier);
		$hold (posedge C &&& D, posedge XR &&& D, 
			 tremoval_XR_C_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFRQX 
`timescale 1ns/10ps
`celldefine
module DFFRQXX4 (Q, XQ, D, XR, C);
	output Q, XQ;
	input D, XR, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire xcr_0;

	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.133541:0.279286:1.23465;
		specparam tpd_XR_Q_negedge_f = 0.133541:0.279286:1.23465;
		specparam tpd_C_Q_posedge_r = 0.447612:0.601317:1.80658;
		specparam tpd_C_Q_posedge_f = 0.382399:0.506546:1.15248;
		specparam tpd_XR_XQ_negedge_r = 0.256521:0.419221:1.8969;
		specparam tpd_XR_XQ_negedge_f = 0.256521:0.419221:1.8969;
		specparam tpd_C_XQ_posedge_r = 0.488275:0.619721:1.8118;
		specparam tpd_C_XQ_posedge_f = 0.558731:0.666074:1.32091;
		specparam tsetup_D_C_XR_posedge_XR_posedge = 0.0967825:0.0977695:0.1233;
		specparam thold_D_C_XR_posedge_XR_posedge = -0.0424496:-0.0524583:-0.0763303;
		specparam tsetup_D_C_XR_negedge_XR_posedge = 0.0967825:0.0977695:0.1233;
		specparam thold_D_C_XR_negedge_XR_posedge = -0.0424496:-0.0524583:-0.0763303;
		specparam trecovery_XR_C_D_posedge_D_posedge = -0.186756:-0.269673:-0.0390992;
		specparam tremoval_XR_C_D_posedge_D_posedge = 0.234301:0.334005:0.797243;
		specparam tpw_XR_negedge = 0.326154:0.417356:2.72095;
		specparam tpw_C_posedge = 0.320358:0.330811:2.72095;
		specparam tpw_C_negedge = 0.320358:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& XR, posedge D &&& XR, 
			 tsetup_D_C_XR_posedge_XR_posedge, 
			 thold_D_C_XR_posedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XR, negedge D &&& XR, 
			 tsetup_D_C_XR_negedge_XR_posedge, 
			 thold_D_C_XR_negedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XR &&& D, posedge C &&& D, 
			 trecovery_XR_C_D_posedge_D_posedge, notifier);
		$hold (posedge C &&& D, posedge XR &&& D, 
			 tremoval_XR_C_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFRQX 
`timescale 1ns/10ps
`celldefine
module DFFRQXXL (Q, XQ, D, XR, C);
	output Q, XQ;
	input D, XR, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire xcr_0;

	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, delayed_D, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XR_Q_negedge_r = 0.112436:0.248288:1.25338;
		specparam tpd_XR_Q_negedge_f = 0.112436:0.248288:1.25338;
		specparam tpd_C_Q_posedge_r = 0.34402:0.486255:1.67951;
		specparam tpd_C_Q_posedge_f = 0.340927:0.459399:1.20583;
		specparam tpd_XR_XQ_negedge_r = 0.210986:0.377491:1.81489;
		specparam tpd_XR_XQ_negedge_f = 0.210986:0.377491:1.81489;
		specparam tpd_C_XQ_posedge_r = 0.413656:0.549087:1.74854;
		specparam tpd_C_XQ_posedge_f = 0.412824:0.527345:1.27613;
		specparam tsetup_D_C_XR_posedge_XR_posedge = 0.148633:0.13402:0.162436;
		specparam thold_D_C_XR_posedge_XR_posedge = -0.0634883:-0.0725889:-0.0995821;
		specparam tsetup_D_C_XR_negedge_XR_posedge = 0.148633:0.13402:0.162436;
		specparam thold_D_C_XR_negedge_XR_posedge = -0.0634883:-0.0725889:-0.0995821;
		specparam trecovery_XR_C_D_posedge_D_posedge = -0.196622:-0.249948:0.00133952;
		specparam tremoval_XR_C_D_posedge_D_posedge = 0.257488:0.356241:0.804677;
		specparam tpw_XR_negedge = 0.304657:0.396376:2.72095;
		specparam tpw_C_posedge = 0.200003:0.330811:2.72095;
		specparam tpw_C_negedge = 0.200003:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& XR, posedge D &&& XR, 
			 tsetup_D_C_XR_posedge_XR_posedge, 
			 thold_D_C_XR_posedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XR, negedge D &&& XR, 
			 tsetup_D_C_XR_negedge_XR_posedge, 
			 thold_D_C_XR_negedge_XR_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XR &&& D, posedge C &&& D, 
			 trecovery_XR_C_D_posedge_D_posedge, notifier);
		$hold (posedge C &&& D, posedge XR &&& D, 
			 tremoval_XR_C_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSQ 
`timescale 1ns/10ps
`celldefine
module DFFSQX1 (Q, D, XS, C);
	output Q;
	input D, XS, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_s, xcr_0;

	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.305769:0.466054:1.9365;
		specparam tpd_XS_Q_negedge_f = 0.305769:0.466054:1.9365;
		specparam tpd_C_Q_posedge_r = 0.310843:0.449603:1.61798;
		specparam tpd_C_Q_posedge_f = 0.351035:0.467668:1.10021;
		specparam tsetup_D_C_XS_posedge_XS_posedge = 0.160711:0.148685:0.231425;
		specparam thold_D_C_XS_posedge_XS_posedge = -0.065216:-0.0821631:-0.152067;
		specparam tsetup_D_C_XS_negedge_XS_posedge = 0.160711:0.148685:0.231425;
		specparam thold_D_C_XS_negedge_XS_posedge = -0.065216:-0.0821631:-0.152067;
		specparam trecovery_XS_C_NTB_D_posedge_NTB_D_posedge = -0.0395406:-0.0614261:0.0630605;
		specparam tremoval_XS_C_NTB_D_posedge_NTB_D_posedge = 0.109041:0.131004:0.108159;
		specparam tpw_XS_negedge = 0.182761:0.330811:2.72095;
		specparam tpw_C_posedge = 0.172749:0.330811:2.72095;
		specparam tpw_C_negedge = 0.172749:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& XS, posedge D &&& XS, 
			 tsetup_D_C_XS_posedge_XS_posedge, 
			 thold_D_C_XS_posedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XS, negedge D &&& XS, 
			 tsetup_D_C_XS_negedge_XS_posedge, 
			 thold_D_C_XS_negedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XS &&& ~D, posedge C &&& ~D, 
			 trecovery_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge C &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSQ 
`timescale 1ns/10ps
`celldefine
module DFFSQX2 (Q, D, XS, C);
	output Q;
	input D, XS, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_s, xcr_0;

	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.324933:0.49081:1.97448;
		specparam tpd_XS_Q_negedge_f = 0.324933:0.49081:1.97448;
		specparam tpd_C_Q_posedge_r = 0.31668:0.460593:1.64296;
		specparam tpd_C_Q_posedge_f = 0.345243:0.468592:1.10066;
		specparam tsetup_D_C_XS_posedge_XS_posedge = 0.132783:0.126459:0.192828;
		specparam thold_D_C_XS_posedge_XS_posedge = -0.0525569:-0.0704805:-0.132192;
		specparam tsetup_D_C_XS_negedge_XS_posedge = 0.132783:0.126459:0.192828;
		specparam thold_D_C_XS_negedge_XS_posedge = -0.0525569:-0.0704805:-0.132192;
		specparam trecovery_XS_C_NTB_D_posedge_NTB_D_posedge = -0.0172306:-0.0395919:0.0962612;
		specparam tremoval_XS_C_NTB_D_posedge_NTB_D_posedge = 0.0834533:0.107112:0.0919956;
		specparam tpw_XS_negedge = 0.185988:0.330811:2.72095;
		specparam tpw_C_posedge = 0.18405:0.330811:2.72095;
		specparam tpw_C_negedge = 0.18405:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& XS, posedge D &&& XS, 
			 tsetup_D_C_XS_posedge_XS_posedge, 
			 thold_D_C_XS_posedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XS, negedge D &&& XS, 
			 tsetup_D_C_XS_negedge_XS_posedge, 
			 thold_D_C_XS_negedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XS &&& ~D, posedge C &&& ~D, 
			 trecovery_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge C &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSQ 
`timescale 1ns/10ps
`celldefine
module DFFSQX4 (Q, D, XS, C);
	output Q;
	input D, XS, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_s, xcr_0;

	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.352648:0.51766:1.99311;
		specparam tpd_XS_Q_negedge_f = 0.352648:0.51766:1.99311;
		specparam tpd_C_Q_posedge_r = 0.356251:0.500504:1.66416;
		specparam tpd_C_Q_posedge_f = 0.37144:0.496696:1.15424;
		specparam tsetup_D_C_XS_posedge_XS_posedge = 0.103375:0.108706:0.17251;
		specparam thold_D_C_XS_posedge_XS_posedge = -0.0464709:-0.06379:-0.12231;
		specparam tsetup_D_C_XS_negedge_XS_posedge = 0.103375:0.108706:0.17251;
		specparam thold_D_C_XS_negedge_XS_posedge = -0.0464709:-0.06379:-0.12231;
		specparam trecovery_XS_C_NTB_D_posedge_NTB_D_posedge = -0.021377:-0.043213:0.106476;
		specparam tremoval_XS_C_NTB_D_posedge_NTB_D_posedge = 0.0882861:0.108768:0.0835624;
		specparam tpw_XS_negedge = 0.203556:0.349169:2.72095;
		specparam tpw_C_posedge = 0.22403:0.330811:2.72095;
		specparam tpw_C_negedge = 0.22403:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& XS, posedge D &&& XS, 
			 tsetup_D_C_XS_posedge_XS_posedge, 
			 thold_D_C_XS_posedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XS, negedge D &&& XS, 
			 tsetup_D_C_XS_negedge_XS_posedge, 
			 thold_D_C_XS_negedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XS &&& ~D, posedge C &&& ~D, 
			 trecovery_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge C &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSQ 
`timescale 1ns/10ps
`celldefine
module DFFSQXL (Q, D, XS, C);
	output Q;
	input D, XS, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_s, xcr_0;

	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.299119:0.455834:1.9095;
		specparam tpd_XS_Q_negedge_f = 0.299119:0.455834:1.9095;
		specparam tpd_C_Q_posedge_r = 0.305861:0.441253:1.59371;
		specparam tpd_C_Q_posedge_f = 0.348052:0.466656:1.21249;
		specparam tsetup_D_C_XS_posedge_XS_posedge = 0.156548:0.147241:0.230363;
		specparam thold_D_C_XS_posedge_XS_posedge = -0.066179:-0.0839041:-0.150338;
		specparam tsetup_D_C_XS_negedge_XS_posedge = 0.156548:0.147241:0.230363;
		specparam thold_D_C_XS_negedge_XS_posedge = -0.066179:-0.0839041:-0.150338;
		specparam trecovery_XS_C_NTB_D_posedge_NTB_D_posedge = -0.0394578:-0.0650193:0.0571623;
		specparam tremoval_XS_C_NTB_D_posedge_NTB_D_posedge = 0.110757:0.134504:0.108656;
		specparam tpw_XS_negedge = 0.176439:0.330811:2.72095;
		specparam tpw_C_posedge = 0.167339:0.330811:2.72095;
		specparam tpw_C_negedge = 0.167339:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& XS, posedge D &&& XS, 
			 tsetup_D_C_XS_posedge_XS_posedge, 
			 thold_D_C_XS_posedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XS, negedge D &&& XS, 
			 tsetup_D_C_XS_negedge_XS_posedge, 
			 thold_D_C_XS_negedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XS &&& ~D, posedge C &&& ~D, 
			 trecovery_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge C &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSQX 
`timescale 1ns/10ps
`celldefine
module DFFSQXX1 (Q, XQ, D, XS, C);
	output Q, XQ;
	input D, XS, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_s;
	wire xcr_0;

	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.324792:0.483814:1.96538;
		specparam tpd_XS_Q_negedge_f = 0.324792:0.483814:1.96538;
		specparam tpd_C_Q_posedge_r = 0.31315:0.452864:1.6362;
		specparam tpd_C_Q_posedge_f = 0.353849:0.472895:1.13252;
		specparam tpd_XS_XQ_negedge_r = 0.139992:0.287007:1.25678;
		specparam tpd_XS_XQ_negedge_f = 0.139992:0.287007:1.25678;
		specparam tpd_C_XQ_posedge_r = 0.470861:0.608118:1.77104;
		specparam tpd_C_XQ_posedge_f = 0.398502:0.508075:1.1364;
		specparam tsetup_D_C_XS_posedge_XS_posedge = 0.161497:0.149523:0.22662;
		specparam thold_D_C_XS_posedge_XS_posedge = -0.0661164:-0.0826409:-0.151674;
		specparam tsetup_D_C_XS_negedge_XS_posedge = 0.161497:0.149523:0.22662;
		specparam thold_D_C_XS_negedge_XS_posedge = -0.0661164:-0.0826409:-0.151674;
		specparam trecovery_XS_C_NTB_D_posedge_NTB_D_posedge = -0.035485:-0.0611488:0.067311;
		specparam tremoval_XS_C_NTB_D_posedge_NTB_D_posedge = 0.105128:0.127503:0.104434;
		specparam tpw_XS_negedge = 0.205948:0.341301:2.72095;
		specparam tpw_C_posedge = 0.18051:0.330811:2.72095;
		specparam tpw_C_negedge = 0.18051:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& XS, posedge D &&& XS, 
			 tsetup_D_C_XS_posedge_XS_posedge, 
			 thold_D_C_XS_posedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XS, negedge D &&& XS, 
			 tsetup_D_C_XS_negedge_XS_posedge, 
			 thold_D_C_XS_negedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XS &&& ~D, posedge C &&& ~D, 
			 trecovery_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge C &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSQX 
`timescale 1ns/10ps
`celldefine
module DFFSQXX2 (Q, XQ, D, XS, C);
	output Q, XQ;
	input D, XS, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_s;
	wire xcr_0;

	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.381139:0.543141:2.03593;
		specparam tpd_XS_Q_negedge_f = 0.381139:0.543141:2.03593;
		specparam tpd_C_Q_posedge_r = 0.319591:0.462225:1.63703;
		specparam tpd_C_Q_posedge_f = 0.348223:0.470499:1.09398;
		specparam tpd_XS_XQ_negedge_r = 0.158558:0.309666:1.28282;
		specparam tpd_XS_XQ_negedge_f = 0.158558:0.309666:1.28282;
		specparam tpd_C_XQ_posedge_r = 0.501494:0.640596:1.78795;
		specparam tpd_C_XQ_posedge_f = 0.436957:0.547639:1.15361;
		specparam tsetup_D_C_XS_posedge_XS_posedge = 0.13154:0.128133:0.196078;
		specparam thold_D_C_XS_posedge_XS_posedge = -0.0542136:-0.0700388:-0.131905;
		specparam tsetup_D_C_XS_negedge_XS_posedge = 0.13154:0.128133:0.196078;
		specparam thold_D_C_XS_negedge_XS_posedge = -0.0542136:-0.0700388:-0.131905;
		specparam trecovery_XS_C_NTB_D_posedge_NTB_D_posedge = -0.0174578:-0.0395367:0.0985814;
		specparam tremoval_XS_C_NTB_D_posedge_NTB_D_posedge = 0.0834533:0.107112:0.0879981;
		specparam tpw_XS_negedge = 0.247865:0.385885:2.72095;
		specparam tpw_C_posedge = 0.200157:0.330811:2.72095;
		specparam tpw_C_negedge = 0.200157:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& XS, posedge D &&& XS, 
			 tsetup_D_C_XS_posedge_XS_posedge, 
			 thold_D_C_XS_posedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XS, negedge D &&& XS, 
			 tsetup_D_C_XS_negedge_XS_posedge, 
			 thold_D_C_XS_negedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XS &&& ~D, posedge C &&& ~D, 
			 trecovery_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge C &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSQX 
`timescale 1ns/10ps
`celldefine
module DFFSQXX4 (Q, XQ, D, XS, C);
	output Q, XQ;
	input D, XS, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_s;
	wire xcr_0;

	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.378176:0.539971:2.02615;
		specparam tpd_XS_Q_negedge_f = 0.378176:0.539971:2.02615;
		specparam tpd_C_Q_posedge_r = 0.3584:0.502686:1.68561;
		specparam tpd_C_Q_posedge_f = 0.372752:0.497094:1.14854;
		specparam tpd_XS_XQ_negedge_r = 0.14752:0.297521:1.28942;
		specparam tpd_XS_XQ_negedge_f = 0.14752:0.297521:1.28942;
		specparam tpd_C_XQ_posedge_r = 0.509901:0.646793:1.8051;
		specparam tpd_C_XQ_posedge_f = 0.468362:0.578758:1.22126;
		specparam tsetup_D_C_XS_posedge_XS_posedge = 0.103164:0.108902:0.171521;
		specparam thold_D_C_XS_posedge_XS_posedge = -0.0465477:-0.063961:-0.121147;
		specparam tsetup_D_C_XS_negedge_XS_posedge = 0.103164:0.108902:0.171521;
		specparam thold_D_C_XS_negedge_XS_posedge = -0.0465477:-0.063961:-0.121147;
		specparam trecovery_XS_C_NTB_D_posedge_NTB_D_posedge = -0.0228594:-0.0429008:0.108798;
		specparam tremoval_XS_C_NTB_D_posedge_NTB_D_posedge = 0.0882861:0.108768:0.0847151;
		specparam tpw_XS_negedge = 0.242438:0.372772:2.72095;
		specparam tpw_C_posedge = 0.241966:0.330811:2.72095;
		specparam tpw_C_negedge = 0.241966:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& XS, posedge D &&& XS, 
			 tsetup_D_C_XS_posedge_XS_posedge, 
			 thold_D_C_XS_posedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XS, negedge D &&& XS, 
			 tsetup_D_C_XS_negedge_XS_posedge, 
			 thold_D_C_XS_negedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XS &&& ~D, posedge C &&& ~D, 
			 trecovery_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge C &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSQX 
`timescale 1ns/10ps
`celldefine
module DFFSQXXL (Q, XQ, D, XS, C);
	output Q, XQ;
	input D, XS, C;
	reg notifier;
	wire delayed_D, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_s;
	wire xcr_0;

	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, delayed_D, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_XS_Q_negedge_r = 0.304458:0.462525:1.92975;
		specparam tpd_XS_Q_negedge_f = 0.304458:0.462525:1.92975;
		specparam tpd_C_Q_posedge_r = 0.30821:0.44438:1.60952;
		specparam tpd_C_Q_posedge_f = 0.348242:0.467391:1.21219;
		specparam tpd_XS_XQ_negedge_r = 0.137487:0.286198:1.33752;
		specparam tpd_XS_XQ_negedge_f = 0.137487:0.286198:1.33752;
		specparam tpd_C_XQ_posedge_r = 0.448098:0.584422:1.75328;
		specparam tpd_C_XQ_posedge_f = 0.379736:0.492169:1.224;
		specparam tsetup_D_C_XS_posedge_XS_posedge = 0.161153:0.150685:0.228655;
		specparam thold_D_C_XS_posedge_XS_posedge = -0.0681163:-0.0824027:-0.151651;
		specparam tsetup_D_C_XS_negedge_XS_posedge = 0.161153:0.150685:0.228655;
		specparam thold_D_C_XS_negedge_XS_posedge = -0.0681163:-0.0824027:-0.151651;
		specparam trecovery_XS_C_NTB_D_posedge_NTB_D_posedge = -0.0349664:-0.0595596:0.0629292;
		specparam tremoval_XS_C_NTB_D_posedge_NTB_D_posedge = 0.107461:0.129641:0.102192;
		specparam tpw_XS_negedge = 0.18568:0.330811:2.72095;
		specparam tpw_C_posedge = 0.171642:0.330811:2.72095;
		specparam tpw_C_negedge = 0.171642:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& XS, posedge D &&& XS, 
			 tsetup_D_C_XS_posedge_XS_posedge, 
			 thold_D_C_XS_posedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& XS, negedge D &&& XS, 
			 tsetup_D_C_XS_negedge_XS_posedge, 
			 thold_D_C_XS_negedge_XS_posedge, notifier,,, delayed_C, delayed_D);
		$recovery (posedge XS &&& ~D, posedge C &&& ~D, 
			 trecovery_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge C &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_C_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSRQ 
`timescale 1ns/10ps
`celldefine
module DFFSRQX1 (Q, D, XR, XS, C);
	output Q;
	input D, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_r, int_fwire_s;
	wire xcr_0;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.125296:0.251163:1.4322;
		specparam tpd_XR_Q_negedge_f = 0.118467:0.25567:1.17835;
		specparam tpd_XS_Q_negedge_r = 0.338698:0.5039:1.97581;
		specparam tpd_XS_Q_negedge_f = 0.338698:0.5039:1.97581;
		specparam tpd_C_Q_posedge_r = 0.352706:0.500023:1.69712;
		specparam tpd_C_Q_posedge_f = 0.369941:0.488278:1.12698;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.141838:0.132694:0.161064;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.0592962:-0.0719715:-0.0878618;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.141838:0.132694:0.161064;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.0592962:-0.0719715:-0.0878618;
		specparam trecovery_XR_C_adacond1_posedge_adacond1_posedge = -0.209339:-0.254351:0.0483951;
		specparam tremoval_XR_C_adacond1_posedge_adacond1_posedge = 0.301162:0.393993:0.846993;
		specparam tpw_XR_negedge = 0.343471:0.43047:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0137302:0.00513585:0.0180789;
		specparam thold_XR_XS_posedge_posedge = 0.0433338:0.0581851:0.131098;
		specparam trecovery_XS_C_adacond2_posedge_adacond2_posedge = -0.0426609:-0.0649763:0.0516036;
		specparam tremoval_XS_C_adacond2_posedge_adacond2_posedge = 0.129085:0.159156:0.143107;
		specparam tsetup_XS_XR_posedge_posedge = 0.0387431:0.0573508:0.177598;
		specparam thold_XS_XR_posedge_posedge = 0.0503677:0.0602465:0.0513411;
		specparam tpw_XS_negedge = 0.204446:0.338678:2.72095;
		specparam tpw_C_posedge = 0.202452:0.330811:2.72095;
		specparam tpw_C_negedge = 0.202452:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge C &&& adacond1, 
			 trecovery_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge C &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge C &&& adacond2, 
			 trecovery_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge C &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSRQ 
`timescale 1ns/10ps
`celldefine
module DFFSRQX2 (Q, D, XR, XS, C);
	output Q;
	input D, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_r, int_fwire_s;
	wire xcr_0;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.140812:0.274052:1.45748;
		specparam tpd_XR_Q_negedge_f = 0.137246:0.28313:1.23504;
		specparam tpd_XS_Q_negedge_r = 0.359567:0.529453:1.98382;
		specparam tpd_XS_Q_negedge_f = 0.359567:0.529453:1.98382;
		specparam tpd_C_Q_posedge_r = 0.358336:0.509944:1.692;
		specparam tpd_C_Q_posedge_f = 0.360998:0.484905:1.11785;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.11965:0.114422:0.141994;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.0498845:-0.0627461:-0.0855237;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.11965:0.114422:0.141994;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.0498845:-0.0627461:-0.0855237;
		specparam trecovery_XR_C_adacond1_posedge_adacond1_posedge = -0.197082:-0.238823:0.101086;
		specparam tremoval_XR_C_adacond1_posedge_adacond1_posedge = 0.296317:0.388196:0.857181;
		specparam tpw_XR_negedge = 0.348695:0.438337:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0175722:0.00551938:0.049485;
		specparam thold_XR_XS_posedge_posedge = 0.030631:0.039973:0.112514;
		specparam trecovery_XS_C_adacond2_posedge_adacond2_posedge = -0.0197775:-0.0416745:0.0895827;
		specparam tremoval_XS_C_adacond2_posedge_adacond2_posedge = 0.105121:0.129953:0.121769;
		specparam tsetup_XS_XR_posedge_posedge = 0.029586:0.0469526:0.175335;
		specparam thold_XS_XR_posedge_posedge = 0.0524681:0.0606506:0.0812654;
		specparam tpw_XS_negedge = 0.212135:0.346546:2.72095;
		specparam tpw_C_posedge = 0.213741:0.330811:2.72095;
		specparam tpw_C_negedge = 0.213741:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge C &&& adacond1, 
			 trecovery_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge C &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge C &&& adacond2, 
			 trecovery_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge C &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSRQ 
`timescale 1ns/10ps
`celldefine
module DFFSRQX4 (Q, D, XR, XS, C);
	output Q;
	input D, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_r, int_fwire_s;
	wire xcr_0;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.142698:0.275152:1.4578;
		specparam tpd_XR_Q_negedge_f = 0.13697:0.283327:1.23838;
		specparam tpd_XS_Q_negedge_r = 0.402774:0.573956:2.04529;
		specparam tpd_XS_Q_negedge_f = 0.402774:0.573956:2.04529;
		specparam tpd_C_Q_posedge_r = 0.41981:0.574046:1.75948;
		specparam tpd_C_Q_posedge_f = 0.403959:0.529793:1.16974;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.0934178:0.0978403:0.125584;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.0434046:-0.0545617:-0.0736478;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.0934178:0.0978403:0.125584;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.0434046:-0.0545617:-0.0736478;
		specparam trecovery_XR_C_adacond1_posedge_adacond1_posedge = -0.208178:-0.277577:-0.00588861;
		specparam tremoval_XR_C_adacond1_posedge_adacond1_posedge = 0.283424:0.379501:0.853428;
		specparam tpw_XR_negedge = 0.364428:0.45145:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0170734:0.0200938:0.108534;
		specparam thold_XR_XS_posedge_posedge = 0.0411993:0.0521995:0.135159;
		specparam trecovery_XS_C_adacond2_posedge_adacond2_posedge = -0.023584:-0.0485482:0.104502;
		specparam tremoval_XS_C_adacond2_posedge_adacond2_posedge = 0.106905:0.132674:0.113314;
		specparam tsetup_XS_XR_posedge_posedge = 0.0150878:0.0179009:0.169524;
		specparam thold_XS_XR_posedge_posedge = 0.0554021:0.0644052:0.14293;
		specparam tpw_XS_negedge = 0.237915:0.37015:2.72095;
		specparam tpw_C_posedge = 0.273323:0.330811:2.72095;
		specparam tpw_C_negedge = 0.273323:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge C &&& adacond1, 
			 trecovery_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge C &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge C &&& adacond2, 
			 trecovery_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge C &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSRQ 
`timescale 1ns/10ps
`celldefine
module DFFSRQXL (Q, D, XR, XS, C);
	output Q;
	input D, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_r, int_fwire_s;
	wire xcr_0;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.122939:0.244693:1.41697;
		specparam tpd_XR_Q_negedge_f = 0.116979:0.254321:1.25978;
		specparam tpd_XS_Q_negedge_r = 0.333007:0.494847:1.95931;
		specparam tpd_XS_Q_negedge_f = 0.333007:0.494847:1.95931;
		specparam tpd_C_Q_posedge_r = 0.348265:0.492258:1.68348;
		specparam tpd_C_Q_posedge_f = 0.36649:0.486779:1.22914;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.140828:0.13252:0.160921;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.0583345:-0.0712161:-0.0905417;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.140828:0.13252:0.160921;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.0583345:-0.0712161:-0.0905417;
		specparam trecovery_XR_C_adacond1_posedge_adacond1_posedge = -0.208329:-0.253051:0.027407;
		specparam tremoval_XR_C_adacond1_posedge_adacond1_posedge = 0.301162:0.393993:0.846993;
		specparam tpw_XR_negedge = 0.345699:0.43047:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.013614:0.00545676:0.00890597;
		specparam thold_XR_XS_posedge_posedge = 0.0524192:0.0645493:0.141016;
		specparam trecovery_XS_C_adacond2_posedge_adacond2_posedge = -0.0414403:-0.0652708:0.0520678;
		specparam tremoval_XS_C_adacond2_posedge_adacond2_posedge = 0.132603:0.159156:0.143107;
		specparam tsetup_XS_XR_posedge_posedge = 0.0386485:0.0624279:0.180058;
		specparam thold_XS_XR_posedge_posedge = 0.050172:0.0606131:0.0565628;
		specparam tpw_XS_negedge = 0.201502:0.336056:2.72095;
		specparam tpw_C_posedge = 0.195209:0.330811:2.72095;
		specparam tpw_C_negedge = 0.195209:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge C &&& adacond1, 
			 trecovery_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge C &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge C &&& adacond2, 
			 trecovery_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge C &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSRQX 
`timescale 1ns/10ps
`celldefine
module DFFSRQXX1 (Q, XQ, D, XR, XS, C);
	output Q, XQ;
	input D, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.125722:0.250861:1.42229;
		specparam tpd_XR_Q_negedge_f = 0.119094:0.255283:1.1742;
		specparam tpd_XS_Q_negedge_r = 0.3452:0.509793:1.97475;
		specparam tpd_XS_Q_negedge_f = 0.3452:0.509793:1.97475;
		specparam tpd_C_Q_posedge_r = 0.360415:0.506319:1.69687;
		specparam tpd_C_Q_posedge_f = 0.374567:0.492104:1.1273;
		specparam tpd_XR_XQ_negedge_r = 0.276998:0.45552:1.90352;
		specparam tpd_XR_XQ_negedge_f = 0.276998:0.45552:1.90352;
		specparam tpd_XS_XQ_negedge_r = 0.152285:0.303473:1.55975;
		specparam tpd_XS_XQ_negedge_f = 0.142612:0.2905:1.31734;
		specparam tpd_C_XQ_posedge_r = 0.494437:0.633843:1.81438;
		specparam tpd_C_XQ_posedge_f = 0.449082:0.562271:1.26139;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.138548:0.131286:0.159223;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.0593177:-0.0720652:-0.0910526;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.138548:0.131286:0.159223;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.0593177:-0.0720652:-0.0910526;
		specparam trecovery_XR_C_adacond1_posedge_adacond1_posedge = -0.213962:-0.258739:0.0317222;
		specparam tremoval_XR_C_adacond1_posedge_adacond1_posedge = 0.300008:0.394516:0.851668;
		specparam tpw_XR_negedge = 0.347218:0.433092:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0129522:0.00211392:-0.00623682;
		specparam thold_XR_XS_posedge_posedge = 0.0566421:0.0771004:0.155663;
		specparam trecovery_XS_C_adacond2_posedge_adacond2_posedge = -0.0426333:-0.0647179:0.0544198;
		specparam tremoval_XS_C_adacond2_posedge_adacond2_posedge = 0.129077:0.155167:0.140127;
		specparam tsetup_XS_XR_posedge_posedge = 0.0576273:0.0896705:0.242069;
		specparam thold_XS_XR_posedge_posedge = 0.0129522:0.00211392:-0.0998228;
		specparam tpw_XS_negedge = 0.217712:0.346546:2.72095;
		specparam tpw_C_posedge = 0.211647:0.330811:2.72095;
		specparam tpw_C_negedge = 0.211647:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge C &&& adacond1, 
			 trecovery_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge C &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge C &&& adacond2, 
			 trecovery_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge C &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSRQX 
`timescale 1ns/10ps
`celldefine
module DFFSRQXX2 (Q, XQ, D, XR, XS, C);
	output Q, XQ;
	input D, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.143546:0.278173:1.47426;
		specparam tpd_XR_Q_negedge_f = 0.139529:0.286067:1.24787;
		specparam tpd_XS_Q_negedge_r = 0.41276:0.581541:2.06433;
		specparam tpd_XS_Q_negedge_f = 0.41276:0.581541:2.06433;
		specparam tpd_C_Q_posedge_r = 0.369768:0.521907:1.71724;
		specparam tpd_C_Q_posedge_f = 0.369411:0.494045:1.13576;
		specparam tpd_XR_XQ_negedge_r = 0.335926:0.520204:2.01944;
		specparam tpd_XR_XQ_negedge_f = 0.335926:0.520204:2.01944;
		specparam tpd_XS_XQ_negedge_r = 0.170168:0.328618:1.6223;
		specparam tpd_XS_XQ_negedge_f = 0.158754:0.311532:1.33496;
		specparam tpd_C_XQ_posedge_r = 0.524865:0.668221:1.85963;
		specparam tpd_C_XQ_posedge_f = 0.493491:0.606839:1.27639;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.116384:0.113712:0.139517;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.0506895:-0.0625388:-0.0802374;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.116384:0.113712:0.139517;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.0506895:-0.0625388:-0.0802374;
		specparam trecovery_XR_C_adacond1_posedge_adacond1_posedge = -0.199241:-0.247237:0.0965627;
		specparam tremoval_XR_C_adacond1_posedge_adacond1_posedge = 0.292555:0.385928:0.852709;
		specparam tpw_XR_negedge = 0.350563:0.44096:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0165701:0.00517811:0.00730609;
		specparam thold_XR_XS_posedge_posedge = 0.0584976:0.0777524:0.156753;
		specparam trecovery_XS_C_adacond2_posedge_adacond2_posedge = -0.0200049:-0.0423289:0.0955577;
		specparam tremoval_XS_C_adacond2_posedge_adacond2_posedge = 0.102768:0.127464:0.117339;
		specparam tsetup_XS_XR_posedge_posedge = 0.0674183:0.100956:0.258687;
		specparam thold_XS_XR_posedge_posedge = 0.0135588:0.00517811:-0.0953804;
		specparam tpw_XS_negedge = 0.26099:0.393753:2.72095;
		specparam tpw_C_posedge = 0.239353:0.330811:2.72095;
		specparam tpw_C_negedge = 0.239353:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge C &&& adacond1, 
			 trecovery_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge C &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge C &&& adacond2, 
			 trecovery_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge C &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSRQX 
`timescale 1ns/10ps
`celldefine
module DFFSRQXX4 (Q, XQ, D, XR, XS, C);
	output Q, XQ;
	input D, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.145147:0.278799:1.47094;
		specparam tpd_XR_Q_negedge_f = 0.138718:0.28533:1.24942;
		specparam tpd_XS_Q_negedge_r = 0.432116:0.601969:2.08302;
		specparam tpd_XS_Q_negedge_f = 0.432116:0.601969:2.08302;
		specparam tpd_C_Q_posedge_r = 0.432832:0.587235:1.78615;
		specparam tpd_C_Q_posedge_f = 0.414608:0.540795:1.18975;
		specparam tpd_XR_XQ_negedge_r = 0.304465:0.478195:1.96462;
		specparam tpd_XR_XQ_negedge_f = 0.304465:0.478195:1.96462;
		specparam tpd_XS_XQ_negedge_r = 0.141556:0.28781:1.51975;
		specparam tpd_XS_XQ_negedge_f = 0.144277:0.291013:1.26544;
		specparam tpd_C_XQ_posedge_r = 0.558376:0.697802:1.88352;
		specparam tpd_C_XQ_posedge_f = 0.548027:0.655861:1.28568;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.0934178:0.0978403:0.12461;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.0427113:-0.0536975:-0.0723908;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.0934178:0.0978403:0.12461;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.0427113:-0.0536975:-0.0723908;
		specparam trecovery_XR_C_adacond1_posedge_adacond1_posedge = -0.207929:-0.281377:-0.0147286;
		specparam tremoval_XR_C_adacond1_posedge_adacond1_posedge = 0.281999:0.377224:0.849831;
		specparam tpw_XR_negedge = 0.368771:0.454073:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0155421:0.00356326:0.0489185;
		specparam thold_XR_XS_posedge_posedge = 0.0475878:0.0631751:0.14288;
		specparam trecovery_XS_C_adacond2_posedge_adacond2_posedge = -0.0239766:-0.0487467:0.11039;
		specparam tremoval_XS_C_adacond2_posedge_adacond2_posedge = 0.106877:0.128705:0.107342;
		specparam tsetup_XS_XR_posedge_posedge = 0.0475575:0.0718987:0.201232;
		specparam thold_XS_XR_posedge_posedge = 0.0144081:0.00365397:-0.0653837;
		specparam tpw_XS_negedge = 0.271157:0.388508:2.72095;
		specparam tpw_C_posedge = 0.302067:0.330811:2.72095;
		specparam tpw_C_negedge = 0.302067:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge C &&& adacond1, 
			 trecovery_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge C &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge C &&& adacond2, 
			 trecovery_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge C &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DFFSRQX 
`timescale 1ns/10ps
`celldefine
module DFFSRQXXL (Q, XQ, D, XR, XS, C);
	output Q, XQ;
	input D, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, delayed_D, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, delayed_D, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_XR_Q_negedge_r = 0.123823:0.2454:1.41335;
		specparam tpd_XR_Q_negedge_f = 0.117329:0.254093:1.2596;
		specparam tpd_XS_Q_negedge_r = 0.339994:0.501587:1.96264;
		specparam tpd_XS_Q_negedge_f = 0.339994:0.501587:1.96264;
		specparam tpd_C_Q_posedge_r = 0.356312:0.499401:1.68525;
		specparam tpd_C_Q_posedge_f = 0.370731:0.490722:1.23632;
		specparam tpd_XR_XQ_negedge_r = 0.258842:0.434224:1.85261;
		specparam tpd_XR_XQ_negedge_f = 0.258842:0.434224:1.85261;
		specparam tpd_XS_XQ_negedge_r = 0.150569:0.297937:1.53785;
		specparam tpd_XS_XQ_negedge_f = 0.138781:0.284598:1.33862;
		specparam tpd_C_XQ_posedge_r = 0.473542:0.611028:1.78343;
		specparam tpd_C_XQ_posedge_f = 0.429649:0.543014:1.28919;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.137468:0.128143:0.158643;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.0615309:-0.070747:-0.0912333;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.137468:0.128143:0.158643;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.0615309:-0.070747:-0.0912333;
		specparam trecovery_XR_C_adacond1_posedge_adacond1_posedge = -0.215054:-0.256778:0.011343;
		specparam tremoval_XR_C_adacond1_posedge_adacond1_posedge = 0.300008:0.394516:0.851668;
		specparam tpw_XR_negedge = 0.349478:0.433092:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0148088:0.00425485:-0.0110367;
		specparam thold_XR_XS_posedge_posedge = 0.0550612:0.0749595:0.146249;
		specparam trecovery_XS_C_adacond2_posedge_adacond2_posedge = -0.0414103:-0.0645228:0.0544713;
		specparam tremoval_XS_C_adacond2_posedge_adacond2_posedge = 0.13073:0.15649:0.13879;
		specparam tsetup_XS_XR_posedge_posedge = 0.0540601:0.0878582:0.225457;
		specparam thold_XS_XR_posedge_posedge = 0.0148088:0.00425485:-0.0870532;
		specparam tpw_XS_negedge = 0.205948:0.341301:2.72095;
		specparam tpw_C_posedge = 0.204571:0.330811:2.72095;
		specparam tpw_C_negedge = 0.204571:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:D)) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:D)) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge C &&& adacond1, 
			 trecovery_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge C &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_C_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge C &&& adacond2, 
			 trecovery_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge C &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_C_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNQ 
`timescale 1ns/10ps
`celldefine
module DLNQX1 (Q, D, XG);
	output Q;
	input D, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ;

	not (int_fwire_clk, delayed_XG);
	altos_latch (int_fwire_IQ, notifier, int_fwire_clk, delayed_D);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.174955:0.310786:1.5525;
		specparam tpd_D_Q_f = 0.225126:0.362146:1.37261;
		specparam tpd_XG_Q_negedge_r = 0.250162:0.421782:1.88175;
		specparam tpd_XG_Q_negedge_f = 0.337202:0.498307:1.50068;
		specparam tsetup_D_XG_posedge_posedge = 0.116202:0.143197:0.396675;
		specparam thold_D_XG_posedge_posedge = -0.082035:-0.106824:-0.275658;
		specparam tsetup_D_XG_negedge_posedge = 0.116202:0.143197:0.396675;
		specparam thold_D_XG_negedge_posedge = -0.082035:-0.106824:-0.275658;
		specparam tpw_XG_negedge = 0.231424:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG, posedge D, 
			 tsetup_D_XG_posedge_posedge, 
			 thold_D_XG_posedge_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG, negedge D, 
			 tsetup_D_XG_negedge_posedge, 
			 thold_D_XG_negedge_posedge, notifier,,, delayed_XG, delayed_D);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNQ 
`timescale 1ns/10ps
`celldefine
module DLNQX2 (Q, D, XG);
	output Q;
	input D, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ;

	not (int_fwire_clk, delayed_XG);
	altos_latch (int_fwire_IQ, notifier, int_fwire_clk, delayed_D);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.136718:0.270797:1.47348;
		specparam tpd_D_Q_f = 0.205205:0.380493:1.96744;
		specparam tpd_XG_Q_negedge_r = 0.202888:0.37702:1.81576;
		specparam tpd_XG_Q_negedge_f = 0.327968:0.530381:2.14693;
		specparam tsetup_D_XG_posedge_posedge = 0.0989476:0.123858:0.378941;
		specparam thold_D_XG_posedge_posedge = -0.0580176:-0.0768271:-0.225033;
		specparam tsetup_D_XG_negedge_posedge = 0.0989476:0.123858:0.378941;
		specparam thold_D_XG_negedge_posedge = -0.0580176:-0.0768271:-0.225033;
		specparam tpw_XG_negedge = 0.194117:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG, posedge D, 
			 tsetup_D_XG_posedge_posedge, 
			 thold_D_XG_posedge_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG, negedge D, 
			 tsetup_D_XG_negedge_posedge, 
			 thold_D_XG_negedge_posedge, notifier,,, delayed_XG, delayed_D);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNQ 
`timescale 1ns/10ps
`celldefine
module DLNQX4 (Q, D, XG);
	output Q;
	input D, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ;

	not (int_fwire_clk, delayed_XG);
	altos_latch (int_fwire_IQ, notifier, int_fwire_clk, delayed_D);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.140576:0.266688:1.45953;
		specparam tpd_D_Q_f = 0.184933:0.307416:1.23176;
		specparam tpd_XG_Q_negedge_r = 0.226647:0.396039:1.85348;
		specparam tpd_XG_Q_negedge_f = 0.360893:0.514117:1.48367;
		specparam tsetup_D_XG_posedge_posedge = 0.0893963:0.106783:0.330301;
		specparam thold_D_XG_posedge_posedge = -0.0577863:-0.0677151:-0.161931;
		specparam tsetup_D_XG_negedge_posedge = 0.0893963:0.106783:0.330301;
		specparam thold_D_XG_negedge_posedge = -0.0577863:-0.0677151:-0.161931;
		specparam tpw_XG_negedge = 0.222912:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG, posedge D, 
			 tsetup_D_XG_posedge_posedge, 
			 thold_D_XG_posedge_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG, negedge D, 
			 tsetup_D_XG_negedge_posedge, 
			 thold_D_XG_negedge_posedge, notifier,,, delayed_XG, delayed_D);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNQ 
`timescale 1ns/10ps
`celldefine
module DLNQXL (Q, D, XG);
	output Q;
	input D, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ;

	not (int_fwire_clk, delayed_XG);
	altos_latch (int_fwire_IQ, notifier, int_fwire_clk, delayed_D);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.174352:0.305116:1.53249;
		specparam tpd_D_Q_f = 0.211998:0.340761:1.32281;
		specparam tpd_XG_Q_negedge_r = 0.24565:0.412334:1.85985;
		specparam tpd_XG_Q_negedge_f = 0.320381:0.473093:1.46253;
		specparam tsetup_D_XG_posedge_posedge = 0.109107:0.140513:0.397708;
		specparam thold_D_XG_posedge_posedge = -0.0807189:-0.105787:-0.285342;
		specparam tsetup_D_XG_negedge_posedge = 0.109107:0.140513:0.397708;
		specparam thold_D_XG_negedge_posedge = -0.0807189:-0.105787:-0.285342;
		specparam tpw_XG_negedge = 0.212269:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG, posedge D, 
			 tsetup_D_XG_posedge_posedge, 
			 thold_D_XG_posedge_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG, negedge D, 
			 tsetup_D_XG_negedge_posedge, 
			 thold_D_XG_negedge_posedge, notifier,,, delayed_XG, delayed_D);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNQX 
`timescale 1ns/10ps
`celldefine
module DLNQXX1 (Q, XQ, D, XG);
	output Q, XQ;
	input D, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;

	not (int_fwire_clk, delayed_XG);
	altos_latch (int_fwire_IQ, notifier, int_fwire_clk, delayed_D);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.174804:0.308827:1.54026;
		specparam tpd_D_Q_f = 0.224573:0.360093:1.36492;
		specparam tpd_XG_Q_negedge_r = 0.250001:0.419871:1.86926;
		specparam tpd_XG_Q_negedge_f = 0.336646:0.496244:1.49353;
		specparam tpd_D_XQ_r = 0.334635:0.466016:1.87488;
		specparam tpd_D_XQ_f = 0.287838:0.396247:1.24142;
		specparam tpd_XG_XQ_negedge_r = 0.44651:0.601991:2.03766;
		specparam tpd_XG_XQ_negedge_f = 0.364519:0.508454:1.58089;
		specparam tsetup_D_XG_posedge_posedge = 0.12901:0.153966:0.400234;
		specparam thold_D_XG_posedge_posedge = -0.0825729:-0.108678:-0.274045;
		specparam tsetup_D_XG_negedge_posedge = 0.12901:0.153966:0.400234;
		specparam thold_D_XG_negedge_posedge = -0.0825729:-0.108678:-0.274045;
		specparam tpw_XG_negedge = 0.253822:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG, posedge D, 
			 tsetup_D_XG_posedge_posedge, 
			 thold_D_XG_posedge_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG, negedge D, 
			 tsetup_D_XG_negedge_posedge, 
			 thold_D_XG_negedge_posedge, notifier,,, delayed_XG, delayed_D);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNQX 
`timescale 1ns/10ps
`celldefine
module DLNQXX2 (Q, XQ, D, XG);
	output Q, XQ;
	input D, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;

	not (int_fwire_clk, delayed_XG);
	altos_latch (int_fwire_IQ, notifier, int_fwire_clk, delayed_D);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.147162:0.27889:1.49415;
		specparam tpd_D_Q_f = 0.188391:0.316934:1.2593;
		specparam tpd_XG_Q_negedge_r = 0.214967:0.385954:1.83651;
		specparam tpd_XG_Q_negedge_f = 0.311212:0.467235:1.43642;
		specparam tpd_D_XQ_r = 0.32276:0.455547:1.83633;
		specparam tpd_D_XQ_f = 0.307246:0.423315:1.21104;
		specparam tpd_XG_XQ_negedge_r = 0.445371:0.60554:2.04467;
		specparam tpd_XG_XQ_negedge_f = 0.378963:0.531669:1.55748;
		specparam tsetup_D_XG_posedge_posedge = 0.11725:0.13858:0.384986;
		specparam thold_D_XG_posedge_posedge = -0.0684901:-0.0949804:-0.257755;
		specparam tsetup_D_XG_negedge_posedge = 0.11725:0.13858:0.384986;
		specparam thold_D_XG_negedge_posedge = -0.0684901:-0.0949804:-0.257755;
		specparam tpw_XG_negedge = 0.221726:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG, posedge D, 
			 tsetup_D_XG_posedge_posedge, 
			 thold_D_XG_posedge_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG, negedge D, 
			 tsetup_D_XG_negedge_posedge, 
			 thold_D_XG_negedge_posedge, notifier,,, delayed_XG, delayed_D);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNQX 
`timescale 1ns/10ps
`celldefine
module DLNQXX4 (Q, XQ, D, XG);
	output Q, XQ;
	input D, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;

	not (int_fwire_clk, delayed_XG);
	altos_latch (int_fwire_IQ, notifier, int_fwire_clk, delayed_D);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.140274:0.265327:1.44667;
		specparam tpd_D_Q_f = 0.184316:0.305801:1.22269;
		specparam tpd_XG_Q_negedge_r = 0.226928:0.395427:1.84753;
		specparam tpd_XG_Q_negedge_f = 0.361487:0.513406:1.48254;
		specparam tpd_D_XQ_r = 0.369609:0.507957:1.87882;
		specparam tpd_D_XQ_f = 0.378912:0.502094:1.24215;
		specparam tpd_XG_XQ_negedge_r = 0.5464:0.71552:2.15993;
		specparam tpd_XG_XQ_negedge_f = 0.471621:0.635173:1.64259;
		specparam tsetup_D_XG_posedge_posedge = 0.103669:0.117476:0.337912;
		specparam thold_D_XG_posedge_posedge = -0.057263:-0.0694589:-0.169847;
		specparam tsetup_D_XG_negedge_posedge = 0.103669:0.117476:0.337912;
		specparam thold_D_XG_negedge_posedge = -0.057263:-0.0694589:-0.169847;
		specparam tpw_XG_negedge = 0.242682:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG, posedge D, 
			 tsetup_D_XG_posedge_posedge, 
			 thold_D_XG_posedge_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG, negedge D, 
			 tsetup_D_XG_negedge_posedge, 
			 thold_D_XG_negedge_posedge, notifier,,, delayed_XG, delayed_D);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNQX 
`timescale 1ns/10ps
`celldefine
module DLNQXXL (Q, XQ, D, XG);
	output Q, XQ;
	input D, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;

	not (int_fwire_clk, delayed_XG);
	altos_latch (int_fwire_IQ, notifier, int_fwire_clk, delayed_D);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.174271:0.304946:1.53946;
		specparam tpd_D_Q_f = 0.211691:0.340346:1.32737;
		specparam tpd_XG_Q_negedge_r = 0.245564:0.412159:1.86677;
		specparam tpd_XG_Q_negedge_f = 0.320086:0.47271:1.4672;
		specparam tpd_D_XQ_r = 0.301306:0.42975:1.8042;
		specparam tpd_D_XQ_f = 0.265345:0.36989:1.20608;
		specparam tpd_XG_XQ_negedge_r = 0.409493:0.561967:1.97974;
		specparam tpd_XG_XQ_negedge_f = 0.338028:0.477924:1.54851;
		specparam tsetup_D_XG_posedge_posedge = 0.114487:0.13956:0.3958;
		specparam thold_D_XG_posedge_posedge = -0.0809769:-0.106824:-0.285467;
		specparam tsetup_D_XG_negedge_posedge = 0.114487:0.13956:0.3958;
		specparam thold_D_XG_negedge_posedge = -0.0809769:-0.106824:-0.285467;
		specparam tpw_XG_negedge = 0.224606:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG, posedge D, 
			 tsetup_D_XG_posedge_posedge, 
			 thold_D_XG_posedge_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG, negedge D, 
			 tsetup_D_XG_negedge_posedge, 
			 thold_D_XG_negedge_posedge, notifier,,, delayed_XG, delayed_D);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNRQ 
`timescale 1ns/10ps
`celldefine
module DLNRQX1 (Q, D, XR, XG);
	output Q;
	input D, XR, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.265348:0.407628:1.68577;
		specparam tpd_D_Q_f = 0.24934:0.397496:1.47017;
		specparam tpd_XR_Q_negedge_r = 0.25602:0.410927:1.73332;
		specparam tpd_XR_Q_negedge_f = 0.180836:0.359751:1.5813;
		specparam tpd_XG_Q_negedge_r = 0.310279:0.499389:1.99266;
		specparam tpd_XG_Q_negedge_f = 0.355218:0.527363:1.61727;
		specparam tsetup_D_XG_XR_posedge_XR_posedge = 0.237529:0.247886:0.538489;
		specparam thold_D_XG_XR_posedge_XR_posedge = -0.164928:-0.183658:-0.419485;
		specparam tsetup_D_XG_XR_negedge_XR_posedge = 0.237529:0.247886:0.538489;
		specparam thold_D_XG_XR_negedge_XR_posedge = -0.164928:-0.183658:-0.419485;
		specparam trecovery_XR_XG_D_posedge_D_posedge = 0.230611:0.254309:0.537496;
		specparam tremoval_XR_XG_D_posedge_D_posedge = -0.152635:-0.18794:-0.437368;
		specparam tpw_XR_negedge = 0.180002:0.330811:2.72095;
		specparam tpw_XG_negedge = 0.290519:0.357037:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& XR, posedge D &&& XR, 
			 tsetup_D_XG_XR_posedge_XR_posedge, 
			 thold_D_XG_XR_posedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XR, negedge D &&& XR, 
			 tsetup_D_XG_XR_negedge_XR_posedge, 
			 thold_D_XG_XR_negedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XR &&& D, posedge XG &&& D, 
			 trecovery_XR_XG_D_posedge_D_posedge, notifier);
		$hold (posedge XG &&& D, posedge XR &&& D, 
			 tremoval_XR_XG_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNRQ 
`timescale 1ns/10ps
`celldefine
module DLNRQX2 (Q, D, XR, XG);
	output Q;
	input D, XR, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.213262:0.34361:1.55385;
		specparam tpd_D_Q_f = 0.218223:0.35551:1.33731;
		specparam tpd_XR_Q_negedge_r = 0.199545:0.34324:1.51893;
		specparam tpd_XR_Q_negedge_f = 0.25422:0.451789:1.78938;
		specparam tpd_XG_Q_negedge_r = 0.268174:0.449804:1.91416;
		specparam tpd_XG_Q_negedge_f = 0.342949:0.506221:1.49925;
		specparam tsetup_D_XG_XR_posedge_XR_posedge = 0.177318:0.18476:0.442162;
		specparam thold_D_XG_XR_posedge_XR_posedge = -0.123878:-0.138214:-0.30247;
		specparam tsetup_D_XG_XR_negedge_XR_posedge = 0.177318:0.18476:0.442162;
		specparam thold_D_XG_XR_negedge_XR_posedge = -0.123878:-0.138214:-0.30247;
		specparam trecovery_XR_XG_D_posedge_D_posedge = 0.165336:0.186173:0.348591;
		specparam tremoval_XR_XG_D_posedge_D_posedge = -0.110236:-0.137369:-0.230254;
		specparam tpw_XR_negedge = 0.256122:0.398998:2.72095;
		specparam tpw_XG_negedge = 0.238982:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& XR, posedge D &&& XR, 
			 tsetup_D_XG_XR_posedge_XR_posedge, 
			 thold_D_XG_XR_posedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XR, negedge D &&& XR, 
			 tsetup_D_XG_XR_negedge_XR_posedge, 
			 thold_D_XG_XR_negedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XR &&& D, posedge XG &&& D, 
			 trecovery_XR_XG_D_posedge_D_posedge, notifier);
		$hold (posedge XG &&& D, posedge XR &&& D, 
			 tremoval_XR_XG_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNRQ 
`timescale 1ns/10ps
`celldefine
module DLNRQX4 (Q, D, XR, XG);
	output Q;
	input D, XR, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.198137:0.328011:1.55059;
		specparam tpd_D_Q_f = 0.20553:0.338042:1.29023;
		specparam tpd_XR_Q_negedge_r = 0.182161:0.324791:1.46124;
		specparam tpd_XR_Q_negedge_f = 0.411445:0.64018:2.18371;
		specparam tpd_XG_Q_negedge_r = 0.232729:0.407849:1.813;
		specparam tpd_XG_Q_negedge_f = 0.32523:0.4804:1.41113;
		specparam tsetup_D_XG_XR_posedge_XR_posedge = 0.147746:0.156466:0.383435;
		specparam thold_D_XG_XR_posedge_XR_posedge = -0.113155:-0.121094:-0.242688;
		specparam tsetup_D_XG_XR_negedge_XR_posedge = 0.147746:0.156466:0.383435;
		specparam thold_D_XG_XR_negedge_XR_posedge = -0.113155:-0.121094:-0.242688;
		specparam trecovery_XR_XG_D_posedge_D_posedge = 0.130979:0.151896:0.259422;
		specparam tremoval_XR_XG_D_posedge_D_posedge = -0.0966076:-0.116348:-0.109099;
		specparam tpw_XR_negedge = 0.378517:0.524288:2.72095;
		specparam tpw_XG_negedge = 0.196369:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& XR, posedge D &&& XR, 
			 tsetup_D_XG_XR_posedge_XR_posedge, 
			 thold_D_XG_XR_posedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XR, negedge D &&& XR, 
			 tsetup_D_XG_XR_negedge_XR_posedge, 
			 thold_D_XG_XR_negedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XR &&& D, posedge XG &&& D, 
			 trecovery_XR_XG_D_posedge_D_posedge, notifier);
		$hold (posedge XG &&& D, posedge XR &&& D, 
			 tremoval_XR_XG_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNRQ 
`timescale 1ns/10ps
`celldefine
module DLNRQXL (Q, D, XR, XG);
	output Q;
	input D, XR, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.257732:0.39333:1.65792;
		specparam tpd_D_Q_f = 0.235822:0.376981:1.44182;
		specparam tpd_XR_Q_negedge_r = 0.248385:0.396546:1.7002;
		specparam tpd_XR_Q_negedge_f = 0.171265:0.342724:1.54813;
		specparam tpd_XG_Q_negedge_r = 0.303664:0.486587:1.97385;
		specparam tpd_XG_Q_negedge_f = 0.342727:0.508255:1.60212;
		specparam tsetup_D_XG_XR_posedge_XR_posedge = 0.215204:0.224735:0.518726;
		specparam thold_D_XG_XR_posedge_XR_posedge = -0.153645:-0.173409:-0.40184;
		specparam tsetup_D_XG_XR_negedge_XR_posedge = 0.215204:0.224735:0.518726;
		specparam thold_D_XG_XR_negedge_XR_posedge = -0.153645:-0.173409:-0.40184;
		specparam trecovery_XR_XG_D_posedge_D_posedge = 0.21004:0.23:0.503992;
		specparam tremoval_XR_XG_D_posedge_D_posedge = -0.143118:-0.176367:-0.415683;
		specparam tpw_XR_negedge = 0.165501:0.330811:2.72095;
		specparam tpw_XG_negedge = 0.268759:0.341301:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& XR, posedge D &&& XR, 
			 tsetup_D_XG_XR_posedge_XR_posedge, 
			 thold_D_XG_XR_posedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XR, negedge D &&& XR, 
			 tsetup_D_XG_XR_negedge_XR_posedge, 
			 thold_D_XG_XR_negedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XR &&& D, posedge XG &&& D, 
			 trecovery_XR_XG_D_posedge_D_posedge, notifier);
		$hold (posedge XG &&& D, posedge XR &&& D, 
			 tremoval_XR_XG_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNRQX 
`timescale 1ns/10ps
`celldefine
module DLNRQXX1 (Q, XQ, D, XR, XG);
	output Q, XQ;
	input D, XR, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.267188:0.407239:1.67703;
		specparam tpd_D_Q_f = 0.245814:0.389167:1.41002;
		specparam tpd_XR_Q_negedge_r = 0.257897:0.410462:1.72494;
		specparam tpd_XR_Q_negedge_f = 0.176261:0.349341:1.51591;
		specparam tpd_XG_Q_negedge_r = 0.314009:0.500853:1.98884;
		specparam tpd_XG_Q_negedge_f = 0.353727:0.521083:1.56243;
		specparam tpd_D_XQ_r = 0.364797:0.495041:1.8552;
		specparam tpd_D_XQ_f = 0.418996:0.515498:1.3326;
		specparam tpd_XR_XQ_negedge_r = 0.296615:0.455035:1.94382;
		specparam tpd_XR_XQ_negedge_f = 0.409932:0.519112:1.38599;
		specparam tpd_XG_XQ_negedge_r = 0.472585:0.627029:2.04151;
		specparam tpd_XG_XQ_negedge_f = 0.466843:0.610636:1.65666;
		specparam tsetup_D_XG_XR_posedge_XR_posedge = 0.258059:0.264808:0.543956;
		specparam thold_D_XG_XR_posedge_XR_posedge = -0.167993:-0.187908:-0.425683;
		specparam tsetup_D_XG_XR_negedge_XR_posedge = 0.258059:0.264808:0.543956;
		specparam thold_D_XG_XR_negedge_XR_posedge = -0.167993:-0.187908:-0.425683;
		specparam trecovery_XR_XG_D_posedge_D_posedge = 0.256285:0.271861:0.563437;
		specparam tremoval_XR_XG_D_posedge_D_posedge = -0.156849:-0.190117:-0.444442;
		specparam tpw_XR_negedge = 0.204616:0.341301:2.72095;
		specparam tpw_XG_negedge = 0.318433:0.375395:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& XR, posedge D &&& XR, 
			 tsetup_D_XG_XR_posedge_XR_posedge, 
			 thold_D_XG_XR_posedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XR, negedge D &&& XR, 
			 tsetup_D_XG_XR_negedge_XR_posedge, 
			 thold_D_XG_XR_negedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XR &&& D, posedge XG &&& D, 
			 trecovery_XR_XG_D_posedge_D_posedge, notifier);
		$hold (posedge XG &&& D, posedge XR &&& D, 
			 tremoval_XR_XG_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNRQX 
`timescale 1ns/10ps
`celldefine
module DLNRQXX2 (Q, XQ, D, XR, XG);
	output Q, XQ;
	input D, XR, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.213857:0.343803:1.55906;
		specparam tpd_D_Q_f = 0.218019:0.354876:1.33481;
		specparam tpd_XR_Q_negedge_r = 0.200144:0.344073:1.5239;
		specparam tpd_XR_Q_negedge_f = 0.253828:0.450385:1.78659;
		specparam tpd_XG_Q_negedge_r = 0.268854:0.450405:1.91991;
		specparam tpd_XG_Q_negedge_f = 0.34294:0.505794:1.49748;
		specparam tpd_D_XQ_r = 0.367238:0.502755:1.90031;
		specparam tpd_D_XQ_f = 0.397924:0.493052:1.17151;
		specparam tpd_XR_XQ_negedge_r = 0.447551:0.612548:2.28369;
		specparam tpd_XR_XQ_negedge_f = 0.384456:0.493171:1.14157;
		specparam tpd_XG_XQ_negedge_r = 0.492033:0.654067:2.09303;
		specparam tpd_XG_XQ_negedge_f = 0.454395:0.600889:1.53863;
		specparam tsetup_D_XG_XR_posedge_XR_posedge = 0.203605:0.206964:0.440724;
		specparam thold_D_XG_XR_posedge_XR_posedge = -0.126776:-0.138342:-0.30416;
		specparam tsetup_D_XG_XR_negedge_XR_posedge = 0.203605:0.206964:0.440724;
		specparam thold_D_XG_XR_negedge_XR_posedge = -0.126776:-0.138342:-0.30416;
		specparam trecovery_XR_XG_D_posedge_D_posedge = 0.194918:0.210948:0.353967;
		specparam tremoval_XR_XG_D_posedge_D_posedge = -0.112822:-0.137438:-0.228548;
		specparam tpw_XR_negedge = 0.299521:0.435715:2.72095;
		specparam tpw_XG_negedge = 0.271939:0.341301:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& XR, posedge D &&& XR, 
			 tsetup_D_XG_XR_posedge_XR_posedge, 
			 thold_D_XG_XR_posedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XR, negedge D &&& XR, 
			 tsetup_D_XG_XR_negedge_XR_posedge, 
			 thold_D_XG_XR_negedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XR &&& D, posedge XG &&& D, 
			 trecovery_XR_XG_D_posedge_D_posedge, notifier);
		$hold (posedge XG &&& D, posedge XR &&& D, 
			 tremoval_XR_XG_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNRQX 
`timescale 1ns/10ps
`celldefine
module DLNRQXX4 (Q, XQ, D, XR, XG);
	output Q, XQ;
	input D, XR, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.202:0.328877:1.52621;
		specparam tpd_D_Q_f = 0.206133:0.332448:1.21571;
		specparam tpd_XR_Q_negedge_r = 0.186021:0.325935:1.4389;
		specparam tpd_XR_Q_negedge_f = 0.410147:0.625695:2.10712;
		specparam tpd_XG_Q_negedge_r = 0.237022:0.408834:1.7889;
		specparam tpd_XG_Q_negedge_f = 0.326519:0.475597:1.33769;
		specparam tpd_D_XQ_r = 0.345896:0.477041:1.8612;
		specparam tpd_D_XQ_f = 0.370664:0.46507:1.15306;
		specparam tpd_XR_XQ_negedge_r = 0.659648:0.815516:2.59048;
		specparam tpd_XR_XQ_negedge_f = 0.354813:0.462196:1.07113;
		specparam tpd_XG_XQ_negedge_r = 0.466183:0.620158:2.01093;
		specparam tpd_XG_XQ_negedge_f = 0.407882:0.546282:1.42139;
		specparam tsetup_D_XG_XR_posedge_XR_posedge = 0.175388:0.17866:0.388224;
		specparam thold_D_XG_XR_posedge_XR_posedge = -0.115805:-0.127172:-0.246322;
		specparam tsetup_D_XG_XR_negedge_XR_posedge = 0.175388:0.17866:0.388224;
		specparam thold_D_XG_XR_negedge_XR_posedge = -0.115805:-0.127172:-0.246322;
		specparam trecovery_XR_XG_D_posedge_D_posedge = 0.163237:0.17802:0.263951;
		specparam tremoval_XR_XG_D_posedge_D_posedge = -0.0980041:-0.121811:-0.114342;
		specparam tpw_XR_negedge = 0.447731:0.581974:2.72095;
		specparam tpw_XG_negedge = 0.224496:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& XR, posedge D &&& XR, 
			 tsetup_D_XG_XR_posedge_XR_posedge, 
			 thold_D_XG_XR_posedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XR, negedge D &&& XR, 
			 tsetup_D_XG_XR_negedge_XR_posedge, 
			 thold_D_XG_XR_negedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XR &&& D, posedge XG &&& D, 
			 trecovery_XR_XG_D_posedge_D_posedge, notifier);
		$hold (posedge XG &&& D, posedge XR &&& D, 
			 tremoval_XR_XG_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNRQX 
`timescale 1ns/10ps
`celldefine
module DLNRQXXL (Q, XQ, D, XR, XG);
	output Q, XQ;
	input D, XR, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.258499:0.393253:1.66277;
		specparam tpd_D_Q_f = 0.236172:0.376566:1.44452;
		specparam tpd_XR_Q_negedge_r = 0.249146:0.39667:1.70524;
		specparam tpd_XR_Q_negedge_f = 0.171763:0.342234:1.55097;
		specparam tpd_XG_Q_negedge_r = 0.304788:0.486898:1.97956;
		specparam tpd_XG_Q_negedge_f = 0.343878:0.508709:1.60693;
		specparam tpd_D_XQ_r = 0.336825:0.467319:1.8307;
		specparam tpd_D_XQ_f = 0.380773:0.476573:1.30995;
		specparam tpd_XR_XQ_negedge_r = 0.274908:0.433082:1.91832;
		specparam tpd_XR_XQ_negedge_f = 0.371686:0.480179:1.35719;
		specparam tpd_XG_XQ_negedge_r = 0.444399:0.599619:2.02696;
		specparam tpd_XG_XQ_negedge_f = 0.428159:0.57158:1.64227;
		specparam tsetup_D_XG_XR_posedge_XR_posedge = 0.225754:0.235287:0.521489;
		specparam thold_D_XG_XR_posedge_XR_posedge = -0.154509:-0.172231:-0.402905;
		specparam tsetup_D_XG_XR_negedge_XR_posedge = 0.225754:0.235287:0.521489;
		specparam thold_D_XG_XR_negedge_XR_posedge = -0.154509:-0.172231:-0.402905;
		specparam trecovery_XR_XG_D_posedge_D_posedge = 0.222794:0.241593:0.514944;
		specparam tremoval_XR_XG_D_posedge_D_posedge = -0.142461:-0.176435:-0.416388;
		specparam tpw_XR_negedge = 0.181022:0.330811:2.72095;
		specparam tpw_XG_negedge = 0.285073:0.349169:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& XR, posedge D &&& XR, 
			 tsetup_D_XG_XR_posedge_XR_posedge, 
			 thold_D_XG_XR_posedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XR, negedge D &&& XR, 
			 tsetup_D_XG_XR_negedge_XR_posedge, 
			 thold_D_XG_XR_negedge_XR_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XR &&& D, posedge XG &&& D, 
			 trecovery_XR_XG_D_posedge_D_posedge, notifier);
		$hold (posedge XG &&& D, posedge XR &&& D, 
			 tremoval_XR_XG_D_posedge_D_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSQ 
`timescale 1ns/10ps
`celldefine
module DLNSQX1 (Q, D, XS, XG);
	output Q;
	input D, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.224975:0.37279:1.66119;
		specparam tpd_D_Q_f = 0.384763:0.542732:1.56628;
		specparam tpd_XS_Q_negedge_r = 0.251586:0.420323:1.88517;
		specparam tpd_XS_Q_negedge_f = 0.411835:0.565723:1.30373;
		specparam tpd_XG_Q_negedge_r = 0.304528:0.486138:1.96991;
		specparam tpd_XG_Q_negedge_f = 0.428263:0.615768:1.69843;
		specparam tsetup_D_XG_XS_posedge_XS_posedge = 0.20263:0.229235:0.518774;
		specparam thold_D_XG_XS_posedge_XS_posedge = -0.130213:-0.168229:-0.413493;
		specparam tsetup_D_XG_XS_negedge_XS_posedge = 0.20263:0.229235:0.518774;
		specparam thold_D_XG_XS_negedge_XS_posedge = -0.130213:-0.168229:-0.413493;
		specparam trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge = 0.301321:0.296325:0.281532;
		specparam tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge = -0.23205:-0.227542:-0.223023;
		specparam tpw_XS_negedge = 0.202704:0.330811:2.72095;
		specparam tpw_XG_negedge = 0.323444:0.354414:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& XS, posedge D &&& XS, 
			 tsetup_D_XG_XS_posedge_XS_posedge, 
			 thold_D_XG_XS_posedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XS, negedge D &&& XS, 
			 tsetup_D_XG_XS_negedge_XS_posedge, 
			 thold_D_XG_XS_negedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XS &&& ~D, posedge XG &&& ~D, 
			 trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge XG &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSQ 
`timescale 1ns/10ps
`celldefine
module DLNSQX2 (Q, D, XS, XG);
	output Q;
	input D, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.175656:0.315497:1.5493;
		specparam tpd_D_Q_f = 0.316693:0.462452:1.42894;
		specparam tpd_XS_Q_negedge_r = 0.345105:0.526849:2.04013;
		specparam tpd_XS_Q_negedge_f = 0.347795:0.496492:1.19882;
		specparam tpd_XG_Q_negedge_r = 0.264364:0.443849:1.93165;
		specparam tpd_XG_Q_negedge_f = 0.391447:0.570567:1.62107;
		specparam tsetup_D_XG_XS_posedge_XS_posedge = 0.149119:0.168711:0.422338;
		specparam thold_D_XG_XS_posedge_XS_posedge = -0.0939881:-0.120844:-0.289149;
		specparam tsetup_D_XG_XS_negedge_XS_posedge = 0.149119:0.168711:0.422338;
		specparam thold_D_XG_XS_negedge_XS_posedge = -0.0939881:-0.120844:-0.289149;
		specparam trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge = 0.214778:0.207407:0.185312;
		specparam tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge = -0.157817:-0.155323:-0.137575;
		specparam tpw_XS_negedge = 0.26736:0.357037:2.72095;
		specparam tpw_XG_negedge = 0.266835:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& XS, posedge D &&& XS, 
			 tsetup_D_XG_XS_posedge_XS_posedge, 
			 thold_D_XG_XS_posedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XS, negedge D &&& XS, 
			 tsetup_D_XG_XS_negedge_XS_posedge, 
			 thold_D_XG_XS_negedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XS &&& ~D, posedge XG &&& ~D, 
			 trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge XG &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSQ 
`timescale 1ns/10ps
`celldefine
module DLNSQX4 (Q, D, XS, XG);
	output Q;
	input D, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.165101:0.300692:1.50379;
		specparam tpd_D_Q_f = 0.309312:0.446356:1.36668;
		specparam tpd_XS_Q_negedge_r = 0.517081:0.712936:2.22494;
		specparam tpd_XS_Q_negedge_f = 0.347379:0.496182:1.19467;
		specparam tpd_XG_Q_negedge_r = 0.221683:0.396142:1.79559;
		specparam tpd_XG_Q_negedge_f = 0.35866:0.525672:1.46769;
		specparam tsetup_D_XG_XS_posedge_XS_posedge = 0.1191:0.143515:0.357185;
		specparam thold_D_XG_XS_posedge_XS_posedge = -0.0859924:-0.107197:-0.218352;
		specparam tsetup_D_XG_XS_negedge_XS_posedge = 0.1191:0.143515:0.357185;
		specparam thold_D_XG_XS_negedge_XS_posedge = -0.0859924:-0.107197:-0.218352;
		specparam trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge = 0.23343:0.230315:0.217533;
		specparam tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge = -0.164595:-0.169711:-0.159202;
		specparam tpw_XS_negedge = 0.345654:0.414734:2.72095;
		specparam tpw_XG_negedge = 0.246347:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& XS, posedge D &&& XS, 
			 tsetup_D_XG_XS_posedge_XS_posedge, 
			 thold_D_XG_XS_posedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XS, negedge D &&& XS, 
			 tsetup_D_XG_XS_negedge_XS_posedge, 
			 thold_D_XG_XS_negedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XS &&& ~D, posedge XG &&& ~D, 
			 trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge XG &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSQ 
`timescale 1ns/10ps
`celldefine
module DLNSQXL (Q, D, XS, XG);
	output Q;
	input D, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.220678:0.364693:1.65993;
		specparam tpd_D_Q_f = 0.358341:0.509275:1.52544;
		specparam tpd_XS_Q_negedge_r = 0.251093:0.417272:1.89811;
		specparam tpd_XS_Q_negedge_f = 0.385245:0.532201:1.26887;
		specparam tpd_XG_Q_negedge_r = 0.29981:0.477938:1.97414;
		specparam tpd_XG_Q_negedge_f = 0.402142:0.582655:1.66411;
		specparam tsetup_D_XG_XS_posedge_XS_posedge = 0.18272:0.213816:0.502696;
		specparam thold_D_XG_XS_posedge_XS_posedge = -0.122967:-0.157351:-0.401331;
		specparam tsetup_D_XG_XS_negedge_XS_posedge = 0.18272:0.213816:0.502696;
		specparam thold_D_XG_XS_negedge_XS_posedge = -0.122967:-0.157351:-0.401331;
		specparam trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge = 0.271242:0.266543:0.25307;
		specparam tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge = -0.20879:-0.204188:-0.19592;
		specparam tpw_XS_negedge = 0.189593:0.330811:2.72095;
		specparam tpw_XG_negedge = 0.295183:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& XS, posedge D &&& XS, 
			 tsetup_D_XG_XS_posedge_XS_posedge, 
			 thold_D_XG_XS_posedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XS, negedge D &&& XS, 
			 tsetup_D_XG_XS_negedge_XS_posedge, 
			 thold_D_XG_XS_negedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XS &&& ~D, posedge XG &&& ~D, 
			 trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge XG &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSQX 
`timescale 1ns/10ps
`celldefine
module DLNSQXX1 (Q, XQ, D, XS, XG);
	output Q, XQ;
	input D, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.218729:0.364007:1.63448;
		specparam tpd_D_Q_f = 0.375322:0.528337:1.54638;
		specparam tpd_XS_Q_negedge_r = 0.247796:0.414721:1.86855;
		specparam tpd_XS_Q_negedge_f = 0.40231:0.551295:1.28566;
		specparam tpd_XG_Q_negedge_r = 0.298057:0.477258:1.94577;
		specparam tpd_XG_Q_negedge_f = 0.418837:0.601488:1.68063;
		specparam tpd_D_XQ_r = 0.508366:0.635093:1.97991;
		specparam tpd_D_XQ_f = 0.364128:0.47816:1.35563;
		specparam tpd_XS_XQ_negedge_r = 0.534831:0.657762:1.75118;
		specparam tpd_XS_XQ_negedge_f = 0.376036:0.525431:1.6016;
		specparam tpd_XG_XQ_negedge_r = 0.551736:0.708188:2.14743;
		specparam tpd_XG_XQ_negedge_f = 0.444932:0.593208:1.67493;
		specparam tsetup_D_XG_XS_posedge_XS_posedge = 0.205621:0.228782:0.509867;
		specparam thold_D_XG_XS_posedge_XS_posedge = -0.124412:-0.161927:-0.403736;
		specparam tsetup_D_XG_XS_negedge_XS_posedge = 0.205621:0.228782:0.509867;
		specparam thold_D_XG_XS_negedge_XS_posedge = -0.124412:-0.161927:-0.403736;
		specparam trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge = 0.350246:0.341963:0.322952;
		specparam tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge = -0.22538:-0.221753:-0.214196;
		specparam tpw_XS_negedge = 0.202704:0.330811:2.72095;
		specparam tpw_XG_negedge = 0.375676:0.401621:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& XS, posedge D &&& XS, 
			 tsetup_D_XG_XS_posedge_XS_posedge, 
			 thold_D_XG_XS_posedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XS, negedge D &&& XS, 
			 tsetup_D_XG_XS_negedge_XS_posedge, 
			 thold_D_XG_XS_negedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XS &&& ~D, posedge XG &&& ~D, 
			 trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge XG &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSQX 
`timescale 1ns/10ps
`celldefine
module DLNSQXX2 (Q, XQ, D, XS, XG);
	output Q, XQ;
	input D, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.174815:0.313364:1.55011;
		specparam tpd_D_Q_f = 0.311234:0.452158:1.39519;
		specparam tpd_XS_Q_negedge_r = 0.344011:0.524419:2.04331;
		specparam tpd_XS_Q_negedge_f = 0.342376:0.486382:1.16709;
		specparam tpd_XG_Q_negedge_r = 0.262755:0.441512:1.93382;
		specparam tpd_XG_Q_negedge_f = 0.386016:0.560368:1.58993;
		specparam tpd_D_XQ_r = 0.476023:0.604312:1.94218;
		specparam tpd_D_XQ_f = 0.344685:0.45773:1.19951;
		specparam tpd_XS_XQ_negedge_r = 0.506719:0.638117:1.7434;
		specparam tpd_XS_XQ_negedge_f = 0.521731:0.66976:1.69672;
		specparam tpd_XG_XQ_negedge_r = 0.55067:0.712258:2.1677;
		specparam tpd_XG_XQ_negedge_f = 0.439024:0.588319:1.58701;
		specparam tsetup_D_XG_XS_posedge_XS_posedge = 0.161356:0.179677:0.420391;
		specparam thold_D_XG_XS_posedge_XS_posedge = -0.0934597:-0.118556:-0.288217;
		specparam tsetup_D_XG_XS_negedge_XS_posedge = 0.161356:0.179677:0.420391;
		specparam thold_D_XG_XS_negedge_XS_posedge = -0.0934597:-0.118556:-0.288217;
		specparam trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge = 0.270622:0.260428:0.228881;
		specparam tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge = -0.155498:-0.152557:-0.134222;
		specparam tpw_XS_negedge = 0.275535:0.362282:2.72095;
		specparam tpw_XG_negedge = 0.322197:0.354414:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& XS, posedge D &&& XS, 
			 tsetup_D_XG_XS_posedge_XS_posedge, 
			 thold_D_XG_XS_posedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XS, negedge D &&& XS, 
			 tsetup_D_XG_XS_negedge_XS_posedge, 
			 thold_D_XG_XS_negedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XS &&& ~D, posedge XG &&& ~D, 
			 trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge XG &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSQX 
`timescale 1ns/10ps
`celldefine
module DLNSQXX4 (Q, XQ, D, XS, XG);
	output Q, XQ;
	input D, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.164822:0.301177:1.5175;
		specparam tpd_D_Q_f = 0.312705:0.453856:1.42451;
		specparam tpd_XS_Q_negedge_r = 0.519428:0.716826:2.2504;
		specparam tpd_XS_Q_negedge_f = 0.352806:0.506264:1.25665;
		specparam tpd_XG_Q_negedge_r = 0.221049:0.396506:1.81015;
		specparam tpd_XG_Q_negedge_f = 0.362144:0.5332:1.52392;
		specparam tpd_D_XQ_r = 0.470296:0.594083:1.91812;
		specparam tpd_D_XQ_f = 0.324854:0.434796:1.14899;
		specparam tpd_XS_XQ_negedge_r = 0.510138:0.646265:1.77871;
		specparam tpd_XS_XQ_negedge_f = 0.72104:0.859651:1.87744;
		specparam tpd_XG_XQ_negedge_r = 0.519718:0.673049:2.04903;
		specparam tpd_XG_XQ_negedge_f = 0.389357:0.532102:1.44484;
		specparam tsetup_D_XG_XS_posedge_XS_posedge = 0.138516:0.155584:0.355174;
		specparam thold_D_XG_XS_posedge_XS_posedge = -0.082272:-0.10741:-0.216169;
		specparam tsetup_D_XG_XS_negedge_XS_posedge = 0.138516:0.155584:0.355174;
		specparam thold_D_XG_XS_negedge_XS_posedge = -0.082272:-0.10741:-0.216169;
		specparam trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge = 0.267968:0.264158:0.251113;
		specparam tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge = -0.172017:-0.175106:-0.165474;
		specparam tpw_XS_negedge = 0.382586:0.44096:2.72095;
		specparam tpw_XG_negedge = 0.283192:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& XS, posedge D &&& XS, 
			 tsetup_D_XG_XS_posedge_XS_posedge, 
			 thold_D_XG_XS_posedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XS, negedge D &&& XS, 
			 tsetup_D_XG_XS_negedge_XS_posedge, 
			 thold_D_XG_XS_negedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XS &&& ~D, posedge XG &&& ~D, 
			 trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge XG &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSQX 
`timescale 1ns/10ps
`celldefine
module DLNSQXXL (Q, XQ, D, XS, XG);
	output Q, XQ;
	input D, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.215939:0.35624:1.62657;
		specparam tpd_D_Q_f = 0.34857:0.491928:1.47924;
		specparam tpd_XS_Q_negedge_r = 0.24855:0.412065:1.87426;
		specparam tpd_XS_Q_negedge_f = 0.375436:0.514804:1.22447;
		specparam tpd_XG_Q_negedge_r = 0.29484:0.469226:1.9458;
		specparam tpd_XG_Q_negedge_f = 0.392361:0.565422:1.6204;
		specparam tpd_D_XQ_r = 0.464441:0.590479:1.91795;
		specparam tpd_D_XQ_f = 0.3275:0.437212:1.29196;
		specparam tpd_XS_XQ_negedge_r = 0.490813:0.613011:1.69518;
		specparam tpd_XS_XQ_negedge_f = 0.349502:0.493329:1.55881;
		specparam tpd_XG_XQ_negedge_r = 0.508061:0.663791:2.0923;
		specparam tpd_XG_XQ_negedge_f = 0.407742:0.551911:1.62371;
		specparam tsetup_D_XG_XS_posedge_XS_posedge = 0.182837:0.206967:0.494431;
		specparam thold_D_XG_XS_posedge_XS_posedge = -0.116332:-0.155111:-0.389559;
		specparam tsetup_D_XG_XS_negedge_XS_posedge = 0.182837:0.206967:0.494431;
		specparam thold_D_XG_XS_negedge_XS_posedge = -0.116332:-0.155111:-0.389559;
		specparam trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge = 0.30615:0.295748:0.276442;
		specparam tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge = -0.197228:-0.196973:-0.187503;
		specparam tpw_XS_negedge = 0.187272:0.330811:2.72095;
		specparam tpw_XG_negedge = 0.329628:0.357037:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& XS, posedge D &&& XS, 
			 tsetup_D_XG_XS_posedge_XS_posedge, 
			 thold_D_XG_XS_posedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& XS, negedge D &&& XS, 
			 tsetup_D_XG_XS_negedge_XS_posedge, 
			 thold_D_XG_XS_negedge_XS_posedge, notifier,,, delayed_XG, delayed_D);
		$recovery (posedge XS &&& ~D, posedge XG &&& ~D, 
			 trecovery_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$hold (posedge XG &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_XG_NTB_D_posedge_NTB_D_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSRQ 
`timescale 1ns/10ps
`celldefine
module DLNSRQX1 (Q, D, XR, XS, XG);
	output Q;
	input D, XR, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_latch_sr_1 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_D_Q_r = 0.297824:0.439661:1.67929;
		specparam tpd_D_Q_f = 0.427047:0.603077:1.68255;
		specparam tpd_XR_Q_negedge_r = 0.289028:0.443359:1.75706;
		specparam tpd_XR_Q_negedge_f = 0.3121:0.485915:1.70925;
		specparam tpd_XS_Q_negedge_r = 0.286777:0.460569:1.96438;
		specparam tpd_XS_Q_negedge_f = 0.446879:0.615684:1.40602;
		specparam tpd_XG_Q_negedge_r = 0.360388:0.549962:2.03205;
		specparam tpd_XG_Q_negedge_f = 0.473152:0.678637:1.81814;
		specparam tsetup_D_XG_adacond0_posedge_adacond0_posedge = 0.269652:0.280733:0.575358;
		specparam thold_D_XG_adacond0_posedge_adacond0_posedge = -0.195476:-0.220499:-0.451468;
		specparam tsetup_D_XG_adacond0_negedge_adacond0_posedge = 0.269652:0.280733:0.575358;
		specparam thold_D_XG_adacond0_negedge_adacond0_posedge = -0.195476:-0.220499:-0.451468;
		specparam trecovery_XR_XG_adacond1_posedge_adacond1_posedge = 0.263562:0.285772:0.59771;
		specparam tremoval_XR_XG_adacond1_posedge_adacond1_posedge = -0.187814:-0.223485:-0.505941;
		specparam tpw_XR_negedge = 0.302114:0.39113:2.72095;
		specparam trecovery_XS_XG_adacond2_posedge_adacond2_posedge = 0.36051:0.352049:0.331539;
		specparam tremoval_XS_XG_adacond2_posedge_adacond2_posedge = -0.248236:-0.242279:-0.235513;
		specparam tsetup_XS_XR_XG_posedge_XG_posedge = 0.332938:0.415919:1.19752;
		specparam thold_XS_XR_XG_posedge_XG_posedge = -0.243575:-0.344204:-0.680956;
		specparam tpw_XS_negedge = 0.236431:0.341301:2.72095;
		specparam tpw_XG_negedge = 0.401748:0.425224:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XG_adacond0_posedge_adacond0_posedge, 
			 thold_D_XG_adacond0_posedge_adacond0_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XG_adacond0_negedge_adacond0_posedge, 
			 thold_D_XG_adacond0_negedge_adacond0_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XR &&& XG, posedge XS &&& XG, 
			 tsetup_XS_XR_XG_posedge_XG_posedge, 
			 thold_XS_XR_XG_posedge_XG_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge XG &&& adacond1, 
			 trecovery_XR_XG_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge XG &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XG_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge XG &&& adacond2, 
			 trecovery_XS_XG_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge XG &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XG_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSRQ 
`timescale 1ns/10ps
`celldefine
module DLNSRQXL (Q, D, XR, XS, XG);
	output Q;
	input D, XR, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_latch_sr_1 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_D_Q_r = 0.340557:0.479607:1.73049;
		specparam tpd_D_Q_f = 0.426428:0.600616:1.68173;
		specparam tpd_XR_Q_negedge_r = 0.332105:0.483798:1.83489;
		specparam tpd_XR_Q_negedge_f = 0.266896:0.424114:1.55819;
		specparam tpd_XS_Q_negedge_r = 0.271821:0.439098:1.94064;
		specparam tpd_XS_Q_negedge_f = 0.443041:0.605685:1.38796;
		specparam tpd_XG_Q_negedge_r = 0.395508:0.583822:2.06983;
		specparam tpd_XG_Q_negedge_f = 0.469992:0.67:1.79729;
		specparam tsetup_D_XG_adacond0_posedge_adacond0_posedge = 0.298652:0.307151:0.600944;
		specparam thold_D_XG_adacond0_posedge_adacond0_posedge = -0.228668:-0.248013:-0.487929;
		specparam tsetup_D_XG_adacond0_negedge_adacond0_posedge = 0.298652:0.307151:0.600944;
		specparam thold_D_XG_adacond0_negedge_adacond0_posedge = -0.228668:-0.248013:-0.487929;
		specparam trecovery_XR_XG_adacond1_posedge_adacond1_posedge = 0.292278:0.31437:0.651615;
		specparam tremoval_XR_XG_adacond1_posedge_adacond1_posedge = -0.220043:-0.252744:-0.571685;
		specparam tpw_XR_negedge = 0.260906:0.346546:2.72095;
		specparam trecovery_XS_XG_adacond2_posedge_adacond2_posedge = 0.358458:0.35032:0.331465;
		specparam tremoval_XS_XG_adacond2_posedge_adacond2_posedge = -0.238733:-0.239525:-0.231229;
		specparam tsetup_XS_XR_XG_posedge_XG_posedge = 0.288615:0.373475:1.12879;
		specparam thold_XS_XR_XG_posedge_XG_posedge = -0.209618:-0.306627:-0.615574;
		specparam tpw_XS_negedge = 0.218496:0.333433:2.72095;
		specparam tpw_XG_negedge = 0.404148:0.427847:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		$setuphold (posedge XG &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XG_adacond0_posedge_adacond0_posedge, 
			 thold_D_XG_adacond0_posedge_adacond0_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XG_adacond0_negedge_adacond0_posedge, 
			 thold_D_XG_adacond0_negedge_adacond0_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XR &&& XG, posedge XS &&& XG, 
			 tsetup_XS_XR_XG_posedge_XG_posedge, 
			 thold_XS_XR_XG_posedge_XG_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge XG &&& adacond1, 
			 trecovery_XR_XG_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge XG &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XG_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge XG &&& adacond2, 
			 trecovery_XS_XG_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge XG &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XG_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSRQX 
`timescale 1ns/10ps
`celldefine
module DLNSRQXX1 (Q, XQ, D, XR, XS, XG);
	output Q, XQ;
	input D, XR, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_latch_sr_1 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_D_Q_r = 0.29523:0.438431:1.69321;
		specparam tpd_D_Q_f = 0.425377:0.604105:1.70527;
		specparam tpd_XR_Q_negedge_r = 0.286406:0.442021:1.77147;
		specparam tpd_XR_Q_negedge_f = 0.309686:0.485814:1.73046;
		specparam tpd_XS_Q_negedge_r = 0.28643:0.461287:1.98331;
		specparam tpd_XS_Q_negedge_f = 0.445974:0.617518:1.43247;
		specparam tpd_XG_Q_negedge_r = 0.357706:0.548667:2.04776;
		specparam tpd_XG_Q_negedge_f = 0.471491:0.679569:1.83973;
		specparam tpd_D_XQ_r = 0.585493:0.719983:2.07704;
		specparam tpd_D_XQ_f = 0.460912:0.564932:1.41504;
		specparam tpd_XR_XQ_negedge_r = 0.463355:0.603083:2.05939;
		specparam tpd_XR_XQ_negedge_f = 0.452299:0.569004:1.49758;
		specparam tpd_XS_XQ_negedge_r = 0.600869:0.73306:1.83551;
		specparam tpd_XS_XQ_negedge_f = 0.42715:0.581234:1.72314;
		specparam tpd_XG_XQ_negedge_r = 0.631512:0.795206:2.24127;
		specparam tpd_XG_XQ_negedge_f = 0.52425:0.676975:1.77676;
		specparam tsetup_D_XG_adacond0_posedge_adacond0_posedge = 0.286209:0.296076:0.570433;
		specparam thold_D_XG_adacond0_posedge_adacond0_posedge = -0.194601:-0.218013:-0.445546;
		specparam tsetup_D_XG_adacond0_negedge_adacond0_posedge = 0.286209:0.296076:0.570433;
		specparam thold_D_XG_adacond0_negedge_adacond0_posedge = -0.194601:-0.218013:-0.445546;
		specparam trecovery_XR_XG_adacond1_posedge_adacond1_posedge = 0.283891:0.30351:0.614101;
		specparam tremoval_XR_XG_adacond1_posedge_adacond1_posedge = -0.184808:-0.221058:-0.499941;
		specparam tpw_XR_negedge = 0.337794:0.419979:2.72095;
		specparam trecovery_XS_XG_adacond2_posedge_adacond2_posedge = 0.397243:0.390853:0.36484;
		specparam tremoval_XS_XG_adacond2_posedge_adacond2_posedge = -0.247741:-0.242692:-0.240556;
		specparam tsetup_XS_XR_XG_posedge_XG_posedge = 0.365864:0.444639:1.19334;
		specparam thold_XS_XR_XG_posedge_XG_posedge = -0.243978:-0.344158:-0.6814;
		specparam tpw_XS_negedge = 0.248143:0.349169:2.72095;
		specparam tpw_XG_negedge = 0.445348:0.467186:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XG_adacond0_posedge_adacond0_posedge, 
			 thold_D_XG_adacond0_posedge_adacond0_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XG_adacond0_negedge_adacond0_posedge, 
			 thold_D_XG_adacond0_negedge_adacond0_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XR &&& XG, posedge XS &&& XG, 
			 tsetup_XS_XR_XG_posedge_XG_posedge, 
			 thold_XS_XR_XG_posedge_XG_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge XG &&& adacond1, 
			 trecovery_XR_XG_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge XG &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XG_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge XG &&& adacond2, 
			 trecovery_XS_XG_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge XG &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XG_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLNSRQX 
`timescale 1ns/10ps
`celldefine
module DLNSRQXXL (Q, XQ, D, XR, XS, XG);
	output Q, XQ;
	input D, XR, XS, XG;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_XG;

	// Function
	wire int_fwire_clk, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s;

	not (int_fwire_clk, delayed_XG);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_latch_sr_1 (int_fwire_IQ, notifier, int_fwire_clk, delayed_D, int_fwire_s, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_D_Q_r = 0.34544:0.483245:1.74043;
		specparam tpd_D_Q_f = 0.430161:0.602153:1.68032;
		specparam tpd_XR_Q_negedge_r = 0.336951:0.487423:1.84686;
		specparam tpd_XR_Q_negedge_f = 0.270037:0.425382:1.55594;
		specparam tpd_XS_Q_negedge_r = 0.275052:0.44172:1.95059;
		specparam tpd_XS_Q_negedge_f = 0.446806:0.60737:1.38665;
		specparam tpd_XG_Q_negedge_r = 0.401694:0.588893:2.08352;
		specparam tpd_XG_Q_negedge_f = 0.475354:0.673481:1.79918;
		specparam tpd_D_XQ_r = 0.575326:0.712236:2.07641;
		specparam tpd_D_XQ_f = 0.477389:0.579823:1.47901;
		specparam tpd_XR_XQ_negedge_r = 0.396431:0.534099:1.94761;
		specparam tpd_XR_XQ_negedge_f = 0.469128:0.584312:1.58914;
		specparam tpd_XS_XQ_negedge_r = 0.586275:0.716874:1.81517;
		specparam tpd_XS_XQ_negedge_f = 0.384639:0.537283:1.7183;
		specparam tpd_XG_XQ_negedge_r = 0.620191:0.783443:2.22232;
		specparam tpd_XG_XQ_negedge_f = 0.534498:0.687148:1.83108;
		specparam tsetup_D_XG_adacond0_posedge_adacond0_posedge = 0.315347:0.321717:0.600809;
		specparam thold_D_XG_adacond0_posedge_adacond0_posedge = -0.231954:-0.249579:-0.487479;
		specparam tsetup_D_XG_adacond0_negedge_adacond0_posedge = 0.315347:0.321717:0.600809;
		specparam thold_D_XG_adacond0_negedge_adacond0_posedge = -0.231954:-0.249579:-0.487479;
		specparam trecovery_XR_XG_adacond1_posedge_adacond1_posedge = 0.311561:0.328613:0.663876;
		specparam tremoval_XR_XG_adacond1_posedge_adacond1_posedge = -0.222138:-0.253768:-0.573466;
		specparam tpw_XR_negedge = 0.283357:0.367527:2.72095;
		specparam trecovery_XS_XG_adacond2_posedge_adacond2_posedge = 0.389561:0.382193:0.354994;
		specparam tremoval_XS_XG_adacond2_posedge_adacond2_posedge = -0.240705:-0.238407:-0.230551;
		specparam tsetup_XS_XR_XG_posedge_XG_posedge = 0.312177:0.39262:1.1306;
		specparam thold_XS_XR_XG_posedge_XG_posedge = -0.209343:-0.308316:-0.618971;
		specparam tpw_XS_negedge = 0.225439:0.333433:2.72095;
		specparam tpw_XG_negedge = 0.439939:0.461941:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XG => (Q+:D)) = ( tpd_XG_Q_negedge_r , tpd_XG_Q_negedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XG => (XQ-:D)) = ( tpd_XG_XQ_negedge_r , tpd_XG_XQ_negedge_f );
		$setuphold (posedge XG &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XG_adacond0_posedge_adacond0_posedge, 
			 thold_D_XG_adacond0_posedge_adacond0_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XG &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XG_adacond0_negedge_adacond0_posedge, 
			 thold_D_XG_adacond0_negedge_adacond0_posedge, notifier,,, delayed_XG, delayed_D);
		$setuphold (posedge XR &&& XG, posedge XS &&& XG, 
			 tsetup_XS_XR_XG_posedge_XG_posedge, 
			 thold_XS_XR_XG_posedge_XG_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, posedge XG &&& adacond1, 
			 trecovery_XR_XG_adacond1_posedge_adacond1_posedge, notifier);
		$hold (posedge XG &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_XG_adacond1_posedge_adacond1_posedge, notifier);
		$recovery (posedge XS &&& adacond2, posedge XG &&& adacond2, 
			 trecovery_XS_XG_adacond2_posedge_adacond2_posedge, notifier);
		$hold (posedge XG &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_XG_adacond2_posedge_adacond2_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (negedge XG, tpw_XG_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLQ 
`timescale 1ns/10ps
`celldefine
module DLQX1 (Q, D, G);
	output Q;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ;

	altos_latch (int_fwire_IQ, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.175115:0.310498:1.54787;
		specparam tpd_D_Q_f = 0.225277:0.361937:1.36986;
		specparam tpd_G_Q_posedge_r = 0.286828:0.435001:1.58996;
		specparam tpd_G_Q_posedge_f = 0.252367:0.389064:1.11818;
		specparam tsetup_D_G_posedge_negedge = 0.00595404:-0.0292038:-0.295642;
		specparam thold_D_G_posedge_negedge = 0.0252636:0.0640491:0.370574;
		specparam tsetup_D_G_negedge_negedge = 0.00595404:-0.0292038:-0.295642;
		specparam thold_D_G_negedge_negedge = 0.0252636:0.0640491:0.370574;
		specparam tpw_G_posedge = 0.189034:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G, posedge D, 
			 tsetup_D_G_posedge_negedge, 
			 thold_D_G_posedge_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 
			 tsetup_D_G_negedge_negedge, 
			 thold_D_G_negedge_negedge, notifier,,, delayed_G, delayed_D);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLQ 
`timescale 1ns/10ps
`celldefine
module DLQX2 (Q, D, G);
	output Q;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ;

	altos_latch (int_fwire_IQ, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.14836:0.28083:1.50065;
		specparam tpd_D_Q_f = 0.190375:0.320889:1.27334;
		specparam tpd_G_Q_posedge_r = 0.268894:0.41564:1.5667;
		specparam tpd_G_Q_posedge_f = 0.217:0.348797:1.0265;
		specparam tsetup_D_G_posedge_negedge = -0.0259022:-0.071555:-0.383769;
		specparam thold_D_G_posedge_negedge = 0.0518333:0.10101:0.469482;
		specparam tsetup_D_G_negedge_negedge = -0.0259022:-0.071555:-0.383769;
		specparam thold_D_G_negedge_negedge = 0.0518333:0.10101:0.469482;
		specparam tpw_G_posedge = 0.153749:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G, posedge D, 
			 tsetup_D_G_posedge_negedge, 
			 thold_D_G_posedge_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 
			 tsetup_D_G_negedge_negedge, 
			 thold_D_G_negedge_negedge, notifier,,, delayed_G, delayed_D);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLQ 
`timescale 1ns/10ps
`celldefine
module DLQX4 (Q, D, G);
	output Q;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ;

	altos_latch (int_fwire_IQ, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.140614:0.264735:1.4407;
		specparam tpd_D_Q_f = 0.183713:0.30546:1.22078;
		specparam tpd_G_Q_posedge_r = 0.304804:0.453846:1.6346;
		specparam tpd_G_Q_posedge_f = 0.226712:0.359174:1.03898;
		specparam tsetup_D_G_posedge_negedge = -0.0837042:-0.146306:-0.572192;
		specparam thold_D_G_posedge_negedge = 0.103687:0.169426:0.647803;
		specparam tsetup_D_G_negedge_negedge = -0.0837042:-0.146306:-0.572192;
		specparam thold_D_G_negedge_negedge = 0.103687:0.169426:0.647803;
		specparam tpw_G_posedge = 0.155073:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G, posedge D, 
			 tsetup_D_G_posedge_negedge, 
			 thold_D_G_posedge_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 
			 tsetup_D_G_negedge_negedge, 
			 thold_D_G_negedge_negedge, notifier,,, delayed_G, delayed_D);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLQ 
`timescale 1ns/10ps
`celldefine
module DLQXL (Q, D, G);
	output Q;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ;

	altos_latch (int_fwire_IQ, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.170811:0.300588:1.52426;
		specparam tpd_D_Q_f = 0.207095:0.334729:1.31296;
		specparam tpd_G_Q_posedge_r = 0.280595:0.421187:1.55507;
		specparam tpd_G_Q_posedge_f = 0.230515:0.35619:1.05644;
		specparam tsetup_D_G_posedge_negedge = -0.00534815:-0.0438087:-0.325306;
		specparam thold_D_G_posedge_negedge = 0.0285558:0.0700903:0.392447;
		specparam tsetup_D_G_negedge_negedge = -0.00534815:-0.0438087:-0.325306;
		specparam thold_D_G_negedge_negedge = 0.0285558:0.0700903:0.392447;
		specparam tpw_G_posedge = 0.163011:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G, posedge D, 
			 tsetup_D_G_posedge_negedge, 
			 thold_D_G_posedge_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 
			 tsetup_D_G_negedge_negedge, 
			 thold_D_G_negedge_negedge, notifier,,, delayed_G, delayed_D);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLQX 
`timescale 1ns/10ps
`celldefine
module DLQXX1 (Q, XQ, D, G);
	output Q, XQ;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ;

	altos_latch (int_fwire_IQ, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.174908:0.308488:1.53371;
		specparam tpd_D_Q_f = 0.224725:0.359833:1.36248;
		specparam tpd_G_Q_posedge_r = 0.286676:0.433034:1.57721;
		specparam tpd_G_Q_posedge_f = 0.251793:0.386846:1.11053;
		specparam tpd_D_XQ_r = 0.334745:0.46547:1.86519;
		specparam tpd_D_XQ_f = 0.288003:0.395799:1.2352;
		specparam tpd_G_XQ_posedge_r = 0.361732:0.492382:1.64633;
		specparam tpd_G_XQ_posedge_f = 0.400545:0.521685:1.28747;
		specparam tsetup_D_G_posedge_negedge = 0.0165576:-0.0201684:-0.270472;
		specparam thold_D_G_posedge_negedge = 0.0251006:0.0622568:0.369723;
		specparam tsetup_D_G_negedge_negedge = 0.0165576:-0.0201684:-0.270472;
		specparam thold_D_G_negedge_negedge = 0.0251006:0.0622568:0.369723;
		specparam tpw_G_posedge = 0.208597:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G, posedge D, 
			 tsetup_D_G_posedge_negedge, 
			 thold_D_G_posedge_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 
			 tsetup_D_G_negedge_negedge, 
			 thold_D_G_negedge_negedge, notifier,,, delayed_G, delayed_D);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLQX 
`timescale 1ns/10ps
`celldefine
module DLQXX2 (Q, XQ, D, G);
	output Q, XQ;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ;

	altos_latch (int_fwire_IQ, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.150162:0.282123:1.50377;
		specparam tpd_D_Q_f = 0.191617:0.321476:1.27479;
		specparam tpd_G_Q_posedge_r = 0.271595:0.418183:1.57285;
		specparam tpd_G_Q_posedge_f = 0.218856:0.350231:1.03201;
		specparam tpd_D_XQ_r = 0.326389:0.45947:1.833;
		specparam tpd_D_XQ_f = 0.312826:0.42903:1.21093;
		specparam tpd_G_XQ_posedge_r = 0.353343:0.488256:1.61945;
		specparam tpd_G_XQ_posedge_f = 0.43506:0.566117:1.28334;
		specparam tsetup_D_G_posedge_negedge = -0.0168739:-0.0585797:-0.350021;
		specparam thold_D_G_posedge_negedge = 0.0515343:0.0997532:0.46415;
		specparam tsetup_D_G_negedge_negedge = -0.0168739:-0.0585797:-0.350021;
		specparam thold_D_G_negedge_negedge = 0.0515343:0.0997532:0.46415;
		specparam tpw_G_posedge = 0.17722:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G, posedge D, 
			 tsetup_D_G_posedge_negedge, 
			 thold_D_G_posedge_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 
			 tsetup_D_G_negedge_negedge, 
			 thold_D_G_negedge_negedge, notifier,,, delayed_G, delayed_D);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLQX 
`timescale 1ns/10ps
`celldefine
module DLQXX4 (Q, XQ, D, G);
	output Q, XQ;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ;

	altos_latch (int_fwire_IQ, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.140332:0.264722:1.44898;
		specparam tpd_D_Q_f = 0.183052:0.304845:1.2232;
		specparam tpd_G_Q_posedge_r = 0.304477:0.453931:1.64383;
		specparam tpd_G_Q_posedge_f = 0.225999:0.358513:1.04199;
		specparam tpd_D_XQ_r = 0.36768:0.506866:1.88454;
		specparam tpd_D_XQ_f = 0.378367:0.501303:1.24385;
		specparam tpd_G_XQ_posedge_r = 0.41132:0.561138:1.72062;
		specparam tpd_G_XQ_posedge_f = 0.543487:0.691489:1.43831;
		specparam tsetup_D_G_posedge_negedge = -0.0783192:-0.13372:-0.528923;
		specparam thold_D_G_posedge_negedge = 0.103582:0.168804:0.647924;
		specparam tsetup_D_G_negedge_negedge = -0.0783192:-0.13372:-0.528923;
		specparam thold_D_G_negedge_negedge = 0.103582:0.168804:0.647924;
		specparam tpw_G_posedge = 0.177244:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G, posedge D, 
			 tsetup_D_G_posedge_negedge, 
			 thold_D_G_posedge_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 
			 tsetup_D_G_negedge_negedge, 
			 thold_D_G_negedge_negedge, notifier,,, delayed_G, delayed_D);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLQX 
`timescale 1ns/10ps
`celldefine
module DLQXXL (Q, XQ, D, G);
	output Q, XQ;
	input D, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ;

	altos_latch (int_fwire_IQ, notifier, delayed_G, delayed_D);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.170789:0.300876:1.53662;
		specparam tpd_D_Q_f = 0.206823:0.334651:1.32085;
		specparam tpd_G_Q_posedge_r = 0.280571:0.421452:1.56869;
		specparam tpd_G_Q_posedge_f = 0.23026:0.356155:1.06406;
		specparam tpd_D_XQ_r = 0.293783:0.423762:1.813;
		specparam tpd_D_XQ_f = 0.259327:0.366444:1.23011;
		specparam tpd_G_XQ_posedge_r = 0.316965:0.445272:1.5907;
		specparam tpd_G_XQ_posedge_f = 0.369892:0.488116:1.27612;
		specparam tsetup_D_G_posedge_negedge = -0.00138782:-0.0363222:-0.311839;
		specparam thold_D_G_posedge_negedge = 0.0276596:0.070816:0.391454;
		specparam tsetup_D_G_negedge_negedge = -0.00138782:-0.0363222:-0.311839;
		specparam thold_D_G_negedge_negedge = 0.0276596:0.070816:0.391454;
		specparam tpw_G_posedge = 0.171085:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G, posedge D, 
			 tsetup_D_G_posedge_negedge, 
			 thold_D_G_posedge_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G, negedge D, 
			 tsetup_D_G_negedge_negedge, 
			 thold_D_G_negedge_negedge, notifier,,, delayed_G, delayed_D);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLRQ 
`timescale 1ns/10ps
`celldefine
module DLRQX1 (Q, D, XR, G);
	output Q;
	input D, XR, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_r;

	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.265077:0.405598:1.66441;
		specparam tpd_D_Q_f = 0.249153:0.395827:1.45513;
		specparam tpd_XR_Q_negedge_r = 0.255774:0.408897:1.71327;
		specparam tpd_XR_Q_negedge_f = 0.180704:0.358152:1.56667;
		specparam tpd_G_Q_posedge_r = 0.342782:0.504553:1.63836;
		specparam tpd_G_Q_posedge_f = 0.271774:0.415052:1.19541;
		specparam tsetup_D_G_XR_posedge_XR_negedge = 0.130628:0.0754806:-0.140092;
		specparam thold_D_G_XR_posedge_XR_negedge = -0.0564556:-0.00773712:0.252945;
		specparam tsetup_D_G_XR_negedge_XR_negedge = 0.130628:0.0754806:-0.140092;
		specparam thold_D_G_XR_negedge_XR_negedge = -0.0564556:-0.00773712:0.252945;
		specparam trecovery_XR_G_D_posedge_D_negedge = 0.13281:0.0912874:-0.0615905;
		specparam tremoval_XR_G_D_posedge_D_negedge = -0.0571787:-0.0235439:0.179137;
		specparam tpw_XR_negedge = 0.180304:0.330811:2.72095;
		specparam tpw_G_posedge = 0.235608:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& XR, posedge D &&& XR, 
			 tsetup_D_G_XR_posedge_XR_negedge, 
			 thold_D_G_XR_posedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XR, negedge D &&& XR, 
			 tsetup_D_G_XR_negedge_XR_negedge, 
			 thold_D_G_XR_negedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XR &&& D, negedge G &&& D, 
			 trecovery_XR_G_D_posedge_D_negedge, notifier);
		$hold (negedge G &&& D, posedge XR &&& D, 
			 tremoval_XR_G_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLRQ 
`timescale 1ns/10ps
`celldefine
module DLRQX2 (Q, D, XR, G);
	output Q;
	input D, XR, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_r;

	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.213482:0.34448:1.56132;
		specparam tpd_D_Q_f = 0.218623:0.356293:1.34274;
		specparam tpd_XR_Q_negedge_r = 0.199746:0.344171:1.52804;
		specparam tpd_XR_Q_negedge_f = 0.254391:0.452611:1.79479;
		specparam tpd_G_Q_posedge_r = 0.319297:0.481343:1.66618;
		specparam tpd_G_Q_posedge_f = 0.252321:0.394184:1.12567;
		specparam tsetup_D_G_XR_posedge_XR_negedge = 0.0341181:-0.0181153:-0.318079;
		specparam thold_D_G_XR_posedge_XR_negedge = 0.00678483:0.0628698:0.412589;
		specparam tsetup_D_G_XR_negedge_XR_negedge = 0.0341181:-0.0181153:-0.318079;
		specparam thold_D_G_XR_negedge_XR_negedge = 0.00678483:0.0628698:0.412589;
		specparam trecovery_XR_G_D_posedge_D_negedge = 0.0264206:-0.0117219:-0.31867;
		specparam tremoval_XR_G_D_posedge_D_negedge = 0.0166526:0.0543451:0.420596;
		specparam tpw_XR_negedge = 0.256122:0.398998:2.72095;
		specparam tpw_G_posedge = 0.190377:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& XR, posedge D &&& XR, 
			 tsetup_D_G_XR_posedge_XR_negedge, 
			 thold_D_G_XR_posedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XR, negedge D &&& XR, 
			 tsetup_D_G_XR_negedge_XR_negedge, 
			 thold_D_G_XR_negedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XR &&& D, negedge G &&& D, 
			 trecovery_XR_G_D_posedge_D_negedge, notifier);
		$hold (negedge G &&& D, posedge XR &&& D, 
			 tremoval_XR_G_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLRQ 
`timescale 1ns/10ps
`celldefine
module DLRQX4 (Q, D, XR, G);
	output Q;
	input D, XR, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_r;

	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.197388:0.325276:1.52766;
		specparam tpd_D_Q_f = 0.204419:0.335219:1.27494;
		specparam tpd_XR_Q_negedge_r = 0.181415:0.322125:1.43695;
		specparam tpd_XR_Q_negedge_f = 0.413066:0.639449:2.1723;
		specparam tpd_G_Q_posedge_r = 0.294545:0.456066:1.66413;
		specparam tpd_G_Q_posedge_f = 0.241304:0.382848:1.1328;
		specparam tsetup_D_G_XR_posedge_XR_negedge = 0.0053268:-0.0441392:-0.319609;
		specparam thold_D_G_XR_posedge_XR_negedge = 0.0160648:0.0701203:0.383047;
		specparam tsetup_D_G_XR_negedge_XR_negedge = 0.0053268:-0.0441392:-0.319609;
		specparam thold_D_G_XR_negedge_XR_negedge = 0.0160648:0.0701203:0.383047;
		specparam trecovery_XR_G_D_posedge_D_negedge = -0.00510892:-0.0412982:-0.379753;
		specparam tremoval_XR_G_D_posedge_D_negedge = 0.0278955:0.0678607:0.447185;
		specparam tpw_XR_negedge = 0.38214:0.525574:2.72095;
		specparam tpw_G_posedge = 0.176397:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& XR, posedge D &&& XR, 
			 tsetup_D_G_XR_posedge_XR_negedge, 
			 thold_D_G_XR_posedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XR, negedge D &&& XR, 
			 tsetup_D_G_XR_negedge_XR_negedge, 
			 thold_D_G_XR_negedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XR &&& D, negedge G &&& D, 
			 trecovery_XR_G_D_posedge_D_negedge, notifier);
		$hold (negedge G &&& D, posedge XR &&& D, 
			 tremoval_XR_G_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLRQ 
`timescale 1ns/10ps
`celldefine
module DLRQXL (Q, D, XR, G);
	output Q;
	input D, XR, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_r;

	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.257385:0.392759:1.65788;
		specparam tpd_D_Q_f = 0.235413:0.376486:1.44138;
		specparam tpd_XR_Q_negedge_r = 0.248036:0.396098:1.70017;
		specparam tpd_XR_Q_negedge_f = 0.170914:0.342354:1.54781;
		specparam tpd_G_Q_posedge_r = 0.338986:0.495779:1.64205;
		specparam tpd_G_Q_posedge_f = 0.25717:0.394804:1.18822;
		specparam tsetup_D_G_XR_posedge_XR_negedge = 0.102983:0.0491269:-0.186764;
		specparam thold_D_G_XR_posedge_XR_negedge = -0.0424812:0.00512869:0.279507;
		specparam tsetup_D_G_XR_negedge_XR_negedge = 0.102983:0.0491269:-0.186764;
		specparam thold_D_G_XR_negedge_XR_negedge = -0.0424812:0.00512869:0.279507;
		specparam trecovery_XR_G_D_posedge_D_negedge = 0.10386:0.0653604:-0.110446;
		specparam tremoval_XR_G_D_posedge_D_negedge = -0.0436621:-0.0108607:0.205956;
		specparam tpw_XR_negedge = 0.165833:0.330811:2.72095;
		specparam tpw_G_posedge = 0.214744:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& XR, posedge D &&& XR, 
			 tsetup_D_G_XR_posedge_XR_negedge, 
			 thold_D_G_XR_posedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XR, negedge D &&& XR, 
			 tsetup_D_G_XR_negedge_XR_negedge, 
			 thold_D_G_XR_negedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XR &&& D, negedge G &&& D, 
			 trecovery_XR_G_D_posedge_D_negedge, notifier);
		$hold (negedge G &&& D, posedge XR &&& D, 
			 tremoval_XR_G_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLRQX 
`timescale 1ns/10ps
`celldefine
module DLRQXX1 (Q, XQ, D, XR, G);
	output Q, XQ;
	input D, XR, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;

	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.266808:0.406716:1.67727;
		specparam tpd_D_Q_f = 0.245546:0.388934:1.41115;
		specparam tpd_XR_Q_negedge_r = 0.257469:0.410067:1.72511;
		specparam tpd_XR_Q_negedge_f = 0.175983:0.349216:1.51681;
		specparam tpd_G_Q_posedge_r = 0.347964:0.509006:1.65525;
		specparam tpd_G_Q_posedge_f = 0.267767:0.407425:1.1484;
		specparam tpd_D_XQ_r = 0.36439:0.495169:1.86388;
		specparam tpd_D_XQ_f = 0.418518:0.515145:1.33855;
		specparam tpd_XR_XQ_negedge_r = 0.296271:0.455222:1.95296;
		specparam tpd_XR_XQ_negedge_f = 0.409428:0.518964:1.3911;
		specparam tpd_G_XQ_posedge_r = 0.386678:0.513783:1.63474;
		specparam tpd_G_XQ_posedge_f = 0.500558:0.618833:1.3272;
		specparam tsetup_D_G_XR_posedge_XR_negedge = 0.156064:0.0996625:-0.117597;
		specparam thold_D_G_XR_posedge_XR_negedge = -0.0565272:-0.00969172:0.252262;
		specparam tsetup_D_G_XR_negedge_XR_negedge = 0.156064:0.0996625:-0.117597;
		specparam thold_D_G_XR_negedge_XR_negedge = -0.0565272:-0.00969172:0.252262;
		specparam trecovery_XR_G_D_posedge_D_negedge = 0.158878:0.114717:-0.034976;
		specparam tremoval_XR_G_D_posedge_D_negedge = -0.0562211:-0.0239849:0.179157;
		specparam tpw_XR_negedge = 0.204616:0.341301:2.72095;
		specparam tpw_G_posedge = 0.269512:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& XR, posedge D &&& XR, 
			 tsetup_D_G_XR_posedge_XR_negedge, 
			 thold_D_G_XR_posedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XR, negedge D &&& XR, 
			 tsetup_D_G_XR_negedge_XR_negedge, 
			 thold_D_G_XR_negedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XR &&& D, negedge G &&& D, 
			 trecovery_XR_G_D_posedge_D_negedge, notifier);
		$hold (negedge G &&& D, posedge XR &&& D, 
			 tremoval_XR_G_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLRQX 
`timescale 1ns/10ps
`celldefine
module DLRQXX2 (Q, XQ, D, XR, G);
	output Q, XQ;
	input D, XR, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;

	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.214151:0.34426:1.55915;
		specparam tpd_D_Q_f = 0.217835:0.353974:1.3269;
		specparam tpd_XR_Q_negedge_r = 0.200425:0.344194:1.52453;
		specparam tpd_XR_Q_negedge_f = 0.253079:0.448785:1.7787;
		specparam tpd_G_Q_posedge_r = 0.320414:0.481934:1.66434;
		specparam tpd_G_Q_posedge_f = 0.251732:0.392098:1.11116;
		specparam tpd_D_XQ_r = 0.367192:0.502306:1.89375;
		specparam tpd_D_XQ_f = 0.397052:0.491247:1.16043;
		specparam tpd_XR_XQ_negedge_r = 0.44707:0.611613:2.27647;
		specparam tpd_XR_XQ_negedge_f = 0.383563:0.491309:1.1293;
		specparam tpd_G_XQ_posedge_r = 0.40124:0.540767:1.70648;
		specparam tpd_G_XQ_posedge_f = 0.504116:0.630422:1.2717;
		specparam tsetup_D_G_XR_posedge_XR_negedge = 0.0627115:0.00841324:-0.274538;
		specparam thold_D_G_XR_posedge_XR_negedge = 0.0086452:0.061037:0.413097;
		specparam tsetup_D_G_XR_negedge_XR_negedge = 0.0627115:0.00841324:-0.274538;
		specparam thold_D_G_XR_negedge_XR_negedge = 0.0086452:0.061037:0.413097;
		specparam trecovery_XR_G_D_posedge_D_negedge = 0.0563019:0.014655:-0.271538;
		specparam tremoval_XR_G_D_posedge_D_negedge = 0.0151134:0.0550784:0.416629;
		specparam tpw_XR_negedge = 0.301681:0.435715:2.72095;
		specparam tpw_G_posedge = 0.218886:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& XR, posedge D &&& XR, 
			 tsetup_D_G_XR_posedge_XR_negedge, 
			 thold_D_G_XR_posedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XR, negedge D &&& XR, 
			 tsetup_D_G_XR_negedge_XR_negedge, 
			 thold_D_G_XR_negedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XR &&& D, negedge G &&& D, 
			 trecovery_XR_G_D_posedge_D_negedge, notifier);
		$hold (negedge G &&& D, posedge XR &&& D, 
			 tremoval_XR_G_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLRQX 
`timescale 1ns/10ps
`celldefine
module DLRQXX4 (Q, XQ, D, XR, G);
	output Q, XQ;
	input D, XR, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;

	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.200572:0.327441:1.52884;
		specparam tpd_D_Q_f = 0.205006:0.331859:1.22626;
		specparam tpd_XR_Q_negedge_r = 0.18459:0.324504:1.43988;
		specparam tpd_XR_Q_negedge_f = 0.40842:0.625734:2.11495;
		specparam tpd_G_Q_posedge_r = 0.297751:0.458149:1.66496;
		specparam tpd_G_Q_posedge_f = 0.241906:0.379486:1.08376;
		specparam tpd_D_XQ_r = 0.344112:0.475659:1.86954;
		specparam tpd_D_XQ_f = 0.363011:0.457456:1.15357;
		specparam tpd_XR_XQ_negedge_r = 0.65782:0.814279:2.59921;
		specparam tpd_XR_XQ_negedge_f = 0.347162:0.454616:1.07051;
		specparam tpd_G_XQ_posedge_r = 0.381236:0.523459:1.75051;
		specparam tpd_G_XQ_posedge_f = 0.460617:0.589453:1.29764;
		specparam tsetup_D_G_XR_posedge_XR_negedge = 0.0292218:-0.0211308:-0.269066;
		specparam thold_D_G_XR_posedge_XR_negedge = 0.0148734:0.0674207:0.375558;
		specparam tsetup_D_G_XR_negedge_XR_negedge = 0.0292218:-0.0211308:-0.269066;
		specparam thold_D_G_XR_negedge_XR_negedge = 0.0148734:0.0674207:0.375558;
		specparam trecovery_XR_G_D_posedge_D_negedge = 0.0190595:-0.017694:-0.325112;
		specparam tremoval_XR_G_D_posedge_D_negedge = 0.0278039:0.0636376:0.439143;
		specparam tpw_XR_negedge = 0.447731:0.581974:2.72095;
		specparam tpw_G_posedge = 0.200412:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& XR, posedge D &&& XR, 
			 tsetup_D_G_XR_posedge_XR_negedge, 
			 thold_D_G_XR_posedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XR, negedge D &&& XR, 
			 tsetup_D_G_XR_negedge_XR_negedge, 
			 thold_D_G_XR_negedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XR &&& D, negedge G &&& D, 
			 trecovery_XR_G_D_posedge_D_negedge, notifier);
		$hold (negedge G &&& D, posedge XR &&& D, 
			 tremoval_XR_G_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLRQX 
`timescale 1ns/10ps
`celldefine
module DLRQXXL (Q, XQ, D, XR, G);
	output Q, XQ;
	input D, XR, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;

	not (int_fwire_r, XR);
	altos_latch_r (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.258266:0.393079:1.66409;
		specparam tpd_D_Q_f = 0.235908:0.376338:1.44521;
		specparam tpd_XR_Q_negedge_r = 0.248926:0.396435:1.71022;
		specparam tpd_XR_Q_negedge_f = 0.171582:0.342115:1.55157;
		specparam tpd_G_Q_posedge_r = 0.339871:0.496152:1.64868;
		specparam tpd_G_Q_posedge_f = 0.257656:0.394654:1.19239;
		specparam tpd_D_XQ_r = 0.336468:0.468131:1.84788;
		specparam tpd_D_XQ_f = 0.380388:0.476824:1.31976;
		specparam tpd_XR_XQ_negedge_r = 0.274584:0.43387:1.9357;
		specparam tpd_XR_XQ_negedge_f = 0.371278:0.480488:1.36766;
		specparam tpd_G_XQ_posedge_r = 0.35823:0.486525:1.62833;
		specparam tpd_G_XQ_posedge_f = 0.462872:0.581144:1.32094;
		specparam tsetup_D_G_XR_posedge_XR_negedge = 0.120039:0.064652:-0.168783;
		specparam thold_D_G_XR_posedge_XR_negedge = -0.0400799:0.00604518:0.281044;
		specparam tsetup_D_G_XR_negedge_XR_negedge = 0.120039:0.064652:-0.168783;
		specparam thold_D_G_XR_negedge_XR_negedge = -0.0400799:0.00604518:0.281044;
		specparam trecovery_XR_G_D_posedge_D_negedge = 0.123301:0.0790473:-0.09051;
		specparam tremoval_XR_G_D_posedge_D_negedge = -0.0414256:-0.0102567:0.207727;
		specparam tpw_XR_negedge = 0.181022:0.330811:2.72095;
		specparam tpw_G_posedge = 0.233278:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& XR, posedge D &&& XR, 
			 tsetup_D_G_XR_posedge_XR_negedge, 
			 thold_D_G_XR_posedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XR, negedge D &&& XR, 
			 tsetup_D_G_XR_negedge_XR_negedge, 
			 thold_D_G_XR_negedge_XR_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XR &&& D, negedge G &&& D, 
			 trecovery_XR_G_D_posedge_D_negedge, notifier);
		$hold (negedge G &&& D, posedge XR &&& D, 
			 tremoval_XR_G_D_posedge_D_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSQ 
`timescale 1ns/10ps
`celldefine
module DLSQX1 (Q, D, XS, G);
	output Q;
	input D, XS, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_s;

	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.210253:0.354984:1.61915;
		specparam tpd_D_Q_f = 0.373012:0.528459:1.56219;
		specparam tpd_XS_Q_negedge_r = 0.242666:0.409821:1.86837;
		specparam tpd_XS_Q_negedge_f = 0.397309:0.546885:1.28609;
		specparam tpd_G_Q_posedge_r = 0.325114:0.475827:1.59788;
		specparam tpd_G_Q_posedge_f = 0.321839:0.47525:1.25595;
		specparam tsetup_D_G_XS_posedge_XS_negedge = 0.0563833:0.0189361:-0.207739;
		specparam thold_D_G_XS_posedge_XS_negedge = 0.000670067:0.0328781:0.321783;
		specparam tsetup_D_G_XS_negedge_XS_negedge = 0.0563833:0.0189361:-0.207739;
		specparam thold_D_G_XS_negedge_XS_negedge = 0.000670067:0.0328781:0.321783;
		specparam trecovery_XS_G_NTB_D_posedge_NTB_D_negedge = 0.351455:0.336972:0.187323;
		specparam tremoval_XS_G_NTB_D_posedge_NTB_D_negedge = -0.258489:-0.253792:-0.0466764;
		specparam tpw_XS_negedge = 0.187272:0.330811:2.72095;
		specparam tpw_G_posedge = 0.277938:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& XS, posedge D &&& XS, 
			 tsetup_D_G_XS_posedge_XS_negedge, 
			 thold_D_G_XS_posedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XS, negedge D &&& XS, 
			 tsetup_D_G_XS_negedge_XS_negedge, 
			 thold_D_G_XS_negedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XS &&& ~D, negedge G &&& ~D, 
			 trecovery_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge G &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSQ 
`timescale 1ns/10ps
`celldefine
module DLSQX2 (Q, D, XS, G);
	output Q;
	input D, XS, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_s;

	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.173361:0.313382:1.55685;
		specparam tpd_D_Q_f = 0.314215:0.459645:1.43648;
		specparam tpd_XS_Q_negedge_r = 0.340896:0.523155:2.04814;
		specparam tpd_XS_Q_negedge_f = 0.344839:0.492916:1.20462;
		specparam tpd_G_Q_posedge_r = 0.315325:0.469479:1.64123;
		specparam tpd_G_Q_posedge_f = 0.274941:0.426189:1.17698;
		specparam tsetup_D_G_XS_posedge_XS_negedge = -0.0223171:-0.0601353:-0.385746;
		specparam thold_D_G_XS_posedge_XS_negedge = 0.0545849:0.0993286:0.484035;
		specparam tsetup_D_G_XS_negedge_XS_negedge = -0.0223171:-0.0601353:-0.385746;
		specparam thold_D_G_XS_negedge_XS_negedge = 0.0545849:0.0993286:0.484035;
		specparam trecovery_XS_G_NTB_D_posedge_NTB_D_negedge = 0.286454:0.280611:0.182153;
		specparam tremoval_XS_G_NTB_D_posedge_NTB_D_negedge = -0.212387:-0.215423:-0.0241151;
		specparam tpw_XS_negedge = 0.253639:0.349169:2.72095;
		specparam tpw_G_posedge = 0.221458:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& XS, posedge D &&& XS, 
			 tsetup_D_G_XS_posedge_XS_negedge, 
			 thold_D_G_XS_posedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XS, negedge D &&& XS, 
			 tsetup_D_G_XS_negedge_XS_negedge, 
			 thold_D_G_XS_negedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XS &&& ~D, negedge G &&& ~D, 
			 trecovery_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge G &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSQ 
`timescale 1ns/10ps
`celldefine
module DLSQX4 (Q, D, XS, G);
	output Q;
	input D, XS, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_s;

	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.163963:0.29962:1.50759;
		specparam tpd_D_Q_f = 0.310674:0.44856:1.37639;
		specparam tpd_XS_Q_negedge_r = 0.516607:0.71333:2.23391;
		specparam tpd_XS_Q_negedge_f = 0.348215:0.497622:1.20058;
		specparam tpd_G_Q_posedge_r = 0.285667:0.440791:1.63903;
		specparam tpd_G_Q_posedge_f = 0.267503:0.417485:1.15846;
		specparam tsetup_D_G_XS_posedge_XS_negedge = -0.0277299:-0.0664665:-0.38226;
		specparam thold_D_G_XS_posedge_XS_negedge = 0.0497156:0.0939785:0.455133;
		specparam tsetup_D_G_XS_negedge_XS_negedge = -0.0277299:-0.0664665:-0.38226;
		specparam thold_D_G_XS_negedge_XS_negedge = 0.0497156:0.0939785:0.455133;
		specparam trecovery_XS_G_NTB_D_posedge_NTB_D_negedge = 0.289677:0.299029:0.304226;
		specparam tremoval_XS_G_NTB_D_posedge_NTB_D_negedge = -0.221104:-0.240739:-0.15682;
		specparam tpw_XS_negedge = 0.345654:0.414734:2.72095;
		specparam tpw_G_posedge = 0.212043:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& XS, posedge D &&& XS, 
			 tsetup_D_G_XS_posedge_XS_negedge, 
			 thold_D_G_XS_posedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XS, negedge D &&& XS, 
			 tsetup_D_G_XS_negedge_XS_negedge, 
			 thold_D_G_XS_negedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XS &&& ~D, negedge G &&& ~D, 
			 trecovery_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge G &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSQ 
`timescale 1ns/10ps
`celldefine
module DLSQXL (Q, D, XS, G);
	output Q;
	input D, XS, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_s;

	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.204153:0.345355:1.61588;
		specparam tpd_D_Q_f = 0.344827:0.494224:1.52349;
		specparam tpd_XS_Q_negedge_r = 0.240179:0.405313:1.87756;
		specparam tpd_XS_Q_negedge_f = 0.368861:0.512469:1.25312;
		specparam tpd_G_Q_posedge_r = 0.319247:0.467022:1.60505;
		specparam tpd_G_Q_posedge_f = 0.293304:0.440884:1.2239;
		specparam tsetup_D_G_XS_posedge_XS_negedge = 0.0335952:0.000717997:-0.252259;
		specparam thold_D_G_XS_posedge_XS_negedge = 0.012346:0.0417806:0.346703;
		specparam tsetup_D_G_XS_negedge_XS_negedge = 0.0335952:0.000717997:-0.252259;
		specparam thold_D_G_XS_negedge_XS_negedge = 0.012346:0.0417806:0.346703;
		specparam trecovery_XS_G_NTB_D_posedge_NTB_D_negedge = 0.318738:0.303841:0.158942;
		specparam tremoval_XS_G_NTB_D_posedge_NTB_D_negedge = -0.231454:-0.229641:-0.0211851;
		specparam tpw_XS_negedge = 0.177373:0.330811:2.72095;
		specparam tpw_G_posedge = 0.24429:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& XS, posedge D &&& XS, 
			 tsetup_D_G_XS_posedge_XS_negedge, 
			 thold_D_G_XS_posedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XS, negedge D &&& XS, 
			 tsetup_D_G_XS_negedge_XS_negedge, 
			 thold_D_G_XS_negedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XS &&& ~D, negedge G &&& ~D, 
			 trecovery_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge G &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSQX 
`timescale 1ns/10ps
`celldefine
module DLSQXX1 (Q, XQ, D, XS, G);
	output Q, XQ;
	input D, XS, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_s;

	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.210772:0.355726:1.6411;
		specparam tpd_D_Q_f = 0.369723:0.522739:1.54506;
		specparam tpd_XS_Q_negedge_r = 0.245606:0.413824:1.89628;
		specparam tpd_XS_Q_negedge_f = 0.393988:0.541133:1.26897;
		specparam tpd_G_Q_posedge_r = 0.325684:0.476693:1.62292;
		specparam tpd_G_Q_posedge_f = 0.318384:0.46936:1.23895;
		specparam tpd_D_XQ_r = 0.504683:0.630651:1.98046;
		specparam tpd_D_XQ_f = 0.353188:0.464228:1.31076;
		specparam tpd_XS_XQ_negedge_r = 0.528454:0.648489:1.73685;
		specparam tpd_XS_XQ_negedge_f = 0.372861:0.519625:1.5776;
		specparam tpd_G_XQ_posedge_r = 0.453359:0.576925:1.70992;
		specparam tpd_G_XQ_posedge_f = 0.469272:0.586754:1.29746;
		specparam tsetup_D_G_XS_posedge_XS_negedge = 0.0763345:0.0371302:-0.178668;
		specparam thold_D_G_XS_posedge_XS_negedge = 0.00257284:0.0333882:0.322503;
		specparam tsetup_D_G_XS_negedge_XS_negedge = 0.0763345:0.0371302:-0.178668;
		specparam thold_D_G_XS_negedge_XS_negedge = 0.00257284:0.0333882:0.322503;
		specparam trecovery_XS_G_NTB_D_posedge_NTB_D_negedge = 0.376811:0.360975:0.18211;
		specparam tremoval_XS_G_NTB_D_posedge_NTB_D_negedge = -0.251962:-0.250782:-0.0434451;
		specparam tpw_XS_negedge = 0.200608:0.330811:2.72095;
		specparam tpw_G_posedge = 0.306654:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& XS, posedge D &&& XS, 
			 tsetup_D_G_XS_posedge_XS_negedge, 
			 thold_D_G_XS_posedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XS, negedge D &&& XS, 
			 tsetup_D_G_XS_negedge_XS_negedge, 
			 thold_D_G_XS_negedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XS &&& ~D, negedge G &&& ~D, 
			 trecovery_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge G &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSQX 
`timescale 1ns/10ps
`celldefine
module DLSQXX2 (Q, XQ, D, XS, G);
	output Q, XQ;
	input D, XS, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_s;

	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.175047:0.313502:1.54682;
		specparam tpd_D_Q_f = 0.312477:0.453545:1.39639;
		specparam tpd_XS_Q_negedge_r = 0.343033:0.523377:2.03853;
		specparam tpd_XS_Q_negedge_f = 0.343069:0.486967:1.16628;
		specparam tpd_G_Q_posedge_r = 0.316957:0.469425:1.63175;
		specparam tpd_G_Q_posedge_f = 0.273267:0.420115:1.1376;
		specparam tpd_D_XQ_r = 0.477525:0.605959:1.9459;
		specparam tpd_D_XQ_f = 0.344925:0.457853:1.19984;
		specparam tpd_XS_XQ_negedge_r = 0.507718:0.638998:1.7451;
		specparam tpd_XS_XQ_negedge_f = 0.520814:0.668881:1.6955;
		specparam tpd_G_XQ_posedge_r = 0.437859:0.572226:1.7171;
		specparam tpd_G_XQ_posedge_f = 0.487479:0.615614:1.28726;
		specparam tsetup_D_G_XS_posedge_XS_negedge = -0.000673088:-0.0397185:-0.340155;
		specparam thold_D_G_XS_posedge_XS_negedge = 0.0526818:0.0976415:0.482339;
		specparam tsetup_D_G_XS_negedge_XS_negedge = -0.000673088:-0.0397185:-0.340155;
		specparam thold_D_G_XS_negedge_XS_negedge = 0.0526818:0.0976415:0.482339;
		specparam trecovery_XS_G_NTB_D_posedge_NTB_D_negedge = 0.326568:0.315163:0.181261;
		specparam tremoval_XS_G_NTB_D_posedge_NTB_D_negedge = -0.213212:-0.215279:-0.0215318;
		specparam tpw_XS_negedge = 0.27597:0.362282:2.72095;
		specparam tpw_G_posedge = 0.257645:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& XS, posedge D &&& XS, 
			 tsetup_D_G_XS_posedge_XS_negedge, 
			 thold_D_G_XS_posedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XS, negedge D &&& XS, 
			 tsetup_D_G_XS_negedge_XS_negedge, 
			 thold_D_G_XS_negedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XS &&& ~D, negedge G &&& ~D, 
			 trecovery_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge G &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSQX 
`timescale 1ns/10ps
`celldefine
module DLSQXX4 (Q, XQ, D, XS, G);
	output Q, XQ;
	input D, XS, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_s;

	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.163953:0.299951:1.51411;
		specparam tpd_D_Q_f = 0.314145:0.455615:1.42965;
		specparam tpd_XS_Q_negedge_r = 0.51893:0.716581:2.25083;
		specparam tpd_XS_Q_negedge_f = 0.35374:0.507291:1.25803;
		specparam tpd_G_Q_posedge_r = 0.285646:0.441135:1.64561;
		specparam tpd_G_Q_posedge_f = 0.270994:0.424425:1.21124;
		specparam tpd_D_XQ_r = 0.471695:0.597746:1.95841;
		specparam tpd_D_XQ_f = 0.322608:0.433836:1.16175;
		specparam tpd_XS_XQ_negedge_r = 0.511037:0.649283:1.81534;
		specparam tpd_XS_XQ_negedge_f = 0.719303:0.859175:1.89425;
		specparam tpd_G_XQ_posedge_r = 0.428381:0.566175:1.77061;
		specparam tpd_G_XQ_posedge_f = 0.444216:0.575825:1.29955;
		specparam tsetup_D_G_XS_posedge_XS_negedge = -0.0158967:-0.0549041:-0.33988;
		specparam thold_D_G_XS_posedge_XS_negedge = 0.0494563:0.0951986:0.456718;
		specparam tsetup_D_G_XS_negedge_XS_negedge = -0.0158967:-0.0549041:-0.33988;
		specparam thold_D_G_XS_negedge_XS_negedge = 0.0494563:0.0951986:0.456718;
		specparam trecovery_XS_G_NTB_D_posedge_NTB_D_negedge = 0.326242:0.332337:0.314328;
		specparam tremoval_XS_G_NTB_D_posedge_NTB_D_negedge = -0.227122:-0.24629:-0.164215;
		specparam tpw_XS_negedge = 0.382586:0.44096:2.72095;
		specparam tpw_G_posedge = 0.244608:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& XS, posedge D &&& XS, 
			 tsetup_D_G_XS_posedge_XS_negedge, 
			 thold_D_G_XS_posedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XS, negedge D &&& XS, 
			 tsetup_D_G_XS_negedge_XS_negedge, 
			 thold_D_G_XS_negedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XS &&& ~D, negedge G &&& ~D, 
			 trecovery_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge G &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSQX 
`timescale 1ns/10ps
`celldefine
module DLSQXXL (Q, XQ, D, XS, G);
	output Q, XQ;
	input D, XS, G;
	reg notifier;
	wire delayed_D, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_s;

	not (int_fwire_s, XS);
	altos_latch_s (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing
	specify
		specparam tpd_D_Q_r = 0.205902:0.34485:1.61595;
		specparam tpd_D_Q_f = 0.341909:0.486013:1.48491;
		specparam tpd_XS_Q_negedge_r = 0.244488:0.408602:1.88495;
		specparam tpd_XS_Q_negedge_f = 0.366091:0.504388:1.21602;
		specparam tpd_G_Q_posedge_r = 0.321042:0.466671:1.6077;
		specparam tpd_G_Q_posedge_f = 0.290438:0.432725:1.1867;
		specparam tpd_D_XQ_r = 0.458482:0.585927:1.93547;
		specparam tpd_D_XQ_f = 0.317155:0.426946:1.28059;
		specparam tpd_XS_XQ_negedge_r = 0.482129:0.603979:1.69786;
		specparam tpd_XS_XQ_negedge_f = 0.346027:0.490753:1.568;
		specparam tpd_G_XQ_posedge_r = 0.406727:0.532443:1.66896;
		specparam tpd_G_XQ_posedge_f = 0.433247:0.550152:1.28229;
		specparam tsetup_D_G_XS_posedge_XS_negedge = 0.0450871:0.0103574:-0.233818;
		specparam thold_D_G_XS_posedge_XS_negedge = 0.0135103:0.0432755:0.348786;
		specparam tsetup_D_G_XS_negedge_XS_negedge = 0.0450871:0.0103574:-0.233818;
		specparam thold_D_G_XS_negedge_XS_negedge = 0.0135103:0.0432755:0.348786;
		specparam trecovery_XS_G_NTB_D_posedge_NTB_D_negedge = 0.333546:0.318097:0.159937;
		specparam tremoval_XS_G_NTB_D_posedge_NTB_D_negedge = -0.227758:-0.225686:-0.0133491;
		specparam tpw_XS_negedge = 0.185624:0.330811:2.72095;
		specparam tpw_G_posedge = 0.25996:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& XS, posedge D &&& XS, 
			 tsetup_D_G_XS_posedge_XS_negedge, 
			 thold_D_G_XS_posedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& XS, negedge D &&& XS, 
			 tsetup_D_G_XS_negedge_XS_negedge, 
			 thold_D_G_XS_negedge_XS_negedge, notifier,,, delayed_G, delayed_D);
		$recovery (posedge XS &&& ~D, negedge G &&& ~D, 
			 trecovery_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$hold (negedge G &&& ~D, posedge XS &&& ~D, 
			 tremoval_XS_G_NTB_D_posedge_NTB_D_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSRQ 
`timescale 1ns/10ps
`celldefine
module DLSRQX1 (Q, D, XR, XS, G);
	output Q;
	input D, XR, XS, G;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_r, int_fwire_s;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_latch_sr_1 (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_D_Q_r = 0.292603:0.433479:1.66272;
		specparam tpd_D_Q_f = 0.420487:0.596986:1.67551;
		specparam tpd_XR_Q_negedge_r = 0.282586:0.435545:1.73889;
		specparam tpd_XR_Q_negedge_f = 0.310198:0.483603:1.70847;
		specparam tpd_XS_Q_negedge_r = 0.286672:0.460262:1.96339;
		specparam tpd_XS_Q_negedge_f = 0.437841:0.60543:1.39192;
		specparam tpd_G_Q_posedge_r = 0.402248:0.563678:1.69948;
		specparam tpd_G_Q_posedge_f = 0.36956:0.543427:1.37137;
		specparam tsetup_D_G_adacond0_posedge_adacond0_negedge = 0.132146:0.0758614:-0.175347;
		specparam thold_D_G_adacond0_posedge_adacond0_negedge = -0.0557058:-0.0100222:0.279119;
		specparam tsetup_D_G_adacond0_negedge_adacond0_negedge = 0.132146:0.0758614:-0.175347;
		specparam thold_D_G_adacond0_negedge_adacond0_negedge = -0.0557058:-0.0100222:0.279119;
		specparam trecovery_XR_G_adacond1_posedge_adacond1_negedge = 0.134114:0.0894544:-0.0625219;
		specparam tremoval_XR_G_adacond1_posedge_adacond1_negedge = -0.0547893:-0.0240397:0.17346;
		specparam tpw_XR_negedge = 0.299241:0.388508:2.72095;
		specparam trecovery_XS_G_adacond2_posedge_adacond2_negedge = 0.400138:0.389532:0.240458;
		specparam tremoval_XS_G_adacond2_posedge_adacond2_negedge = -0.287639:-0.287514:-0.100199;
		specparam tsetup_XS_XR_NTB_G_posedge_NTB_G_posedge = 0.329546:0.413446:1.20162;
		specparam thold_XS_XR_NTB_G_posedge_NTB_G_posedge = -0.241182:-0.344204:-0.680956;
		specparam tpw_XS_negedge = 0.239024:0.346546:2.72095;
		specparam tpw_G_posedge = 0.339927:0.330811:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_G_adacond0_posedge_adacond0_negedge, 
			 thold_D_G_adacond0_posedge_adacond0_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_G_adacond0_negedge_adacond0_negedge, 
			 thold_D_G_adacond0_negedge_adacond0_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (posedge XR &&& ~G, posedge XS &&& ~G, 
			 tsetup_XS_XR_NTB_G_posedge_NTB_G_posedge, 
			 thold_XS_XR_NTB_G_posedge_NTB_G_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge G &&& adacond1, 
			 trecovery_XR_G_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge G &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_G_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge G &&& adacond2, 
			 trecovery_XS_G_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge G &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_G_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSRQ 
`timescale 1ns/10ps
`celldefine
module DLSRQXL (Q, D, XR, XS, G);
	output Q;
	input D, XR, XS, G;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_r, int_fwire_s;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_latch_sr_1 (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s, int_fwire_r);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_D_Q_r = 0.341778:0.484527:1.76001;
		specparam tpd_D_Q_f = 0.432673:0.612076:1.71389;
		specparam tpd_XR_Q_negedge_r = 0.332971:0.488311:1.86595;
		specparam tpd_XR_Q_negedge_f = 0.271925:0.433331:1.59066;
		specparam tpd_XS_Q_negedge_r = 0.275321:0.445423:1.9773;
		specparam tpd_XS_Q_negedge_f = 0.44843:0.615266:1.41498;
		specparam tpd_G_Q_posedge_r = 0.44257:0.607784:1.78122;
		specparam tpd_G_Q_posedge_f = 0.379169:0.553059:1.39777;
		specparam tsetup_D_G_adacond0_posedge_adacond0_negedge = 0.172559:0.115817:-0.13042;
		specparam thold_D_G_adacond0_posedge_adacond0_negedge = -0.0985889:-0.0476679:0.22308;
		specparam tsetup_D_G_adacond0_negedge_adacond0_negedge = 0.172559:0.115817:-0.13042;
		specparam thold_D_G_adacond0_negedge_adacond0_negedge = -0.0985889:-0.0476679:0.22308;
		specparam trecovery_XR_G_adacond1_posedge_adacond1_negedge = 0.179701:0.132176:0.0134744;
		specparam tremoval_XR_G_adacond1_posedge_adacond1_negedge = -0.105257:-0.0647052:0.0824715;
		specparam tpw_XR_negedge = 0.268237:0.354414:2.72095;
		specparam trecovery_XS_G_adacond2_posedge_adacond2_negedge = 0.413296:0.403016:0.241338;
		specparam tremoval_XS_G_adacond2_posedge_adacond2_negedge = -0.292958:-0.293085:-0.100878;
		specparam tsetup_XS_XR_NTB_G_posedge_NTB_G_posedge = 0.299034:0.381042:1.13023;
		specparam thold_XS_XR_NTB_G_posedge_NTB_G_posedge = -0.212915:-0.313008:-0.626523;
		specparam tpw_XS_negedge = 0.222625:0.338678:2.72095;
		specparam tpw_G_posedge = 0.355632:0.346546:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		$setuphold (negedge G &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_G_adacond0_posedge_adacond0_negedge, 
			 thold_D_G_adacond0_posedge_adacond0_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_G_adacond0_negedge_adacond0_negedge, 
			 thold_D_G_adacond0_negedge_adacond0_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (posedge XR &&& ~G, posedge XS &&& ~G, 
			 tsetup_XS_XR_NTB_G_posedge_NTB_G_posedge, 
			 thold_XS_XR_NTB_G_posedge_NTB_G_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge G &&& adacond1, 
			 trecovery_XR_G_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge G &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_G_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge G &&& adacond2, 
			 trecovery_XS_G_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge G &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_G_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSRQX 
`timescale 1ns/10ps
`celldefine
module DLSRQXX1 (Q, XQ, D, XR, XS, G);
	output Q, XQ;
	input D, XR, XS, G;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire int_fwire_s;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_latch_sr_1 (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_D_Q_r = 0.288954:0.430954:1.66424;
		specparam tpd_D_Q_f = 0.418986:0.598448:1.70177;
		specparam tpd_XR_Q_negedge_r = 0.278962:0.432978:1.73995;
		specparam tpd_XR_Q_negedge_f = 0.308728:0.485269:1.73503;
		specparam tpd_XS_Q_negedge_r = 0.284448:0.458919:1.96873;
		specparam tpd_XS_Q_negedge_f = 0.436265:0.606841:1.41818;
		specparam tpd_G_Q_posedge_r = 0.398769:0.561358:1.70222;
		specparam tpd_G_Q_posedge_f = 0.368019:0.545044:1.39768;
		specparam tpd_D_XQ_r = 0.566989:0.700805:2.04877;
		specparam tpd_D_XQ_f = 0.450721:0.554705:1.4106;
		specparam tpd_XR_XQ_negedge_r = 0.451725:0.589175:2.03515;
		specparam tpd_XR_XQ_negedge_f = 0.441003:0.55725:1.49003;
		specparam tpd_XS_XQ_negedge_r = 0.579611:0.709306:1.79898;
		specparam tpd_XS_XQ_negedge_f = 0.422519:0.576233:1.73142;
		specparam tpd_G_XQ_posedge_r = 0.515956:0.647051:1.77436;
		specparam tpd_G_XQ_posedge_f = 0.56138:0.686919:1.45492;
		specparam tsetup_D_G_adacond0_posedge_adacond0_negedge = 0.154681:0.0965796:-0.148732;
		specparam thold_D_G_adacond0_posedge_adacond0_negedge = -0.05439:-0.00921542:0.286406;
		specparam tsetup_D_G_adacond0_negedge_adacond0_negedge = 0.154681:0.0965796:-0.148732;
		specparam thold_D_G_adacond0_negedge_adacond0_negedge = -0.05439:-0.00921542:0.286406;
		specparam trecovery_XR_G_adacond1_posedge_adacond1_negedge = 0.152171:0.108505:-0.0380577;
		specparam tremoval_XR_G_adacond1_posedge_adacond1_negedge = -0.052918:-0.0202574:0.179103;
		specparam tpw_XR_negedge = 0.329376:0.412111:2.72095;
		specparam trecovery_XS_G_adacond2_posedge_adacond2_negedge = 0.427405:0.417675:0.240336;
		specparam tremoval_XS_G_adacond2_posedge_adacond2_negedge = -0.29048:-0.287653:-0.0991129;
		specparam tsetup_XS_XR_NTB_G_posedge_NTB_G_posedge = 0.358388:0.43743:1.19678;
		specparam thold_XS_XR_NTB_G_posedge_NTB_G_posedge = -0.239981:-0.344158:-0.682655;
		specparam tpw_XS_negedge = 0.248143:0.349169:2.72095;
		specparam tpw_G_posedge = 0.373598:0.362282:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_G_adacond0_posedge_adacond0_negedge, 
			 thold_D_G_adacond0_posedge_adacond0_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_G_adacond0_negedge_adacond0_negedge, 
			 thold_D_G_adacond0_negedge_adacond0_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (posedge XR &&& ~G, posedge XS &&& ~G, 
			 tsetup_XS_XR_NTB_G_posedge_NTB_G_posedge, 
			 thold_XS_XR_NTB_G_posedge_NTB_G_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge G &&& adacond1, 
			 trecovery_XR_G_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge G &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_G_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge G &&& adacond2, 
			 trecovery_XS_G_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge G &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_G_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLSRQX 
`timescale 1ns/10ps
`celldefine
module DLSRQXXL (Q, XQ, D, XR, XS, G);
	output Q, XQ;
	input D, XR, XS, G;
	reg notifier;
	wire delayed_D, delayed_XR, delayed_XS, delayed_G;

	// Function
	wire int_fwire_IQ, int_fwire_IXQ, int_fwire_r;
	wire int_fwire_s;

	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_latch_sr_1 (int_fwire_IQ, notifier, delayed_G, delayed_D, int_fwire_s, int_fwire_r);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire D__bar;


	// Additional timing gates
	and (adacond0, XR, XS);
	and (adacond1, D, XS);
	not (D__bar, D);
	and (adacond2, D__bar, XR);

	specify
		specparam tpd_D_Q_r = 0.342958:0.483317:1.74403;
		specparam tpd_D_Q_f = 0.434076:0.610816:1.7048;
		specparam tpd_XR_Q_negedge_r = 0.334148:0.487079:1.85029;
		specparam tpd_XR_Q_negedge_f = 0.273228:0.432458:1.58137;
		specparam tpd_XS_Q_negedge_r = 0.276352:0.444718:1.96214;
		specparam tpd_XS_Q_negedge_f = 0.449808:0.614193:1.40598;
		specparam tpd_G_Q_posedge_r = 0.44393:0.606711:1.76623;
		specparam tpd_G_Q_posedge_f = 0.380571:0.551992:1.38858;
		specparam tpd_D_XQ_r = 0.573375:0.709048:2.06447;
		specparam tpd_D_XQ_f = 0.46884:0.567479:1.43637;
		specparam tpd_XR_XQ_negedge_r = 0.394722:0.53024:1.93719;
		specparam tpd_XR_XQ_negedge_f = 0.460308:0.571554:1.5461;
		specparam tpd_XS_XQ_negedge_r = 0.583758:0.712136:1.79914;
		specparam tpd_XS_XQ_negedge_f = 0.380352:0.529028:1.68759;
		specparam tpd_G_XQ_posedge_r = 0.519588:0.650092:1.77684;
		specparam tpd_G_XQ_posedge_f = 0.570757:0.69244:1.46769;
		specparam tsetup_D_G_adacond0_posedge_adacond0_negedge = 0.193013:0.131459:-0.112614;
		specparam thold_D_G_adacond0_posedge_adacond0_negedge = -0.0989919:-0.048042:0.223332;
		specparam tsetup_D_G_adacond0_negedge_adacond0_negedge = 0.193013:0.131459:-0.112614;
		specparam thold_D_G_adacond0_negedge_adacond0_negedge = -0.0989919:-0.048042:0.223332;
		specparam trecovery_XR_G_adacond1_posedge_adacond1_negedge = 0.19357:0.147944:0.0311824;
		specparam tremoval_XR_G_adacond1_posedge_adacond1_negedge = -0.103166:-0.0666591:0.0826137;
		specparam tpw_XR_negedge = 0.285077:0.37015:2.72095;
		specparam trecovery_XS_G_adacond2_posedge_adacond2_negedge = 0.435572:0.421428:0.240907;
		specparam tremoval_XS_G_adacond2_posedge_adacond2_negedge = -0.291822:-0.290285:-0.102117;
		specparam tsetup_XS_XR_NTB_G_posedge_NTB_G_posedge = 0.31568:0.395368:1.12735;
		specparam thold_XS_XR_NTB_G_posedge_NTB_G_posedge = -0.214334:-0.312232:-0.626628;
		specparam tpw_XS_negedge = 0.22751:0.338678:2.72095;
		specparam tpw_G_posedge = 0.381089:0.367527:2.72095;

		(D => Q) = ( tpd_D_Q_r , tpd_D_Q_f );
		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge G => (Q+:D)) = ( tpd_G_Q_posedge_r , tpd_G_Q_posedge_f );
		(D => XQ) = ( tpd_D_XQ_r , tpd_D_XQ_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge G => (XQ-:D)) = ( tpd_G_XQ_posedge_r , tpd_G_XQ_posedge_f );
		$setuphold (negedge G &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_G_adacond0_posedge_adacond0_negedge, 
			 thold_D_G_adacond0_posedge_adacond0_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (negedge G &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_G_adacond0_negedge_adacond0_negedge, 
			 thold_D_G_adacond0_negedge_adacond0_negedge, notifier,,, delayed_G, delayed_D);
		$setuphold (posedge XR &&& ~G, posedge XS &&& ~G, 
			 tsetup_XS_XR_NTB_G_posedge_NTB_G_posedge, 
			 thold_XS_XR_NTB_G_posedge_NTB_G_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond1, negedge G &&& adacond1, 
			 trecovery_XR_G_adacond1_posedge_adacond1_negedge, notifier);
		$hold (negedge G &&& adacond1, posedge XR &&& adacond1, 
			 tremoval_XR_G_adacond1_posedge_adacond1_negedge, notifier);
		$recovery (posedge XS &&& adacond2, negedge G &&& adacond2, 
			 trecovery_XS_G_adacond2_posedge_adacond2_negedge, notifier);
		$hold (negedge G &&& adacond2, posedge XS &&& adacond2, 
			 tremoval_XS_G_adacond2_posedge_adacond2_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge G, tpw_G_posedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: DLY1X1 
`timescale 1ns/10ps
`celldefine
module DLY1X1 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.167486:0.292718:1.46904;
		specparam tpd_A_Y_f = 0.172232:0.311331:1.61508;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: DLY2X1 
`timescale 1ns/10ps
`celldefine
module DLY2X1 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.384961:0.528768:1.76654;
		specparam tpd_A_Y_f = 0.377025:0.539444:1.89446;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: DLY3X1 
`timescale 1ns/10ps
`celldefine
module DLY3X1 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.591084:0.746823:2.01245;
		specparam tpd_A_Y_f = 0.556758:0.733458:2.12282;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: DLY4X1 
`timescale 1ns/10ps
`celldefine
module DLY4X1 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.908661:1.07652:2.35827;
		specparam tpd_A_Y_f = 0.820781:1.01104:2.42864;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: ENO 
`timescale 1ns/10ps
`celldefine
module ENOX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	and (int_fwire_0, C, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0621553:0.196194:1.73205;
		specparam tpd_A_Y_f = 0.0476174:0.144253:1.24337;
		specparam tpd_B_Y_r = 0.0847983:0.199018:1.55301;
		specparam tpd_B_Y_f = 0.0675662:0.17281:1.31402;
		specparam tpd_C_Y_r = 0.129466:0.214384:0.792363;
		specparam tpd_C_Y_f = 0.164295:0.280985:1.20163;
		specparam tpd_D_Y_r = 0.137611:0.211788:0.757275;
		specparam tpd_D_Y_f = 0.178473:0.299396:1.26105;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: ENO 
`timescale 1ns/10ps
`celldefine
module ENOXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	and (int_fwire_0, C, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0878802:0.224907:1.79633;
		specparam tpd_A_Y_f = 0.0580272:0.142941:1.09711;
		specparam tpd_B_Y_r = 0.118387:0.238668:1.6226;
		specparam tpd_B_Y_f = 0.0878563:0.182251:1.21126;
		specparam tpd_C_Y_r = 0.158502:0.23534:0.732617;
		specparam tpd_C_Y_f = 0.225914:0.346637:1.32783;
		specparam tpd_D_Y_r = 0.173563:0.239815:0.70759;
		specparam tpd_D_Y_f = 0.243718:0.366889:1.38706;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: EOR 
`timescale 1ns/10ps
`celldefine
module EORX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	not (B__bar, B);
	and (int_fwire_0, B__bar, D);
	and (int_fwire_1, B__bar, C);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D);
	and (int_fwire_3, A__bar, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.050624:0.182485:1.69289;
		specparam tpd_A_Y_f = 0.0582798:0.174424:1.5378;
		specparam tpd_B_Y_r = 0.0621934:0.195386:1.70675;
		specparam tpd_B_Y_f = 0.0679338:0.173423:1.45038;
		specparam tpd_C_Y_r = 0.15285:0.265491:1.25443;
		specparam tpd_C_Y_f = 0.180877:0.28639:1.11666;
		specparam tpd_D_Y_r = 0.171337:0.294491:1.35626;
		specparam tpd_D_Y_f = 0.205291:0.294952:1.06349;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: EOR 
`timescale 1ns/10ps
`celldefine
module EORXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1, int_fwire_2, int_fwire_3;

	not (B__bar, B);
	and (int_fwire_0, B__bar, D);
	and (int_fwire_1, B__bar, C);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D);
	and (int_fwire_3, A__bar, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0826786:0.220732:1.78896;
		specparam tpd_A_Y_f = 0.0619157:0.141433:1.03588;
		specparam tpd_B_Y_r = 0.100073:0.235576:1.78559;
		specparam tpd_B_Y_f = 0.0720464:0.138671:0.931678;
		specparam tpd_C_Y_r = 0.241434:0.345997:1.32926;
		specparam tpd_C_Y_f = 0.166972:0.255084:0.882269;
		specparam tpd_D_Y_r = 0.266879:0.37787:1.41945;
		specparam tpd_D_Y_f = 0.191106:0.266118:0.839839;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: FAD1 
`timescale 1ns/10ps
`celldefine
module FAD1X1 (CO, SO, A, B, CI);
	output CO, SO;
	input A, B, CI;

	// Function
	wire A__bar, B__bar, CI__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6;

	and (int_fwire_0, B, CI);
	and (int_fwire_1, A, CI);
	and (int_fwire_2, A, B);
	or (CO, int_fwire_2, int_fwire_1, int_fwire_0);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_3, A__bar, B__bar, CI);
	not (CI__bar, CI);
	and (int_fwire_4, A__bar, B, CI__bar);
	and (int_fwire_5, A, B__bar, CI__bar);
	and (int_fwire_6, A, B, CI);
	or (SO, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3);

	// Timing
	specify
		specparam tpd_A_CO_r = 0.189865:0.346561:1.655;
		specparam tpd_A_CO_f = 0.257513:0.450782:2.08124;
		specparam tpd_B_CO_r = 0.183531:0.325904:1.57764;
		specparam tpd_B_CO_f = 0.275114:0.455007:1.97103;
		specparam tpd_CI_CO_r = 0.16967:0.327506:1.61596;
		specparam tpd_CI_CO_f = 0.215592:0.425873:2.04678;
		specparam tpd_A_SO_posedge_r = 0.206133:0.346067:1.61542;
		specparam tpd_A_SO_posedge_f = 0.322489:0.493913:1.92579;
		specparam tpd_A_SO_negedge_r = 0.369679:0.525274:2.05511;
		specparam tpd_A_SO_negedge_f = 0.334074:0.503889:1.70679;
		specparam tpd_B_SO_posedge_r = 0.212515:0.340483:1.53957;
		specparam tpd_B_SO_posedge_f = 0.345823:0.514547:1.82944;
		specparam tpd_B_SO_negedge_r = 0.408505:0.55335:1.95064;
		specparam tpd_B_SO_negedge_f = 0.32855:0.486283:1.62605;
		specparam tpd_CI_SO_posedge_r = 0.21075:0.361761:1.67159;
		specparam tpd_CI_SO_posedge_f = 0.272908:0.455706:1.96989;
		specparam tpd_CI_SO_negedge_r = 0.383232:0.539922:2.02397;
		specparam tpd_CI_SO_negedge_f = 0.326472:0.47992:1.63369;

		(A => CO) = ( tpd_A_CO_r , tpd_A_CO_f );
		(B => CO) = ( tpd_B_CO_r , tpd_B_CO_f );
		(CI => CO) = ( tpd_CI_CO_r , tpd_CI_CO_f );
		(posedge A => (SO:A)) = ( tpd_A_SO_posedge_r , tpd_A_SO_posedge_f );
		(negedge A => (SO:A)) = ( tpd_A_SO_negedge_r , tpd_A_SO_negedge_f );
		(posedge B => (SO:B)) = ( tpd_B_SO_posedge_r , tpd_B_SO_posedge_f );
		(negedge B => (SO:B)) = ( tpd_B_SO_negedge_r , tpd_B_SO_negedge_f );
		(posedge CI => (SO:CI)) = ( tpd_CI_SO_posedge_r , tpd_CI_SO_posedge_f );
		(negedge CI => (SO:CI)) = ( tpd_CI_SO_negedge_r , tpd_CI_SO_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: FAD1 
`timescale 1ns/10ps
`celldefine
module FAD1XL (CO, SO, A, B, CI);
	output CO, SO;
	input A, B, CI;

	// Function
	wire A__bar, B__bar, CI__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6;

	and (int_fwire_0, B, CI);
	and (int_fwire_1, A, CI);
	and (int_fwire_2, A, B);
	or (CO, int_fwire_2, int_fwire_1, int_fwire_0);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_3, A__bar, B__bar, CI);
	not (CI__bar, CI);
	and (int_fwire_4, A__bar, B, CI__bar);
	and (int_fwire_5, A, B__bar, CI__bar);
	and (int_fwire_6, A, B, CI);
	or (SO, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3);

	// Timing
	specify
		specparam tpd_A_CO_r = 0.237698:0.393572:1.65814;
		specparam tpd_A_CO_f = 0.385893:0.600649:2.48374;
		specparam tpd_B_CO_r = 0.240839:0.380538:1.55757;
		specparam tpd_B_CO_f = 0.406735:0.611896:2.34661;
		specparam tpd_CI_CO_r = 0.212938:0.370624:1.6142;
		specparam tpd_CI_CO_f = 0.307316:0.537013:2.40574;
		specparam tpd_A_SO_posedge_r = 0.250044:0.387542:1.59968;
		specparam tpd_A_SO_posedge_f = 0.472477:0.673504:2.38066;
		specparam tpd_A_SO_negedge_r = 0.532019:0.692907:2.35432;
		specparam tpd_A_SO_negedge_f = 0.452066:0.631372:1.96629;
		specparam tpd_B_SO_posedge_r = 0.257241:0.379862:1.50684;
		specparam tpd_B_SO_posedge_f = 0.498791:0.698404:2.27843;
		specparam tpd_B_SO_negedge_r = 0.555607:0.706934:2.21559;
		specparam tpd_B_SO_negedge_f = 0.445563:0.608935:1.85778;
		specparam tpd_CI_SO_posedge_r = 0.255252:0.408077:1.68368;
		specparam tpd_CI_SO_posedge_f = 0.406335:0.613962:2.43551;
		specparam tpd_CI_SO_negedge_r = 0.513775:0.678664:2.28668;
		specparam tpd_CI_SO_negedge_f = 0.446356:0.61204:1.89231;

		(A => CO) = ( tpd_A_CO_r , tpd_A_CO_f );
		(B => CO) = ( tpd_B_CO_r , tpd_B_CO_f );
		(CI => CO) = ( tpd_CI_CO_r , tpd_CI_CO_f );
		(posedge A => (SO:A)) = ( tpd_A_SO_posedge_r , tpd_A_SO_posedge_f );
		(negedge A => (SO:A)) = ( tpd_A_SO_negedge_r , tpd_A_SO_negedge_f );
		(posedge B => (SO:B)) = ( tpd_B_SO_posedge_r , tpd_B_SO_posedge_f );
		(negedge B => (SO:B)) = ( tpd_B_SO_negedge_r , tpd_B_SO_negedge_f );
		(posedge CI => (SO:CI)) = ( tpd_CI_SO_posedge_r , tpd_CI_SO_posedge_f );
		(negedge CI => (SO:CI)) = ( tpd_CI_SO_negedge_r , tpd_CI_SO_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: GA_AND2 
`timescale 1ns/10ps
`celldefine
module GA_AND2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	and (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.112389:0.238182:1.41292;
		specparam tpd_A_Y_f = 0.0992548:0.219382:1.14724;
		specparam tpd_B_Y_r = 0.122777:0.237215:1.37378;
		specparam tpd_B_Y_f = 0.113155:0.239825:1.21196;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_AND3 
`timescale 1ns/10ps
`celldefine
module GA_AND3 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	and (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.138649:0.282398:1.55632;
		specparam tpd_A_Y_f = 0.10064:0.233611:1.21821;
		specparam tpd_B_Y_r = 0.15681:0.288864:1.52979;
		specparam tpd_B_Y_f = 0.11482:0.253393:1.27956;
		specparam tpd_C_Y_r = 0.166956:0.290088:1.47794;
		specparam tpd_C_Y_f = 0.124008:0.266712:1.32627;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_AOI21 
`timescale 1ns/10ps
`celldefine
module GA_AOI21 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1;

	not (C__bar, C);
	not (A__bar, A);
	and (int_fwire_0, A__bar, C__bar);
	not (B__bar, B);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0944651:0.23074:1.77537;
		specparam tpd_A_Y_f = 0.0330363:0.0966387:0.764161;
		specparam tpd_B_Y_r = 0.117736:0.239415:1.60429;
		specparam tpd_B_Y_f = 0.0662446:0.158045:1.05932;
		specparam tpd_C_Y_r = 0.140567:0.26229:1.61075;
		specparam tpd_C_Y_f = 0.0773713:0.158523:0.977469;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_AOI211 
`timescale 1ns/10ps
`celldefine
module GA_AOI211 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, D__bar);
	not (C__bar, C);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.138443:0.26751:1.75751;
		specparam tpd_A_Y_f = 0.0357636:0.0900617:0.568741;
		specparam tpd_B_Y_r = 0.208681:0.32109:1.68134;
		specparam tpd_B_Y_f = 0.0432963:0.106216:0.576951;
		specparam tpd_C_Y_r = 0.215834:0.331246:1.53412;
		specparam tpd_C_Y_f = 0.0707506:0.155408:0.821354;
		specparam tpd_D_Y_r = 0.251741:0.367789:1.55792;
		specparam tpd_D_Y_f = 0.0820782:0.155117:0.756258;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_AOI22 
`timescale 1ns/10ps
`celldefine
module GA_AOI22 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2, int_fwire_3;

	not (D__bar, D);
	not (B__bar, B);
	and (int_fwire_0, B__bar, D__bar);
	not (C__bar, C);
	and (int_fwire_1, B__bar, C__bar);
	not (A__bar, A);
	and (int_fwire_2, A__bar, D__bar);
	and (int_fwire_3, A__bar, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0915408:0.226336:1.75362;
		specparam tpd_A_Y_f = 0.0467752:0.128565:1.019;
		specparam tpd_B_Y_r = 0.114769:0.248117:1.76386;
		specparam tpd_B_Y_f = 0.0577792:0.130912:0.939415;
		specparam tpd_C_Y_r = 0.155258:0.279891:1.62949;
		specparam tpd_C_Y_f = 0.0876289:0.180243:1.08533;
		specparam tpd_D_Y_r = 0.177218:0.30191:1.63395;
		specparam tpd_D_Y_f = 0.0986491:0.180548:1.00115;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_BUF1 
`timescale 1ns/10ps
`celldefine
module GA_BUF1 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0803561:0.194611:1.30144;
		specparam tpd_A_Y_f = 0.0910007:0.207701:1.15341;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_BUF2 
`timescale 1ns/10ps
`celldefine
module GA_BUF2 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0793888:0.207333:1.3512;
		specparam tpd_A_Y_f = 0.0980582:0.231034:1.21515;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_BUF3 
`timescale 1ns/10ps
`celldefine
module GA_BUF3 (Y, A);
	output Y;
	input A;

	// Function
	buf (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0924664:0.228766:1.39927;
		specparam tpd_A_Y_f = 0.11853:0.260249:1.28789;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_INV1 
`timescale 1ns/10ps
`celldefine
module GA_INV1 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0331168:0.175595:1.79224;
		specparam tpd_A_Y_f = 0.0258209:0.123408:1.29238;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_INV2 
`timescale 1ns/10ps
`celldefine
module GA_INV2 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0296568:0.17147:1.78212;
		specparam tpd_A_Y_f = 0.0228558:0.11689:1.25606;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_INV3 
`timescale 1ns/10ps
`celldefine
module GA_INV3 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0306664:0.172553:1.78175;
		specparam tpd_A_Y_f = 0.0235072:0.11693:1.24676;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_INV4 
`timescale 1ns/10ps
`celldefine
module GA_INV4 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0295339:0.172133:1.79245;
		specparam tpd_A_Y_f = 0.0227694:0.11751:1.26423;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_NAND2 
`timescale 1ns/10ps
`celldefine
module GA_NAND2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0391302:0.178205:1.7518;
		specparam tpd_A_Y_f = 0.0407234:0.164492:1.64096;
		specparam tpd_B_Y_r = 0.0506362:0.194251:1.79262;
		specparam tpd_B_Y_f = 0.0510956:0.160396:1.5119;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_NAND3 
`timescale 1ns/10ps
`celldefine
module GA_NAND3 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0480221:0.172038:1.53663;
		specparam tpd_A_Y_f = 0.0641664:0.190756:1.70603;
		specparam tpd_B_Y_r = 0.0603792:0.188384:1.57458;
		specparam tpd_B_Y_f = 0.0823095:0.19607:1.62228;
		specparam tpd_C_Y_r = 0.0677823:0.198408:1.58844;
		specparam tpd_C_Y_f = 0.0925232:0.196653:1.50263;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_NAND4 
`timescale 1ns/10ps
`celldefine
module GA_NAND4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0567308:0.167513:1.32002;
		specparam tpd_A_Y_f = 0.0944483:0.214606:1.67457;
		specparam tpd_B_Y_r = 0.0700056:0.184079:1.35739;
		specparam tpd_B_Y_f = 0.121161:0.229601:1.6162;
		specparam tpd_C_Y_r = 0.0784567:0.194686:1.37311;
		specparam tpd_C_Y_f = 0.13926:0.23941:1.52276;
		specparam tpd_D_Y_r = 0.0816699:0.199214:1.36655;
		specparam tpd_D_Y_f = 0.14982:0.247905:1.45192;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_NOR2 
`timescale 1ns/10ps
`celldefine
module GA_NOR2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0620126:0.200455:1.7668;
		specparam tpd_A_Y_f = 0.0299098:0.0926656:0.794071;
		specparam tpd_B_Y_r = 0.0940771:0.214027:1.61256;
		specparam tpd_B_Y_f = 0.035988:0.107701:0.793488;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_NOR3 
`timescale 1ns/10ps
`celldefine
module GA_NOR3 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.101699:0.234387:1.75252;
		specparam tpd_A_Y_f = 0.0355421:0.0893575:0.571417;
		specparam tpd_B_Y_r = 0.172909:0.287441:1.67735;
		specparam tpd_B_Y_f = 0.0428696:0.105385:0.57939;
		specparam tpd_C_Y_r = 0.201678:0.314427:1.55091;
		specparam tpd_C_Y_f = 0.0418995:0.111895:0.604772;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_NOR4 
`timescale 1ns/10ps
`celldefine
module GA_NOR4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.148071:0.275973:1.74924;
		specparam tpd_A_Y_f = 0.0412576:0.0931306:0.443083;
		specparam tpd_B_Y_r = 0.258066:0.365342:1.72535;
		specparam tpd_B_Y_f = 0.049258:0.109257:0.456098;
		specparam tpd_C_Y_r = 0.323844:0.432258:1.64906;
		specparam tpd_C_Y_f = 0.0491629:0.116358:0.483635;
		specparam tpd_D_Y_r = 0.351364:0.458678:1.56951;
		specparam tpd_D_Y_f = 0.049117:0.121061:0.527682;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_OAI21 
`timescale 1ns/10ps
`celldefine
module GA_OAI21 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0;

	not (C__bar, C);
	not (B__bar, B);
	and (int_fwire_0, B__bar, C__bar);
	not (A__bar, A);
	or (Y, A__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.045229:0.147433:1.21395;
		specparam tpd_A_Y_f = 0.0611276:0.151951:1.05923;
		specparam tpd_B_Y_r = 0.110684:0.244931:1.78166;
		specparam tpd_B_Y_f = 0.061433:0.133149:0.913636;
		specparam tpd_C_Y_r = 0.1405:0.258583:1.61057;
		specparam tpd_C_Y_f = 0.0790078:0.159155:0.97355;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_OAI211 
`timescale 1ns/10ps
`celldefine
module GA_OAI211 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0494433:0.149574:1.17379;
		specparam tpd_A_Y_f = 0.0928736:0.194019:1.29022;
		specparam tpd_B_Y_r = 0.0620773:0.167194:1.21214;
		specparam tpd_B_Y_f = 0.111652:0.199966:1.20239;
		specparam tpd_C_Y_r = 0.139554:0.271367:1.77719;
		specparam tpd_C_Y_f = 0.100806:0.178341:1.03204;
		specparam tpd_D_Y_r = 0.168724:0.286455:1.60921;
		specparam tpd_D_Y_f = 0.128447:0.211941:1.10054;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_OAI22 
`timescale 1ns/10ps
`celldefine
module GA_OAI22 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0874837:0.215328:1.65425;
		specparam tpd_A_Y_f = 0.070138:0.158885:1.00494;
		specparam tpd_B_Y_r = 0.128738:0.241594:1.49733;
		specparam tpd_B_Y_f = 0.0929489:0.184293:1.04392;
		specparam tpd_C_Y_r = 0.138133:0.266197:1.73457;
		specparam tpd_C_Y_f = 0.0939393:0.172389:0.910545;
		specparam tpd_D_Y_r = 0.167425:0.280203:1.5703;
		specparam tpd_D_Y_f = 0.113393:0.192562:0.939053;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_OR2 
`timescale 1ns/10ps
`celldefine
module GA_OR2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0866586:0.204434:1.26716;
		specparam tpd_A_Y_f = 0.150998:0.288294:1.36218;
		specparam tpd_B_Y_r = 0.0965313:0.22295:1.3314;
		specparam tpd_B_Y_f = 0.18255:0.302612:1.31184;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GA_OR3 
`timescale 1ns/10ps
`celldefine
module GA_OR3 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.083584:0.210411:1.26898;
		specparam tpd_A_Y_f = 0.203997:0.367876:1.60895;
		specparam tpd_B_Y_r = 0.0941384:0.22774:1.32184;
		specparam tpd_B_Y_f = 0.274984:0.421115:1.5947;
		specparam tpd_C_Y_r = 0.0966004:0.237524:1.3786;
		specparam tpd_C_Y_f = 0.303792:0.44812:1.51296;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GEN2 
`timescale 1ns/10ps
`celldefine
module GEN2X1 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, B, D, E);
	and (int_fwire_1, B, C);
	or (Y, A, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0840938:0.224963:1.34169;
		specparam tpd_A_Y_f = 0.235028:0.41931:1.90064;
		specparam tpd_B_Y_r = 0.212715:0.36955:1.71654;
		specparam tpd_B_Y_f = 0.210579:0.367513:1.61937;
		specparam tpd_C_Y_r = 0.16583:0.302135:1.47155;
		specparam tpd_C_Y_f = 0.330746:0.49973:1.87755;
		specparam tpd_D_Y_r = 0.247375:0.39667:1.70172;
		specparam tpd_D_Y_f = 0.348902:0.515039:1.74206;
		specparam tpd_E_Y_r = 0.254403:0.390192:1.6033;
		specparam tpd_E_Y_f = 0.371142:0.541731:1.79526;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GEN2 
`timescale 1ns/10ps
`celldefine
module GEN2XL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, B, D, E);
	and (int_fwire_1, B, C);
	or (Y, A, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.103629:0.246153:1.33112;
		specparam tpd_A_Y_f = 0.334057:0.54875:2.35781;
		specparam tpd_B_Y_r = 0.246965:0.407969:1.73606;
		specparam tpd_B_Y_f = 0.287437:0.469595:2.00476;
		specparam tpd_C_Y_r = 0.200963:0.334281:1.45854;
		specparam tpd_C_Y_f = 0.460833:0.661289:2.32467;
		specparam tpd_D_Y_r = 0.29453:0.44639:1.71751;
		specparam tpd_D_Y_f = 0.485443:0.684585:2.19069;
		specparam tpd_E_Y_r = 0.30269:0.437932:1.60058;
		specparam tpd_E_Y_f = 0.515426:0.72016:2.25347;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GEN3 
`timescale 1ns/10ps
`celldefine
module GEN3X1 (Y, A, B, C, D, E, F, G);
	output Y;
	input A, B, C, D, E, F, G;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	and (int_fwire_0, B, D, F, G);
	and (int_fwire_1, B, D, E);
	and (int_fwire_2, B, C);
	or (Y, A, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0889656:0.24029:1.39785;
		specparam tpd_A_Y_f = 0.331874:0.524545:1.98023;
		specparam tpd_B_Y_r = 0.305244:0.476503:1.93249;
		specparam tpd_B_Y_f = 0.210185:0.363802:1.50761;
		specparam tpd_C_Y_r = 0.198448:0.343687:1.53224;
		specparam tpd_C_Y_f = 0.476532:0.652479:1.98875;
		specparam tpd_D_Y_r = 0.363002:0.52368:1.90152;
		specparam tpd_D_Y_f = 0.378841:0.540394:1.64824;
		specparam tpd_E_Y_r = 0.28951:0.436824:1.61734;
		specparam tpd_E_Y_f = 0.565559:0.74333:1.96714;
		specparam tpd_F_Y_r = 0.397811:0.556652:1.85088;
		specparam tpd_F_Y_f = 0.572836:0.747233:1.86102;
		specparam tpd_G_Y_r = 0.406144:0.554935:1.753;
		specparam tpd_G_Y_f = 0.603765:0.783229:1.91947;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
	endspecify
endmodule
`endcelldefine

// type: GEN3 
`timescale 1ns/10ps
`celldefine
module GEN3XL (Y, A, B, C, D, E, F, G);
	output Y;
	input A, B, C, D, E, F, G;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	and (int_fwire_0, B, D, F, G);
	and (int_fwire_1, B, D, E);
	and (int_fwire_2, B, C);
	or (Y, A, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.109477:0.264577:1.41342;
		specparam tpd_A_Y_f = 0.523828:0.766343:2.69868;
		specparam tpd_B_Y_r = 0.33405:0.515597:1.96855;
		specparam tpd_B_Y_f = 0.299531:0.489012:2.04042;
		specparam tpd_C_Y_r = 0.242885:0.38602:1.52838;
		specparam tpd_C_Y_f = 0.733154:0.959427:2.72227;
		specparam tpd_D_Y_r = 0.413304:0.581646:1.92847;
		specparam tpd_D_Y_f = 0.549397:0.752964:2.27651;
		specparam tpd_E_Y_r = 0.346397:0.497173:1.6397;
		specparam tpd_E_Y_f = 0.846561:1.07412:2.70862;
		specparam tpd_F_Y_r = 0.470287:0.639001:1.91011;
		specparam tpd_F_Y_f = 0.858278:1.08378:2.61283;
		specparam tpd_G_Y_r = 0.478177:0.631822:1.79576;
		specparam tpd_G_Y_f = 0.894995:1.12685:2.67707;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
	endspecify
endmodule
`endcelldefine

// type: HAD1 
`timescale 1ns/10ps
`celldefine
module HAD1X1 (CO, SO, A, B);
	output CO, SO;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	and (CO, A, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (SO, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_CO_r = 0.093761:0.224303:1.40473;
		specparam tpd_A_CO_f = 0.0966431:0.243877:1.49553;
		specparam tpd_B_CO_r = 0.101894:0.220967:1.36211;
		specparam tpd_B_CO_f = 0.110002:0.263852:1.55902;
		specparam tpd_A_SO_posedge_r = 0.0961328:0.231365:1.37493;
		specparam tpd_A_SO_posedge_f = 0.134929:0.305743:1.66577;
		specparam tpd_A_SO_negedge_r = 0.136597:0.293844:1.62958;
		specparam tpd_A_SO_negedge_f = 0.137334:0.293382:1.35429;
		specparam tpd_B_SO_posedge_r = 0.151956:0.302525:1.54751;
		specparam tpd_B_SO_posedge_f = 0.194393:0.377639:1.77088;
		specparam tpd_B_SO_negedge_r = 0.212819:0.371533:1.76848;
		specparam tpd_B_SO_negedge_f = 0.201064:0.343973:1.36067;

		(A => CO) = ( tpd_A_CO_r , tpd_A_CO_f );
		(B => CO) = ( tpd_B_CO_r , tpd_B_CO_f );
		(posedge A => (SO:A)) = ( tpd_A_SO_posedge_r , tpd_A_SO_posedge_f );
		(negedge A => (SO:A)) = ( tpd_A_SO_negedge_r , tpd_A_SO_negedge_f );
		(posedge B => (SO:B)) = ( tpd_B_SO_posedge_r , tpd_B_SO_posedge_f );
		(negedge B => (SO:B)) = ( tpd_B_SO_negedge_r , tpd_B_SO_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: HAD1 
`timescale 1ns/10ps
`celldefine
module HAD1XL (CO, SO, A, B);
	output CO, SO;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	and (CO, A, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (SO, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_CO_r = 0.103497:0.233025:1.36985;
		specparam tpd_A_CO_f = 0.131575:0.305822:1.85654;
		specparam tpd_B_CO_r = 0.111942:0.229086:1.32504;
		specparam tpd_B_CO_f = 0.150498:0.329717:1.92639;
		specparam tpd_A_SO_posedge_r = 0.107826:0.245845:1.41895;
		specparam tpd_A_SO_posedge_f = 0.139428:0.314794:1.77335;
		specparam tpd_A_SO_negedge_r = 0.161464:0.329593:1.6993;
		specparam tpd_A_SO_negedge_f = 0.155265:0.320122:1.49793;
		specparam tpd_B_SO_posedge_r = 0.211961:0.364168:1.65921;
		specparam tpd_B_SO_posedge_f = 0.202506:0.391859:1.89789;
		specparam tpd_B_SO_negedge_r = 0.242284:0.405394:1.81742;
		specparam tpd_B_SO_negedge_f = 0.250388:0.399934:1.55567;

		(A => CO) = ( tpd_A_CO_r , tpd_A_CO_f );
		(B => CO) = ( tpd_B_CO_r , tpd_B_CO_f );
		(posedge A => (SO:A)) = ( tpd_A_SO_posedge_r , tpd_A_SO_posedge_f );
		(negedge A => (SO:A)) = ( tpd_A_SO_negedge_r , tpd_A_SO_negedge_f );
		(posedge B => (SO:B)) = ( tpd_B_SO_posedge_r , tpd_B_SO_posedge_f );
		(negedge B => (SO:B)) = ( tpd_B_SO_negedge_r , tpd_B_SO_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX1 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0271877:0.166065:1.76444;
		specparam tpd_A_Y_f = 0.0302736:0.172223:1.83456;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX12 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.178452:0.334779:1.77654;
		specparam tpd_A_Y_f = 0.152808:0.263743:0.88022;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX16 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.178307:0.333818:1.7507;
		specparam tpd_A_Y_f = 0.170371:0.287554:0.961082;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX2 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0253146:0.163266:1.75581;
		specparam tpd_A_Y_f = 0.027049:0.164844:1.7739;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX20 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.185999:0.341975:1.74467;
		specparam tpd_A_Y_f = 0.187922:0.308966:0.971819;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX24 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.211601:0.371176:1.82888;
		specparam tpd_A_Y_f = 0.180324:0.299991:0.950213;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX3 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0259091:0.166424:1.77724;
		specparam tpd_A_Y_f = 0.0230836:0.135292:1.468;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX30 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.22372:0.38486:1.84092;
		specparam tpd_A_Y_f = 0.199075:0.322846:0.978895;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX36 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.234823:0.398641:1.86699;
		specparam tpd_A_Y_f = 0.217262:0.345204:1.01712;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX4 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0258887:0.166516:1.77769;
		specparam tpd_A_Y_f = 0.0226206:0.133148:1.44944;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX6 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0262289:0.167181:1.78181;
		specparam tpd_A_Y_f = 0.022627:0.131664:1.43278;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVX8 (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0261023:0.167261:1.78308;
		specparam tpd_A_Y_f = 0.0223497:0.130266:1.42016;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: INV 
`timescale 1ns/10ps
`celldefine
module INVXL (Y, A);
	output Y;
	input A;

	// Function
	not (Y, A);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0343997:0.178848:1.81416;
		specparam tpd_A_Y_f = 0.0287987:0.134807:1.40089;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
	endspecify
endmodule
`endcelldefine

// type: MAJ3 
`timescale 1ns/10ps
`celldefine
module MAJ3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	and (int_fwire_0, B, C);
	and (int_fwire_1, A, C);
	and (int_fwire_2, A, B);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.133086:0.276913:1.48268;
		specparam tpd_A_Y_f = 0.149527:0.336995:1.75832;
		specparam tpd_B_Y_r = 0.154926:0.300579:1.54581;
		specparam tpd_B_Y_f = 0.185603:0.353628:1.75452;
		specparam tpd_C_Y_r = 0.149699:0.281969:1.48696;
		specparam tpd_C_Y_f = 0.204011:0.357167:1.67342;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: MAJ3 
`timescale 1ns/10ps
`celldefine
module MAJ3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	and (int_fwire_0, B, C);
	and (int_fwire_1, A, C);
	and (int_fwire_2, A, B);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.166188:0.312916:1.49822;
		specparam tpd_A_Y_f = 0.216582:0.427845:2.13857;
		specparam tpd_B_Y_r = 0.191502:0.337095:1.56565;
		specparam tpd_B_Y_f = 0.288897:0.482654:2.19181;
		specparam tpd_C_Y_r = 0.195181:0.328045:1.49295;
		specparam tpd_C_Y_f = 0.310169:0.493145:2.08095;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2A 
`timescale 1ns/10ps
`celldefine
module MUX2AX1 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D0__bar, int_fwire_0, int_fwire_1;
	wire S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	not (D0__bar, D0);
	and (int_fwire_1, D0__bar, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.193745:0.319913:1.54039;
		specparam tpd_D0_Y_f = 0.260499:0.435641:1.93078;
		specparam tpd_D1_Y_r = 0.153742:0.28757:1.49803;
		specparam tpd_D1_Y_f = 0.212042:0.388917:1.97313;
		specparam tpd_S_Y_posedge_r = 0.146032:0.294992:1.56078;
		specparam tpd_S_Y_posedge_f = 0.198551:0.369753:1.92069;
		specparam tpd_S_Y_negedge_r = 0.169845:0.309066:1.60212;
		specparam tpd_S_Y_negedge_f = 0.244314:0.409997:1.81802;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2A 
`timescale 1ns/10ps
`celldefine
module MUX2AX2 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D0__bar, int_fwire_0, int_fwire_1;
	wire S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	not (D0__bar, D0);
	and (int_fwire_1, D0__bar, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.202014:0.336496:1.6141;
		specparam tpd_D0_Y_f = 0.274442:0.448972:1.78606;
		specparam tpd_D1_Y_r = 0.164713:0.308402:1.56063;
		specparam tpd_D1_Y_f = 0.242386:0.42216:1.89821;
		specparam tpd_S_Y_posedge_r = 0.155098:0.312443:1.61456;
		specparam tpd_S_Y_posedge_f = 0.227579:0.402781:1.85586;
		specparam tpd_S_Y_negedge_r = 0.176387:0.324778:1.68918;
		specparam tpd_S_Y_negedge_f = 0.25722:0.419708:1.64932;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2A 
`timescale 1ns/10ps
`celldefine
module MUX2AX4 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D0__bar, int_fwire_0, int_fwire_1;
	wire S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	not (D0__bar, D0);
	and (int_fwire_1, D0__bar, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.250533:0.390784:1.66019;
		specparam tpd_D0_Y_f = 0.340844:0.501957:1.53378;
		specparam tpd_D1_Y_r = 0.224594:0.375469:1.67361;
		specparam tpd_D1_Y_f = 0.278794:0.439863:1.60421;
		specparam tpd_S_Y_posedge_r = 0.213833:0.377632:1.71872;
		specparam tpd_S_Y_posedge_f = 0.28991:0.454054:1.64764;
		specparam tpd_S_Y_negedge_r = 0.22441:0.379635:1.73365;
		specparam tpd_S_Y_negedge_f = 0.30456:0.452755:1.37369;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2A 
`timescale 1ns/10ps
`celldefine
module MUX2AXL (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D0__bar, int_fwire_0, int_fwire_1;
	wire S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	not (D0__bar, D0);
	and (int_fwire_1, D0__bar, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.226749:0.357924:1.65609;
		specparam tpd_D0_Y_f = 0.294678:0.444921:1.57601;
		specparam tpd_D1_Y_r = 0.195432:0.32044:1.49605;
		specparam tpd_D1_Y_f = 0.264578:0.431182:1.79159;
		specparam tpd_S_Y_posedge_r = 0.186472:0.330604:1.57746;
		specparam tpd_S_Y_posedge_f = 0.247278:0.407989:1.73367;
		specparam tpd_S_Y_negedge_r = 0.200689:0.346272:1.72699;
		specparam tpd_S_Y_negedge_f = 0.282409:0.423754:1.46793;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2B 
`timescale 1ns/10ps
`celldefine
module MUX2BX1 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D1__bar, int_fwire_0, int_fwire_1;
	wire S__bar;

	not (D1__bar, D1);
	and (int_fwire_0, D1__bar, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.156743:0.288676:1.48318;
		specparam tpd_D0_Y_f = 0.22165:0.391619:1.94838;
		specparam tpd_D1_Y_r = 0.206624:0.370004:1.77938;
		specparam tpd_D1_Y_f = 0.18055:0.310899:1.55991;
		specparam tpd_S_Y_posedge_r = 0.140744:0.272746:1.45292;
		specparam tpd_S_Y_posedge_f = 0.197303:0.38251:2.00945;
		specparam tpd_S_Y_negedge_r = 0.206821:0.365472:1.72371;
		specparam tpd_S_Y_negedge_f = 0.172699:0.314177:1.60875;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2B 
`timescale 1ns/10ps
`celldefine
module MUX2BX2 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D1__bar, int_fwire_0, int_fwire_1;
	wire S__bar;

	not (D1__bar, D1);
	and (int_fwire_0, D1__bar, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.175243:0.319615:1.56694;
		specparam tpd_D0_Y_f = 0.260202:0.441368:1.98873;
		specparam tpd_D1_Y_r = 0.22476:0.398891:1.83933;
		specparam tpd_D1_Y_f = 0.199259:0.336374:1.55354;
		specparam tpd_S_Y_posedge_r = 0.156298:0.299257:1.52023;
		specparam tpd_S_Y_posedge_f = 0.23591:0.43196:2.07598;
		specparam tpd_S_Y_negedge_r = 0.224768:0.395963:1.78611;
		specparam tpd_S_Y_negedge_f = 0.190722:0.339188:1.60189;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2B 
`timescale 1ns/10ps
`celldefine
module MUX2BX4 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D1__bar, int_fwire_0, int_fwire_1;
	wire S__bar;

	not (D1__bar, D1);
	and (int_fwire_0, D1__bar, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.234367:0.388612:1.67017;
		specparam tpd_D0_Y_f = 0.342723:0.511802:1.76;
		specparam tpd_D1_Y_r = 0.28463:0.467922:1.89817;
		specparam tpd_D1_Y_f = 0.23897:0.36399:1.23396;
		specparam tpd_S_Y_posedge_r = 0.21527:0.369813:1.63265;
		specparam tpd_S_Y_posedge_f = 0.319186:0.502026:1.87509;
		specparam tpd_S_Y_negedge_r = 0.282739:0.462983:1.84341;
		specparam tpd_S_Y_negedge_f = 0.230318:0.367035:1.27903;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2B 
`timescale 1ns/10ps
`celldefine
module MUX2BXL (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D1__bar, int_fwire_0, int_fwire_1;
	wire S__bar;

	not (D1__bar, D1);
	and (int_fwire_0, D1__bar, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.212995:0.336488:1.48437;
		specparam tpd_D0_Y_f = 0.288382:0.443118:1.75047;
		specparam tpd_D1_Y_r = 0.282361:0.452835:1.9903;
		specparam tpd_D1_Y_f = 0.215036:0.31978:1.17294;
		specparam tpd_S_Y_posedge_r = 0.189718:0.312762:1.43454;
		specparam tpd_S_Y_posedge_f = 0.258624:0.425221:1.84186;
		specparam tpd_S_Y_negedge_r = 0.284537:0.453001:1.93689;
		specparam tpd_S_Y_negedge_f = 0.205738:0.32224:1.2225;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2I 
`timescale 1ns/10ps
`celldefine
module MUX2IX1 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D0__bar, D1__bar, int_fwire_0;
	wire int_fwire_1, S__bar;

	not (D1__bar, D1);
	and (int_fwire_0, D1__bar, S);
	not (S__bar, S);
	not (D0__bar, D0);
	and (int_fwire_1, D0__bar, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.088133:0.211569:1.46149;
		specparam tpd_D0_Y_f = 0.0818684:0.177844:1.1409;
		specparam tpd_D1_Y_r = 0.0942601:0.220206:1.51958;
		specparam tpd_D1_Y_f = 0.0799352:0.177223:1.15335;
		specparam tpd_S_Y_posedge_r = 0.0802948:0.187095:1.21442;
		specparam tpd_S_Y_posedge_f = 0.0812873:0.182542:0.977584;
		specparam tpd_S_Y_negedge_r = 0.0577521:0.180109:1.23335;
		specparam tpd_S_Y_negedge_f = 0.0464318:0.138141:0.997869;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2I 
`timescale 1ns/10ps
`celldefine
module MUX2IX2 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D0__bar, D1__bar, int_fwire_0;
	wire int_fwire_1, S__bar;

	not (D1__bar, D1);
	and (int_fwire_0, D1__bar, S);
	not (S__bar, S);
	not (D0__bar, D0);
	and (int_fwire_1, D0__bar, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.0874973:0.211435:1.47423;
		specparam tpd_D0_Y_f = 0.0861972:0.187153:1.21194;
		specparam tpd_D1_Y_r = 0.0909967:0.214958:1.47538;
		specparam tpd_D1_Y_f = 0.0824142:0.184779:1.2104;
		specparam tpd_S_Y_posedge_r = 0.0918677:0.20092:1.21476;
		specparam tpd_S_Y_posedge_f = 0.0967116:0.205459:1.07361;
		specparam tpd_S_Y_negedge_r = 0.0560801:0.185423:1.29165;
		specparam tpd_S_Y_negedge_f = 0.0476195:0.146629:1.05934;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2I 
`timescale 1ns/10ps
`celldefine
module MUX2IX4 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D0__bar, D1__bar, int_fwire_0;
	wire int_fwire_1, S__bar;

	not (D1__bar, D1);
	and (int_fwire_0, D1__bar, S);
	not (S__bar, S);
	not (D0__bar, D0);
	and (int_fwire_1, D0__bar, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.077394:0.200809:1.46743;
		specparam tpd_D0_Y_f = 0.0774617:0.178039:1.20809;
		specparam tpd_D1_Y_r = 0.0840456:0.206562:1.47339;
		specparam tpd_D1_Y_f = 0.0702539:0.173006:1.20565;
		specparam tpd_S_Y_posedge_r = 0.110753:0.223002:1.28634;
		specparam tpd_S_Y_posedge_f = 0.119354:0.233345:1.13938;
		specparam tpd_S_Y_negedge_r = 0.0555898:0.191417:1.33592;
		specparam tpd_S_Y_negedge_f = 0.0474188:0.149251:1.09366;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2I 
`timescale 1ns/10ps
`celldefine
module MUX2IXL (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire D0__bar, D1__bar, int_fwire_0;
	wire int_fwire_1, S__bar;

	not (D1__bar, D1);
	and (int_fwire_0, D1__bar, S);
	not (S__bar, S);
	not (D0__bar, D0);
	and (int_fwire_1, D0__bar, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.108274:0.237153:1.54653;
		specparam tpd_D0_Y_f = 0.103839:0.191519:1.10795;
		specparam tpd_D1_Y_r = 0.111202:0.241203:1.56324;
		specparam tpd_D1_Y_f = 0.0963027:0.178851:1.02195;
		specparam tpd_S_Y_posedge_r = 0.0780264:0.179335:1.12004;
		specparam tpd_S_Y_posedge_f = 0.0949219:0.200213:1.07623;
		specparam tpd_S_Y_negedge_r = 0.0751844:0.196608:1.28109;
		specparam tpd_S_Y_negedge_f = 0.0522259:0.132933:0.903439;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2 
`timescale 1ns/10ps
`celldefine
module MUX2X1 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire int_fwire_0, int_fwire_1, S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.146771:0.297478:1.54008;
		specparam tpd_D0_Y_f = 0.174415:0.368962:1.98046;
		specparam tpd_D1_Y_r = 0.145654:0.297372:1.53978;
		specparam tpd_D1_Y_f = 0.180238:0.375011:1.99153;
		specparam tpd_S_Y_posedge_r = 0.10682:0.249486:1.43256;
		specparam tpd_S_Y_posedge_f = 0.150232:0.33832:1.96643;
		specparam tpd_S_Y_negedge_r = 0.159248:0.331953:1.75318;
		specparam tpd_S_Y_negedge_f = 0.155374:0.333366:1.61677;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2 
`timescale 1ns/10ps
`celldefine
module MUX2X2 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire int_fwire_0, int_fwire_1, S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.144228:0.300942:1.56686;
		specparam tpd_D0_Y_f = 0.169737:0.359398:1.84919;
		specparam tpd_D1_Y_r = 0.142059:0.29827:1.53064;
		specparam tpd_D1_Y_f = 0.202839:0.406792:1.97817;
		specparam tpd_S_Y_posedge_r = 0.110453:0.260227:1.46416;
		specparam tpd_S_Y_posedge_f = 0.158379:0.346238:1.88872;
		specparam tpd_S_Y_negedge_r = 0.160581:0.338809:1.76809;
		specparam tpd_S_Y_negedge_f = 0.171375:0.35939:1.5578;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2 
`timescale 1ns/10ps
`celldefine
module MUX2X4 (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire int_fwire_0, int_fwire_1, S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.17831:0.347675:1.6714;
		specparam tpd_D0_Y_f = 0.217741:0.416404:1.88595;
		specparam tpd_D1_Y_r = 0.177062:0.346063:1.64168;
		specparam tpd_D1_Y_f = 0.258013:0.470958:2.02102;
		specparam tpd_S_Y_posedge_r = 0.146918:0.31041:1.58173;
		specparam tpd_S_Y_posedge_f = 0.211144:0.409411:1.95259;
		specparam tpd_S_Y_negedge_r = 0.18993:0.378828:1.83548;
		specparam tpd_S_Y_negedge_f = 0.223194:0.42037:1.58408;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX2 
`timescale 1ns/10ps
`celldefine
module MUX2XL (Y, D0, D1, S);
	output Y;
	input D0, D1, S;

	// Function
	wire int_fwire_0, int_fwire_1, S__bar;

	and (int_fwire_0, D1, S);
	not (S__bar, S);
	and (int_fwire_1, D0, S__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.180428:0.319123:1.50187;
		specparam tpd_D0_Y_f = 0.201218:0.389631:1.91518;
		specparam tpd_D1_Y_r = 0.178202:0.317266:1.50132;
		specparam tpd_D1_Y_f = 0.199046:0.386159:1.90484;
		specparam tpd_S_Y_posedge_r = 0.132804:0.270008:1.40317;
		specparam tpd_S_Y_posedge_f = 0.169936:0.350148:1.86268;
		specparam tpd_S_Y_negedge_r = 0.179033:0.348488:1.77243;
		specparam tpd_S_Y_negedge_f = 0.159985:0.323405:1.41551;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(posedge S => (Y:S)) = ( tpd_S_Y_posedge_r , tpd_S_Y_posedge_f );
		(negedge S => (Y:S)) = ( tpd_S_Y_negedge_r , tpd_S_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX3I 
`timescale 1ns/10ps
`celldefine
module MUX3IX1 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire D0__bar, D1__bar, D2__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	not (D2__bar, D2);
	and (int_fwire_0, D2__bar, S1);
	not (S1__bar, S1);
	not (D1__bar, D1);
	and (int_fwire_1, D1__bar, S0, S1__bar);
	not (S0__bar, S0);
	not (D0__bar, D0);
	and (int_fwire_2, D0__bar, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.361593:0.519075:1.97075;
		specparam tpd_D0_Y_f = 0.30012:0.448299:1.82457;
		specparam tpd_D1_Y_r = 0.343176:0.491888:1.86305;
		specparam tpd_D1_Y_f = 0.310603:0.462269:1.89171;
		specparam tpd_D2_Y_r = 0.205757:0.346511:1.65431;
		specparam tpd_D2_Y_f = 0.189756:0.335327:1.68931;
		specparam tpd_S0_Y_posedge_r = 0.333474:0.480766:1.63651;
		specparam tpd_S0_Y_posedge_f = 0.314143:0.484173:2.01521;
		specparam tpd_S0_Y_negedge_r = 0.351534:0.507849:2.00739;
		specparam tpd_S0_Y_negedge_f = 0.280667:0.429718:1.80492;
		specparam tpd_S1_Y_posedge_r = 0.202432:0.343505:1.47513;
		specparam tpd_S1_Y_posedge_f = 0.226017:0.392757:1.89811;
		specparam tpd_S1_Y_negedge_r = 0.228282:0.385611:1.89199;
		specparam tpd_S1_Y_negedge_f = 0.161787:0.302599:1.51406;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX3I 
`timescale 1ns/10ps
`celldefine
module MUX3IX2 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire D0__bar, D1__bar, D2__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	not (D2__bar, D2);
	and (int_fwire_0, D2__bar, S1);
	not (S1__bar, S1);
	not (D1__bar, D1);
	and (int_fwire_1, D1__bar, S0, S1__bar);
	not (S0__bar, S0);
	not (D0__bar, D0);
	and (int_fwire_2, D0__bar, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.382328:0.546903:2.01892;
		specparam tpd_D0_Y_f = 0.316416:0.466565:1.80086;
		specparam tpd_D1_Y_r = 0.363311:0.519127:1.90947;
		specparam tpd_D1_Y_f = 0.327319:0.481082:1.86763;
		specparam tpd_D2_Y_r = 0.221398:0.368176:1.6988;
		specparam tpd_D2_Y_f = 0.203005:0.350746:1.66354;
		specparam tpd_S0_Y_posedge_r = 0.353774:0.507984:1.68062;
		specparam tpd_S0_Y_posedge_f = 0.330468:0.50255:1.98772;
		specparam tpd_S0_Y_negedge_r = 0.372263:0.536017:2.05584;
		specparam tpd_S0_Y_negedge_f = 0.297436:0.448468:1.78338;
		specparam tpd_S1_Y_posedge_r = 0.218011:0.365038:1.51398;
		specparam tpd_S1_Y_posedge_f = 0.242382:0.411076:1.87;
		specparam tpd_S1_Y_negedge_r = 0.247862:0.411891:1.93906;
		specparam tpd_S1_Y_negedge_f = 0.175061:0.317993:1.48962;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX3I 
`timescale 1ns/10ps
`celldefine
module MUX3IX4 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire D0__bar, D1__bar, D2__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	not (D2__bar, D2);
	and (int_fwire_0, D2__bar, S1);
	not (S1__bar, S1);
	not (D1__bar, D1);
	and (int_fwire_1, D1__bar, S0, S1__bar);
	not (S0__bar, S0);
	not (D0__bar, D0);
	and (int_fwire_2, D0__bar, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.42313:0.594593:2.06734;
		specparam tpd_D0_Y_f = 0.351585:0.505979:1.80146;
		specparam tpd_D1_Y_r = 0.403424:0.565988:1.95778;
		specparam tpd_D1_Y_f = 0.363375:0.521313:1.86919;
		specparam tpd_D2_Y_r = 0.253378:0.406898:1.74074;
		specparam tpd_D2_Y_f = 0.233554:0.386119:1.66209;
		specparam tpd_S0_Y_posedge_r = 0.393827:0.554973:1.72486;
		specparam tpd_S0_Y_posedge_f = 0.365836:0.542216:1.98372;
		specparam tpd_S0_Y_negedge_r = 0.41347:0.584091:2.10645;
		specparam tpd_S0_Y_negedge_f = 0.333497:0.488733:1.78838;
		specparam tpd_S1_Y_posedge_r = 0.249942:0.403461:1.54989;
		specparam tpd_S1_Y_posedge_f = 0.277888:0.450867:1.86564;
		specparam tpd_S1_Y_negedge_r = 0.287431:0.458164:1.98547;
		specparam tpd_S1_Y_negedge_f = 0.205642:0.353332:1.48989;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX3I 
`timescale 1ns/10ps
`celldefine
module MUX3IXL (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire D0__bar, D1__bar, D2__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	not (D2__bar, D2);
	and (int_fwire_0, D2__bar, S1);
	not (S1__bar, S1);
	not (D1__bar, D1);
	and (int_fwire_1, D1__bar, S0, S1__bar);
	not (S0__bar, S0);
	not (D0__bar, D0);
	and (int_fwire_2, D0__bar, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.392725:0.553686:2.08751;
		specparam tpd_D0_Y_f = 0.348998:0.48065:1.59448;
		specparam tpd_D1_Y_r = 0.390736:0.551721:2.08412;
		specparam tpd_D1_Y_f = 0.341132:0.472522:1.57871;
		specparam tpd_D2_Y_r = 0.251488:0.408313:1.87352;
		specparam tpd_D2_Y_f = 0.224045:0.35213:1.37688;
		specparam tpd_S0_Y_posedge_r = 0.356333:0.500478:1.68685;
		specparam tpd_S0_Y_posedge_f = 0.347318:0.498739:1.74221;
		specparam tpd_S0_Y_negedge_r = 0.365128:0.51739:2.02075;
		specparam tpd_S0_Y_negedge_f = 0.304314:0.432327:1.50749;
		specparam tpd_S1_Y_posedge_r = 0.221839:0.359096:1.49435;
		specparam tpd_S1_Y_posedge_f = 0.240911:0.390651:1.62366;
		specparam tpd_S1_Y_negedge_r = 0.214709:0.372197:1.88346;
		specparam tpd_S1_Y_negedge_f = 0.183431:0.306314:1.24117;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX3 
`timescale 1ns/10ps
`celldefine
module MUX3X1 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	and (int_fwire_0, D2, S1);
	not (S1__bar, S1);
	and (int_fwire_1, D1, S0, S1__bar);
	not (S0__bar, S0);
	and (int_fwire_2, D0, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.234071:0.39592:1.6793;
		specparam tpd_D0_Y_f = 0.294475:0.518906:2.22486;
		specparam tpd_D1_Y_r = 0.244435:0.412284:1.75376;
		specparam tpd_D1_Y_f = 0.274066:0.485397:2.09936;
		specparam tpd_D2_Y_r = 0.131003:0.276932:1.53485;
		specparam tpd_D2_Y_f = 0.151466:0.329704:1.85623;
		specparam tpd_S0_Y_posedge_r = 0.214119:0.379145:1.6762;
		specparam tpd_S0_Y_posedge_f = 0.285065:0.509018:2.27339;
		specparam tpd_S0_Y_negedge_r = 0.248656:0.432851:1.85246;
		specparam tpd_S0_Y_negedge_f = 0.265905:0.476508:1.8548;
		specparam tpd_S1_Y_posedge_r = 0.102868:0.243498:1.36445;
		specparam tpd_S1_Y_posedge_f = 0.165772:0.38351:2.13963;
		specparam tpd_S1_Y_negedge_r = 0.161219:0.341678:1.73747;
		specparam tpd_S1_Y_negedge_f = 0.14832:0.32652:1.65303;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX3 
`timescale 1ns/10ps
`celldefine
module MUX3X2 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	and (int_fwire_0, D2, S1);
	not (S1__bar, S1);
	and (int_fwire_1, D1, S0, S1__bar);
	not (S0__bar, S0);
	and (int_fwire_2, D0, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.257757:0.429236:1.73343;
		specparam tpd_D0_Y_f = 0.332245:0.56126:2.20259;
		specparam tpd_D1_Y_r = 0.269511:0.44696:1.8087;
		specparam tpd_D1_Y_f = 0.309433:0.525311:2.0713;
		specparam tpd_D2_Y_r = 0.14644:0.302515:1.57906;
		specparam tpd_D2_Y_f = 0.173364:0.359478:1.81883;
		specparam tpd_S0_Y_posedge_r = 0.239502:0.414269:1.7413;
		specparam tpd_S0_Y_posedge_f = 0.323812:0.552594:2.25206;
		specparam tpd_S0_Y_negedge_r = 0.271661:0.465418:1.89176;
		specparam tpd_S0_Y_negedge_f = 0.30039:0.515538:1.82186;
		specparam tpd_S1_Y_posedge_r = 0.12083:0.275356:1.44489;
		specparam tpd_S1_Y_posedge_f = 0.207628:0.433301:2.13043;
		specparam tpd_S1_Y_negedge_r = 0.181669:0.373999:1.78121;
		specparam tpd_S1_Y_negedge_f = 0.167358:0.354735:1.60292;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX3 
`timescale 1ns/10ps
`celldefine
module MUX3X4 (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	and (int_fwire_0, D2, S1);
	not (S1__bar, S1);
	and (int_fwire_1, D1, S0, S1__bar);
	not (S0__bar, S0);
	and (int_fwire_2, D0, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.314617:0.498117:1.83759;
		specparam tpd_D0_Y_f = 0.432078:0.673692:2.37368;
		specparam tpd_D1_Y_r = 0.328992:0.518582:1.91344;
		specparam tpd_D1_Y_f = 0.408941:0.638401:2.24657;
		specparam tpd_D2_Y_r = 0.187029:0.356581:1.66765;
		specparam tpd_D2_Y_f = 0.234558:0.436839:1.95153;
		specparam tpd_S0_Y_posedge_r = 0.299833:0.486523:1.86291;
		specparam tpd_S0_Y_posedge_f = 0.424711:0.666157:2.42034;
		specparam tpd_S0_Y_negedge_r = 0.327401:0.532939:1.97051;
		specparam tpd_S0_Y_negedge_f = 0.397603:0.625944:1.9829;
		specparam tpd_S1_Y_posedge_r = 0.164118:0.33268:1.58197;
		specparam tpd_S1_Y_posedge_f = 0.319276:0.558084:2.31141;
		specparam tpd_S1_Y_negedge_r = 0.236022:0.441986:1.86901;
		specparam tpd_S1_Y_negedge_f = 0.225338:0.428624:1.72459;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX3 
`timescale 1ns/10ps
`celldefine
module MUX3XL (Y, D0, D1, D2, S0, S1);
	output Y;
	input D0, D1, D2, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire S0__bar, S1__bar;

	and (int_fwire_0, D2, S1);
	not (S1__bar, S1);
	and (int_fwire_1, D1, S0, S1__bar);
	not (S0__bar, S0);
	and (int_fwire_2, D0, S0__bar, S1__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.283902:0.435404:1.71239;
		specparam tpd_D0_Y_f = 0.31108:0.5074:1.94546;
		specparam tpd_D1_Y_r = 0.275761:0.426273:1.68927;
		specparam tpd_D1_Y_f = 0.309034:0.504608:1.9414;
		specparam tpd_D2_Y_r = 0.165812:0.303359:1.49519;
		specparam tpd_D2_Y_f = 0.184215:0.349805:1.66957;
		specparam tpd_S0_Y_posedge_r = 0.243826:0.393302:1.62741;
		specparam tpd_S0_Y_posedge_f = 0.291199:0.482068:1.93154;
		specparam tpd_S0_Y_negedge_r = 0.286559:0.459683:1.85438;
		specparam tpd_S0_Y_negedge_f = 0.280141:0.461015:1.55183;
		specparam tpd_S1_Y_posedge_r = 0.129178:0.260057:1.3297;
		specparam tpd_S1_Y_posedge_f = 0.163276:0.343364:1.78785;
		specparam tpd_S1_Y_negedge_r = 0.182261:0.352639:1.74377;
		specparam tpd_S1_Y_negedge_f = 0.157966:0.305477:1.29027;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX4I 
`timescale 1ns/10ps
`celldefine
module MUX4IX1 (Y, D0, D1, D2, D3, S0, S1);
	output Y;
	input D0, D1, D2, D3, S0, S1;

	// Function
	wire D0__bar, D1__bar, D2__bar;
	wire D3__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2, int_fwire_3, S0__bar;
	wire S1__bar;

	not (D3__bar, D3);
	and (int_fwire_0, D3__bar, S0, S1);
	not (S0__bar, S0);
	not (D2__bar, D2);
	and (int_fwire_1, D2__bar, S0__bar, S1);
	not (S1__bar, S1);
	not (D1__bar, D1);
	and (int_fwire_2, D1__bar, S0, S1__bar);
	not (D0__bar, D0);
	and (int_fwire_3, D0__bar, S0__bar, S1__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.392481:0.549672:2.00446;
		specparam tpd_D0_Y_f = 0.31198:0.454161:1.77692;
		specparam tpd_D1_Y_r = 0.398374:0.555029:2.01041;
		specparam tpd_D1_Y_f = 0.318213:0.459285:1.77388;
		specparam tpd_D2_Y_r = 0.380328:0.537939:1.9975;
		specparam tpd_D2_Y_f = 0.295626:0.436671:1.74047;
		specparam tpd_D3_Y_r = 0.382757:0.538546:1.97775;
		specparam tpd_D3_Y_f = 0.305527:0.450679:1.79128;
		specparam tpd_S0_Y_posedge_r = 0.386458:0.542026:1.8226;
		specparam tpd_S0_Y_posedge_f = 0.324991:0.484714:1.8741;
		specparam tpd_S0_Y_negedge_r = 0.389232:0.544641:2.00882;
		specparam tpd_S0_Y_negedge_f = 0.299334:0.446051:1.77328;
		specparam tpd_S1_Y_posedge_r = 0.261456:0.411416:1.63238;
		specparam tpd_S1_Y_posedge_f = 0.217329:0.367015:1.70899;
		specparam tpd_S1_Y_negedge_r = 0.243819:0.39619:1.84588;
		specparam tpd_S1_Y_negedge_f = 0.18941:0.332717:1.55259;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(D3 => Y) = ( tpd_D3_Y_r , tpd_D3_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX4I 
`timescale 1ns/10ps
`celldefine
module MUX4IX2 (Y, D0, D1, D2, D3, S0, S1);
	output Y;
	input D0, D1, D2, D3, S0, S1;

	// Function
	wire D0__bar, D1__bar, D2__bar;
	wire D3__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2, int_fwire_3, S0__bar;
	wire S1__bar;

	not (D3__bar, D3);
	and (int_fwire_0, D3__bar, S0, S1);
	not (S0__bar, S0);
	not (D2__bar, D2);
	and (int_fwire_1, D2__bar, S0__bar, S1);
	not (S1__bar, S1);
	not (D1__bar, D1);
	and (int_fwire_2, D1__bar, S0, S1__bar);
	not (D0__bar, D0);
	and (int_fwire_3, D0__bar, S0__bar, S1__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.416828:0.5804:2.03259;
		specparam tpd_D0_Y_f = 0.330669:0.474292:1.73774;
		specparam tpd_D1_Y_r = 0.423198:0.586056:2.03938;
		specparam tpd_D1_Y_f = 0.337109:0.479595:1.73493;
		specparam tpd_D2_Y_r = 0.404316:0.567469:2.02195;
		specparam tpd_D2_Y_f = 0.313055:0.455198:1.69959;
		specparam tpd_D3_Y_r = 0.408135:0.569878:2.0038;
		specparam tpd_D3_Y_f = 0.3241:0.470746:1.75287;
		specparam tpd_S0_Y_posedge_r = 0.411164:0.573134:1.84954;
		specparam tpd_S0_Y_posedge_f = 0.343719:0.504813:1.83169;
		specparam tpd_S0_Y_negedge_r = 0.413451:0.574955:2.04081;
		specparam tpd_S0_Y_negedge_f = 0.31884:0.467347:1.73627;
		specparam tpd_S1_Y_posedge_r = 0.285357:0.441002:1.65726;
		specparam tpd_S1_Y_posedge_f = 0.236249:0.387083:1.66328;
		specparam tpd_S1_Y_negedge_r = 0.2672:0.42529:1.87603;
		specparam tpd_S1_Y_negedge_f = 0.207945:0.352383:1.51342;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(D3 => Y) = ( tpd_D3_Y_r , tpd_D3_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX4I 
`timescale 1ns/10ps
`celldefine
module MUX4IX4 (Y, D0, D1, D2, D3, S0, S1);
	output Y;
	input D0, D1, D2, D3, S0, S1;

	// Function
	wire D0__bar, D1__bar, D2__bar;
	wire D3__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2, int_fwire_3, S0__bar;
	wire S1__bar;

	not (D3__bar, D3);
	and (int_fwire_0, D3__bar, S0, S1);
	not (S0__bar, S0);
	not (D2__bar, D2);
	and (int_fwire_1, D2__bar, S0__bar, S1);
	not (S1__bar, S1);
	not (D1__bar, D1);
	and (int_fwire_2, D1__bar, S0, S1__bar);
	not (D0__bar, D0);
	and (int_fwire_3, D0__bar, S0__bar, S1__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.470602:0.64257:2.12079;
		specparam tpd_D0_Y_f = 0.370356:0.519032:1.74419;
		specparam tpd_D1_Y_r = 0.473188:0.645033:2.12596;
		specparam tpd_D1_Y_f = 0.378374:0.525949:1.74211;
		specparam tpd_D2_Y_r = 0.453296:0.625922:2.10902;
		specparam tpd_D2_Y_f = 0.353177:0.500528:1.70638;
		specparam tpd_D3_Y_r = 0.456685:0.626952:2.08569;
		specparam tpd_D3_Y_f = 0.364642:0.516636:1.76393;
		specparam tpd_S0_Y_posedge_r = 0.46152:0.632729:1.93442;
		specparam tpd_S0_Y_posedge_f = 0.384511:0.550799:1.83589;
		specparam tpd_S0_Y_negedge_r = 0.467362:0.638367:2.13788;
		specparam tpd_S0_Y_negedge_f = 0.359872:0.513186:1.74787;
		specparam tpd_S1_Y_posedge_r = 0.334202:0.498764:1.73761;
		specparam tpd_S1_Y_posedge_f = 0.277368:0.433421:1.66714;
		specparam tpd_S1_Y_negedge_r = 0.31699:0.48413:1.96816;
		specparam tpd_S1_Y_negedge_f = 0.248308:0.397664:1.52288;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(D3 => Y) = ( tpd_D3_Y_r , tpd_D3_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX4I 
`timescale 1ns/10ps
`celldefine
module MUX4IXL (Y, D0, D1, D2, D3, S0, S1);
	output Y;
	input D0, D1, D2, D3, S0, S1;

	// Function
	wire D0__bar, D1__bar, D2__bar;
	wire D3__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_2, int_fwire_3, S0__bar;
	wire S1__bar;

	not (D3__bar, D3);
	and (int_fwire_0, D3__bar, S0, S1);
	not (S0__bar, S0);
	not (D2__bar, D2);
	and (int_fwire_1, D2__bar, S0__bar, S1);
	not (S1__bar, S1);
	not (D1__bar, D1);
	and (int_fwire_2, D1__bar, S0, S1__bar);
	not (D0__bar, D0);
	and (int_fwire_3, D0__bar, S0__bar, S1__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.401762:0.562077:2.08819;
		specparam tpd_D0_Y_f = 0.349409:0.471346:1.48279;
		specparam tpd_D1_Y_r = 0.415949:0.576012:2.10973;
		specparam tpd_D1_Y_f = 0.358559:0.480885:1.49221;
		specparam tpd_D2_Y_r = 0.392232:0.552777:2.08293;
		specparam tpd_D2_Y_f = 0.331658:0.452945:1.4479;
		specparam tpd_D3_Y_r = 0.393865:0.552938:2.06137;
		specparam tpd_D3_Y_f = 0.347707:0.472557:1.50833;
		specparam tpd_S0_Y_posedge_r = 0.394102:0.543689:1.80381;
		specparam tpd_S0_Y_posedge_f = 0.382556:0.531658:1.73589;
		specparam tpd_S0_Y_negedge_r = 0.409862:0.567071:2.12829;
		specparam tpd_S0_Y_negedge_f = 0.327583:0.451225:1.45764;
		specparam tpd_S1_Y_posedge_r = 0.246668:0.391936:1.56168;
		specparam tpd_S1_Y_posedge_f = 0.245624:0.387533:1.5211;
		specparam tpd_S1_Y_negedge_r = 0.234494:0.392349:1.91161;
		specparam tpd_S1_Y_negedge_f = 0.196085:0.317162:1.19888;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(D3 => Y) = ( tpd_D3_Y_r , tpd_D3_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX4 
`timescale 1ns/10ps
`celldefine
module MUX4X1 (Y, D0, D1, D2, D3, S0, S1);
	output Y;
	input D0, D1, D2, D3, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, S0__bar, S1__bar;

	and (int_fwire_0, D3, S0, S1);
	not (S0__bar, S0);
	and (int_fwire_1, D2, S0__bar, S1);
	not (S1__bar, S1);
	and (int_fwire_2, D1, S0, S1__bar);
	and (int_fwire_3, D0, S0__bar, S1__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.246955:0.407896:1.6891;
		specparam tpd_D0_Y_f = 0.317917:0.539465:2.11309;
		specparam tpd_D1_Y_r = 0.252454:0.413936:1.68751;
		specparam tpd_D1_Y_f = 0.32364:0.5447:2.11947;
		specparam tpd_D2_Y_r = 0.231458:0.388944:1.64842;
		specparam tpd_D2_Y_f = 0.307195:0.526398:2.09781;
		specparam tpd_D3_Y_r = 0.240709:0.404031:1.7021;
		specparam tpd_D3_Y_f = 0.309364:0.527398:2.07967;
		specparam tpd_S0_Y_posedge_r = 0.233539:0.400697:1.69829;
		specparam tpd_S0_Y_posedge_f = 0.314366:0.534513:2.14431;
		specparam tpd_S0_Y_negedge_r = 0.259909:0.438474:1.76888;
		specparam tpd_S0_Y_negedge_f = 0.311737:0.531933:1.90743;
		specparam tpd_S1_Y_posedge_r = 0.124915:0.285287:1.4659;
		specparam tpd_S1_Y_posedge_f = 0.173234:0.384695:1.96366;
		specparam tpd_S1_Y_negedge_r = 0.152185:0.320912:1.60554;
		specparam tpd_S1_Y_negedge_f = 0.189606:0.39965:1.70013;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(D3 => Y) = ( tpd_D3_Y_r , tpd_D3_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX4 
`timescale 1ns/10ps
`celldefine
module MUX4X2 (Y, D0, D1, D2, D3, S0, S1);
	output Y;
	input D0, D1, D2, D3, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, S0__bar, S1__bar;

	and (int_fwire_0, D3, S0, S1);
	not (S0__bar, S0);
	and (int_fwire_1, D2, S0__bar, S1);
	not (S1__bar, S1);
	and (int_fwire_2, D1, S0, S1__bar);
	and (int_fwire_3, D0, S0__bar, S1__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.276669:0.447684:1.75065;
		specparam tpd_D0_Y_f = 0.364849:0.59211:2.11933;
		specparam tpd_D1_Y_r = 0.283655:0.45525:1.74984;
		specparam tpd_D1_Y_f = 0.371985:0.598847:2.12871;
		specparam tpd_D2_Y_r = 0.259755:0.427467:1.71014;
		specparam tpd_D2_Y_f = 0.354041:0.579265:2.10604;
		specparam tpd_D3_Y_r = 0.270331:0.443989:1.76384;
		specparam tpd_D3_Y_f = 0.355946:0.580051:2.08856;
		specparam tpd_S0_Y_posedge_r = 0.265073:0.442769:1.78064;
		specparam tpd_S0_Y_posedge_f = 0.361762:0.587601:2.14962;
		specparam tpd_S0_Y_negedge_r = 0.289067:0.477703:1.81628;
		specparam tpd_S0_Y_negedge_f = 0.358885:0.584374:1.91306;
		specparam tpd_S1_Y_posedge_r = 0.155138:0.328478:1.57812;
		specparam tpd_S1_Y_posedge_f = 0.224962:0.444568:1.98529;
		specparam tpd_S1_Y_negedge_r = 0.180384:0.362462:1.66661;
		specparam tpd_S1_Y_negedge_f = 0.238761:0.455239:1.71146;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(D3 => Y) = ( tpd_D3_Y_r , tpd_D3_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX4 
`timescale 1ns/10ps
`celldefine
module MUX4X4 (Y, D0, D1, D2, D3, S0, S1);
	output Y;
	input D0, D1, D2, D3, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, S0__bar, S1__bar;

	and (int_fwire_0, D3, S0, S1);
	not (S0__bar, S0);
	and (int_fwire_1, D2, S0__bar, S1);
	not (S1__bar, S1);
	and (int_fwire_2, D1, S0, S1__bar);
	and (int_fwire_3, D0, S0__bar, S1__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.358126:0.537487:1.86396;
		specparam tpd_D0_Y_f = 0.478186:0.698878:2.09635;
		specparam tpd_D1_Y_r = 0.368655:0.548374:1.86588;
		specparam tpd_D1_Y_f = 0.486158:0.706344:2.10616;
		specparam tpd_D2_Y_r = 0.338795:0.515175:1.81859;
		specparam tpd_D2_Y_f = 0.466729:0.686162:2.08334;
		specparam tpd_D3_Y_r = 0.352317:0.534608:1.88053;
		specparam tpd_D3_Y_f = 0.468867:0.687213:2.06525;
		specparam tpd_S0_Y_posedge_r = 0.350731:0.536852:1.9273;
		specparam tpd_S0_Y_posedge_f = 0.475823:0.695161:2.12131;
		specparam tpd_S0_Y_negedge_r = 0.369804:0.566854:1.90528;
		specparam tpd_S0_Y_negedge_f = 0.472232:0.690341:1.88834;
		specparam tpd_S1_Y_posedge_r = 0.23934:0.419573:1.76003;
		specparam tpd_S1_Y_posedge_f = 0.355475:0.567733:1.96769;
		specparam tpd_S1_Y_negedge_r = 0.263527:0.454855:1.76986;
		specparam tpd_S1_Y_negedge_f = 0.360949:0.571264:1.71936;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(D3 => Y) = ( tpd_D3_Y_r , tpd_D3_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: MUX4 
`timescale 1ns/10ps
`celldefine
module MUX4XL (Y, D0, D1, D2, D3, S0, S1);
	output Y;
	input D0, D1, D2, D3, S0, S1;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, S0__bar, S1__bar;

	and (int_fwire_0, D3, S0, S1);
	not (S0__bar, S0);
	and (int_fwire_1, D2, S0__bar, S1);
	not (S1__bar, S1);
	and (int_fwire_2, D1, S0, S1__bar);
	and (int_fwire_3, D0, S0__bar, S1__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_D0_Y_r = 0.287414:0.443513:1.7382;
		specparam tpd_D0_Y_f = 0.305542:0.496769:1.75665;
		specparam tpd_D1_Y_r = 0.295999:0.45396:1.74992;
		specparam tpd_D1_Y_f = 0.318773:0.510549:1.77968;
		specparam tpd_D2_Y_r = 0.270293:0.423945:1.69957;
		specparam tpd_D2_Y_f = 0.297841:0.487012:1.74312;
		specparam tpd_D3_Y_r = 0.285709:0.444936:1.76348;
		specparam tpd_D3_Y_f = 0.299429:0.487313:1.72009;
		specparam tpd_S0_Y_posedge_r = 0.264967:0.424377:1.72243;
		specparam tpd_S0_Y_posedge_f = 0.313532:0.501844:1.80356;
		specparam tpd_S0_Y_negedge_r = 0.320475:0.504063:1.97309;
		specparam tpd_S0_Y_negedge_f = 0.296614:0.479316:1.44228;
		specparam tpd_S1_Y_posedge_r = 0.133953:0.287526:1.45116;
		specparam tpd_S1_Y_posedge_f = 0.153522:0.325453:1.55836;
		specparam tpd_S1_Y_negedge_r = 0.183485:0.359442:1.75972;
		specparam tpd_S1_Y_negedge_f = 0.160534:0.326002:1.17011;

		(D0 => Y) = ( tpd_D0_Y_r , tpd_D0_Y_f );
		(D1 => Y) = ( tpd_D1_Y_r , tpd_D1_Y_f );
		(D2 => Y) = ( tpd_D2_Y_r , tpd_D2_Y_f );
		(D3 => Y) = ( tpd_D3_Y_r , tpd_D3_Y_f );
		(posedge S0 => (Y:S0)) = ( tpd_S0_Y_posedge_r , tpd_S0_Y_posedge_f );
		(negedge S0 => (Y:S0)) = ( tpd_S0_Y_negedge_r , tpd_S0_Y_negedge_f );
		(posedge S1 => (Y:S1)) = ( tpd_S1_Y_posedge_r , tpd_S1_Y_posedge_f );
		(negedge S1 => (Y:S1)) = ( tpd_S1_Y_negedge_r , tpd_S1_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: NAND21 
`timescale 1ns/10ps
`celldefine
module NAND21X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0369237:0.179306:1.79608;
		specparam tpd_A_Y_f = 0.0331829:0.145117:1.48718;
		specparam tpd_B_Y_r = 0.0968204:0.214622:1.30022;
		specparam tpd_B_Y_f = 0.0902441:0.207341:1.23147;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND21 
`timescale 1ns/10ps
`celldefine
module NAND21X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0341597:0.177411:1.79957;
		specparam tpd_A_Y_f = 0.0299401:0.13679:1.42932;
		specparam tpd_B_Y_r = 0.11768:0.246862:1.36922;
		specparam tpd_B_Y_f = 0.108933:0.237989:1.27297;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND21 
`timescale 1ns/10ps
`celldefine
module NAND21X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0353118:0.178097:1.79307;
		specparam tpd_A_Y_f = 0.0303968:0.135965:1.40793;
		specparam tpd_B_Y_r = 0.13985:0.276562:1.45998;
		specparam tpd_B_Y_f = 0.125309:0.259111:1.29892;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND21 
`timescale 1ns/10ps
`celldefine
module NAND21XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0476585:0.193992:1.83423;
		specparam tpd_A_Y_f = 0.0420413:0.151581:1.46283;
		specparam tpd_B_Y_r = 0.108023:0.217418:1.24338;
		specparam tpd_B_Y_f = 0.112147:0.239095:1.35507;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND2 
`timescale 1ns/10ps
`celldefine
module NAND2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0363799:0.178516:1.79229;
		specparam tpd_A_Y_f = 0.0335035:0.147957:1.51834;
		specparam tpd_B_Y_r = 0.0460732:0.190334:1.80471;
		specparam tpd_B_Y_f = 0.0407814:0.143227:1.40461;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND2 
`timescale 1ns/10ps
`celldefine
module NAND2X12 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.156114:0.304945:1.68579;
		specparam tpd_A_Y_f = 0.14857:0.246576:0.854549;
		specparam tpd_B_Y_r = 0.168111:0.321783:1.73451;
		specparam tpd_B_Y_f = 0.155506:0.247364:0.833162;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND2 
`timescale 1ns/10ps
`celldefine
module NAND2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0339929:0.177086:1.80008;
		specparam tpd_A_Y_f = 0.02994:0.13722:1.43596;
		specparam tpd_B_Y_r = 0.0439513:0.188892:1.80717;
		specparam tpd_B_Y_f = 0.0370959:0.134791:1.33795;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND2 
`timescale 1ns/10ps
`celldefine
module NAND2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0352986:0.178117:1.79568;
		specparam tpd_A_Y_f = 0.0309545:0.138554:1.43548;
		specparam tpd_B_Y_r = 0.045791:0.190846:1.80753;
		specparam tpd_B_Y_f = 0.0384427:0.134785:1.32317;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND2 
`timescale 1ns/10ps
`celldefine
module NAND2X6 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.161143:0.310316:1.67415;
		specparam tpd_A_Y_f = 0.148436:0.248465:0.864075;
		specparam tpd_B_Y_r = 0.174169:0.32756:1.73638;
		specparam tpd_B_Y_f = 0.155525:0.245018:0.821267;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND2 
`timescale 1ns/10ps
`celldefine
module NAND2X8 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.133369:0.278246:1.65255;
		specparam tpd_A_Y_f = 0.147473:0.240939:0.797882;
		specparam tpd_B_Y_r = 0.145712:0.295483:1.70588;
		specparam tpd_B_Y_f = 0.154695:0.243187:0.780008;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND2 
`timescale 1ns/10ps
`celldefine
module NAND2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.04834:0.194519:1.83429;
		specparam tpd_A_Y_f = 0.0434157:0.155552:1.50011;
		specparam tpd_B_Y_r = 0.0590563:0.20611:1.84698;
		specparam tpd_B_Y_f = 0.0516174:0.150471:1.37647;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND31 
`timescale 1ns/10ps
`celldefine
module NAND31X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0442936:0.182587:1.73856;
		specparam tpd_A_Y_f = 0.048354:0.175387:1.69927;
		specparam tpd_B_Y_r = 0.0558006:0.196205:1.75407;
		specparam tpd_B_Y_f = 0.0625339:0.177861:1.61939;
		specparam tpd_C_Y_r = 0.113758:0.228246:1.25683;
		specparam tpd_C_Y_f = 0.12039:0.249411:1.48621;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND31 
`timescale 1ns/10ps
`celldefine
module NAND31X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0441336:0.18697:1.78891;
		specparam tpd_A_Y_f = 0.0405804:0.153615:1.51373;
		specparam tpd_B_Y_r = 0.0572978:0.201546:1.8026;
		specparam tpd_B_Y_f = 0.0540131:0.157993:1.44721;
		specparam tpd_C_Y_r = 0.140514:0.26689:1.36885;
		specparam tpd_C_Y_f = 0.131643:0.261764:1.38649;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND31 
`timescale 1ns/10ps
`celldefine
module NAND31X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0491097:0.193914:1.81162;
		specparam tpd_A_Y_f = 0.0348728:0.12634:1.22252;
		specparam tpd_B_Y_r = 0.0671081:0.212483:1.83169;
		specparam tpd_B_Y_f = 0.0475944:0.130849:1.1505;
		specparam tpd_C_Y_r = 0.166245:0.295811:1.41741;
		specparam tpd_C_Y_f = 0.134472:0.252727:1.16438;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND31 
`timescale 1ns/10ps
`celldefine
module NAND31XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0490223:0.188414:1.74681;
		specparam tpd_A_Y_f = 0.0542615:0.180903:1.7015;
		specparam tpd_B_Y_r = 0.0607068:0.201809:1.76125;
		specparam tpd_B_Y_f = 0.0687094:0.183566:1.61823;
		specparam tpd_C_Y_r = 0.124567:0.232862:1.1758;
		specparam tpd_C_Y_f = 0.149382:0.294473:1.64951;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND32 
`timescale 1ns/10ps
`celldefine
module NAND32X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.036746:0.178476:1.78454;
		specparam tpd_A_Y_f = 0.0326991:0.142463:1.45799;
		specparam tpd_B_Y_r = 0.105186:0.225021:1.27313;
		specparam tpd_B_Y_f = 0.131929:0.261223:1.35277;
		specparam tpd_C_Y_r = 0.117721:0.243499:1.32608;
		specparam tpd_C_Y_f = 0.154512:0.268048:1.31157;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND32 
`timescale 1ns/10ps
`celldefine
module NAND32X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0338892:0.177196:1.80139;
		specparam tpd_A_Y_f = 0.0295395:0.135884:1.42224;
		specparam tpd_B_Y_r = 0.127648:0.259528:1.36469;
		specparam tpd_B_Y_f = 0.17026:0.310002:1.43982;
		specparam tpd_C_Y_r = 0.138339:0.272357:1.40295;
		specparam tpd_C_Y_f = 0.192662:0.31563:1.38118;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND32 
`timescale 1ns/10ps
`celldefine
module NAND32X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0353493:0.17844:1.79704;
		specparam tpd_A_Y_f = 0.0303078:0.135551:1.40392;
		specparam tpd_B_Y_r = 0.1494:0.286287:1.42199;
		specparam tpd_B_Y_f = 0.205631:0.348281:1.49896;
		specparam tpd_C_Y_r = 0.158757:0.295815:1.45055;
		specparam tpd_C_Y_f = 0.227867:0.354069:1.42724;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND32 
`timescale 1ns/10ps
`celldefine
module NAND32XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.048958:0.200646:1.91116;
		specparam tpd_A_Y_f = 0.0418138:0.154106:1.50123;
		specparam tpd_B_Y_r = 0.10948:0.228113:1.33836;
		specparam tpd_B_Y_f = 0.141852:0.273757:1.45787;
		specparam tpd_C_Y_r = 0.120329:0.246251:1.394;
		specparam tpd_C_Y_f = 0.16652:0.282623:1.41508;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND3 
`timescale 1ns/10ps
`celldefine
module NAND3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0442228:0.181897:1.73171;
		specparam tpd_A_Y_f = 0.0484702:0.175409:1.69909;
		specparam tpd_B_Y_r = 0.0557624:0.195614:1.74566;
		specparam tpd_B_Y_f = 0.0628692:0.178157:1.62044;
		specparam tpd_C_Y_r = 0.0632644:0.204766:1.75662;
		specparam tpd_C_Y_f = 0.0704792:0.176512:1.51137;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND3 
`timescale 1ns/10ps
`celldefine
module NAND3X12 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.235878:0.399485:1.881;
		specparam tpd_A_Y_f = 0.218681:0.354519:1.45412;
		specparam tpd_B_Y_r = 0.252327:0.417492:1.93215;
		specparam tpd_B_Y_f = 0.232033:0.356671:1.41979;
		specparam tpd_C_Y_r = 0.265714:0.431316:1.9725;
		specparam tpd_C_Y_f = 0.23894:0.352543:1.35655;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND3 
`timescale 1ns/10ps
`celldefine
module NAND3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0442016:0.186334:1.77932;
		specparam tpd_A_Y_f = 0.0407098:0.153311:1.50836;
		specparam tpd_B_Y_r = 0.0573544:0.200936:1.79299;
		specparam tpd_B_Y_f = 0.0543523:0.157789:1.44221;
		specparam tpd_C_Y_r = 0.0666801:0.211805:1.80617;
		specparam tpd_C_Y_f = 0.0617624:0.156219:1.33366;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND3 
`timescale 1ns/10ps
`celldefine
module NAND3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0491927:0.192372:1.78866;
		specparam tpd_A_Y_f = 0.0348162:0.124716:1.20106;
		specparam tpd_B_Y_r = 0.067401:0.211225:1.80907;
		specparam tpd_B_Y_f = 0.0477234:0.129375:1.12959;
		specparam tpd_C_Y_r = 0.0811905:0.226882:1.82783;
		specparam tpd_C_Y_f = 0.0550142:0.127564:1.01007;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND3 
`timescale 1ns/10ps
`celldefine
module NAND3X8 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.20341:0.364338:1.82378;
		specparam tpd_A_Y_f = 0.19854:0.331982:1.41364;
		specparam tpd_B_Y_r = 0.21965:0.382682:1.87923;
		specparam tpd_B_Y_f = 0.212124:0.334949:1.38337;
		specparam tpd_C_Y_r = 0.232729:0.396291:1.91953;
		specparam tpd_C_Y_f = 0.219324:0.332255:1.32947;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND3 
`timescale 1ns/10ps
`celldefine
module NAND3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0498037:0.188719:1.74065;
		specparam tpd_A_Y_f = 0.0550147:0.18141:1.69992;
		specparam tpd_B_Y_r = 0.0619856:0.202664:1.75532;
		specparam tpd_B_Y_f = 0.0706336:0.185609:1.62147;
		specparam tpd_C_Y_r = 0.0693494:0.211321:1.76679;
		specparam tpd_C_Y_f = 0.0776555:0.182856:1.50851;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND41 
`timescale 1ns/10ps
`celldefine
module NAND41X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0526785:0.190254:1.71938;
		specparam tpd_A_Y_f = 0.0554245:0.177923:1.65304;
		specparam tpd_B_Y_r = 0.0668037:0.205292:1.73591;
		specparam tpd_B_Y_f = 0.0743687:0.186134:1.59285;
		specparam tpd_C_Y_r = 0.0776813:0.217781:1.75217;
		specparam tpd_C_Y_f = 0.0876384:0.190211:1.4928;
		specparam tpd_D_Y_r = 0.134346:0.246776:1.23866;
		specparam tpd_D_Y_f = 0.144625:0.271096:1.48284;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND41 
`timescale 1ns/10ps
`celldefine
module NAND41X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0545984:0.196107:1.77622;
		specparam tpd_A_Y_f = 0.0544324:0.176034:1.64199;
		specparam tpd_B_Y_r = 0.0691854:0.210931:1.78765;
		specparam tpd_B_Y_f = 0.0737485:0.186491:1.60048;
		specparam tpd_C_Y_r = 0.0806369:0.223085:1.79523;
		specparam tpd_C_Y_f = 0.0875237:0.191542:1.50743;
		specparam tpd_D_Y_r = 0.162358:0.286643:1.3419;
		specparam tpd_D_Y_f = 0.168368:0.307159:1.57077;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND41 
`timescale 1ns/10ps
`celldefine
module NAND41X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.181755:0.334915:1.7339;
		specparam tpd_A_Y_f = 0.221849:0.325921:0.954192;
		specparam tpd_B_Y_r = 0.200535:0.356329:1.79885;
		specparam tpd_B_Y_f = 0.242469:0.336544:0.939228;
		specparam tpd_C_Y_r = 0.215341:0.372111:1.84596;
		specparam tpd_C_Y_f = 0.256372:0.342773:0.903161;
		specparam tpd_D_Y_r = 0.273192:0.403011:1.62882;
		specparam tpd_D_Y_f = 0.309813:0.417581:1.0799;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND41 
`timescale 1ns/10ps
`celldefine
module NAND41XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0617464:0.201706:1.74877;
		specparam tpd_A_Y_f = 0.0557174:0.165549:1.46765;
		specparam tpd_B_Y_r = 0.0829248:0.22528:1.81661;
		specparam tpd_B_Y_f = 0.0757375:0.174973:1.40515;
		specparam tpd_C_Y_r = 0.098635:0.242391:1.84288;
		specparam tpd_C_Y_f = 0.089596:0.180494:1.30671;
		specparam tpd_D_Y_r = 0.162978:0.272765:1.23991;
		specparam tpd_D_Y_f = 0.165904:0.294903:1.45019;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND42 
`timescale 1ns/10ps
`celldefine
module NAND42X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.044302:0.182819:1.74281;
		specparam tpd_A_Y_f = 0.0483787:0.17538:1.6991;
		specparam tpd_B_Y_r = 0.0552086:0.195781:1.75635;
		specparam tpd_B_Y_f = 0.0614998:0.176764:1.61805;
		specparam tpd_C_Y_r = 0.122448:0.239695:1.23943;
		specparam tpd_C_Y_f = 0.1658:0.307093:1.64372;
		specparam tpd_D_Y_r = 0.135399:0.258687:1.29473;
		specparam tpd_D_Y_f = 0.190156:0.315838:1.59744;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND42 
`timescale 1ns/10ps
`celldefine
module NAND42X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0440899:0.186926:1.78959;
		specparam tpd_A_Y_f = 0.0403612:0.152803:1.50593;
		specparam tpd_B_Y_r = 0.0572446:0.201574:1.80337;
		specparam tpd_B_Y_f = 0.0536004:0.156842:1.43814;
		specparam tpd_C_Y_r = 0.150635:0.278847:1.35778;
		specparam tpd_C_Y_f = 0.192095:0.329739:1.54904;
		specparam tpd_D_Y_r = 0.161079:0.291717:1.39615;
		specparam tpd_D_Y_f = 0.214378:0.335291:1.49177;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND42 
`timescale 1ns/10ps
`celldefine
module NAND42X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0491705:0.193799:1.80894;
		specparam tpd_A_Y_f = 0.0347529:0.125598:1.21394;
		specparam tpd_B_Y_r = 0.0672482:0.212464:1.82914;
		specparam tpd_B_Y_f = 0.0474157:0.130066:1.14181;
		specparam tpd_C_Y_r = 0.176557:0.306948:1.4007;
		specparam tpd_C_Y_f = 0.200862:0.324158:1.33424;
		specparam tpd_D_Y_r = 0.187698:0.319876:1.44251;
		specparam tpd_D_Y_f = 0.224749:0.330862:1.2622;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND42 
`timescale 1ns/10ps
`celldefine
module NAND42XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.049644:0.189986:1.76022;
		specparam tpd_A_Y_f = 0.0544148:0.18091:1.70049;
		specparam tpd_B_Y_r = 0.0608462:0.202808:1.77366;
		specparam tpd_B_Y_f = 0.0681278:0.182975:1.61764;
		specparam tpd_C_Y_r = 0.120969:0.231656:1.16824;
		specparam tpd_C_Y_f = 0.182949:0.32791:1.72265;
		specparam tpd_D_Y_r = 0.132826:0.250373:1.23003;
		specparam tpd_D_Y_f = 0.208:0.336414:1.66357;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND43 
`timescale 1ns/10ps
`celldefine
module NAND43X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.036631:0.178429:1.78509;
		specparam tpd_A_Y_f = 0.0326441:0.142689:1.4623;
		specparam tpd_B_Y_r = 0.106747:0.2282:1.22005;
		specparam tpd_B_Y_f = 0.188022:0.333978:1.56339;
		specparam tpd_C_Y_r = 0.120312:0.247004:1.27241;
		specparam tpd_C_Y_f = 0.243439:0.3714:1.54659;
		specparam tpd_D_Y_r = 0.126252:0.259171:1.33439;
		specparam tpd_D_Y_f = 0.266304:0.390447:1.46321;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND43 
`timescale 1ns/10ps
`celldefine
module NAND43X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0339402:0.177233:1.80116;
		specparam tpd_A_Y_f = 0.029616:0.136009:1.42321;
		specparam tpd_B_Y_r = 0.124895:0.257085:1.30576;
		specparam tpd_B_Y_f = 0.245547:0.398137:1.6613;
		specparam tpd_C_Y_r = 0.138039:0.272505:1.34966;
		specparam tpd_C_Y_f = 0.300974:0.438339:1.63189;
		specparam tpd_D_Y_r = 0.144452:0.282291:1.40012;
		specparam tpd_D_Y_f = 0.322128:0.454499:1.53724;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND43 
`timescale 1ns/10ps
`celldefine
module NAND43X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0353484:0.17815:1.79348;
		specparam tpd_A_Y_f = 0.0303439:0.135518:1.40359;
		specparam tpd_B_Y_r = 0.14405:0.28278:1.38933;
		specparam tpd_B_Y_f = 0.294277:0.448151:1.72677;
		specparam tpd_C_Y_r = 0.156914:0.296122:1.42728;
		specparam tpd_C_Y_f = 0.350381:0.490551:1.68894;
		specparam tpd_D_Y_r = 0.163991:0.305507:1.4733;
		specparam tpd_D_Y_f = 0.371644:0.506857:1.58722;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND43 
`timescale 1ns/10ps
`celldefine
module NAND43XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar;

	not (A__bar, A);
	or (Y, A__bar, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0467029:0.198725:1.91375;
		specparam tpd_A_Y_f = 0.0401133:0.151593:1.49249;
		specparam tpd_B_Y_r = 0.111592:0.236274:1.34595;
		specparam tpd_B_Y_f = 0.170322:0.310821:1.54733;
		specparam tpd_C_Y_r = 0.125072:0.256535:1.40383;
		specparam tpd_C_Y_f = 0.221708:0.343875:1.53455;
		specparam tpd_D_Y_r = 0.132246:0.271037:1.47076;
		specparam tpd_D_Y_f = 0.244106:0.363077:1.45252;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND4 
`timescale 1ns/10ps
`celldefine
module NAND4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0527094:0.189613:1.711;
		specparam tpd_A_Y_f = 0.0556509:0.178089:1.6522;
		specparam tpd_B_Y_r = 0.066806:0.204809:1.72819;
		specparam tpd_B_Y_f = 0.074925:0.186614:1.59332;
		specparam tpd_C_Y_r = 0.0777808:0.217277:1.74369;
		specparam tpd_C_Y_f = 0.0884205:0.191075:1.49484;
		specparam tpd_D_Y_r = 0.0860171:0.227417:1.75755;
		specparam tpd_D_Y_f = 0.096743:0.196724:1.42119;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND4 
`timescale 1ns/10ps
`celldefine
module NAND4X12 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.194446:0.34958:1.77091;
		specparam tpd_A_Y_f = 0.205016:0.306314:0.925155;
		specparam tpd_B_Y_r = 0.211579:0.368914:1.82186;
		specparam tpd_B_Y_f = 0.224074:0.318091:0.924995;
		specparam tpd_C_Y_r = 0.225603:0.38395:1.86453;
		specparam tpd_C_Y_f = 0.237621:0.323595:0.891872;
		specparam tpd_D_Y_r = 0.233125:0.391907:1.88987;
		specparam tpd_D_Y_f = 0.245498:0.327848:0.854699;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND4 
`timescale 1ns/10ps
`celldefine
module NAND4X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0544292:0.197584:1.79905;
		specparam tpd_A_Y_f = 0.054425:0.178301:1.6763;
		specparam tpd_B_Y_r = 0.0690925:0.2123:1.8096;
		specparam tpd_B_Y_f = 0.0741155:0.189175:1.63655;
		specparam tpd_C_Y_r = 0.0803465:0.224142:1.81621;
		specparam tpd_C_Y_f = 0.0881147:0.194479:1.54456;
		specparam tpd_D_Y_r = 0.0862532:0.22987:1.79428;
		specparam tpd_D_Y_f = 0.0963975:0.199881:1.47193;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND4 
`timescale 1ns/10ps
`celldefine
module NAND4X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.179817:0.334168:1.74504;
		specparam tpd_A_Y_f = 0.215882:0.318374:0.922564;
		specparam tpd_B_Y_r = 0.196475:0.353365:1.80399;
		specparam tpd_B_Y_f = 0.23435:0.327376:0.907913;
		specparam tpd_C_Y_r = 0.210614:0.368796:1.85264;
		specparam tpd_C_Y_f = 0.247332:0.33172:0.868785;
		specparam tpd_D_Y_r = 0.222665:0.381728:1.89439;
		specparam tpd_D_Y_f = 0.254913:0.335147:0.821933;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND4 
`timescale 1ns/10ps
`celldefine
module NAND4X8 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.169397:0.322197:1.73278;
		specparam tpd_A_Y_f = 0.205684:0.308422:0.929851;
		specparam tpd_B_Y_r = 0.186392:0.341699:1.78605;
		specparam tpd_B_Y_f = 0.224883:0.320571:0.930315;
		specparam tpd_C_Y_r = 0.20093:0.357423:1.83289;
		specparam tpd_C_Y_f = 0.238446:0.326103:0.899043;
		specparam tpd_D_Y_r = 0.210501:0.367852:1.86516;
		specparam tpd_D_Y_f = 0.246219:0.330293:0.861272;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND4 
`timescale 1ns/10ps
`celldefine
module NAND4XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0642859:0.204929:1.76488;
		specparam tpd_A_Y_f = 0.0576382:0.168503:1.48206;
		specparam tpd_B_Y_r = 0.085895:0.228527:1.82495;
		specparam tpd_B_Y_f = 0.0788475:0.17899:1.42029;
		specparam tpd_C_Y_r = 0.101666:0.245331:1.84449;
		specparam tpd_C_Y_f = 0.0937075:0.186178:1.32638;
		specparam tpd_D_Y_r = 0.107253:0.250532:1.81457;
		specparam tpd_D_Y_f = 0.100646:0.189111:1.24649;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND5 
`timescale 1ns/10ps
`celldefine
module NAND5X1 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.144991:0.287568:1.62546;
		specparam tpd_A_Y_f = 0.167798:0.303225:1.44421;
		specparam tpd_B_Y_r = 0.15986:0.30868:1.69868;
		specparam tpd_B_Y_f = 0.175411:0.302581:1.4048;
		specparam tpd_C_Y_r = 0.169263:0.315279:1.6448;
		specparam tpd_C_Y_f = 0.217748:0.3586:1.54254;
		specparam tpd_D_Y_r = 0.183042:0.33372:1.71105;
		specparam tpd_D_Y_f = 0.230803:0.362213:1.51464;
		specparam tpd_E_Y_r = 0.195663:0.348979:1.76036;
		specparam tpd_E_Y_f = 0.238271:0.361131:1.46187;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND5 
`timescale 1ns/10ps
`celldefine
module NAND5X2 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.155735:0.303562:1.64677;
		specparam tpd_A_Y_f = 0.194754:0.341906:1.51426;
		specparam tpd_B_Y_r = 0.170947:0.32488:1.71886;
		specparam tpd_B_Y_f = 0.202375:0.341233:1.47469;
		specparam tpd_C_Y_r = 0.181401:0.333494:1.67522;
		specparam tpd_C_Y_f = 0.245743:0.397842:1.60767;
		specparam tpd_D_Y_r = 0.194824:0.351009:1.73343;
		specparam tpd_D_Y_f = 0.258592:0.401688:1.58236;
		specparam tpd_E_Y_r = 0.206364:0.364622:1.77811;
		specparam tpd_E_Y_f = 0.266086:0.400544:1.53278;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND5 
`timescale 1ns/10ps
`celldefine
module NAND5X4 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.191823:0.349454:1.72786;
		specparam tpd_A_Y_f = 0.254883:0.393804:1.28596;
		specparam tpd_B_Y_r = 0.207505:0.370905:1.79767;
		specparam tpd_B_Y_f = 0.262514:0.393621:1.24837;
		specparam tpd_C_Y_r = 0.212481:0.371846:1.7335;
		specparam tpd_C_Y_f = 0.305849:0.450992:1.38922;
		specparam tpd_D_Y_r = 0.229189:0.392773:1.80216;
		specparam tpd_D_Y_f = 0.318839:0.454276:1.35758;
		specparam tpd_E_Y_r = 0.241658:0.408036:1.85354;
		specparam tpd_E_Y_f = 0.32636:0.453141:1.30512;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND5 
`timescale 1ns/10ps
`celldefine
module NAND5XL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.18718:0.342596:1.79259;
		specparam tpd_A_Y_f = 0.201486:0.325328:1.22083;
		specparam tpd_B_Y_r = 0.204974:0.3626:1.86325;
		specparam tpd_B_Y_f = 0.209044:0.320604:1.17022;
		specparam tpd_C_Y_r = 0.187224:0.338102:1.73806;
		specparam tpd_C_Y_f = 0.23497:0.357687:1.27143;
		specparam tpd_D_Y_r = 0.205795:0.360278:1.80734;
		specparam tpd_D_Y_f = 0.249542:0.363099:1.24619;
		specparam tpd_E_Y_r = 0.216294:0.372388:1.84889;
		specparam tpd_E_Y_f = 0.256272:0.361395:1.19816;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND6 
`timescale 1ns/10ps
`celldefine
module NAND6X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.156302:0.301408:1.62881;
		specparam tpd_A_Y_f = 0.198588:0.340811:1.53578;
		specparam tpd_B_Y_r = 0.172555:0.322377:1.70119;
		specparam tpd_B_Y_f = 0.212616:0.345201:1.50453;
		specparam tpd_C_Y_r = 0.183954:0.337138:1.75257;
		specparam tpd_C_Y_f = 0.220161:0.343626:1.4506;
		specparam tpd_D_Y_r = 0.168079:0.31368:1.64011;
		specparam tpd_D_Y_f = 0.217994:0.358376:1.53688;
		specparam tpd_E_Y_r = 0.183784:0.334103:1.71217;
		specparam tpd_E_Y_f = 0.230379:0.361188:1.50515;
		specparam tpd_F_Y_r = 0.195933:0.349379:1.76318;
		specparam tpd_F_Y_f = 0.237986:0.359972:1.45044;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND6 
`timescale 1ns/10ps
`celldefine
module NAND6X2 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.168069:0.318424:1.65321;
		specparam tpd_A_Y_f = 0.22735:0.381375:1.61217;
		specparam tpd_B_Y_r = 0.184636:0.339758:1.72416;
		specparam tpd_B_Y_f = 0.241393:0.385702:1.58122;
		specparam tpd_C_Y_r = 0.196395:0.354358:1.77507;
		specparam tpd_C_Y_f = 0.248959:0.384176:1.52812;
		specparam tpd_D_Y_r = 0.180569:0.332417:1.67345;
		specparam tpd_D_Y_f = 0.246752:0.398371:1.60574;
		specparam tpd_E_Y_r = 0.193246:0.349279:1.73023;
		specparam tpd_E_Y_f = 0.259052:0.401649:1.57966;
		specparam tpd_F_Y_r = 0.206785:0.365212:1.78305;
		specparam tpd_F_Y_f = 0.266469:0.400207:1.52555;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND6 
`timescale 1ns/10ps
`celldefine
module NAND6X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.204561:0.363698:1.72103;
		specparam tpd_A_Y_f = 0.287586:0.433069:1.3798;
		specparam tpd_B_Y_r = 0.22163:0.38489:1.79124;
		specparam tpd_B_Y_f = 0.301618:0.437712:1.35059;
		specparam tpd_C_Y_r = 0.234127:0.400037:1.84021;
		specparam tpd_C_Y_f = 0.309194:0.436337:1.29956;
		specparam tpd_D_Y_r = 0.214901:0.374724:1.73618;
		specparam tpd_D_Y_f = 0.307029:0.450688:1.37405;
		specparam tpd_E_Y_r = 0.227813:0.39131:1.79162;
		specparam tpd_E_Y_f = 0.31933:0.45386:1.34771;
		specparam tpd_F_Y_r = 0.241861:0.407568:1.84313;
		specparam tpd_F_Y_f = 0.326723:0.452399:1.29426;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND6 
`timescale 1ns/10ps
`celldefine
module NAND6XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.180159:0.33027:1.71749;
		specparam tpd_A_Y_f = 0.213541:0.338852:1.28521;
		specparam tpd_B_Y_r = 0.198326:0.351885:1.78685;
		specparam tpd_B_Y_f = 0.227513:0.343532:1.25859;
		specparam tpd_C_Y_r = 0.211486:0.366189:1.83537;
		specparam tpd_C_Y_f = 0.234581:0.341065:1.20512;
		specparam tpd_D_Y_r = 0.19155:0.342258:1.73505;
		specparam tpd_D_Y_f = 0.233945:0.356969:1.27836;
		specparam tpd_E_Y_r = 0.206201:0.359648:1.78858;
		specparam tpd_E_Y_f = 0.246506:0.360681:1.25765;
		specparam tpd_F_Y_r = 0.219591:0.37498:1.83959;
		specparam tpd_F_Y_f = 0.253203:0.357875:1.20348;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND8 
`timescale 1ns/10ps
`celldefine
module NAND8X1 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire G__bar, H__bar;

	not (H__bar, H);
	not (G__bar, G);
	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar, G__bar, H__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.156191:0.297235:1.63921;
		specparam tpd_A_Y_f = 0.178633:0.298668:1.29107;
		specparam tpd_B_Y_r = 0.168965:0.315562:1.69991;
		specparam tpd_B_Y_f = 0.186177:0.299215:1.26093;
		specparam tpd_C_Y_r = 0.173846:0.316452:1.66625;
		specparam tpd_C_Y_f = 0.204228:0.324016:1.30137;
		specparam tpd_D_Y_r = 0.185953:0.333982:1.72352;
		specparam tpd_D_Y_f = 0.211025:0.323281:1.27076;
		specparam tpd_E_Y_r = 0.166824:0.307844:1.65362;
		specparam tpd_E_Y_f = 0.185463:0.302027:1.29226;
		specparam tpd_F_Y_r = 0.181039:0.327709:1.72212;
		specparam tpd_F_Y_f = 0.193654:0.302891:1.25815;
		specparam tpd_G_Y_r = 0.183925:0.32528:1.67219;
		specparam tpd_G_Y_f = 0.211983:0.328767:1.31117;
		specparam tpd_H_Y_r = 0.196066:0.342949:1.73242;
		specparam tpd_H_Y_f = 0.218721:0.32753:1.27562;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND8 
`timescale 1ns/10ps
`celldefine
module NAND8X2 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire G__bar, H__bar;

	not (H__bar, H);
	not (G__bar, G);
	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar, G__bar, H__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.173071:0.31835:1.67093;
		specparam tpd_A_Y_f = 0.208958:0.333754:1.2887;
		specparam tpd_B_Y_r = 0.186115:0.336953:1.73075;
		specparam tpd_B_Y_f = 0.216549:0.334484:1.25925;
		specparam tpd_C_Y_r = 0.190583:0.33736:1.69644;
		specparam tpd_C_Y_f = 0.234428:0.359083:1.29828;
		specparam tpd_D_Y_r = 0.202881:0.354896:1.7525;
		specparam tpd_D_Y_f = 0.241174:0.358331:1.268;
		specparam tpd_E_Y_r = 0.191166:0.33602:1.69545;
		specparam tpd_E_Y_f = 0.224329:0.347391:1.30043;
		specparam tpd_F_Y_r = 0.205918:0.356162:1.75772;
		specparam tpd_F_Y_f = 0.232647:0.348997:1.27316;
		specparam tpd_G_Y_r = 0.205085:0.349285:1.6993;
		specparam tpd_G_Y_f = 0.248974:0.372124:1.31872;
		specparam tpd_H_Y_r = 0.217413:0.36706:1.75856;
		specparam tpd_H_Y_f = 0.255755:0.370645:1.28368;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND8 
`timescale 1ns/10ps
`celldefine
module NAND8X4 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire G__bar, H__bar;

	not (H__bar, H);
	not (G__bar, G);
	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar, G__bar, H__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.197132:0.343336:1.66784;
		specparam tpd_A_Y_f = 0.249931:0.375743:1.27955;
		specparam tpd_B_Y_r = 0.210452:0.362029:1.72679;
		specparam tpd_B_Y_f = 0.25749:0.376365:1.25167;
		specparam tpd_C_Y_r = 0.214936:0.362588:1.69247;
		specparam tpd_C_Y_f = 0.275261:0.401084:1.28922;
		specparam tpd_D_Y_r = 0.227381:0.380025:1.7471;
		specparam tpd_D_Y_f = 0.28204:0.400531:1.25961;
		specparam tpd_E_Y_r = 0.210555:0.357363:1.72558;
		specparam tpd_E_Y_f = 0.254336:0.3762:1.27458;
		specparam tpd_F_Y_r = 0.225447:0.37731:1.78848;
		specparam tpd_F_Y_f = 0.262591:0.37765:1.24686;
		specparam tpd_G_Y_r = 0.226095:0.372088:1.73167;
		specparam tpd_G_Y_f = 0.280236:0.403186:1.29776;
		specparam tpd_H_Y_r = 0.238481:0.389759:1.78971;
		specparam tpd_H_Y_f = 0.286986:0.401692:1.26341;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NAND8 
`timescale 1ns/10ps
`celldefine
module NAND8XL (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire G__bar, H__bar;

	not (H__bar, H);
	not (G__bar, G);
	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar, G__bar, H__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.194462:0.346593:1.76712;
		specparam tpd_A_Y_f = 0.220416:0.349437:1.411;
		specparam tpd_B_Y_r = 0.206839:0.361267:1.80944;
		specparam tpd_B_Y_f = 0.229243:0.349018:1.38614;
		specparam tpd_C_Y_r = 0.211258:0.365243:1.80097;
		specparam tpd_C_Y_f = 0.24491:0.371962:1.40697;
		specparam tpd_D_Y_r = 0.228444:0.384013:1.86262;
		specparam tpd_D_Y_f = 0.252842:0.369305:1.36751;
		specparam tpd_E_Y_r = 0.206631:0.358496:1.77778;
		specparam tpd_E_Y_f = 0.228595:0.354905:1.42153;
		specparam tpd_F_Y_r = 0.219041:0.373143:1.8216;
		specparam tpd_F_Y_f = 0.237407:0.354063:1.39279;
		specparam tpd_G_Y_r = 0.228192:0.381885:1.81898;
		specparam tpd_G_Y_f = 0.255577:0.380225:1.4226;
		specparam tpd_H_Y_r = 0.238688:0.393487:1.84932;
		specparam tpd_H_Y_f = 0.264579:0.379946:1.40308;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR21 
`timescale 1ns/10ps
`celldefine
module NOR21X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0452212:0.178722:1.71547;
		specparam tpd_A_Y_f = 0.0336338:0.122738:1.14665;
		specparam tpd_B_Y_r = 0.113169:0.225335:1.28274;
		specparam tpd_B_Y_f = 0.0937775:0.185509:0.868629;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR21 
`timescale 1ns/10ps
`celldefine
module NOR21X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0400234:0.173007:1.70882;
		specparam tpd_A_Y_f = 0.0299807:0.117879:1.13407;
		specparam tpd_B_Y_r = 0.127452:0.250092:1.33912;
		specparam tpd_B_Y_f = 0.114088:0.218741:0.937435;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR21 
`timescale 1ns/10ps
`celldefine
module NOR21X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0564243:0.197735:1.78614;
		specparam tpd_A_Y_f = 0.0241394:0.074861:0.67546;
		specparam tpd_B_Y_r = 0.170853:0.301828:1.44623;
		specparam tpd_B_Y_f = 0.119343:0.214317:0.732486;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR21 
`timescale 1ns/10ps
`celldefine
module NOR21XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0526015:0.189201:1.74806;
		specparam tpd_A_Y_f = 0.033507:0.112826:1.01772;
		specparam tpd_B_Y_r = 0.131558:0.241378:1.24393;
		specparam tpd_B_Y_f = 0.117889:0.222229:0.951887;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR2 
`timescale 1ns/10ps
`celldefine
module NOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0450189:0.177684:1.70946;
		specparam tpd_A_Y_f = 0.0350241:0.129544:1.21214;
		specparam tpd_B_Y_r = 0.0671472:0.180965:1.53768;
		specparam tpd_B_Y_f = 0.0484813:0.15098:1.2322;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR2 
`timescale 1ns/10ps
`celldefine
module NOR2X12 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.19653:0.343344:1.72912;
		specparam tpd_A_Y_f = 0.149333:0.258451:0.906189;
		specparam tpd_B_Y_r = 0.219523:0.348897:1.6515;
		specparam tpd_B_Y_f = 0.167923:0.287249:1.01208;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR2 
`timescale 1ns/10ps
`celldefine
module NOR2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0397965:0.172648:1.70869;
		specparam tpd_A_Y_f = 0.0300511:0.119329:1.15086;
		specparam tpd_B_Y_r = 0.0623603:0.176009:1.53134;
		specparam tpd_B_Y_f = 0.0418246:0.141109:1.17643;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR2 
`timescale 1ns/10ps
`celldefine
module NOR2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0603716:0.201629:1.79211;
		specparam tpd_A_Y_f = 0.0239972:0.072441:0.643516;
		specparam tpd_B_Y_r = 0.0854657:0.203929:1.62065;
		specparam tpd_B_Y_f = 0.0278012:0.0860657:0.664585;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR2 
`timescale 1ns/10ps
`celldefine
module NOR2X6 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.21638:0.363412:1.77029;
		specparam tpd_A_Y_f = 0.152058:0.260502:0.890837;
		specparam tpd_B_Y_r = 0.238949:0.36856:1.69881;
		specparam tpd_B_Y_f = 0.165716:0.278847:0.956893;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR2 
`timescale 1ns/10ps
`celldefine
module NOR2X8 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.169695:0.311158:1.66776;
		specparam tpd_A_Y_f = 0.148397:0.252553:0.830113;
		specparam tpd_B_Y_r = 0.193611:0.319076:1.60928;
		specparam tpd_B_Y_f = 0.163255:0.276471:0.912182;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR2 
`timescale 1ns/10ps
`celldefine
module NOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0510306:0.187651:1.75147;
		specparam tpd_A_Y_f = 0.0330074:0.11333:1.03433;
		specparam tpd_B_Y_r = 0.0754936:0.193394:1.58302;
		specparam tpd_B_Y_f = 0.0438202:0.133432:1.05483;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR31 
`timescale 1ns/10ps
`celldefine
module NOR31X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0678054:0.200161:1.69877;
		specparam tpd_A_Y_f = 0.0367728:0.105676:0.811912;
		specparam tpd_B_Y_r = 0.122379:0.236197:1.6165;
		specparam tpd_B_Y_f = 0.0479864:0.124294:0.812382;
		specparam tpd_C_Y_r = 0.191711:0.303253:1.34667;
		specparam tpd_C_Y_f = 0.0993477:0.177889:0.657292;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR31 
`timescale 1ns/10ps
`celldefine
module NOR31X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0655288:0.198978:1.7075;
		specparam tpd_A_Y_f = 0.0341738:0.0985087:0.763025;
		specparam tpd_B_Y_r = 0.121916:0.237931:1.62745;
		specparam tpd_B_Y_f = 0.0490334:0.126613:0.830221;
		specparam tpd_C_Y_r = 0.20859:0.328737:1.39675;
		specparam tpd_C_Y_f = 0.125633:0.216796:0.758807;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR31 
`timescale 1ns/10ps
`celldefine
module NOR31X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.250983:0.399905:1.87978;
		specparam tpd_A_Y_f = 0.165279:0.276954:0.85964;
		specparam tpd_B_Y_r = 0.306818:0.43807:1.85716;
		specparam tpd_B_Y_f = 0.179826:0.296774:0.921056;
		specparam tpd_C_Y_r = 0.376462:0.505574:1.69363;
		specparam tpd_C_Y_f = 0.241544:0.357063:1.09152;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR31 
`timescale 1ns/10ps
`celldefine
module NOR31XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0811547:0.215325:1.74239;
		specparam tpd_A_Y_f = 0.0373949:0.0991483:0.710501;
		specparam tpd_B_Y_r = 0.143016:0.25935:1.66471;
		specparam tpd_B_Y_f = 0.0479749:0.117824:0.715926;
		specparam tpd_C_Y_r = 0.214733:0.318662:1.27013;
		specparam tpd_C_Y_f = 0.125617:0.218885:0.80318;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR32 
`timescale 1ns/10ps
`celldefine
module NOR32X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0453249:0.178535:1.7126;
		specparam tpd_A_Y_f = 0.0337776:0.12315:1.14887;
		specparam tpd_B_Y_r = 0.119331:0.224826:1.21888;
		specparam tpd_B_Y_f = 0.11328:0.217599:1.02283;
		specparam tpd_C_Y_r = 0.126659:0.225219:1.19802;
		specparam tpd_C_Y_f = 0.123128:0.232396:1.05992;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR32 
`timescale 1ns/10ps
`celldefine
module NOR32X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.042635:0.175694:1.7098;
		specparam tpd_A_Y_f = 0.0311192:0.119077:1.13029;
		specparam tpd_B_Y_r = 0.131834:0.246091:1.26609;
		specparam tpd_B_Y_f = 0.128216:0.238829:1.02851;
		specparam tpd_C_Y_r = 0.139199:0.244064:1.23648;
		specparam tpd_C_Y_f = 0.139853:0.253845:1.07062;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR32 
`timescale 1ns/10ps
`celldefine
module NOR32X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0595595:0.201143:1.79241;
		specparam tpd_A_Y_f = 0.0238991:0.0723083:0.644193;
		specparam tpd_B_Y_r = 0.170893:0.292831:1.36454;
		specparam tpd_B_Y_f = 0.131881:0.230973:0.820526;
		specparam tpd_C_Y_r = 0.178277:0.289168:1.3295;
		specparam tpd_C_Y_f = 0.143117:0.244782:0.860593;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR32 
`timescale 1ns/10ps
`celldefine
module NOR32XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0521745:0.189078:1.751;
		specparam tpd_A_Y_f = 0.0327735:0.110108:0.994741;
		specparam tpd_B_Y_r = 0.15175:0.263982:1.26359;
		specparam tpd_B_Y_f = 0.137078:0.247027:1.00358;
		specparam tpd_C_Y_r = 0.15932:0.259532:1.21571;
		specparam tpd_C_Y_f = 0.154076:0.267545:1.06977;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR3 
`timescale 1ns/10ps
`celldefine
module NOR3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0613759:0.192069:1.67952;
		specparam tpd_A_Y_f = 0.0380098:0.113605:0.906773;
		specparam tpd_B_Y_r = 0.112193:0.225601:1.591;
		specparam tpd_B_Y_f = 0.0513497:0.134085:0.911;
		specparam tpd_C_Y_r = 0.13162:0.238846:1.43979;
		specparam tpd_C_Y_f = 0.0553384:0.149129:0.965659;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR3 
`timescale 1ns/10ps
`celldefine
module NOR3X12 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.359916:0.510431:2.04416;
		specparam tpd_A_Y_f = 0.182737:0.30272:0.951737;
		specparam tpd_B_Y_r = 0.41584:0.551538:2.006;
		specparam tpd_B_Y_f = 0.195971:0.317799:0.998134;
		specparam tpd_C_Y_r = 0.437756:0.568232:1.90598;
		specparam tpd_C_Y_f = 0.203442:0.327204:1.04808;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR3 
`timescale 1ns/10ps
`celldefine
module NOR3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0552302:0.187584:1.69216;
		specparam tpd_A_Y_f = 0.0333434:0.103495:0.845729;
		specparam tpd_B_Y_r = 0.110665:0.22647:1.60405;
		specparam tpd_B_Y_f = 0.0466642:0.128268:0.878182;
		specparam tpd_C_Y_r = 0.132165:0.243684:1.46675;
		specparam tpd_C_Y_f = 0.0469369:0.139009:0.907435;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR3 
`timescale 1ns/10ps
`celldefine
module NOR3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.250004:0.399404:1.8901;
		specparam tpd_A_Y_f = 0.16397:0.275773:0.863997;
		specparam tpd_B_Y_r = 0.305989:0.437645:1.86713;
		specparam tpd_B_Y_f = 0.178504:0.295568:0.925502;
		specparam tpd_C_Y_r = 0.32757:0.454854:1.77606;
		specparam tpd_C_Y_f = 0.186148:0.307988:0.989582;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR3 
`timescale 1ns/10ps
`celldefine
module NOR3X8 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.377715:0.50468:1.82203;
		specparam tpd_A_Y_f = 0.199603:0.324561:1.04107;
		specparam tpd_B_Y_r = 0.355863:0.487434:1.91778;
		specparam tpd_B_Y_f = 0.192361:0.314502:0.988523;
		specparam tpd_C_Y_r = 0.299226:0.44685:1.95028;
		specparam tpd_C_Y_f = 0.178712:0.298324:0.939204;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR3 
`timescale 1ns/10ps
`celldefine
module NOR3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0797301:0.213362:1.73456;
		specparam tpd_A_Y_f = 0.0369858:0.0991208:0.721491;
		specparam tpd_B_Y_r = 0.135287:0.250566:1.64802;
		specparam tpd_B_Y_f = 0.0474725:0.117484:0.729664;
		specparam tpd_C_Y_r = 0.157279:0.268157:1.50216;
		specparam tpd_C_Y_f = 0.0512064:0.134142:0.806419;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR41 
`timescale 1ns/10ps
`celldefine
module NOR41X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.066574:0.196202:1.65099;
		specparam tpd_A_Y_f = 0.0482185:0.119239:0.808886;
		specparam tpd_B_Y_r = 0.154516:0.266055:1.61402;
		specparam tpd_B_Y_f = 0.073817:0.154613:0.863813;
		specparam tpd_C_Y_r = 0.206701:0.317772:1.52966;
		specparam tpd_C_Y_f = 0.0859865:0.174242:0.924644;
		specparam tpd_D_Y_r = 0.295485:0.41539:1.46772;
		specparam tpd_D_Y_f = 0.168626:0.264412:0.865263;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR41 
`timescale 1ns/10ps
`celldefine
module NOR41X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0637195:0.193499:1.65073;
		specparam tpd_A_Y_f = 0.0358257:0.0967811:0.667006;
		specparam tpd_B_Y_r = 0.148375:0.258801:1.61065;
		specparam tpd_B_Y_f = 0.0485913:0.120066:0.683082;
		specparam tpd_C_Y_r = 0.20062:0.310827:1.52453;
		specparam tpd_C_Y_f = 0.0499872:0.130781:0.711921;
		specparam tpd_D_Y_r = 0.292746:0.412299:1.45419;
		specparam tpd_D_Y_f = 0.127623:0.21438:0.688774;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR41 
`timescale 1ns/10ps
`celldefine
module NOR41X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.222275:0.375397:1.86932;
		specparam tpd_A_Y_f = 0.177837:0.287531:0.856014;
		specparam tpd_B_Y_r = 0.316644:0.446868:1.86466;
		specparam tpd_B_Y_f = 0.211702:0.328028:0.973955;
		specparam tpd_C_Y_r = 0.368935:0.498759:1.81081;
		specparam tpd_C_Y_f = 0.235004:0.353008:1.06719;
		specparam tpd_D_Y_r = 0.457875:0.596639:1.83543;
		specparam tpd_D_Y_f = 0.329064:0.453142:1.21545;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR41 
`timescale 1ns/10ps
`celldefine
module NOR41XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0945481:0.225068:1.7029;
		specparam tpd_A_Y_f = 0.0388689:0.0926071:0.539688;
		specparam tpd_B_Y_r = 0.186153:0.295566:1.67157;
		specparam tpd_B_Y_f = 0.0489544:0.111032:0.54597;
		specparam tpd_C_Y_r = 0.247081:0.357743:1.59343;
		specparam tpd_C_Y_f = 0.0496348:0.120387:0.574109;
		specparam tpd_D_Y_r = 0.319702:0.420793:1.3244;
		specparam tpd_D_Y_f = 0.128784:0.217028:0.733344;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR42 
`timescale 1ns/10ps
`celldefine
module NOR42X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0701947:0.203145:1.70861;
		specparam tpd_A_Y_f = 0.0360842:0.102425:0.77753;
		specparam tpd_B_Y_r = 0.126009:0.240396:1.62562;
		specparam tpd_B_Y_f = 0.0465618:0.120395:0.776714;
		specparam tpd_C_Y_r = 0.197662:0.300433:1.26744;
		specparam tpd_C_Y_f = 0.112546:0.199263:0.75351;
		specparam tpd_D_Y_r = 0.20453:0.299723:1.23822;
		specparam tpd_D_Y_f = 0.124383:0.216711:0.802976;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR42 
`timescale 1ns/10ps
`celldefine
module NOR42X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0556466:0.18794:1.69194;
		specparam tpd_A_Y_f = 0.0334612:0.10366:0.844913;
		specparam tpd_B_Y_r = 0.110829:0.226932:1.60329;
		specparam tpd_B_Y_f = 0.0470781:0.128646:0.87919;
		specparam tpd_C_Y_r = 0.199056:0.310811:1.30714;
		specparam tpd_C_Y_f = 0.139873:0.239051:0.874884;
		specparam tpd_D_Y_r = 0.20555:0.306695:1.26796;
		specparam tpd_D_Y_f = 0.151705:0.253923:0.922855;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR42 
`timescale 1ns/10ps
`celldefine
module NOR42X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.253137:0.401064:1.88079;
		specparam tpd_A_Y_f = 0.165586:0.275974:0.833955;
		specparam tpd_B_Y_r = 0.309813:0.440149:1.85845;
		specparam tpd_B_Y_f = 0.179959:0.29529:0.893236;
		specparam tpd_C_Y_r = 0.381265:0.500633:1.61584;
		specparam tpd_C_Y_f = 0.25365:0.374262:1.15836;
		specparam tpd_D_Y_r = 0.388766:0.501148:1.59085;
		specparam tpd_D_Y_f = 0.266232:0.392059:1.21214;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR42 
`timescale 1ns/10ps
`celldefine
module NOR42XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar;

	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0823573:0.216344:1.7469;
		specparam tpd_A_Y_f = 0.0372378:0.0984363:0.705954;
		specparam tpd_B_Y_r = 0.139277:0.255154:1.66259;
		specparam tpd_B_Y_f = 0.0470316:0.115555:0.707256;
		specparam tpd_C_Y_r = 0.240568:0.350246:1.32953;
		specparam tpd_C_Y_f = 0.149511:0.247942:0.868671;
		specparam tpd_D_Y_r = 0.248136:0.346001:1.28351;
		specparam tpd_D_Y_f = 0.166351:0.267496:0.931888;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR43 
`timescale 1ns/10ps
`celldefine
module NOR43X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0456908:0.179215:1.7142;
		specparam tpd_A_Y_f = 0.0337963:0.121649:1.12796;
		specparam tpd_B_Y_r = 0.14672:0.25889:1.29366;
		specparam tpd_B_Y_f = 0.120336:0.22594:0.983448;
		specparam tpd_C_Y_r = 0.160676:0.263558:1.27385;
		specparam tpd_C_Y_f = 0.133883:0.244082:1.03603;
		specparam tpd_D_Y_r = 0.167984:0.263162:1.22922;
		specparam tpd_D_Y_f = 0.143993:0.257508:1.07899;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR43 
`timescale 1ns/10ps
`celldefine
module NOR43X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0399632:0.174136:1.72159;
		specparam tpd_A_Y_f = 0.0297146:0.116373:1.12006;
		specparam tpd_B_Y_r = 0.156524:0.276619:1.34481;
		specparam tpd_B_Y_f = 0.136299:0.24903:1.03025;
		specparam tpd_C_Y_r = 0.170113:0.279501:1.31686;
		specparam tpd_C_Y_f = 0.149782:0.265721:1.08035;
		specparam tpd_D_Y_r = 0.177063:0.276634:1.2621;
		specparam tpd_D_Y_f = 0.160109:0.278387:1.12338;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR43 
`timescale 1ns/10ps
`celldefine
module NOR43X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.060196:0.201677:1.79261;
		specparam tpd_A_Y_f = 0.0240363:0.0725274:0.644104;
		specparam tpd_B_Y_r = 0.210313:0.335711:1.45947;
		specparam tpd_B_Y_f = 0.142022:0.241715:0.827057;
		specparam tpd_C_Y_r = 0.22463:0.338872:1.43;
		specparam tpd_C_Y_f = 0.154928:0.257137:0.872597;
		specparam tpd_D_Y_r = 0.232241:0.337599:1.38044;
		specparam tpd_D_Y_f = 0.164916:0.267815:0.905228;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR43 
`timescale 1ns/10ps
`celldefine
module NOR43XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar;

	not (A__bar, A);
	and (Y, A__bar, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0538216:0.190336:1.74866;
		specparam tpd_A_Y_f = 0.0334478:0.111246:0.99715;
		specparam tpd_B_Y_r = 0.163963:0.278056:1.31289;
		specparam tpd_B_Y_f = 0.133238:0.240017:0.96918;
		specparam tpd_C_Y_r = 0.17874:0.283728:1.29228;
		specparam tpd_C_Y_f = 0.148835:0.259334:1.02495;
		specparam tpd_D_Y_r = 0.186115:0.282936:1.24857;
		specparam tpd_D_Y_f = 0.158705:0.27118:1.06274;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR4 
`timescale 1ns/10ps
`celldefine
module NOR4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0683157:0.197138:1.64045;
		specparam tpd_A_Y_f = 0.0489304:0.119925:0.806047;
		specparam tpd_B_Y_r = 0.154269:0.264726:1.60008;
		specparam tpd_B_Y_f = 0.0741228:0.154623:0.859973;
		specparam tpd_C_Y_r = 0.206976:0.316992:1.51477;
		specparam tpd_C_Y_f = 0.0865853:0.174718:0.921832;
		specparam tpd_D_Y_r = 0.22882:0.336665:1.4096;
		specparam tpd_D_Y_f = 0.0958717:0.200916:1.09859;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR4 
`timescale 1ns/10ps
`celldefine
module NOR4X12 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.309492:0.463498:2.00315;
		specparam tpd_A_Y_f = 0.190826:0.303262:0.901796;
		specparam tpd_B_Y_r = 0.403042:0.537768:1.99063;
		specparam tpd_B_Y_f = 0.224354:0.339506:1.00698;
		specparam tpd_C_Y_r = 0.455847:0.590015:1.92958;
		specparam tpd_C_Y_f = 0.249595:0.364986:1.09708;
		specparam tpd_D_Y_r = 0.477662:0.609566:1.82449;
		specparam tpd_D_Y_f = 0.275154:0.400954:1.27088;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR4 
`timescale 1ns/10ps
`celldefine
module NOR4X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0680747:0.197911:1.65024;
		specparam tpd_A_Y_f = 0.0371272:0.098979:0.669072;
		specparam tpd_B_Y_r = 0.154017:0.263778:1.60987;
		specparam tpd_B_Y_f = 0.0501368:0.122189:0.685631;
		specparam tpd_C_Y_r = 0.20646:0.31578:1.52354;
		specparam tpd_C_Y_f = 0.0520281:0.133174:0.716275;
		specparam tpd_D_Y_r = 0.231092:0.339744:1.44115;
		specparam tpd_D_Y_f = 0.051252:0.140587:0.767801;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR4 
`timescale 1ns/10ps
`celldefine
module NOR4X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.202575:0.35187:1.77509;
		specparam tpd_A_Y_f = 0.177931:0.297198:0.944242;
		specparam tpd_B_Y_r = 0.298446:0.430159:1.79768;
		specparam tpd_B_Y_f = 0.211056:0.336769:1.05067;
		specparam tpd_C_Y_r = 0.353822:0.485436:1.7626;
		specparam tpd_C_Y_f = 0.231522:0.359183:1.13438;
		specparam tpd_D_Y_r = 0.379673:0.511329:1.71606;
		specparam tpd_D_Y_f = 0.247264:0.377762:1.22358;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR4 
`timescale 1ns/10ps
`celldefine
module NOR4X8 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.261637:0.414149:1.93342;
		specparam tpd_A_Y_f = 0.188834:0.302031:0.903045;
		specparam tpd_B_Y_r = 0.356283:0.487988:1.91584;
		specparam tpd_B_Y_f = 0.226981:0.344362:1.02961;
		specparam tpd_C_Y_r = 0.410346:0.541665:1.8626;
		specparam tpd_C_Y_f = 0.250437:0.367962:1.11171;
		specparam tpd_D_Y_r = 0.432501:0.562248:1.77719;
		specparam tpd_D_Y_f = 0.259282:0.386589:1.23249;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR4 
`timescale 1ns/10ps
`celldefine
module NOR4XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0940893:0.22443:1.69747;
		specparam tpd_A_Y_f = 0.0389739:0.0930858:0.546174;
		specparam tpd_B_Y_r = 0.184535:0.29385:1.6662;
		specparam tpd_B_Y_f = 0.0492475:0.111844:0.554155;
		specparam tpd_C_Y_r = 0.244416:0.354638:1.58528;
		specparam tpd_C_Y_f = 0.0500877:0.122042:0.587022;
		specparam tpd_D_Y_r = 0.266378:0.37411:1.49263;
		specparam tpd_D_Y_f = 0.0519196:0.132546:0.662525;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR5 
`timescale 1ns/10ps
`celldefine
module NOR5X1 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.182255:0.329708:1.72794;
		specparam tpd_A_Y_f = 0.147564:0.286588:1.48615;
		specparam tpd_B_Y_r = 0.205874:0.336918:1.66782;
		specparam tpd_B_Y_f = 0.162018:0.307886:1.55962;
		specparam tpd_C_Y_r = 0.238357:0.39054:1.8861;
		specparam tpd_C_Y_f = 0.158723:0.300593:1.45367;
		specparam tpd_D_Y_r = 0.29461:0.428558:1.86287;
		specparam tpd_D_Y_f = 0.172926:0.320079:1.5128;
		specparam tpd_E_Y_r = 0.317869:0.448333:1.77259;
		specparam tpd_E_Y_f = 0.180373:0.332443:1.57846;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR5 
`timescale 1ns/10ps
`celldefine
module NOR5X2 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.191079:0.342638:1.73601;
		specparam tpd_A_Y_f = 0.160385:0.305146:1.49843;
		specparam tpd_B_Y_r = 0.214708:0.349802:1.67698;
		specparam tpd_B_Y_f = 0.17499:0.326211:1.57025;
		specparam tpd_C_Y_r = 0.246876:0.402981:1.89262;
		specparam tpd_C_Y_f = 0.170921:0.318454:1.46428;
		specparam tpd_D_Y_r = 0.30307:0.441126:1.86978;
		specparam tpd_D_Y_f = 0.185308:0.33794:1.52219;
		specparam tpd_E_Y_r = 0.326322:0.46095:1.77999;
		specparam tpd_E_Y_f = 0.193239:0.350641:1.58783;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR5 
`timescale 1ns/10ps
`celldefine
module NOR5X4 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.224075:0.380382:1.76296;
		specparam tpd_A_Y_f = 0.189773:0.323436:1.21428;
		specparam tpd_B_Y_r = 0.247593:0.387364:1.7094;
		specparam tpd_B_Y_f = 0.204608:0.344706:1.28394;
		specparam tpd_C_Y_r = 0.282076:0.442384:1.91826;
		specparam tpd_C_Y_f = 0.199657:0.336322:1.17904;
		specparam tpd_D_Y_r = 0.33839:0.480616:1.89729;
		specparam tpd_D_Y_f = 0.214158:0.355824:1.2371;
		specparam tpd_E_Y_r = 0.361522:0.500524:1.80856;
		specparam tpd_E_Y_f = 0.222816:0.368944:1.30161;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR5 
`timescale 1ns/10ps
`celldefine
module NOR5XL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.218009:0.368255:1.78541;
		specparam tpd_A_Y_f = 0.16331:0.279831:1.14362;
		specparam tpd_B_Y_r = 0.243089:0.377337:1.73844;
		specparam tpd_B_Y_f = 0.173644:0.29698:1.20157;
		specparam tpd_C_Y_r = 0.298966:0.453204:1.97871;
		specparam tpd_C_Y_f = 0.190389:0.316617:1.16604;
		specparam tpd_D_Y_r = 0.360474:0.497439:1.95243;
		specparam tpd_D_Y_f = 0.204828:0.3358:1.22781;
		specparam tpd_E_Y_r = 0.385187:0.519338:1.86426;
		specparam tpd_E_Y_f = 0.211888:0.347074:1.28536;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR6 
`timescale 1ns/10ps
`celldefine
module NOR6X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.205676:0.358222:1.72182;
		specparam tpd_A_Y_f = 0.158186:0.30001:1.4905;
		specparam tpd_B_Y_r = 0.231058:0.368667:1.67638;
		specparam tpd_B_Y_f = 0.171861:0.319807:1.55266;
		specparam tpd_C_Y_r = 0.220111:0.373504:1.74629;
		specparam tpd_C_Y_f = 0.171705:0.315128:1.50317;
		specparam tpd_D_Y_r = 0.242673:0.379663:1.68641;
		specparam tpd_D_Y_f = 0.18623:0.335972:1.57472;
		specparam tpd_E_Y_r = 0.222112:0.376309:1.76162;
		specparam tpd_E_Y_f = 0.173522:0.314493:1.47011;
		specparam tpd_F_Y_r = 0.247486:0.385329:1.69072;
		specparam tpd_F_Y_f = 0.190966:0.341233:1.56548;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR6 
`timescale 1ns/10ps
`celldefine
module NOR6X2 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.218896:0.379041:1.76532;
		specparam tpd_A_Y_f = 0.171855:0.322375:1.54669;
		specparam tpd_B_Y_r = 0.244244:0.389508:1.72047;
		specparam tpd_B_Y_f = 0.185696:0.34201:1.60823;
		specparam tpd_C_Y_r = 0.232489:0.393487:1.78805;
		specparam tpd_C_Y_f = 0.185001:0.337015:1.55722;
		specparam tpd_D_Y_r = 0.25506:0.39951:1.72811;
		specparam tpd_D_Y_f = 0.199669:0.357755:1.62845;
		specparam tpd_E_Y_r = 0.234171:0.395942:1.80222;
		specparam tpd_E_Y_f = 0.1868:0.335991:1.52303;
		specparam tpd_F_Y_r = 0.258691:0.403744:1.73079;
		specparam tpd_F_Y_f = 0.204067:0.362451:1.61519;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR6 
`timescale 1ns/10ps
`celldefine
module NOR6X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.260795:0.427598:1.81179;
		specparam tpd_A_Y_f = 0.200176:0.3387:1.25425;
		specparam tpd_B_Y_r = 0.286175:0.438064:1.77058;
		specparam tpd_B_Y_f = 0.214142:0.358357:1.31333;
		specparam tpd_C_Y_r = 0.274146:0.441702:1.83368;
		specparam tpd_C_Y_f = 0.212726:0.352941:1.26359;
		specparam tpd_D_Y_r = 0.296757:0.4479:1.77583;
		specparam tpd_D_Y_f = 0.227551:0.373901:1.3338;
		specparam tpd_E_Y_r = 0.275322:0.443808:1.8514;
		specparam tpd_E_Y_f = 0.213652:0.350013:1.22077;
		specparam tpd_F_Y_r = 0.299843:0.451534:1.77854;
		specparam tpd_F_Y_f = 0.231315:0.376812:1.3152;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR6 
`timescale 1ns/10ps
`celldefine
module NOR6XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.237823:0.390668:1.81303;
		specparam tpd_A_Y_f = 0.162147:0.278891:1.12906;
		specparam tpd_B_Y_r = 0.26234:0.398409:1.75279;
		specparam tpd_B_Y_f = 0.174015:0.2972:1.19369;
		specparam tpd_C_Y_r = 0.250574:0.405696:1.85931;
		specparam tpd_C_Y_f = 0.17249:0.287329:1.10269;
		specparam tpd_D_Y_r = 0.275638:0.412696:1.78296;
		specparam tpd_D_Y_f = 0.186914:0.310463:1.19062;
		specparam tpd_E_Y_r = 0.257214:0.410552:1.83373;
		specparam tpd_E_Y_f = 0.188687:0.309872:1.16423;
		specparam tpd_F_Y_r = 0.281973:0.418548:1.7784;
		specparam tpd_F_Y_f = 0.19844:0.324142:1.21221;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR8 
`timescale 1ns/10ps
`celldefine
module NOR8X1 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire G__bar, H__bar;

	not (H__bar, H);
	not (G__bar, G);
	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar, G__bar, H__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.204221:0.346445:1.73721;
		specparam tpd_A_Y_f = 0.152832:0.2509:0.905013;
		specparam tpd_B_Y_r = 0.228741:0.35441:1.6745;
		specparam tpd_B_Y_f = 0.168286:0.273762:0.985186;
		specparam tpd_C_Y_r = 0.2029:0.344563:1.73579;
		specparam tpd_C_Y_f = 0.156941:0.2525:0.889932;
		specparam tpd_D_Y_r = 0.225745:0.350294:1.66476;
		specparam tpd_D_Y_f = 0.173615:0.278278:0.983988;
		specparam tpd_E_Y_r = 0.228871:0.370144:1.75338;
		specparam tpd_E_Y_f = 0.17116:0.268125:0.92554;
		specparam tpd_F_Y_r = 0.251425:0.376002:1.69328;
		specparam tpd_F_Y_f = 0.18509:0.288797:0.998495;
		specparam tpd_G_Y_r = 0.227484:0.368456:1.75736;
		specparam tpd_G_Y_f = 0.174519:0.268177:0.903315;
		specparam tpd_H_Y_r = 0.250256:0.374148:1.68581;
		specparam tpd_H_Y_f = 0.191348:0.294229:0.998253;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR8 
`timescale 1ns/10ps
`celldefine
module NOR8X2 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire G__bar, H__bar;

	not (H__bar, H);
	not (G__bar, G);
	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar, G__bar, H__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.21159:0.356128:1.74978;
		specparam tpd_A_Y_f = 0.166576:0.267967:0.888503;
		specparam tpd_B_Y_r = 0.2373:0.365626:1.68937;
		specparam tpd_B_Y_f = 0.182801:0.291447:0.968933;
		specparam tpd_C_Y_r = 0.206412:0.34991:1.74016;
		specparam tpd_C_Y_f = 0.166965:0.264489:0.86409;
		specparam tpd_D_Y_r = 0.229267:0.355938:1.67167;
		specparam tpd_D_Y_f = 0.183926:0.290732:0.957352;
		specparam tpd_E_Y_r = 0.243199:0.387756:1.77502;
		specparam tpd_E_Y_f = 0.187241:0.285308:0.911725;
		specparam tpd_F_Y_r = 0.26579:0.393591:1.71842;
		specparam tpd_F_Y_f = 0.201245:0.305967:0.983018;
		specparam tpd_G_Y_r = 0.240735:0.384862:1.77723;
		specparam tpd_G_Y_f = 0.189346:0.283973:0.886109;
		specparam tpd_H_Y_r = 0.263501:0.390405:1.70617;
		specparam tpd_H_Y_f = 0.206368:0.310176:0.980143;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR8 
`timescale 1ns/10ps
`celldefine
module NOR8X4 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire G__bar, H__bar;

	not (H__bar, H);
	not (G__bar, G);
	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar, G__bar, H__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.266101:0.408358:1.79394;
		specparam tpd_A_Y_f = 0.185221:0.270007:0.638235;
		specparam tpd_B_Y_r = 0.292278:0.419307:1.73967;
		specparam tpd_B_Y_f = 0.201035:0.292488:0.71254;
		specparam tpd_C_Y_r = 0.261064:0.403208:1.78903;
		specparam tpd_C_Y_f = 0.186056:0.267471:0.612511;
		specparam tpd_D_Y_r = 0.283827:0.40919:1.72162;
		specparam tpd_D_Y_f = 0.203113:0.293356:0.703626;
		specparam tpd_E_Y_r = 0.287876:0.43218:1.81374;
		specparam tpd_E_Y_f = 0.193783:0.27519:0.639543;
		specparam tpd_F_Y_r = 0.31056:0.438101:1.75561;
		specparam tpd_F_Y_f = 0.207945:0.295824:0.709661;
		specparam tpd_G_Y_r = 0.284865:0.428805:1.81482;
		specparam tpd_G_Y_f = 0.194937:0.273009:0.613063;
		specparam tpd_H_Y_r = 0.307628:0.434398:1.74493;
		specparam tpd_H_Y_f = 0.212084:0.299214:0.705583;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: NOR8 
`timescale 1ns/10ps
`celldefine
module NOR8XL (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire G__bar, H__bar;

	not (H__bar, H);
	not (G__bar, G);
	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (Y, A__bar, B__bar, C__bar, D__bar, E__bar, F__bar, G__bar, H__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.243071:0.390201:1.83761;
		specparam tpd_A_Y_f = 0.177733:0.262643:0.707431;
		specparam tpd_B_Y_r = 0.267985:0.397283:1.75625;
		specparam tpd_B_Y_f = 0.195224:0.2921:0.821007;
		specparam tpd_C_Y_r = 0.244494:0.389696:1.80942;
		specparam tpd_C_Y_f = 0.195183:0.285616:0.766151;
		specparam tpd_D_Y_r = 0.269163:0.398207:1.75795;
		specparam tpd_D_Y_f = 0.206287:0.303353:0.825504;
		specparam tpd_E_Y_r = 0.271337:0.418251:1.86113;
		specparam tpd_E_Y_f = 0.197561:0.281364:0.743777;
		specparam tpd_F_Y_r = 0.296096:0.425609:1.77487;
		specparam tpd_F_Y_f = 0.217147:0.313385:0.865721;
		specparam tpd_G_Y_r = 0.269051:0.413853:1.83276;
		specparam tpd_G_Y_f = 0.212333:0.299076:0.783527;
		specparam tpd_H_Y_r = 0.293625:0.422561:1.78086;
		specparam tpd_H_Y_f = 0.223409:0.316844:0.842784;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA21 
`timescale 1ns/10ps
`celldefine
module OA21X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, A, C);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.116433:0.261758:1.53939;
		specparam tpd_A_Y_f = 0.0933217:0.264313:1.76164;
		specparam tpd_B_Y_r = 0.110957:0.237301:1.39275;
		specparam tpd_B_Y_f = 0.170747:0.351615:1.98021;
		specparam tpd_C_Y_r = 0.136261:0.272882:1.50309;
		specparam tpd_C_Y_f = 0.192845:0.356706:1.88481;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA21 
`timescale 1ns/10ps
`celldefine
module OA21X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, A, C);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.181623:0.343752:1.68724;
		specparam tpd_A_Y_f = 0.134896:0.302776:1.4759;
		specparam tpd_B_Y_r = 0.171888:0.319367:1.53973;
		specparam tpd_B_Y_f = 0.266155:0.440888:1.76282;
		specparam tpd_C_Y_r = 0.200879:0.354793:1.63979;
		specparam tpd_C_Y_f = 0.287891:0.446358:1.63602;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA21 
`timescale 1ns/10ps
`celldefine
module OA21XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire int_fwire_0, int_fwire_1;

	and (int_fwire_0, A, C);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.132224:0.271231:1.47431;
		specparam tpd_A_Y_f = 0.118274:0.284694:1.62304;
		specparam tpd_B_Y_r = 0.133967:0.256713:1.34191;
		specparam tpd_B_Y_f = 0.250428:0.424057:1.92147;
		specparam tpd_C_Y_r = 0.160124:0.29183:1.45375;
		specparam tpd_C_Y_f = 0.279432:0.438587:1.80138;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA2222 
`timescale 1ns/10ps
`celldefine
module OA2222X1 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;
	wire int_fwire_9, int_fwire_10, int_fwire_11;
	wire int_fwire_12, int_fwire_13, int_fwire_14;
	wire int_fwire_15;

	and (int_fwire_0, B, D, F, H);
	and (int_fwire_1, B, D, F, G);
	and (int_fwire_2, B, D, E, H);
	and (int_fwire_3, B, D, E, G);
	and (int_fwire_4, B, C, F, H);
	and (int_fwire_5, B, C, F, G);
	and (int_fwire_6, B, C, E, H);
	and (int_fwire_7, B, C, E, G);
	and (int_fwire_8, A, D, F, H);
	and (int_fwire_9, A, D, F, G);
	and (int_fwire_10, A, D, E, H);
	and (int_fwire_11, A, D, E, G);
	and (int_fwire_12, A, C, F, H);
	and (int_fwire_13, A, C, F, G);
	and (int_fwire_14, A, C, E, H);
	and (int_fwire_15, A, C, E, G);
	or (Y, int_fwire_15, int_fwire_14, int_fwire_13, int_fwire_12, int_fwire_11, int_fwire_10, int_fwire_9, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.149116:0.284029:1.46762;
		specparam tpd_A_Y_f = 0.182753:0.325479:1.3738;
		specparam tpd_B_Y_r = 0.17148:0.309552:1.55145;
		specparam tpd_B_Y_f = 0.208649:0.333531:1.28418;
		specparam tpd_C_Y_r = 0.17107:0.298899:1.4782;
		specparam tpd_C_Y_f = 0.224002:0.369521:1.45205;
		specparam tpd_D_Y_r = 0.19077:0.318853:1.53246;
		specparam tpd_D_Y_f = 0.249586:0.378837:1.35708;
		specparam tpd_E_Y_r = 0.171975:0.304953:1.47593;
		specparam tpd_E_Y_f = 0.210539:0.343652:1.36807;
		specparam tpd_F_Y_r = 0.192772:0.328961:1.56205;
		specparam tpd_F_Y_f = 0.235425:0.350551:1.27699;
		specparam tpd_G_Y_r = 0.19351:0.319182:1.47978;
		specparam tpd_G_Y_f = 0.257348:0.392168:1.45217;
		specparam tpd_H_Y_r = 0.212062:0.337871:1.53255;
		specparam tpd_H_Y_f = 0.285205:0.404461:1.36325;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA2222 
`timescale 1ns/10ps
`celldefine
module OA2222X4 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;
	wire int_fwire_9, int_fwire_10, int_fwire_11;
	wire int_fwire_12, int_fwire_13, int_fwire_14;
	wire int_fwire_15;

	and (int_fwire_0, B, D, F, H);
	and (int_fwire_1, B, D, F, G);
	and (int_fwire_2, B, D, E, H);
	and (int_fwire_3, B, D, E, G);
	and (int_fwire_4, B, C, F, H);
	and (int_fwire_5, B, C, F, G);
	and (int_fwire_6, B, C, E, H);
	and (int_fwire_7, B, C, E, G);
	and (int_fwire_8, A, D, F, H);
	and (int_fwire_9, A, D, F, G);
	and (int_fwire_10, A, D, E, H);
	and (int_fwire_11, A, D, E, G);
	and (int_fwire_12, A, C, F, H);
	and (int_fwire_13, A, C, F, G);
	and (int_fwire_14, A, C, E, H);
	and (int_fwire_15, A, C, E, G);
	or (Y, int_fwire_15, int_fwire_14, int_fwire_13, int_fwire_12, int_fwire_11, int_fwire_10, int_fwire_9, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.210749:0.353493:1.62023;
		specparam tpd_A_Y_f = 0.252428:0.37395:1.23212;
		specparam tpd_B_Y_r = 0.23472:0.377914:1.69758;
		specparam tpd_B_Y_f = 0.277766:0.382705:1.10995;
		specparam tpd_C_Y_r = 0.237514:0.37178:1.62845;
		specparam tpd_C_Y_f = 0.290516:0.41449:1.2987;
		specparam tpd_D_Y_r = 0.253032:0.384927:1.65314;
		specparam tpd_D_Y_f = 0.315768:0.424999:1.18209;
		specparam tpd_E_Y_r = 0.234317:0.377171:1.63885;
		specparam tpd_E_Y_f = 0.275046:0.391922:1.24281;
		specparam tpd_F_Y_r = 0.255246:0.399059:1.71421;
		specparam tpd_F_Y_f = 0.299048:0.399222:1.11928;
		specparam tpd_G_Y_r = 0.260786:0.395496:1.64087;
		specparam tpd_G_Y_f = 0.323981:0.442915:1.32946;
		specparam tpd_H_Y_r = 0.273791:0.406269:1.66226;
		specparam tpd_H_Y_f = 0.347863:0.452419:1.2141;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA2222 
`timescale 1ns/10ps
`celldefine
module OA2222XL (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;
	wire int_fwire_9, int_fwire_10, int_fwire_11;
	wire int_fwire_12, int_fwire_13, int_fwire_14;
	wire int_fwire_15;

	and (int_fwire_0, B, D, F, H);
	and (int_fwire_1, B, D, F, G);
	and (int_fwire_2, B, D, E, H);
	and (int_fwire_3, B, D, E, G);
	and (int_fwire_4, B, C, F, H);
	and (int_fwire_5, B, C, F, G);
	and (int_fwire_6, B, C, E, H);
	and (int_fwire_7, B, C, E, G);
	and (int_fwire_8, A, D, F, H);
	and (int_fwire_9, A, D, F, G);
	and (int_fwire_10, A, D, E, H);
	and (int_fwire_11, A, D, E, G);
	and (int_fwire_12, A, C, F, H);
	and (int_fwire_13, A, C, F, G);
	and (int_fwire_14, A, C, E, H);
	and (int_fwire_15, A, C, E, G);
	or (Y, int_fwire_15, int_fwire_14, int_fwire_13, int_fwire_12, int_fwire_11, int_fwire_10, int_fwire_9, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.165546:0.301186:1.4459;
		specparam tpd_A_Y_f = 0.222921:0.363628:1.45055;
		specparam tpd_B_Y_r = 0.184909:0.320715:1.50978;
		specparam tpd_B_Y_f = 0.253314:0.377995:1.34888;
		specparam tpd_C_Y_r = 0.193106:0.321114:1.46818;
		specparam tpd_C_Y_f = 0.281822:0.425184:1.50751;
		specparam tpd_D_Y_r = 0.213361:0.338644:1.49778;
		specparam tpd_D_Y_f = 0.335721:0.471402:1.42854;
		specparam tpd_E_Y_r = 0.189632:0.322595:1.45451;
		specparam tpd_E_Y_f = 0.244328:0.379381:1.44649;
		specparam tpd_F_Y_r = 0.211859:0.346342:1.53775;
		specparam tpd_F_Y_f = 0.27467:0.393404:1.33854;
		specparam tpd_G_Y_r = 0.205511:0.326122:1.41403;
		specparam tpd_G_Y_f = 0.305972:0.441061:1.52323;
		specparam tpd_H_Y_r = 0.24298:0.369428:1.54366;
		specparam tpd_H_Y_f = 0.360104:0.486482:1.40923;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA222 
`timescale 1ns/10ps
`celldefine
module OA222X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7;

	and (int_fwire_0, B, D, F);
	and (int_fwire_1, B, D, E);
	and (int_fwire_2, B, C, F);
	and (int_fwire_3, B, C, E);
	and (int_fwire_4, A, D, F);
	and (int_fwire_5, A, D, E);
	and (int_fwire_6, A, C, F);
	and (int_fwire_7, A, C, E);
	or (Y, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.198295:0.360025:1.66806;
		specparam tpd_A_Y_f = 0.183312:0.405586:2.05364;
		specparam tpd_B_Y_r = 0.235157:0.400689:1.78044;
		specparam tpd_B_Y_f = 0.205766:0.409951:1.93879;
		specparam tpd_C_Y_r = 0.245761:0.39798:1.67367;
		specparam tpd_C_Y_f = 0.245631:0.471348:2.17225;
		specparam tpd_D_Y_r = 0.285996:0.444936:1.78157;
		specparam tpd_D_Y_f = 0.270767:0.481321:2.04846;
		specparam tpd_E_Y_r = 0.267507:0.414718:1.62977;
		specparam tpd_E_Y_f = 0.272708:0.501956:2.23064;
		specparam tpd_F_Y_r = 0.305026:0.459119:1.72179;
		specparam tpd_F_Y_f = 0.295107:0.509724:2.10239;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA222 
`timescale 1ns/10ps
`celldefine
module OA222X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7;

	and (int_fwire_0, B, D, F);
	and (int_fwire_1, B, D, E);
	and (int_fwire_2, B, C, F);
	and (int_fwire_3, B, C, E);
	and (int_fwire_4, A, D, F);
	and (int_fwire_5, A, D, E);
	and (int_fwire_6, A, C, F);
	and (int_fwire_7, A, C, E);
	or (Y, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.282413:0.458797:1.86002;
		specparam tpd_A_Y_f = 0.272907:0.479412:1.86267;
		specparam tpd_B_Y_r = 0.322356:0.502416:1.96226;
		specparam tpd_B_Y_f = 0.295005:0.484753:1.72276;
		specparam tpd_C_Y_r = 0.329096:0.497234:1.84867;
		specparam tpd_C_Y_f = 0.33574:0.546218:1.9736;
		specparam tpd_D_Y_r = 0.372638:0.546681:1.95249;
		specparam tpd_D_Y_f = 0.360719:0.557586:1.82996;
		specparam tpd_E_Y_r = 0.348987:0.510522:1.77383;
		specparam tpd_E_Y_f = 0.361363:0.574263:2.02511;
		specparam tpd_F_Y_r = 0.391248:0.559703:1.87456;
		specparam tpd_F_Y_f = 0.383714:0.583018:1.87661;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA222 
`timescale 1ns/10ps
`celldefine
module OA222XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7;

	and (int_fwire_0, B, D, F);
	and (int_fwire_1, B, D, E);
	and (int_fwire_2, B, C, F);
	and (int_fwire_3, B, C, E);
	and (int_fwire_4, A, D, F);
	and (int_fwire_5, A, D, E);
	and (int_fwire_6, A, C, F);
	and (int_fwire_7, A, C, E);
	or (Y, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.227198:0.383635:1.64031;
		specparam tpd_A_Y_f = 0.234078:0.436378:1.91738;
		specparam tpd_B_Y_r = 0.266729:0.424142:1.74762;
		specparam tpd_B_Y_f = 0.267924:0.455712:1.79552;
		specparam tpd_C_Y_r = 0.289739:0.437026:1.67378;
		specparam tpd_C_Y_f = 0.329759:0.539124:2.08856;
		specparam tpd_D_Y_r = 0.329355:0.479825:1.76611;
		specparam tpd_D_Y_f = 0.362968:0.561486:1.95203;
		specparam tpd_E_Y_r = 0.313128:0.45543:1.63116;
		specparam tpd_E_Y_f = 0.376534:0.59061:2.17079;
		specparam tpd_F_Y_r = 0.35626:0.504237:1.73186;
		specparam tpd_F_Y_f = 0.406495:0.610635:2.02311;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA22 
`timescale 1ns/10ps
`celldefine
module OA22X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	and (int_fwire_0, B, D);
	and (int_fwire_1, B, C);
	and (int_fwire_2, A, D);
	and (int_fwire_3, A, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.122047:0.268657:1.47837;
		specparam tpd_A_Y_f = 0.156244:0.357474:1.98996;
		specparam tpd_B_Y_r = 0.149324:0.302337:1.59377;
		specparam tpd_B_Y_f = 0.178901:0.361541:1.88867;
		specparam tpd_C_Y_r = 0.150691:0.288563:1.47582;
		specparam tpd_C_Y_f = 0.209902:0.416727:2.10516;
		specparam tpd_D_Y_r = 0.179577:0.324967:1.58228;
		specparam tpd_D_Y_f = 0.232032:0.421283:1.98669;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA22 
`timescale 1ns/10ps
`celldefine
module OA22X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	and (int_fwire_0, B, D);
	and (int_fwire_1, B, C);
	and (int_fwire_2, A, D);
	and (int_fwire_3, A, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.185135:0.349184:1.64822;
		specparam tpd_A_Y_f = 0.249276:0.43882:1.7848;
		specparam tpd_B_Y_r = 0.215757:0.383703:1.75451;
		specparam tpd_B_Y_f = 0.271298:0.443603:1.65517;
		specparam tpd_C_Y_r = 0.213618:0.367927:1.62167;
		specparam tpd_C_Y_f = 0.301838:0.495423:1.88638;
		specparam tpd_D_Y_r = 0.245985:0.406708:1.72215;
		specparam tpd_D_Y_f = 0.323677:0.50159:1.74371;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA22 
`timescale 1ns/10ps
`celldefine
module OA22XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	and (int_fwire_0, B, D);
	and (int_fwire_1, B, C);
	and (int_fwire_2, A, D);
	and (int_fwire_3, A, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.139611:0.281786:1.42571;
		specparam tpd_A_Y_f = 0.212239:0.405374:1.93746;
		specparam tpd_B_Y_r = 0.168208:0.315751:1.54176;
		specparam tpd_B_Y_f = 0.242132:0.418537:1.81922;
		specparam tpd_C_Y_r = 0.180865:0.315302:1.44481;
		specparam tpd_C_Y_f = 0.31389:0.514362:2.12031;
		specparam tpd_D_Y_r = 0.211791:0.352415:1.55141;
		specparam tpd_D_Y_f = 0.342722:0.530151:1.97861;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA33 
`timescale 1ns/10ps
`celldefine
module OA33X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;

	and (int_fwire_0, C, F);
	and (int_fwire_1, C, E);
	and (int_fwire_2, C, D);
	and (int_fwire_3, B, F);
	and (int_fwire_4, B, E);
	and (int_fwire_5, B, D);
	and (int_fwire_6, A, F);
	and (int_fwire_7, A, E);
	and (int_fwire_8, A, D);
	or (Y, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0999207:0.225412:1.35125;
		specparam tpd_A_Y_f = 0.170884:0.299962:1.26501;
		specparam tpd_B_Y_r = 0.112569:0.244986:1.41002;
		specparam tpd_B_Y_f = 0.221322:0.332249:1.25387;
		specparam tpd_C_Y_r = 0.118043:0.257598:1.47195;
		specparam tpd_C_Y_f = 0.243171:0.350089:1.17633;
		specparam tpd_D_Y_r = 0.124192:0.249474:1.35986;
		specparam tpd_D_Y_f = 0.197006:0.321115:1.28801;
		specparam tpd_E_Y_r = 0.137777:0.270115:1.42387;
		specparam tpd_E_Y_f = 0.253492:0.359786:1.2824;
		specparam tpd_F_Y_r = 0.142196:0.280772:1.48288;
		specparam tpd_F_Y_f = 0.274538:0.376235:1.20485;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA33 
`timescale 1ns/10ps
`celldefine
module OA33X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;

	and (int_fwire_0, C, F);
	and (int_fwire_1, C, E);
	and (int_fwire_2, C, D);
	and (int_fwire_3, B, F);
	and (int_fwire_4, B, E);
	and (int_fwire_5, B, D);
	and (int_fwire_6, A, F);
	and (int_fwire_7, A, E);
	and (int_fwire_8, A, D);
	or (Y, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.139392:0.278355:1.44553;
		specparam tpd_A_Y_f = 0.265207:0.379391:1.20743;
		specparam tpd_B_Y_r = 0.156767:0.299054:1.51505;
		specparam tpd_B_Y_f = 0.314582:0.413624:1.15494;
		specparam tpd_C_Y_r = 0.175158:0.321996:1.61219;
		specparam tpd_C_Y_f = 0.334447:0.428115:1.03324;
		specparam tpd_D_Y_r = 0.169524:0.310141:1.48535;
		specparam tpd_D_Y_f = 0.284983:0.393862:1.21152;
		specparam tpd_E_Y_r = 0.182004:0.32426:1.52669;
		specparam tpd_E_Y_f = 0.340897:0.435699:1.17778;
		specparam tpd_F_Y_r = 0.188053:0.332971:1.57467;
		specparam tpd_F_Y_f = 0.36382:0.454469:1.08138;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA33 
`timescale 1ns/10ps
`celldefine
module OA33XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;

	and (int_fwire_0, C, F);
	and (int_fwire_1, C, E);
	and (int_fwire_2, C, D);
	and (int_fwire_3, B, F);
	and (int_fwire_4, B, E);
	and (int_fwire_5, B, D);
	and (int_fwire_6, A, F);
	and (int_fwire_7, A, E);
	and (int_fwire_8, A, D);
	or (Y, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.109248:0.23422:1.33988;
		specparam tpd_A_Y_f = 0.188766:0.31382:1.24091;
		specparam tpd_B_Y_r = 0.122062:0.253361:1.39949;
		specparam tpd_B_Y_f = 0.244126:0.351272:1.22485;
		specparam tpd_C_Y_r = 0.129492:0.26817:1.4719;
		specparam tpd_C_Y_f = 0.266065:0.369359:1.13616;
		specparam tpd_D_Y_r = 0.135286:0.259385:1.34704;
		specparam tpd_D_Y_f = 0.210918:0.329244:1.24634;
		specparam tpd_E_Y_r = 0.14847:0.278995:1.40849;
		specparam tpd_E_Y_f = 0.272803:0.374326:1.23654;
		specparam tpd_F_Y_r = 0.152102:0.288257:1.46345;
		specparam tpd_F_Y_f = 0.295427:0.393274:1.1577;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA44 
`timescale 1ns/10ps
`celldefine
module OA44X1 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;
	wire int_fwire_9, int_fwire_10, int_fwire_11;
	wire int_fwire_12, int_fwire_13, int_fwire_14;
	wire int_fwire_15;

	and (int_fwire_0, D, H);
	and (int_fwire_1, D, G);
	and (int_fwire_2, D, F);
	and (int_fwire_3, D, E);
	and (int_fwire_4, C, H);
	and (int_fwire_5, C, G);
	and (int_fwire_6, C, F);
	and (int_fwire_7, C, E);
	and (int_fwire_8, B, H);
	and (int_fwire_9, B, G);
	and (int_fwire_10, B, F);
	and (int_fwire_11, B, E);
	and (int_fwire_12, A, H);
	and (int_fwire_13, A, G);
	and (int_fwire_14, A, F);
	and (int_fwire_15, A, E);
	or (Y, int_fwire_15, int_fwire_14, int_fwire_13, int_fwire_12, int_fwire_11, int_fwire_10, int_fwire_9, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.106089:0.238997:1.42208;
		specparam tpd_A_Y_f = 0.134278:0.271032:1.26631;
		specparam tpd_B_Y_r = 0.136949:0.27936:1.52421;
		specparam tpd_B_Y_f = 0.22779:0.350554:1.31905;
		specparam tpd_C_Y_r = 0.15348:0.302034:1.60944;
		specparam tpd_C_Y_f = 0.28307:0.406221:1.29687;
		specparam tpd_D_Y_r = 0.163848:0.319842:1.70079;
		specparam tpd_D_Y_f = 0.308925:0.432086:1.25138;
		specparam tpd_E_Y_r = 0.129549:0.262041:1.43143;
		specparam tpd_E_Y_f = 0.163581:0.29387:1.28237;
		specparam tpd_F_Y_r = 0.160019:0.301976:1.53695;
		specparam tpd_F_Y_f = 0.258409:0.374099:1.33376;
		specparam tpd_G_Y_r = 0.175481:0.322561:1.62219;
		specparam tpd_G_Y_f = 0.313782:0.429564:1.31133;
		specparam tpd_H_Y_r = 0.184586:0.33807:1.71032;
		specparam tpd_H_Y_f = 0.339608:0.455435:1.26549;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA44 
`timescale 1ns/10ps
`celldefine
module OA44X4 (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;
	wire int_fwire_9, int_fwire_10, int_fwire_11;
	wire int_fwire_12, int_fwire_13, int_fwire_14;
	wire int_fwire_15;

	and (int_fwire_0, D, H);
	and (int_fwire_1, D, G);
	and (int_fwire_2, D, F);
	and (int_fwire_3, D, E);
	and (int_fwire_4, C, H);
	and (int_fwire_5, C, G);
	and (int_fwire_6, C, F);
	and (int_fwire_7, C, E);
	and (int_fwire_8, B, H);
	and (int_fwire_9, B, G);
	and (int_fwire_10, B, F);
	and (int_fwire_11, B, E);
	and (int_fwire_12, A, H);
	and (int_fwire_13, A, G);
	and (int_fwire_14, A, F);
	and (int_fwire_15, A, E);
	or (Y, int_fwire_15, int_fwire_14, int_fwire_13, int_fwire_12, int_fwire_11, int_fwire_10, int_fwire_9, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.149291:0.293498:1.53993;
		specparam tpd_A_Y_f = 0.180446:0.295181:1.02644;
		specparam tpd_B_Y_r = 0.181216:0.327553:1.62485;
		specparam tpd_B_Y_f = 0.279077:0.376964:1.05417;
		specparam tpd_C_Y_r = 0.202151:0.349093:1.70101;
		specparam tpd_C_Y_f = 0.334503:0.431785:1.01585;
		specparam tpd_D_Y_r = 0.21923:0.371617:1.79287;
		specparam tpd_D_Y_f = 0.360295:0.457421:0.961279;
		specparam tpd_E_Y_r = 0.175081:0.319002:1.55627;
		specparam tpd_E_Y_f = 0.19719:0.306803:1.02994;
		specparam tpd_F_Y_r = 0.205071:0.351755:1.64221;
		specparam tpd_F_Y_f = 0.295842:0.389053:1.05879;
		specparam tpd_G_Y_r = 0.223709:0.372198:1.71793;
		specparam tpd_G_Y_f = 0.35128:0.443889:1.02106;
		specparam tpd_H_Y_r = 0.237901:0.390841:1.80318;
		specparam tpd_H_Y_f = 0.377193:0.469528:0.967553;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OA44 
`timescale 1ns/10ps
`celldefine
module OA44XL (Y, A, B, C, D, E, F, G, H);
	output Y;
	input A, B, C, D, E, F, G, H;

	// Function
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3, int_fwire_4, int_fwire_5;
	wire int_fwire_6, int_fwire_7, int_fwire_8;
	wire int_fwire_9, int_fwire_10, int_fwire_11;
	wire int_fwire_12, int_fwire_13, int_fwire_14;
	wire int_fwire_15;

	and (int_fwire_0, D, H);
	and (int_fwire_1, D, G);
	and (int_fwire_2, D, F);
	and (int_fwire_3, D, E);
	and (int_fwire_4, C, H);
	and (int_fwire_5, C, G);
	and (int_fwire_6, C, F);
	and (int_fwire_7, C, E);
	and (int_fwire_8, B, H);
	and (int_fwire_9, B, G);
	and (int_fwire_10, B, F);
	and (int_fwire_11, B, E);
	and (int_fwire_12, A, H);
	and (int_fwire_13, A, G);
	and (int_fwire_14, A, F);
	and (int_fwire_15, A, E);
	or (Y, int_fwire_15, int_fwire_14, int_fwire_13, int_fwire_12, int_fwire_11, int_fwire_10, int_fwire_9, int_fwire_8, int_fwire_7, int_fwire_6, int_fwire_5, int_fwire_4, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.108997:0.235974:1.31909;
		specparam tpd_A_Y_f = 0.215694:0.350078:1.35513;
		specparam tpd_B_Y_r = 0.121396:0.254073:1.36805;
		specparam tpd_B_Y_f = 0.308194:0.420752:1.368;
		specparam tpd_C_Y_r = 0.127215:0.265604:1.4208;
		specparam tpd_C_Y_f = 0.367665:0.480896:1.3237;
		specparam tpd_D_Y_r = 0.125924:0.268975:1.46035;
		specparam tpd_D_Y_f = 0.388917:0.499495:1.25976;
		specparam tpd_E_Y_r = 0.134775:0.260763:1.32763;
		specparam tpd_E_Y_f = 0.242478:0.370023:1.37129;
		specparam tpd_F_Y_r = 0.147246:0.278901:1.37989;
		specparam tpd_F_Y_f = 0.338471:0.444145:1.38746;
		specparam tpd_G_Y_r = 0.152292:0.289487:1.43187;
		specparam tpd_G_Y_f = 0.400437:0.50713:1.34608;
		specparam tpd_H_Y_r = 0.150753:0.291846:1.46613;
		specparam tpd_H_Y_f = 0.423025:0.527567:1.28516;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
		(G => Y) = ( tpd_G_Y_r , tpd_G_Y_f );
		(H => Y) = ( tpd_H_Y_r , tpd_H_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI211 
`timescale 1ns/10ps
`celldefine
module OAI211X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0445534:0.143012:1.171;
		specparam tpd_A_Y_f = 0.079694:0.180881:1.28399;
		specparam tpd_B_Y_r = 0.0539987:0.157231:1.20626;
		specparam tpd_B_Y_f = 0.0922087:0.18084:1.1935;
		specparam tpd_C_Y_r = 0.120568:0.252902:1.76401;
		specparam tpd_C_Y_f = 0.0886755:0.168617:1.07559;
		specparam tpd_D_Y_r = 0.142629:0.258722:1.60276;
		specparam tpd_D_Y_f = 0.106229:0.186708:1.07008;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI211 
`timescale 1ns/10ps
`celldefine
module OAI211X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.161298:0.309643:1.62245;
		specparam tpd_A_Y_f = 0.273228:0.395129:1.30427;
		specparam tpd_B_Y_r = 0.17197:0.3234:1.67695;
		specparam tpd_B_Y_f = 0.286267:0.39554:1.25759;
		specparam tpd_C_Y_r = 0.265203:0.413937:1.89388;
		specparam tpd_C_Y_f = 0.2721:0.373215:1.11099;
		specparam tpd_D_Y_r = 0.287442:0.420644:1.80415;
		specparam tpd_D_Y_f = 0.300664:0.402586:1.17097;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI211 
`timescale 1ns/10ps
`celldefine
module OAI211XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0660331:0.171829:1.21665;
		specparam tpd_A_Y_f = 0.109556:0.199892:1.17479;
		specparam tpd_B_Y_r = 0.0785899:0.187633:1.24999;
		specparam tpd_B_Y_f = 0.125761:0.203741:1.09232;
		specparam tpd_C_Y_r = 0.195327:0.325447:1.83449;
		specparam tpd_C_Y_f = 0.124505:0.196463:0.938191;
		specparam tpd_D_Y_r = 0.224612:0.343489:1.67648;
		specparam tpd_D_Y_f = 0.152827:0.229169:1.00019;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21A 
`timescale 1ns/10ps
`celldefine
module OAI21AX1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire B__bar, C__bar, int_fwire_0;

	not (C__bar, C);
	not (B__bar, B);
	and (int_fwire_0, B__bar, C__bar);
	or (Y, A, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0860116:0.167784:0.744815;
		specparam tpd_A_Y_f = 0.11961:0.22228:1.03632;
		specparam tpd_B_Y_r = 0.0868471:0.22189:1.75867;
		specparam tpd_B_Y_f = 0.0612548:0.141646:1.07492;
		specparam tpd_C_Y_r = 0.109621:0.226312:1.58183;
		specparam tpd_C_Y_f = 0.0803753:0.168032:1.13455;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21A 
`timescale 1ns/10ps
`celldefine
module OAI21AX4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire B__bar, C__bar, int_fwire_0;

	not (C__bar, C);
	not (B__bar, B);
	and (int_fwire_0, B__bar, C__bar);
	or (Y, A, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.208091:0.340345:1.53935;
		specparam tpd_A_Y_f = 0.283349:0.409329:1.26763;
		specparam tpd_B_Y_r = 0.234337:0.382262:1.8276;
		specparam tpd_B_Y_f = 0.209581:0.315488:1.02863;
		specparam tpd_C_Y_r = 0.25905:0.390071:1.72623;
		specparam tpd_C_Y_f = 0.239779:0.351509:1.14012;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21A 
`timescale 1ns/10ps
`celldefine
module OAI21AXL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire B__bar, C__bar, int_fwire_0;

	not (C__bar, C);
	not (B__bar, B);
	and (int_fwire_0, B__bar, C__bar);
	or (Y, A, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.104901:0.181388:0.73487;
		specparam tpd_A_Y_f = 0.124787:0.219252:0.927098;
		specparam tpd_B_Y_r = 0.142574:0.277107:1.83271;
		specparam tpd_B_Y_f = 0.0785269:0.149418:0.902674;
		specparam tpd_C_Y_r = 0.171764:0.292698:1.66546;
		specparam tpd_C_Y_f = 0.0978236:0.174024:0.941295;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21BB 
`timescale 1ns/10ps
`celldefine
module OAI21BBX1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire C__bar, int_fwire_0;

	not (C__bar, C);
	and (int_fwire_0, A, B);
	or (Y, int_fwire_0, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.104485:0.222714:1.26722;
		specparam tpd_A_Y_f = 0.101828:0.245438:1.58615;
		specparam tpd_B_Y_r = 0.111876:0.218996:1.22889;
		specparam tpd_B_Y_f = 0.109902:0.258415:1.63303;
		specparam tpd_C_Y_r = 0.0420488:0.18119:1.73184;
		specparam tpd_C_Y_f = 0.0505881:0.172874:1.69706;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21BB 
`timescale 1ns/10ps
`celldefine
module OAI21BBX4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire C__bar, int_fwire_0;

	not (C__bar, C);
	and (int_fwire_0, A, B);
	or (Y, int_fwire_0, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.218936:0.347881:1.56644;
		specparam tpd_A_Y_f = 0.249062:0.368752:1.11874;
		specparam tpd_B_Y_r = 0.226414:0.343983:1.52129;
		specparam tpd_B_Y_f = 0.257384:0.381643:1.17197;
		specparam tpd_C_Y_r = 0.154211:0.302265:1.65239;
		specparam tpd_C_Y_f = 0.195227:0.291728:0.930577;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21BB 
`timescale 1ns/10ps
`celldefine
module OAI21BBXL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire C__bar, int_fwire_0;

	not (C__bar, C);
	and (int_fwire_0, A, B);
	or (Y, int_fwire_0, C__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.130844:0.243786:1.22769;
		specparam tpd_A_Y_f = 0.12995:0.269633:1.47684;
		specparam tpd_B_Y_r = 0.139776:0.241123:1.19041;
		specparam tpd_B_Y_f = 0.145176:0.28965:1.53742;
		specparam tpd_C_Y_r = 0.0619719:0.209112:1.84253;
		specparam tpd_C_Y_f = 0.0573175:0.153881:1.3695;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21B 
`timescale 1ns/10ps
`celldefine
module OAI21BX1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, int_fwire_0;

	not (B__bar, B);
	and (int_fwire_0, B__bar, C);
	not (A__bar, A);
	or (Y, A__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.037836:0.135885:1.18201;
		specparam tpd_A_Y_f = 0.0439711:0.124742:0.939784;
		specparam tpd_B_Y_r = 0.09955:0.234614:1.77572;
		specparam tpd_B_Y_f = 0.0473718:0.109193:0.793318;
		specparam tpd_C_Y_r = 0.175327:0.289802:1.31998;
		specparam tpd_C_Y_f = 0.118169:0.208601:0.823039;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21B 
`timescale 1ns/10ps
`celldefine
module OAI21BX4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, int_fwire_0;

	not (B__bar, B);
	and (int_fwire_0, B__bar, C);
	not (A__bar, A);
	or (Y, A__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.174132:0.323272:1.66756;
		specparam tpd_A_Y_f = 0.203057:0.317846:1.03176;
		specparam tpd_B_Y_r = 0.258754:0.411287:1.89765;
		specparam tpd_B_Y_f = 0.193471:0.291547:0.871692;
		specparam tpd_C_Y_r = 0.330825:0.462123:1.65779;
		specparam tpd_C_Y_f = 0.275655:0.39228:1.13843;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21B 
`timescale 1ns/10ps
`celldefine
module OAI21BXL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, int_fwire_0;

	not (B__bar, B);
	and (int_fwire_0, B__bar, C);
	not (A__bar, A);
	or (Y, A__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0522803:0.157951:1.2355;
		specparam tpd_A_Y_f = 0.0638104:0.144267:0.921053;
		specparam tpd_B_Y_r = 0.149763:0.283722:1.8504;
		specparam tpd_B_Y_f = 0.0689994:0.129458:0.760807;
		specparam tpd_C_Y_r = 0.234816:0.342812:1.35335;
		specparam tpd_C_Y_f = 0.138674:0.225192:0.831518;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21 
`timescale 1ns/10ps
`celldefine
module OAI21X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0;

	not (C__bar, C);
	not (B__bar, B);
	and (int_fwire_0, B__bar, C__bar);
	not (A__bar, A);
	or (Y, A__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0343626:0.129732:1.16925;
		specparam tpd_A_Y_f = 0.0608064:0.166012:1.29505;
		specparam tpd_B_Y_r = 0.0832859:0.217923:1.74222;
		specparam tpd_B_Y_f = 0.0599254:0.144509:1.11629;
		specparam tpd_C_Y_r = 0.105072:0.221162:1.5629;
		specparam tpd_C_Y_f = 0.0803565:0.17453:1.2009;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21 
`timescale 1ns/10ps
`celldefine
module OAI21X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0;

	not (C__bar, C);
	not (B__bar, B);
	and (int_fwire_0, B__bar, C__bar);
	not (A__bar, A);
	or (Y, A__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.172046:0.318561:1.62938;
		specparam tpd_A_Y_f = 0.207825:0.322496:1.03741;
		specparam tpd_B_Y_r = 0.256555:0.407253:1.86207;
		specparam tpd_B_Y_f = 0.199469:0.297817:0.878639;
		specparam tpd_C_Y_r = 0.27868:0.411088:1.75574;
		specparam tpd_C_Y_f = 0.227907:0.333293:0.994972;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI21 
`timescale 1ns/10ps
`celldefine
module OAI21XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0;

	not (C__bar, C);
	not (B__bar, B);
	and (int_fwire_0, B__bar, C__bar);
	not (A__bar, A);
	or (Y, A__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0465642:0.151968:1.24439;
		specparam tpd_A_Y_f = 0.0595293:0.140703:0.938314;
		specparam tpd_B_Y_r = 0.131842:0.268319:1.84279;
		specparam tpd_B_Y_f = 0.063564:0.12386:0.774955;
		specparam tpd_C_Y_r = 0.161292:0.282362:1.674;
		specparam tpd_C_Y_f = 0.0802831:0.14839:0.830302;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI221 
`timescale 1ns/10ps
`celldefine
module OAI221X1 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.106817:0.234734:1.69806;
		specparam tpd_A_Y_f = 0.13309:0.236352:1.44432;
		specparam tpd_B_Y_r = 0.130524:0.242216:1.53097;
		specparam tpd_B_Y_f = 0.158671:0.259318:1.42817;
		specparam tpd_C_Y_r = 0.128264:0.256918:1.7104;
		specparam tpd_C_Y_f = 0.150257:0.248721:1.33575;
		specparam tpd_D_Y_r = 0.150683:0.26379:1.53693;
		specparam tpd_D_Y_f = 0.176998:0.273965:1.33761;
		specparam tpd_E_Y_r = 0.0433444:0.138681:1.12363;
		specparam tpd_E_Y_f = 0.127268:0.237939:1.51036;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI221 
`timescale 1ns/10ps
`celldefine
module OAI221X4 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.283721:0.433048:1.90244;
		specparam tpd_A_Y_f = 0.318154:0.423981:1.15499;
		specparam tpd_B_Y_r = 0.3077:0.441681:1.81106;
		specparam tpd_B_Y_f = 0.347282:0.452052:1.208;
		specparam tpd_C_Y_r = 0.310515:0.460074:1.96278;
		specparam tpd_C_Y_f = 0.335016:0.436205:1.10451;
		specparam tpd_D_Y_r = 0.333277:0.467536:1.85443;
		specparam tpd_D_Y_f = 0.365942:0.467164:1.1578;
		specparam tpd_E_Y_r = 0.176435:0.326208:1.65529;
		specparam tpd_E_Y_f = 0.314597:0.429775:1.25832;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI221 
`timescale 1ns/10ps
`celldefine
module OAI221XL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1;

	not (E__bar, E);
	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0, E__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.203397:0.328491:1.79488;
		specparam tpd_A_Y_f = 0.139399:0.220181:1.0488;
		specparam tpd_B_Y_r = 0.235647:0.349002:1.63807;
		specparam tpd_B_Y_f = 0.161646:0.240373:1.05271;
		specparam tpd_C_Y_r = 0.253058:0.377568:1.83485;
		specparam tpd_C_Y_f = 0.163217:0.236606:0.92763;
		specparam tpd_D_Y_r = 0.281514:0.395595:1.66864;
		specparam tpd_D_Y_f = 0.188141:0.262044:0.961863;
		specparam tpd_E_Y_r = 0.0644317:0.168395:1.18726;
		specparam tpd_E_Y_f = 0.110756:0.193506:1.015;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI222 
`timescale 1ns/10ps
`celldefine
module OAI222X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	not (F__bar, F);
	not (E__bar, E);
	and (int_fwire_0, E__bar, F__bar);
	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_1, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_2, A__bar, B__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.248765:0.397252:1.84037;
		specparam tpd_A_Y_f = 0.280496:0.385537:1.15474;
		specparam tpd_B_Y_r = 0.272487:0.403502:1.72638;
		specparam tpd_B_Y_f = 0.32287:0.429399:1.26886;
		specparam tpd_C_Y_r = 0.303597:0.450291:1.93767;
		specparam tpd_C_Y_f = 0.328613:0.425117:1.1541;
		specparam tpd_D_Y_r = 0.329029:0.460381:1.81354;
		specparam tpd_D_Y_f = 0.375174:0.474993:1.26636;
		specparam tpd_E_Y_r = 0.327227:0.473273:1.97276;
		specparam tpd_E_Y_f = 0.360643:0.454669:1.14197;
		specparam tpd_F_Y_r = 0.349393:0.481483:1.85986;
		specparam tpd_F_Y_f = 0.394527:0.489512:1.19973;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI222 
`timescale 1ns/10ps
`celldefine
module OAI222X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	not (F__bar, F);
	not (E__bar, E);
	and (int_fwire_0, E__bar, F__bar);
	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_1, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_2, A__bar, B__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.275766:0.427777:1.87979;
		specparam tpd_A_Y_f = 0.330438:0.443428:1.2122;
		specparam tpd_B_Y_r = 0.299502:0.433729:1.76355;
		specparam tpd_B_Y_f = 0.373764:0.487981:1.32439;
		specparam tpd_C_Y_r = 0.328205:0.477544:1.96944;
		specparam tpd_C_Y_f = 0.378641:0.483043:1.2143;
		specparam tpd_D_Y_r = 0.353623:0.488004:1.84213;
		specparam tpd_D_Y_f = 0.427015:0.534678:1.32549;
		specparam tpd_E_Y_r = 0.353729:0.502829:2.00685;
		specparam tpd_E_Y_f = 0.410026:0.511576:1.19404;
		specparam tpd_F_Y_r = 0.37606:0.510906:1.88851;
		specparam tpd_F_Y_f = 0.446308:0.549217:1.25696;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI222 
`timescale 1ns/10ps
`celldefine
module OAI222XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;

	not (F__bar, F);
	not (E__bar, E);
	and (int_fwire_0, E__bar, F__bar);
	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_1, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_2, A__bar, B__bar);
	or (Y, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.125379:0.246704:1.60093;
		specparam tpd_A_Y_f = 0.124762:0.209164:1.03007;
		specparam tpd_B_Y_r = 0.155167:0.259409:1.41624;
		specparam tpd_B_Y_f = 0.161444:0.245237:1.12159;
		specparam tpd_C_Y_r = 0.242023:0.360866:1.74853;
		specparam tpd_C_Y_f = 0.199725:0.273239:1.003;
		specparam tpd_D_Y_r = 0.272158:0.378791:1.57841;
		specparam tpd_D_Y_f = 0.236994:0.314754:1.09756;
		specparam tpd_E_Y_r = 0.294436:0.413305:1.78898;
		specparam tpd_E_Y_f = 0.233512:0.306993:0.968705;
		specparam tpd_F_Y_r = 0.325408:0.433742:1.62949;
		specparam tpd_F_Y_f = 0.263952:0.337444:1.00625;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22A 
`timescale 1ns/10ps
`celldefine
module OAI22AX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0648143:0.193996:1.65372;
		specparam tpd_A_Y_f = 0.0624424:0.157888:1.13665;
		specparam tpd_B_Y_r = 0.0883501:0.197216:1.4691;
		specparam tpd_B_Y_f = 0.0856934:0.186357:1.21875;
		specparam tpd_C_Y_r = 0.112545:0.243618:1.7312;
		specparam tpd_C_Y_f = 0.0899102:0.175659:1.04361;
		specparam tpd_D_Y_r = 0.186882:0.300713:1.32955;
		specparam tpd_D_Y_f = 0.161331:0.253203:0.949485;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22A 
`timescale 1ns/10ps
`celldefine
module OAI22AX4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.228452:0.378259:1.82866;
		specparam tpd_A_Y_f = 0.217056:0.332272:1.00046;
		specparam tpd_B_Y_r = 0.251456:0.382622:1.72109;
		specparam tpd_B_Y_f = 0.246894:0.365781:1.118;
		specparam tpd_C_Y_r = 0.285161:0.436059:1.95048;
		specparam tpd_C_Y_f = 0.244337:0.350283:0.983637;
		specparam tpd_D_Y_r = 0.35918:0.493005:1.72857;
		specparam tpd_D_Y_f = 0.322651:0.433485:1.11805;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22A 
`timescale 1ns/10ps
`celldefine
module OAI22AXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.103841:0.233467:1.71014;
		specparam tpd_A_Y_f = 0.0691392:0.146488:0.84228;
		specparam tpd_B_Y_r = 0.138768:0.251823:1.54029;
		specparam tpd_B_Y_f = 0.0885873:0.168046:0.87716;
		specparam tpd_C_Y_r = 0.178751:0.306782:1.79759;
		specparam tpd_C_Y_f = 0.0983033:0.168597:0.796341;
		specparam tpd_D_Y_r = 0.256173:0.355487:1.23774;
		specparam tpd_D_Y_f = 0.182111:0.27516:0.914827;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22B 
`timescale 1ns/10ps
`celldefine
module OAI22BX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, C__bar, int_fwire_0;
	wire int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0712202:0.202383:1.6843;
		specparam tpd_A_Y_f = 0.0654238:0.158936:1.10442;
		specparam tpd_B_Y_r = 0.144235:0.250366:1.2247;
		specparam tpd_B_Y_f = 0.137622:0.231345:0.943301;
		specparam tpd_C_Y_r = 0.106837:0.237325:1.72372;
		specparam tpd_C_Y_f = 0.085897:0.169257:1.02487;
		specparam tpd_D_Y_r = 0.178239:0.28554:1.26745;
		specparam tpd_D_Y_f = 0.15495:0.246742:0.937465;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22B 
`timescale 1ns/10ps
`celldefine
module OAI22BX4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, C__bar, int_fwire_0;
	wire int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.2395:0.391551:1.85579;
		specparam tpd_A_Y_f = 0.223392:0.345949:1.11797;
		specparam tpd_B_Y_r = 0.3131:0.440546:1.60762;
		specparam tpd_B_Y_f = 0.301087:0.424216:1.27711;
		specparam tpd_C_Y_r = 0.280538:0.432926:1.93881;
		specparam tpd_C_Y_f = 0.244519:0.356992:1.10563;
		specparam tpd_D_Y_r = 0.352054:0.480802:1.6539;
		specparam tpd_D_Y_f = 0.318761:0.43978:1.2768;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22B 
`timescale 1ns/10ps
`celldefine
module OAI22BXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, C__bar, int_fwire_0;
	wire int_fwire_1;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.102383:0.22752:1.63607;
		specparam tpd_A_Y_f = 0.0668085:0.141331:0.789869;
		specparam tpd_B_Y_r = 0.19846:0.295799:1.10818;
		specparam tpd_B_Y_f = 0.16549:0.260029:0.892339;
		specparam tpd_C_Y_r = 0.194854:0.322388:1.81603;
		specparam tpd_C_Y_f = 0.102305:0.172877:0.786889;
		specparam tpd_D_Y_r = 0.272045:0.370594:1.24952;
		specparam tpd_D_Y_f = 0.178553:0.268959:0.873043;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22C 
`timescale 1ns/10ps
`celldefine
module OAI22CX1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire C__bar, D__bar, int_fwire_0;
	wire int_fwire_1;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.107627:0.19114:0.714005;
		specparam tpd_A_Y_f = 0.159565:0.278744:1.19617;
		specparam tpd_B_Y_r = 0.115567:0.189254:0.690348;
		specparam tpd_B_Y_f = 0.170826:0.291746:1.2339;
		specparam tpd_C_Y_r = 0.116129:0.233424:1.58798;
		specparam tpd_C_Y_f = 0.0799821:0.167651:1.1046;
		specparam tpd_D_Y_r = 0.0911799:0.226567:1.76503;
		specparam tpd_D_Y_f = 0.0599013:0.13788:1.02161;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22C 
`timescale 1ns/10ps
`celldefine
module OAI22CX4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire C__bar, D__bar, int_fwire_0;
	wire int_fwire_1;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.235216:0.362417:1.50278;
		specparam tpd_A_Y_f = 0.315769:0.449675:1.34174;
		specparam tpd_B_Y_r = 0.243116:0.36048:1.47483;
		specparam tpd_B_Y_f = 0.327227:0.463356:1.38325;
		specparam tpd_C_Y_r = 0.272003:0.403543:1.76837;
		specparam tpd_C_Y_f = 0.233844:0.338695:0.99961;
		specparam tpd_D_Y_r = 0.247258:0.396693:1.87819;
		specparam tpd_D_Y_f = 0.205346:0.303373:0.884113;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22C 
`timescale 1ns/10ps
`celldefine
module OAI22CXL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire C__bar, D__bar, int_fwire_0;
	wire int_fwire_1;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.14194:0.224255:0.783241;
		specparam tpd_A_Y_f = 0.15188:0.256665:0.988886;
		specparam tpd_B_Y_r = 0.151111:0.222145:0.756273;
		specparam tpd_B_Y_f = 0.159939:0.266956:1.0162;
		specparam tpd_C_Y_r = 0.179323:0.301736:1.71623;
		specparam tpd_C_Y_f = 0.0797992:0.151591:0.838652;
		specparam tpd_D_Y_r = 0.149359:0.285511:1.88583;
		specparam tpd_D_Y_f = 0.0648262:0.129232:0.785579;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22 
`timescale 1ns/10ps
`celldefine
module OAI22X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0639271:0.195074:1.68082;
		specparam tpd_A_Y_f = 0.0627943:0.160742:1.17431;
		specparam tpd_B_Y_r = 0.0874623:0.198459:1.49949;
		specparam tpd_B_Y_f = 0.0864608:0.189139:1.25557;
		specparam tpd_C_Y_r = 0.11123:0.242983:1.73701;
		specparam tpd_C_Y_f = 0.0911244:0.179336:1.07689;
		specparam tpd_D_Y_r = 0.134289:0.248813:1.55733;
		specparam tpd_D_Y_f = 0.116292:0.210497:1.16773;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22 
`timescale 1ns/10ps
`celldefine
module OAI22X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.228942:0.377896:1.80473;
		specparam tpd_A_Y_f = 0.21979:0.334357:0.997305;
		specparam tpd_B_Y_r = 0.251907:0.381579:1.69775;
		specparam tpd_B_Y_f = 0.250025:0.367877:1.11438;
		specparam tpd_C_Y_r = 0.283797:0.433036:1.92135;
		specparam tpd_C_Y_f = 0.24719:0.352866:0.982184;
		specparam tpd_D_Y_r = 0.306736:0.438658:1.79828;
		specparam tpd_D_Y_f = 0.279946:0.389565:1.09144;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI22 
`timescale 1ns/10ps
`celldefine
module OAI22XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0, int_fwire_1;

	not (D__bar, D);
	not (C__bar, C);
	and (int_fwire_0, C__bar, D__bar);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.103071:0.233732:1.72771;
		specparam tpd_A_Y_f = 0.0687191:0.150484:0.903117;
		specparam tpd_B_Y_r = 0.135331:0.24946:1.55049;
		specparam tpd_B_Y_f = 0.0944091:0.181381:0.99764;
		specparam tpd_C_Y_r = 0.197796:0.326591:1.82546;
		specparam tpd_C_Y_f = 0.110441:0.182803:0.827308;
		specparam tpd_D_Y_r = 0.227156:0.342301:1.65784;
		specparam tpd_D_Y_f = 0.131547:0.20525:0.865764;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI2B11 
`timescale 1ns/10ps
`celldefine
module OAI2B11X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.04493:0.14392:1.17675;
		specparam tpd_A_Y_f = 0.0931114:0.201509:1.42295;
		specparam tpd_B_Y_r = 0.0535003:0.156568:1.20095;
		specparam tpd_B_Y_f = 0.108338:0.205391:1.34564;
		specparam tpd_C_Y_r = 0.121343:0.253771:1.76161;
		specparam tpd_C_Y_f = 0.100299:0.187865:1.18134;
		specparam tpd_D_Y_r = 0.19278:0.307766:1.3515;
		specparam tpd_D_Y_f = 0.173905:0.277985:1.17197;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI2B11 
`timescale 1ns/10ps
`celldefine
module OAI2B11X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.168341:0.317166:1.64409;
		specparam tpd_A_Y_f = 0.269668:0.383287:1.1593;
		specparam tpd_B_Y_r = 0.178668:0.33063:1.69017;
		specparam tpd_B_Y_f = 0.28474:0.387443:1.12846;
		specparam tpd_C_Y_r = 0.28188:0.430052:1.92493;
		specparam tpd_C_Y_f = 0.267949:0.363003:0.968206;
		specparam tpd_D_Y_r = 0.353158:0.48391:1.70573;
		specparam tpd_D_Y_f = 0.350085:0.460554:1.14515;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI2B11 
`timescale 1ns/10ps
`celldefine
module OAI2B11XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0;

	not (C__bar, C);
	and (int_fwire_0, C__bar, D);
	not (B__bar, B);
	not (A__bar, A);
	or (Y, A__bar, B__bar, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0601613:0.164346:1.19995;
		specparam tpd_A_Y_f = 0.0979968:0.186521:1.11798;
		specparam tpd_B_Y_r = 0.073068:0.181397:1.2396;
		specparam tpd_B_Y_f = 0.113325:0.18856:1.03083;
		specparam tpd_C_Y_r = 0.189989:0.321284:1.84166;
		specparam tpd_C_Y_f = 0.115298:0.184569:0.886557;
		specparam tpd_D_Y_r = 0.261105:0.369301:1.37364;
		specparam tpd_D_Y_f = 0.179174:0.261763:0.918612;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI31 
`timescale 1ns/10ps
`celldefine
module OAI31X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C__bar);
	or (Y, int_fwire_0, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.281374:0.425357:1.95661;
		specparam tpd_A_Y_f = 0.172252:0.266617:0.861069;
		specparam tpd_B_Y_r = 0.333386:0.461816:1.908;
		specparam tpd_B_Y_f = 0.197092:0.294855:0.944024;
		specparam tpd_C_Y_r = 0.355769:0.479996:1.79804;
		specparam tpd_C_Y_f = 0.214264:0.316852:1.0276;
		specparam tpd_D_Y_r = 0.140191:0.280588:1.59668;
		specparam tpd_D_Y_f = 0.19259:0.307425:1.10656;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI31 
`timescale 1ns/10ps
`celldefine
module OAI31X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C__bar);
	or (Y, int_fwire_0, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.306345:0.451502:1.96742;
		specparam tpd_A_Y_f = 0.215448:0.318195:0.898151;
		specparam tpd_B_Y_r = 0.358082:0.488963:1.92624;
		specparam tpd_B_Y_f = 0.2395:0.342889:0.957381;
		specparam tpd_C_Y_r = 0.380473:0.507244:1.81666;
		specparam tpd_C_Y_f = 0.259781:0.366326:1.03886;
		specparam tpd_D_Y_r = 0.153216:0.296869:1.60058;
		specparam tpd_D_Y_f = 0.238399:0.359885:1.13982;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI31 
`timescale 1ns/10ps
`celldefine
module OAI31XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, int_fwire_0;

	not (D__bar, D);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C__bar);
	or (Y, int_fwire_0, D__bar);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.132412:0.259484:1.73153;
		specparam tpd_A_Y_f = 0.0904959:0.166248:0.970612;
		specparam tpd_B_Y_r = 0.192:0.306921:1.64206;
		specparam tpd_B_Y_f = 0.126856:0.207824:1.05492;
		specparam tpd_C_Y_r = 0.214388:0.325346:1.50265;
		specparam tpd_C_Y_f = 0.147674:0.237097:1.1478;
		specparam tpd_D_Y_r = 0.0392254:0.120447:0.926416;
		specparam tpd_D_Y_f = 0.112803:0.212806:1.23302;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI32 
`timescale 1ns/10ps
`celldefine
module OAI32X1 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1;

	not (E__bar, E);
	not (D__bar, D);
	and (int_fwire_0, D__bar, E__bar);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0934645:0.219029:1.64867;
		specparam tpd_A_Y_f = 0.074924:0.160171:0.930478;
		specparam tpd_B_Y_r = 0.14847:0.256018:1.55199;
		specparam tpd_B_Y_f = 0.0988842:0.185045:0.972365;
		specparam tpd_C_Y_r = 0.170854:0.273579:1.40576;
		specparam tpd_C_Y_f = 0.113557:0.203041:1.03624;
		specparam tpd_D_Y_r = 0.119624:0.226967:1.37017;
		specparam tpd_D_Y_f = 0.109632:0.189945:0.888969;
		specparam tpd_E_Y_r = 0.144569:0.233804:1.18474;
		specparam tpd_E_Y_f = 0.140426:0.221785:0.961868;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI32 
`timescale 1ns/10ps
`celldefine
module OAI32X4 (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1;

	not (E__bar, E);
	not (D__bar, D);
	and (int_fwire_0, D__bar, E__bar);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.304702:0.455235:1.99111;
		specparam tpd_A_Y_f = 0.234113:0.35196:1.01624;
		specparam tpd_B_Y_r = 0.359878:0.493515:1.94107;
		specparam tpd_B_Y_f = 0.260831:0.378194:1.09362;
		specparam tpd_C_Y_r = 0.382607:0.511785:1.8311;
		specparam tpd_C_Y_f = 0.283333:0.401507:1.17871;
		specparam tpd_D_Y_r = 0.298996:0.450776:1.97405;
		specparam tpd_D_Y_f = 0.27714:0.386421:1.07754;
		specparam tpd_E_Y_r = 0.323928:0.458425:1.8564;
		specparam tpd_E_Y_f = 0.309953:0.420844:1.16473;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI32 
`timescale 1ns/10ps
`celldefine
module OAI32XL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, int_fwire_0;
	wire int_fwire_1;

	not (E__bar, E);
	not (D__bar, D);
	and (int_fwire_0, D__bar, E__bar);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.125909:0.250713:1.69191;
		specparam tpd_A_Y_f = 0.0837998:0.161188:0.803591;
		specparam tpd_B_Y_r = 0.195185:0.303808:1.60434;
		specparam tpd_B_Y_f = 0.110505:0.188041:0.852097;
		specparam tpd_C_Y_r = 0.221984:0.328363:1.47246;
		specparam tpd_C_Y_f = 0.125871:0.205701:0.91798;
		specparam tpd_D_Y_r = 0.166762:0.27364:1.44083;
		specparam tpd_D_Y_f = 0.130152:0.201656:0.77891;
		specparam tpd_E_Y_r = 0.195702:0.286804:1.2602;
		specparam tpd_E_Y_f = 0.163098:0.234408:0.848718;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI33 
`timescale 1ns/10ps
`celldefine
module OAI33X1 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	and (int_fwire_0, D__bar, E__bar, F__bar);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.373012:0.517366:2.06582;
		specparam tpd_A_Y_f = 0.288523:0.398102:1.18028;
		specparam tpd_B_Y_r = 0.42516:0.557707:2.02427;
		specparam tpd_B_Y_f = 0.309514:0.415662:1.20119;
		specparam tpd_C_Y_r = 0.44843:0.5775:1.92038;
		specparam tpd_C_Y_f = 0.330261:0.436047:1.24774;
		specparam tpd_D_Y_r = 0.280218:0.427171:1.93153;
		specparam tpd_D_Y_f = 0.246142:0.362766:1.16809;
		specparam tpd_E_Y_r = 0.337155:0.468176:1.89929;
		specparam tpd_E_Y_f = 0.274855:0.388602:1.22556;
		specparam tpd_F_Y_r = 0.360521:0.487868:1.80532;
		specparam tpd_F_Y_f = 0.296132:0.408307:1.28283;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI33 
`timescale 1ns/10ps
`celldefine
module OAI33X4 (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	and (int_fwire_0, D__bar, E__bar, F__bar);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.399545:0.547193:2.10375;
		specparam tpd_A_Y_f = 0.331553:0.446109:1.18777;
		specparam tpd_B_Y_r = 0.451605:0.587645:2.05953;
		specparam tpd_B_Y_f = 0.352:0.463167:1.20628;
		specparam tpd_C_Y_r = 0.47488:0.607671:1.95556;
		specparam tpd_C_Y_f = 0.373785:0.484431:1.25182;
		specparam tpd_D_Y_r = 0.306582:0.456407:1.97384;
		specparam tpd_D_Y_f = 0.288496:0.409559:1.17584;
		specparam tpd_E_Y_r = 0.363455:0.497829:1.93711;
		specparam tpd_E_Y_f = 0.317259:0.435839:1.2306;
		specparam tpd_F_Y_r = 0.386806:0.517449:1.84253;
		specparam tpd_F_Y_f = 0.339649:0.45674:1.28743;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OAI33 
`timescale 1ns/10ps
`celldefine
module OAI33XL (Y, A, B, C, D, E, F);
	output Y;
	input A, B, C, D, E, F;

	// Function
	wire A__bar, B__bar, C__bar;
	wire D__bar, E__bar, F__bar;
	wire int_fwire_0, int_fwire_1;

	not (F__bar, F);
	not (E__bar, E);
	not (D__bar, D);
	and (int_fwire_0, D__bar, E__bar, F__bar);
	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_1, A__bar, B__bar, C__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.291173:0.400133:1.69712;
		specparam tpd_A_Y_f = 0.155511:0.228249:0.768595;
		specparam tpd_B_Y_r = 0.3538:0.452549:1.62322;
		specparam tpd_B_Y_f = 0.173187:0.240605:0.742791;
		specparam tpd_C_Y_r = 0.381354:0.479068:1.50189;
		specparam tpd_C_Y_f = 0.186767:0.2534:0.765709;
		specparam tpd_D_Y_r = 0.147387:0.261045:1.56019;
		specparam tpd_D_Y_f = 0.102875:0.183482:0.774086;
		specparam tpd_E_Y_r = 0.216453:0.314943:1.48133;
		specparam tpd_E_Y_f = 0.1283:0.203487:0.79359;
		specparam tpd_F_Y_r = 0.244104:0.340717:1.35961;
		specparam tpd_F_Y_f = 0.141809:0.215214:0.822524;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
		(E => Y) = ( tpd_E_Y_r , tpd_E_Y_f );
		(F => Y) = ( tpd_F_Y_r , tpd_F_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR2 
`timescale 1ns/10ps
`celldefine
module OR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0781907:0.2019:1.26602;
		specparam tpd_A_Y_f = 0.17604:0.33628:1.58767;
		specparam tpd_B_Y_r = 0.0843741:0.21286:1.30572;
		specparam tpd_B_Y_f = 0.204266:0.348033:1.527;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR2 
`timescale 1ns/10ps
`celldefine
module OR2X12 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.240939:0.375327:1.58149;
		specparam tpd_A_Y_f = 0.261004:0.381922:1.20248;
		specparam tpd_B_Y_r = 0.260101:0.402687:1.67337;
		specparam tpd_B_Y_f = 0.282689:0.387449:1.13428;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR2 
`timescale 1ns/10ps
`celldefine
module OR2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.112587:0.254885:1.45676;
		specparam tpd_A_Y_f = 0.159395:0.308503:1.37557;
		specparam tpd_B_Y_r = 0.125312:0.269143:1.49625;
		specparam tpd_B_Y_f = 0.183701:0.31698:1.3166;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR2 
`timescale 1ns/10ps
`celldefine
module OR2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.139183:0.291444:1.53598;
		specparam tpd_A_Y_f = 0.210355:0.368162:1.4941;
		specparam tpd_B_Y_r = 0.150296:0.301794:1.56678;
		specparam tpd_B_Y_f = 0.234636:0.377332:1.4182;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR2 
`timescale 1ns/10ps
`celldefine
module OR2X6 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.16296:0.330396:1.6738;
		specparam tpd_A_Y_f = 0.272855:0.447306:1.73053;
		specparam tpd_B_Y_r = 0.181266:0.349793:1.73414;
		specparam tpd_B_Y_f = 0.29498:0.454208:1.6242;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR2 
`timescale 1ns/10ps
`celldefine
module OR2X8 (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.195804:0.370601:1.76562;
		specparam tpd_A_Y_f = 0.337783:0.518757:1.85126;
		specparam tpd_B_Y_r = 0.215207:0.391435:1.82322;
		specparam tpd_B_Y_f = 0.359795:0.526226:1.72987;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR2 
`timescale 1ns/10ps
`celldefine
module OR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	or (Y, A, B);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.110837:0.240935:1.32942;
		specparam tpd_A_Y_f = 0.230603:0.41151:1.91;
		specparam tpd_B_Y_r = 0.1338:0.271834:1.43624;
		specparam tpd_B_Y_f = 0.263811:0.430446:1.80824;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR3 
`timescale 1ns/10ps
`celldefine
module OR3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.10265:0.2329:1.32771;
		specparam tpd_A_Y_f = 0.195042:0.344601:1.43471;
		specparam tpd_B_Y_r = 0.117687:0.252272:1.38334;
		specparam tpd_B_Y_f = 0.25676:0.38963:1.41653;
		specparam tpd_C_Y_r = 0.124564:0.265838:1.44709;
		specparam tpd_C_Y_f = 0.282111:0.412717:1.33248;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR3 
`timescale 1ns/10ps
`celldefine
module OR3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0869291:0.22267:1.38058;
		specparam tpd_A_Y_f = 0.153863:0.302257:1.35918;
		specparam tpd_B_Y_r = 0.100284:0.241509:1.43395;
		specparam tpd_B_Y_f = 0.202049:0.332817:1.3474;
		specparam tpd_C_Y_r = 0.106997:0.255683:1.49956;
		specparam tpd_C_Y_f = 0.222619:0.348442:1.26527;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR3 
`timescale 1ns/10ps
`celldefine
module OR3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0764281:0.203068:1.30175;
		specparam tpd_A_Y_f = 0.141547:0.29056:1.37255;
		specparam tpd_B_Y_r = 0.091981:0.228276:1.38343;
		specparam tpd_B_Y_f = 0.192399:0.322099:1.34987;
		specparam tpd_C_Y_r = 0.0989502:0.244844:1.46271;
		specparam tpd_C_Y_f = 0.213034:0.337899:1.26408;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR3 
`timescale 1ns/10ps
`celldefine
module OR3X6 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.147259:0.311155:1.58084;
		specparam tpd_A_Y_f = 0.40312:0.590876:2.0082;
		specparam tpd_B_Y_r = 0.160662:0.324511:1.61314;
		specparam tpd_B_Y_f = 0.458318:0.634732:1.95373;
		specparam tpd_C_Y_r = 0.175245:0.342433:1.68336;
		specparam tpd_C_Y_f = 0.479603:0.651271:1.83258;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR3 
`timescale 1ns/10ps
`celldefine
module OR3X8 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.174001:0.346676:1.68356;
		specparam tpd_A_Y_f = 0.503139:0.699562:2.18522;
		specparam tpd_B_Y_r = 0.187148:0.358785:1.71402;
		specparam tpd_B_Y_f = 0.55825:0.744575:2.12039;
		specparam tpd_C_Y_r = 0.208278:0.383673:1.79841;
		specparam tpd_C_Y_f = 0.579717:0.761059:1.98823;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR3 
`timescale 1ns/10ps
`celldefine
module OR3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	or (Y, A, B, C);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.109529:0.238001:1.28982;
		specparam tpd_A_Y_f = 0.260401:0.446428:1.95726;
		specparam tpd_B_Y_r = 0.12569:0.257406:1.34368;
		specparam tpd_B_Y_f = 0.330133:0.500398:1.928;
		specparam tpd_C_Y_r = 0.132768:0.270499:1.40669;
		specparam tpd_C_Y_f = 0.359137:0.528814:1.84051;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR4 
`timescale 1ns/10ps
`celldefine
module OR4X1 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	or (Y, A, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.121578:0.265252:1.42233;
		specparam tpd_A_Y_f = 0.253587:0.415831:1.58817;
		specparam tpd_B_Y_r = 0.131543:0.273769:1.42688;
		specparam tpd_B_Y_f = 0.354748:0.50084:1.61717;
		specparam tpd_C_Y_r = 0.138837:0.284757:1.47207;
		specparam tpd_C_Y_f = 0.411157:0.556741:1.56645;
		specparam tpd_D_Y_r = 0.140074:0.291582:1.51897;
		specparam tpd_D_Y_f = 0.434942:0.580023:1.50168;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR4 
`timescale 1ns/10ps
`celldefine
module OR4X2 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	or (Y, A, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0870281:0.223772:1.33776;
		specparam tpd_A_Y_f = 0.182953:0.366846:1.72583;
		specparam tpd_B_Y_r = 0.106799:0.244756:1.36779;
		specparam tpd_B_Y_f = 0.286877:0.447635:1.76461;
		specparam tpd_C_Y_r = 0.115585:0.260676:1.43629;
		specparam tpd_C_Y_f = 0.330416:0.48869:1.70777;
		specparam tpd_D_Y_r = 0.116218:0.27605:1.55394;
		specparam tpd_D_Y_f = 0.347872:0.502993:1.5951;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR4 
`timescale 1ns/10ps
`celldefine
module OR4X4 (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	or (Y, A, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.122638:0.28049:1.55351;
		specparam tpd_A_Y_f = 0.201262:0.381071:1.65496;
		specparam tpd_B_Y_r = 0.156973:0.31103:1.6022;
		specparam tpd_B_Y_f = 0.293261:0.452838:1.67686;
		specparam tpd_C_Y_r = 0.177214:0.334819:1.68176;
		specparam tpd_C_Y_f = 0.332928:0.489277:1.61608;
		specparam tpd_D_Y_r = 0.18433:0.353804:1.80423;
		specparam tpd_D_Y_f = 0.349103:0.501559:1.50924;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: OR4 
`timescale 1ns/10ps
`celldefine
module OR4XL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;

	// Function
	or (Y, A, B, C, D);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.125766:0.262697:1.36268;
		specparam tpd_A_Y_f = 0.27716:0.472306:2.01047;
		specparam tpd_B_Y_r = 0.147551:0.286639:1.41738;
		specparam tpd_B_Y_f = 0.392959:0.570275:2.02653;
		specparam tpd_C_Y_r = 0.152589:0.293688:1.44638;
		specparam tpd_C_Y_f = 0.454728:0.632131:1.98598;
		specparam tpd_D_Y_r = 0.148749:0.294207:1.4753;
		specparam tpd_D_Y_f = 0.479496:0.656658:1.93211;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(B => Y) = ( tpd_B_Y_r , tpd_B_Y_f );
		(C => Y) = ( tpd_C_Y_r , tpd_C_Y_f );
		(D => Y) = ( tpd_D_Y_r , tpd_D_Y_f );
	endspecify
endmodule
`endcelldefine

// type: SDFFNQ 
`timescale 1ns/10ps
`celldefine
module SDFFNQX1 (Q, D, SIN, SMC, XC);
	output Q;
	input D, SIN, SMC, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_XC_Q_negedge_r = 0.39382:0.558434:1.9964;
		specparam tpd_XC_Q_negedge_f = 0.298435:0.433777:1.33051;
		specparam tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = 0.181297:0.142984:-0.096976;
		specparam thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = -0.0318175:-0.00402285:0.232134;
		specparam tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = 0.181297:0.142984:-0.096976;
		specparam thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = -0.0318175:-0.00402285:0.232134;
		specparam tsetup_SIN_XC_SMC_posedge_SMC_negedge = 0.177272:0.140831:-0.101136;
		specparam thold_SIN_XC_SMC_posedge_SMC_negedge = -0.0297552:-0.00276833:0.235566;
		specparam tsetup_SIN_XC_SMC_negedge_SMC_negedge = 0.177272:0.140831:-0.101136;
		specparam thold_SIN_XC_SMC_negedge_SMC_negedge = -0.0297552:-0.00276833:0.235566;
		specparam tsetup_SMC_XC_adacond0_posedge_adacond0_negedge = 0.412731:0.374569:0.0903628;
		specparam thold_SMC_XC_adacond0_posedge_adacond0_negedge = -0.0051941:0.00664365:0.234925;
		specparam tsetup_SMC_XC_adacond0_negedge_adacond0_negedge = 0.412731:0.374569:0.0903628;
		specparam thold_SMC_XC_adacond0_negedge_adacond0_negedge = -0.0051941:0.00664365:0.234925;
		specparam tpw_XC_posedge = 0.225451:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.225451:0.330811:2.72095;

		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_posedge_SMC_negedge, 
			 thold_SIN_XC_SMC_posedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_negedge_SMC_negedge, 
			 thold_SIN_XC_SMC_negedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_posedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_negedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNQ 
`timescale 1ns/10ps
`celldefine
module SDFFNQX2 (Q, D, SIN, SMC, XC);
	output Q;
	input D, SIN, SMC, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_XC_Q_negedge_r = 0.376874:0.543549:1.99079;
		specparam tpd_XC_Q_negedge_f = 0.312041:0.45483:1.34774;
		specparam tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = 0.161309:0.122633:-0.112638;
		specparam thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = -0.0340213:-0.00842307:0.225867;
		specparam tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = 0.161309:0.122633:-0.112638;
		specparam thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = -0.0340213:-0.00842307:0.225867;
		specparam tsetup_SIN_XC_SMC_posedge_SMC_negedge = 0.157092:0.120396:-0.114673;
		specparam thold_SIN_XC_SMC_posedge_SMC_negedge = -0.0300146:-0.00729639:0.226227;
		specparam tsetup_SIN_XC_SMC_negedge_SMC_negedge = 0.157092:0.120396:-0.114673;
		specparam thold_SIN_XC_SMC_negedge_SMC_negedge = -0.0300146:-0.00729639:0.226227;
		specparam tsetup_SMC_XC_adacond0_posedge_adacond0_negedge = 0.409177:0.378846:0.0876238;
		specparam thold_SMC_XC_adacond0_posedge_adacond0_negedge = -0.00997581:0.00270369:0.227324;
		specparam tsetup_SMC_XC_adacond0_negedge_adacond0_negedge = 0.409177:0.378846:0.0876238;
		specparam thold_SMC_XC_adacond0_negedge_adacond0_negedge = -0.00997581:0.00270369:0.227324;
		specparam tpw_XC_posedge = 0.223117:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.223117:0.330811:2.72095;

		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_posedge_SMC_negedge, 
			 thold_SIN_XC_SMC_posedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_negedge_SMC_negedge, 
			 thold_SIN_XC_SMC_negedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_posedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_negedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNQ 
`timescale 1ns/10ps
`celldefine
module SDFFNQX4 (Q, D, SIN, SMC, XC);
	output Q;
	input D, SIN, SMC, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_XC_Q_negedge_r = 0.395424:0.559758:2.0059;
		specparam tpd_XC_Q_negedge_f = 0.324439:0.463185:1.35765;
		specparam tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = 0.138312:0.102489:-0.15292;
		specparam thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = -0.0193172:0.00809103:0.256835;
		specparam tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = 0.138312:0.102489:-0.15292;
		specparam thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = -0.0193172:0.00809103:0.256835;
		specparam tsetup_SIN_XC_SMC_posedge_SMC_negedge = 0.135612:0.0989325:-0.155464;
		specparam thold_SIN_XC_SMC_posedge_SMC_negedge = -0.0178311:0.010455:0.257631;
		specparam tsetup_SIN_XC_SMC_negedge_SMC_negedge = 0.135612:0.0989325:-0.155464;
		specparam thold_SIN_XC_SMC_negedge_SMC_negedge = -0.0178311:0.010455:0.257631;
		specparam tsetup_SMC_XC_adacond0_posedge_adacond0_negedge = 0.37779:0.339881:0.0401127;
		specparam thold_SMC_XC_adacond0_posedge_adacond0_negedge = 0.00407935:0.0189965:0.261801;
		specparam tsetup_SMC_XC_adacond0_negedge_adacond0_negedge = 0.37779:0.339881:0.0401127;
		specparam thold_SMC_XC_adacond0_negedge_adacond0_negedge = 0.00407935:0.0189965:0.261801;
		specparam tpw_XC_posedge = 0.205113:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.205113:0.330811:2.72095;

		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_posedge_SMC_negedge, 
			 thold_SIN_XC_SMC_posedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_negedge_SMC_negedge, 
			 thold_SIN_XC_SMC_negedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_posedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_negedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNQ 
`timescale 1ns/10ps
`celldefine
module SDFFNQXL (Q, D, SIN, SMC, XC);
	output Q;
	input D, SIN, SMC, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_XC_Q_negedge_r = 0.380018:0.545634:1.99351;
		specparam tpd_XC_Q_negedge_f = 0.298283:0.454416:1.71501;
		specparam tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = 0.188545:0.147739:-0.096307;
		specparam thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = -0.0295605:-0.00301483:0.233643;
		specparam tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = 0.188545:0.147739:-0.096307;
		specparam thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = -0.0295605:-0.00301483:0.233643;
		specparam tsetup_SIN_XC_SMC_posedge_SMC_negedge = 0.184741:0.145004:-0.0964851;
		specparam thold_SIN_XC_SMC_posedge_SMC_negedge = -0.0301572:-0.0035809:0.2328;
		specparam tsetup_SIN_XC_SMC_negedge_SMC_negedge = 0.184741:0.145004:-0.0964851;
		specparam thold_SIN_XC_SMC_negedge_SMC_negedge = -0.0301572:-0.0035809:0.2328;
		specparam tsetup_SMC_XC_adacond0_posedge_adacond0_negedge = 0.413439:0.379683:0.103611;
		specparam thold_SMC_XC_adacond0_posedge_adacond0_negedge = -0.00612201:0.00639249:0.236611;
		specparam tsetup_SMC_XC_adacond0_negedge_adacond0_negedge = 0.413439:0.379683:0.103611;
		specparam thold_SMC_XC_adacond0_negedge_adacond0_negedge = -0.00612201:0.00639249:0.236611;
		specparam tpw_XC_posedge = 0.225451:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.225451:0.330811:2.72095;

		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_posedge_SMC_negedge, 
			 thold_SIN_XC_SMC_posedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_negedge_SMC_negedge, 
			 thold_SIN_XC_SMC_negedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_posedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_negedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNQX 
`timescale 1ns/10ps
`celldefine
module SDFFNQXX1 (Q, XQ, D, SIN, SMC, XC);
	output Q, XQ;
	input D, SIN, SMC, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_XC_Q_negedge_r = 0.420114:0.590624:2.0335;
		specparam tpd_XC_Q_negedge_f = 0.318528:0.459758:1.36331;
		specparam tpd_XC_XQ_negedge_r = 0.403258:0.554305:1.99798;
		specparam tpd_XC_XQ_negedge_f = 0.481177:0.608746:1.57432;
		specparam tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = 0.181306:0.140973:-0.0998537;
		specparam thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = -0.0318803:-0.00464519:0.231037;
		specparam tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = 0.181306:0.140973:-0.0998537;
		specparam thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = -0.0318803:-0.00464519:0.231037;
		specparam tsetup_SIN_XC_SMC_posedge_SMC_negedge = 0.17752:0.139143:-0.10155;
		specparam thold_SIN_XC_SMC_posedge_SMC_negedge = -0.0294416:-0.00356046:0.235221;
		specparam tsetup_SIN_XC_SMC_negedge_SMC_negedge = 0.17752:0.139143:-0.10155;
		specparam thold_SIN_XC_SMC_negedge_SMC_negedge = -0.0294416:-0.00356046:0.235221;
		specparam tsetup_SMC_XC_adacond0_posedge_adacond0_negedge = 0.408152:0.373383:0.0904478;
		specparam thold_SMC_XC_adacond0_posedge_adacond0_negedge = -0.00789479:0.0061157:0.235523;
		specparam tsetup_SMC_XC_adacond0_negedge_adacond0_negedge = 0.408152:0.373383:0.0904478;
		specparam thold_SMC_XC_adacond0_negedge_adacond0_negedge = -0.00789479:0.0061157:0.235523;
		specparam tpw_XC_posedge = 0.222841:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.222841:0.330811:2.72095;

		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_posedge_SMC_negedge, 
			 thold_SIN_XC_SMC_posedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_negedge_SMC_negedge, 
			 thold_SIN_XC_SMC_negedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_posedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_negedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNQX 
`timescale 1ns/10ps
`celldefine
module SDFFNQXX2 (Q, XQ, D, SIN, SMC, XC);
	output Q, XQ;
	input D, SIN, SMC, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_XC_Q_negedge_r = 0.398494:0.57003:2.01639;
		specparam tpd_XC_Q_negedge_f = 0.336031:0.487082:1.38908;
		specparam tpd_XC_XQ_negedge_r = 0.416753:0.564042:2.01254;
		specparam tpd_XC_XQ_negedge_f = 0.479264:0.603995:1.4944;
		specparam tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = 0.160448:0.12137:-0.115949;
		specparam thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = -0.0346472:-0.00889441:0.226525;
		specparam tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = 0.160448:0.12137:-0.115949;
		specparam thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = -0.0346472:-0.00889441:0.226525;
		specparam tsetup_SIN_XC_SMC_posedge_SMC_negedge = 0.155445:0.119226:-0.11653;
		specparam thold_SIN_XC_SMC_posedge_SMC_negedge = -0.0338525:-0.00489441:0.225727;
		specparam tsetup_SIN_XC_SMC_negedge_SMC_negedge = 0.155445:0.119226:-0.11653;
		specparam thold_SIN_XC_SMC_negedge_SMC_negedge = -0.0338525:-0.00489441:0.225727;
		specparam tsetup_SMC_XC_adacond0_posedge_adacond0_negedge = 0.407062:0.374846:0.0845696;
		specparam thold_SMC_XC_adacond0_posedge_adacond0_negedge = -0.0111611:0.00290174:0.225248;
		specparam tsetup_SMC_XC_adacond0_negedge_adacond0_negedge = 0.407062:0.374846:0.0845696;
		specparam thold_SMC_XC_adacond0_negedge_adacond0_negedge = -0.0111611:0.00290174:0.225248;
		specparam tpw_XC_posedge = 0.220506:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.220506:0.330811:2.72095;

		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_posedge_SMC_negedge, 
			 thold_SIN_XC_SMC_posedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_negedge_SMC_negedge, 
			 thold_SIN_XC_SMC_negedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_posedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_negedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNQX 
`timescale 1ns/10ps
`celldefine
module SDFFNQXX4 (Q, XQ, D, SIN, SMC, XC);
	output Q, XQ;
	input D, SIN, SMC, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_XC_Q_negedge_r = 0.407542:0.574983:2.03226;
		specparam tpd_XC_Q_negedge_f = 0.337061:0.480442:1.38401;
		specparam tpd_XC_XQ_negedge_r = 0.443623:0.591977:2.04093;
		specparam tpd_XC_XQ_negedge_f = 0.529645:0.659111:1.56143;
		specparam tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = 0.137862:0.101979:-0.152163;
		specparam thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = -0.0194248:0.00761044:0.257671;
		specparam tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = 0.137862:0.101979:-0.152163;
		specparam thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = -0.0194248:0.00761044:0.257671;
		specparam tsetup_SIN_XC_SMC_posedge_SMC_negedge = 0.135292:0.0986474:-0.155214;
		specparam thold_SIN_XC_SMC_posedge_SMC_negedge = -0.0172466:0.010826:0.25714;
		specparam tsetup_SIN_XC_SMC_negedge_SMC_negedge = 0.135292:0.0986474:-0.155214;
		specparam thold_SIN_XC_SMC_negedge_SMC_negedge = -0.0172466:0.010826:0.25714;
		specparam tsetup_SMC_XC_adacond0_posedge_adacond0_negedge = 0.374008:0.340326:0.0390933;
		specparam thold_SMC_XC_adacond0_posedge_adacond0_negedge = 0.00216569:0.0195385:0.263093;
		specparam tsetup_SMC_XC_adacond0_negedge_adacond0_negedge = 0.374008:0.340326:0.0390933;
		specparam thold_SMC_XC_adacond0_negedge_adacond0_negedge = 0.00216569:0.0195385:0.263093;
		specparam tpw_XC_posedge = 0.204843:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.204843:0.330811:2.72095;

		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_posedge_SMC_negedge, 
			 thold_SIN_XC_SMC_posedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_negedge_SMC_negedge, 
			 thold_SIN_XC_SMC_negedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_posedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_negedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNQX 
`timescale 1ns/10ps
`celldefine
module SDFFNQXXL (Q, XQ, D, SIN, SMC, XC);
	output Q, XQ;
	input D, SIN, SMC, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	altos_dff_err (xcr_0, int_fwire_clk, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_XC_Q_negedge_r = 0.400083:0.5699:2.01984;
		specparam tpd_XC_Q_negedge_f = 0.316963:0.478451:1.74362;
		specparam tpd_XC_XQ_negedge_r = 0.368012:0.520674:1.96424;
		specparam tpd_XC_XQ_negedge_f = 0.477939:0.627343:1.91326;
		specparam tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = 0.186736:0.147057:-0.0959722;
		specparam thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge = -0.032855:-0.00373139:0.230545;
		specparam tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = 0.186736:0.147057:-0.0959722;
		specparam thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge = -0.032855:-0.00373139:0.230545;
		specparam tsetup_SIN_XC_SMC_posedge_SMC_negedge = 0.180677:0.1436:-0.0988507;
		specparam thold_SIN_XC_SMC_posedge_SMC_negedge = -0.030686:-0.00247381:0.232229;
		specparam tsetup_SIN_XC_SMC_negedge_SMC_negedge = 0.180677:0.1436:-0.0988507;
		specparam thold_SIN_XC_SMC_negedge_SMC_negedge = -0.030686:-0.00247381:0.232229;
		specparam tsetup_SMC_XC_adacond0_posedge_adacond0_negedge = 0.412326:0.378238:0.100394;
		specparam thold_SMC_XC_adacond0_posedge_adacond0_negedge = -0.00732769:0.00592385:0.236115;
		specparam tsetup_SMC_XC_adacond0_negedge_adacond0_negedge = 0.412326:0.378238:0.100394;
		specparam thold_SMC_XC_adacond0_negedge_adacond0_negedge = -0.00732769:0.00592385:0.236115;
		specparam tpw_XC_posedge = 0.225451:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.225451:0.330811:2.72095;

		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_posedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, 
			 thold_D_XC_NTB_SMC_negedge_NTB_SMC_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_posedge_SMC_negedge, 
			 thold_SIN_XC_SMC_posedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_XC_SMC_negedge_SMC_negedge, 
			 thold_SIN_XC_SMC_negedge_SMC_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_posedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_XC_adacond0_negedge_adacond0_negedge, 
			 thold_SMC_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_SMC);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNRQ 
`timescale 1ns/10ps
`celldefine
module SDFFNRQX1 (Q, D, SIN, SMC, XR, XC);
	output Q;
	input D, SIN, SMC, XR, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.117997:0.255151:1.18539;
		specparam tpd_XR_Q_negedge_f = 0.117997:0.255151:1.18539;
		specparam tpd_XC_Q_negedge_r = 0.406857:0.577884:2.09376;
		specparam tpd_XC_Q_negedge_f = 0.333588:0.474466:1.45942;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.117406:0.0729789:-0.241249;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0145518:0.0187614:0.327225;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.117406:0.0729789:-0.241249;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0145518:0.0187614:0.327225;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.11845:0.0786512:-0.214226;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0133343:0.0151287:0.299611;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.11845:0.0786512:-0.214226;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0133343:0.0151287:0.299611;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.387665:0.343235:-0.0466536;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00762769:0.0306112:0.328733;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.387665:0.343235:-0.0466536;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00762769:0.0306112:0.328733;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.280418:-0.34852:-0.584737;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.373364:0.497293:1.26997;
		specparam tpw_XR_negedge = 0.299592:0.396376:2.72095;
		specparam tpw_XC_posedge = 0.212676:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.212676:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNRQ 
`timescale 1ns/10ps
`celldefine
module SDFFNRQX2 (Q, D, SIN, SMC, XR, XC);
	output Q;
	input D, SIN, SMC, XR, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.132545:0.276436:1.20675;
		specparam tpd_XR_Q_negedge_f = 0.132545:0.276436:1.20675;
		specparam tpd_XC_Q_negedge_r = 0.395612:0.567068:2.0063;
		specparam tpd_XC_Q_negedge_f = 0.315784:0.456766:1.33909;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.141487:0.103775:-0.13256;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0374726:-0.00784446:0.229408;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.141487:0.103775:-0.13256;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0374726:-0.00784446:0.229408;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.145848:0.111688:-0.103881;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0374581:-0.0128847:0.198493;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.145848:0.111688:-0.103881;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0374581:-0.0128847:0.198493;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.409:0.374511:0.0656407;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.015538:-0.000387797:0.233924;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.409:0.374511:0.0656407;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.015538:-0.000387797:0.233924;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.251828:-0.310228:-0.389255;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.35322:0.470607:1.17034;
		specparam tpw_XR_negedge = 0.297484:0.396376:2.72095;
		specparam tpw_XC_posedge = 0.236171:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.236171:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNRQ 
`timescale 1ns/10ps
`celldefine
module SDFFNRQX4 (Q, D, SIN, SMC, XR, XC);
	output Q;
	input D, SIN, SMC, XR, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.150486:0.301475:1.28076;
		specparam tpd_XR_Q_negedge_f = 0.150486:0.301475:1.28076;
		specparam tpd_XC_Q_negedge_r = 0.448787:0.623313:2.08167;
		specparam tpd_XC_Q_negedge_f = 0.352598:0.493989:1.37944;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.117893:0.0845049:-0.186623;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0190135:0.00878387:0.276241;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.117893:0.0845049:-0.186623;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0190135:0.00878387:0.276241;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.151188:0.117359:-0.0907684;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0392104:-0.0167149:0.182033;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.151188:0.117359:-0.0907684;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0392104:-0.0167149:0.182033;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.407925:0.367031:0.0272388;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0151376:-0.00118614:0.217747;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.407925:0.367031:0.0272388;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0151376:-0.00118614:0.217747;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.26777:-0.347534:-0.487143;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.341701:0.460769:1.16139;
		specparam tpw_XR_negedge = 0.30786:0.404243:2.72095;
		specparam tpw_XC_posedge = 0.23617:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.23617:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNRQ 
`timescale 1ns/10ps
`celldefine
module SDFFNRQXL (Q, D, SIN, SMC, XR, XC);
	output Q;
	input D, SIN, SMC, XR, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.112835:0.248534:1.2316;
		specparam tpd_XR_Q_negedge_f = 0.112835:0.248534:1.2316;
		specparam tpd_XC_Q_negedge_r = 0.404601:0.573849:2.0958;
		specparam tpd_XC_Q_negedge_f = 0.330221:0.471769:1.53717;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.116513:0.0721333:-0.240769;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0125936:0.0209139:0.326865;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.116513:0.0721333:-0.240769;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0125936:0.0209139:0.326865;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.11597:0.0776653:-0.215333;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.01416:0.016:0.303247;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.11597:0.0776653:-0.215333;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.01416:0.016:0.303247;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.388796:0.344891:-0.0488149;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00928778:0.0318152:0.334716;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.388796:0.344891:-0.0488149;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00928778:0.0318152:0.334716;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.284003:-0.350572:-0.597336;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.375874:0.500357:1.27584;
		specparam tpw_XR_negedge = 0.299393:0.396376:2.72095;
		specparam tpw_XC_posedge = 0.215285:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.215285:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNRQX 
`timescale 1ns/10ps
`celldefine
module SDFFNRQXX1 (Q, XQ, D, SIN, SMC, XR, XC);
	output Q, XQ;
	input D, SIN, SMC, XR, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.120941:0.258836:1.19431;
		specparam tpd_XR_Q_negedge_f = 0.120941:0.258836:1.19431;
		specparam tpd_XC_Q_negedge_r = 0.414531:0.585177:2.1002;
		specparam tpd_XC_Q_negedge_f = 0.339704:0.481039:1.46926;
		specparam tpd_XR_XQ_negedge_r = 0.218156:0.383243:1.81514;
		specparam tpd_XR_XQ_negedge_f = 0.218156:0.383243:1.81514;
		specparam tpd_XC_XQ_negedge_r = 0.411229:0.565962:2.07597;
		specparam tpd_XC_XQ_negedge_f = 0.496938:0.638969:1.7736;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.11707:0.0727988:-0.238426;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0121889:0.018403:0.326036;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.11707:0.0727988:-0.238426;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0121889:0.018403:0.326036;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.116285:0.077595:-0.212966;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0132984:0.0175781:0.297704;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.116285:0.077595:-0.212966;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0132984:0.0175781:0.297704;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.386538:0.343583:-0.0489116;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00858191:0.029344:0.327149;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.386538:0.343583:-0.0489116;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00858191:0.029344:0.327149;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.286388:-0.351017:-0.576392;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.375319:0.497293:1.26723;
		specparam tpw_XR_negedge = 0.299393:0.396376:2.72095;
		specparam tpw_XC_posedge = 0.212675:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.212675:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNRQX 
`timescale 1ns/10ps
`celldefine
module SDFFNRQXX2 (Q, XQ, D, SIN, SMC, XR, XC);
	output Q, XQ;
	input D, SIN, SMC, XR, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.1369:0.281209:1.21913;
		specparam tpd_XR_Q_negedge_f = 0.1369:0.281209:1.21913;
		specparam tpd_XC_Q_negedge_r = 0.405976:0.577207:2.02068;
		specparam tpd_XC_Q_negedge_f = 0.324829:0.466489:1.35331;
		specparam tpd_XR_XQ_negedge_r = 0.262783:0.430197:1.90644;
		specparam tpd_XR_XQ_negedge_f = 0.262783:0.430197:1.90644;
		specparam tpd_XC_XQ_negedge_r = 0.423393:0.574265:2.02126;
		specparam tpd_XC_XQ_negedge_f = 0.522444:0.658946:1.67516;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.141974:0.104874:-0.133317;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0339959:-0.00674935:0.228545;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.141974:0.104874:-0.133317;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0339959:-0.00674935:0.228545;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.14585:0.111773:-0.103451;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0377879:-0.0149708:0.195789;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.14585:0.111773:-0.103451;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0377879:-0.0149708:0.195789;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.408717:0.374155:0.062031;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0143497:0.000702672:0.23143;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.408717:0.374155:0.062031;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0143497:0.000702672:0.23143;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.252904:-0.314492:-0.389193;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.350834:0.468329:1.16862;
		specparam tpw_XR_negedge = 0.299153:0.398998:2.72095;
		specparam tpw_XC_posedge = 0.23617:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.23617:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNRQX 
`timescale 1ns/10ps
`celldefine
module SDFFNRQXX4 (Q, XQ, D, SIN, SMC, XR, XC);
	output Q, XQ;
	input D, SIN, SMC, XR, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.153074:0.303309:1.28525;
		specparam tpd_XR_Q_negedge_f = 0.153074:0.303309:1.28525;
		specparam tpd_XC_Q_negedge_r = 0.460249:0.633075:2.09029;
		specparam tpd_XC_Q_negedge_f = 0.364137:0.505689:1.39312;
		specparam tpd_XR_XQ_negedge_r = 0.274403:0.437365:1.96173;
		specparam tpd_XR_XQ_negedge_f = 0.274403:0.437365:1.96173;
		specparam tpd_XC_XQ_negedge_r = 0.46226:0.612564:2.06528;
		specparam tpd_XC_XQ_negedge_f = 0.568616:0.702572:1.7203;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.117893:0.0845049:-0.185222;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0183008:0.0101609:0.27343;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.117893:0.0845049:-0.185222;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0183008:0.0101609:0.27343;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.150149:0.116501:-0.0880648;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0415802:-0.0180146:0.181237;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.150149:0.116501:-0.0880648;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0415802:-0.0180146:0.181237;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.406192:0.366531:0.0227404;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0164422:-0.00264082:0.217707;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.406192:0.366531:0.0227404;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0164422:-0.00264082:0.217707;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.270364:-0.352674:-0.491779;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.337959:0.458501:1.15778;
		specparam tpw_XR_negedge = 0.309858:0.404243:2.72095;
		specparam tpw_XC_posedge = 0.23617:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.23617:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNRQX 
`timescale 1ns/10ps
`celldefine
module SDFFNRQXXL (Q, XQ, D, SIN, SMC, XR, XC);
	output Q, XQ;
	input D, SIN, SMC, XR, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.115487:0.252567:1.24512;
		specparam tpd_XR_Q_negedge_f = 0.115487:0.252567:1.24512;
		specparam tpd_XC_Q_negedge_r = 0.412285:0.582046:2.1087;
		specparam tpd_XC_Q_negedge_f = 0.335614:0.477963:1.55066;
		specparam tpd_XR_XQ_negedge_r = 0.208901:0.373065:1.80086;
		specparam tpd_XR_XQ_negedge_f = 0.208901:0.373065:1.80086;
		specparam tpd_XC_XQ_negedge_r = 0.402297:0.557962:2.08862;
		specparam tpd_XC_XQ_negedge_f = 0.480073:0.613855:1.66939;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.116277:0.0720983:-0.240641;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0135443:0.0202944:0.329342;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.116277:0.0720983:-0.240641;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0135443:0.0202944:0.329342;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.11615:0.0776181:-0.21551;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0134058:0.0156733:0.30103;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.11615:0.0776181:-0.21551;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0134058:0.0156733:0.30103;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.388793:0.344651:-0.0488731;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00834329:0.0311663:0.333381;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.388793:0.344651:-0.0488731;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00834329:0.0311663:0.333381;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.284574:-0.353344:-0.593567;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.376217:0.500357:1.2731;
		specparam tpw_XR_negedge = 0.299393:0.396376:2.72095;
		specparam tpw_XC_posedge = 0.215285:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.215285:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSQ 
`timescale 1ns/10ps
`celldefine
module SDFFNSQX1 (Q, D, SIN, SMC, XS, XC);
	output Q;
	input D, SIN, SMC, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.283523:0.440581:1.88179;
		specparam tpd_XS_Q_negedge_f = 0.283523:0.440581:1.88179;
		specparam tpd_XC_Q_negedge_r = 0.367405:0.530877:2.04294;
		specparam tpd_XC_Q_negedge_f = 0.342541:0.481865:1.48748;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.128864:0.0860965:-0.239117;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0145555:0.018804:0.326636;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.128864:0.0860965:-0.239117;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0145555:0.018804:0.326636;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.130733:0.0911194:-0.209254;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0136765:0.0153779:0.300362;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.130733:0.0911194:-0.209254;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0136765:0.0153779:0.300362;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.422514:0.374989:0.000433442;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00652012:0.0296277:0.334215;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.422514:0.374989:0.000433442;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00652012:0.0296277:0.334215;
		specparam trecovery_XS_XC_adacond3_posedge_adacond3_negedge = -0.0284091:-0.0809647:-0.340475;
		specparam tremoval_XS_XC_adacond3_posedge_adacond3_negedge = 0.0936737:0.146813:0.511944;
		specparam tpw_XS_negedge = 0.167109:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.243432:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.243432:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XS &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSQ 
`timescale 1ns/10ps
`celldefine
module SDFFNSQX2 (Q, D, SIN, SMC, XS, XC);
	output Q;
	input D, SIN, SMC, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.292207:0.453362:1.8978;
		specparam tpd_XS_Q_negedge_f = 0.292207:0.453362:1.8978;
		specparam tpd_XC_Q_negedge_r = 0.348785:0.51183:1.9598;
		specparam tpd_XC_Q_negedge_f = 0.322173:0.462352:1.37978;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.150328:0.11503:-0.127124;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0386008:-0.0115722:0.228615;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.150328:0.11503:-0.127124;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0386008:-0.0115722:0.228615;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.155463:0.12047:-0.0990417;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0393243:-0.0141972:0.196901;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.155463:0.12047:-0.0990417;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0393243:-0.0141972:0.196901;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.444151:0.403158:0.108949;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0147908:-0.00274728:0.23121;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.444151:0.403158:0.108949;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0147908:-0.00274728:0.23121;
		specparam trecovery_XS_XC_adacond3_posedge_adacond3_negedge = -0.00517927:-0.0483933:-0.202113;
		specparam tremoval_XS_XC_adacond3_posedge_adacond3_negedge = 0.0657853:0.116917:0.401542;
		specparam tpw_XS_negedge = 0.176647:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.272118:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.272118:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XS &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSQ 
`timescale 1ns/10ps
`celldefine
module SDFFNSQX4 (Q, D, SIN, SMC, XS, XC);
	output Q;
	input D, SIN, SMC, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.338118:0.500498:1.96268;
		specparam tpd_XS_Q_negedge_f = 0.338118:0.500498:1.96268;
		specparam tpd_XC_Q_negedge_r = 0.398955:0.564246:2.01758;
		specparam tpd_XC_Q_negedge_f = 0.368592:0.508149:1.39391;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.129796:0.09337:-0.179632;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0208084:0.00764877:0.273976;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.129796:0.09337:-0.179632;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0208084:0.00764877:0.273976;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.13994:0.107186:-0.12714;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0284969:-0.00377366:0.219574;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.13994:0.107186:-0.12714;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0284969:-0.00377366:0.219574;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.450713:0.407221:0.0772966;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.00792889:0.00894586:0.259106;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.450713:0.407221:0.0772966;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.00792889:0.00894586:0.259106;
		specparam trecovery_XS_XC_adacond3_posedge_adacond3_negedge = -0.0120819:-0.0567113:-0.205724;
		specparam tremoval_XS_XC_adacond3_posedge_adacond3_negedge = 0.0657756:0.115209:0.394607;
		specparam tpw_XS_negedge = 0.193243:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.267198:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.267198:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XS &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSQ 
`timescale 1ns/10ps
`celldefine
module SDFFNSQXL (Q, D, SIN, SMC, XS, XC);
	output Q;
	input D, SIN, SMC, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.281461:0.437219:1.88947;
		specparam tpd_XS_Q_negedge_f = 0.281461:0.437219:1.88947;
		specparam tpd_XC_Q_negedge_r = 0.36787:0.530436:2.05547;
		specparam tpd_XC_Q_negedge_f = 0.344449:0.485989:1.57784;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.129062:0.0828979:-0.238213;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0152373:0.0195576:0.327949;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.129062:0.0828979:-0.238213;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0152373:0.0195576:0.327949;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.131512:0.0885733:-0.209134;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0156079:0.0144014:0.301564;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.131512:0.0885733:-0.209134;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0156079:0.0144014:0.301564;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.422325:0.37773:-0.000648077;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00557936:0.0294192:0.3347;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.422325:0.37773:-0.000648077;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00557936:0.0294192:0.3347;
		specparam trecovery_XS_XC_adacond3_posedge_adacond3_negedge = -0.0334553:-0.0807263:-0.353999;
		specparam tremoval_XS_XC_adacond3_posedge_adacond3_negedge = 0.0965598:0.151716:0.521111;
		specparam tpw_XS_negedge = 0.166101:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.248648:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.248648:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XS &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSQX 
`timescale 1ns/10ps
`celldefine
module SDFFNSQXX1 (Q, XQ, D, SIN, SMC, XS, XC);
	output Q, XQ;
	input D, SIN, SMC, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.310975:0.465271:1.90833;
		specparam tpd_XS_Q_negedge_f = 0.310975:0.465271:1.90833;
		specparam tpd_XC_Q_negedge_r = 0.370314:0.532611:2.03385;
		specparam tpd_XC_Q_negedge_f = 0.346129:0.485231:1.48477;
		specparam tpd_XS_XQ_negedge_r = 0.138501:0.296523:1.42415;
		specparam tpd_XS_XQ_negedge_f = 0.138501:0.296523:1.42415;
		specparam tpd_XC_XQ_negedge_r = 0.451147:0.613326:2.13799;
		specparam tpd_XC_XQ_negedge_f = 0.457223:0.603389:1.7496;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.127902:0.0854827:-0.235986;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0133587:0.0191078:0.327416;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.127902:0.0854827:-0.235986;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0133587:0.0191078:0.327416;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.128146:0.086476:-0.208377;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0157148:0.0156457:0.302103;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.128146:0.086476:-0.208377;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0157148:0.0156457:0.302103;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.418204:0.374757:-0.00150111;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.0048931:0.0282678:0.333008;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.418204:0.374757:-0.00150111;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.0048931:0.0282678:0.333008;
		specparam trecovery_XS_XC_adacond3_posedge_adacond3_negedge = -0.0313127:-0.0810126:-0.346363;
		specparam tremoval_XS_XC_adacond3_posedge_adacond3_negedge = 0.0939231:0.148059:0.509469;
		specparam tpw_XS_negedge = 0.195289:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.243432:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.243432:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XS &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSQX 
`timescale 1ns/10ps
`celldefine
module SDFFNSQXX2 (Q, XQ, D, SIN, SMC, XS, XC);
	output Q, XQ;
	input D, SIN, SMC, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.353877:0.512872:1.98541;
		specparam tpd_XS_Q_negedge_f = 0.353877:0.512872:1.98541;
		specparam tpd_XC_Q_negedge_r = 0.355794:0.517779:1.95676;
		specparam tpd_XC_Q_negedge_f = 0.332946:0.473945:1.38793;
		specparam tpd_XS_XQ_negedge_r = 0.150125:0.310889:1.42522;
		specparam tpd_XS_XQ_negedge_f = 0.150125:0.310889:1.42522;
		specparam tpd_XC_XQ_negedge_r = 0.467464:0.628179:2.07196;
		specparam tpd_XC_XQ_negedge_f = 0.471847:0.614531:1.65152;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.151572:0.115249:-0.130462;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0366727:-0.00836982:0.228099;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.151572:0.115249:-0.130462;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0366727:-0.00836982:0.228099;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.152391:0.11965:-0.0998945;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0396984:-0.0143536:0.197873;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.152391:0.11965:-0.0998945;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0396984:-0.0143536:0.197873;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.44348:0.404726:0.102671;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0138611:0.00125029:0.23621;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.44348:0.404726:0.102671;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0138611:0.00125029:0.23621;
		specparam trecovery_XS_XC_adacond3_posedge_adacond3_negedge = -0.00835176:-0.0478806:-0.199963;
		specparam tremoval_XS_XC_adacond3_posedge_adacond3_negedge = 0.0686684:0.115209:0.399478;
		specparam tpw_XS_negedge = 0.230151:0.364904:2.72095;
		specparam tpw_XC_posedge = 0.269808:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.269808:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XS &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSQX 
`timescale 1ns/10ps
`celldefine
module SDFFNSQXX4 (Q, XQ, D, SIN, SMC, XS, XC);
	output Q, XQ;
	input D, SIN, SMC, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.385337:0.547208:2.04263;
		specparam tpd_XS_Q_negedge_f = 0.385337:0.547208:2.04263;
		specparam tpd_XC_Q_negedge_r = 0.404858:0.569202:2.02551;
		specparam tpd_XC_Q_negedge_f = 0.377168:0.516721:1.4029;
		specparam tpd_XS_XQ_negedge_r = 0.143993:0.302387:1.40141;
		specparam tpd_XS_XQ_negedge_f = 0.143993:0.302387:1.40141;
		specparam tpd_XC_XQ_negedge_r = 0.511349:0.669796:2.10975;
		specparam tpd_XC_XQ_negedge_f = 0.510276:0.647404:1.65762;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.129305:0.0899764:-0.184737;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0188175:0.0112882:0.276413;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.129305:0.0899764:-0.184737;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0188175:0.0112882:0.276413;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.160847:0.128473:-0.0841409;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.042864:-0.0182718:0.178366;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.160847:0.128473:-0.0841409;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.042864:-0.0182718:0.178366;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.441604:0.399344:0.0723006;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0167798:-0.0045637:0.216237;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.441604:0.399344:0.0723006;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0167798:-0.0045637:0.216237;
		specparam trecovery_XS_XC_adacond3_posedge_adacond3_negedge = -0.0155788:-0.0568729:-0.204908;
		specparam tremoval_XS_XC_adacond3_posedge_adacond3_negedge = 0.06365:0.111806:0.394012;
		specparam tpw_XS_negedge = 0.245991:0.375395:2.72095;
		specparam tpw_XC_posedge = 0.269512:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.269512:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XS &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSQX 
`timescale 1ns/10ps
`celldefine
module SDFFNSQXXL (Q, XQ, D, SIN, SMC, XS, XC);
	output Q, XQ;
	input D, SIN, SMC, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.296553:0.450771:1.8944;
		specparam tpd_XS_Q_negedge_f = 0.296553:0.450771:1.8944;
		specparam tpd_XC_Q_negedge_r = 0.368853:0.531207:2.05096;
		specparam tpd_XC_Q_negedge_f = 0.348305:0.491367:1.59808;
		specparam tpd_XS_XQ_negedge_r = 0.132855:0.277929:1.29801;
		specparam tpd_XS_XQ_negedge_f = 0.132855:0.277929:1.29801;
		specparam tpd_XC_XQ_negedge_r = 0.449135:0.6085:2.13091;
		specparam tpd_XC_XQ_negedge_f = 0.444875:0.581296:1.6408;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.128945:0.0828525:-0.238127;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.014253:0.0183067:0.330975;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.128945:0.0828525:-0.238127;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.014253:0.0183067:0.330975;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.131224:0.0886027:-0.209047;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0168116:0.0132913:0.301548;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.131224:0.0886027:-0.209047;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0168116:0.0132913:0.301548;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.421911:0.377631:-0.000808775;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00665724:0.0291639:0.336646;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.421911:0.377631:-0.000808775;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00665724:0.0291639:0.336646;
		specparam trecovery_XS_XC_adacond3_posedge_adacond3_negedge = -0.0335087:-0.0849473:-0.353769;
		specparam tremoval_XS_XC_adacond3_posedge_adacond3_negedge = 0.0965598:0.151716:0.521111;
		specparam tpw_XS_negedge = 0.181784:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.248648:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.248648:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$recovery (posedge XS &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_XC_adacond3_posedge_adacond3_negedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSRQ 
`timescale 1ns/10ps
`celldefine
module SDFFNSRQX1 (Q, D, SIN, SMC, XR, XS, XC);
	output Q;
	input D, SIN, SMC, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.12662:0.253098:1.44589;
		specparam tpd_XR_Q_negedge_f = 0.119076:0.256301:1.19483;
		specparam tpd_XS_Q_negedge_r = 0.327456:0.492203:1.95435;
		specparam tpd_XS_Q_negedge_f = 0.327456:0.492203:1.95435;
		specparam tpd_XC_Q_negedge_r = 0.409356:0.581057:2.10184;
		specparam tpd_XC_Q_negedge_f = 0.351386:0.491105:1.48795;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.132236:0.0924068:-0.229457;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0144046:0.0199125:0.326195;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.132236:0.0924068:-0.229457;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0144046:0.0199125:0.326195;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.136665:0.0955038:-0.19942;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0180761:0.0142104:0.300157;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.136665:0.0955038:-0.19942;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0180761:0.0142104:0.300157;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.427115:0.382247:0.00397949;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00585711:0.0293909:0.328615;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.427115:0.382247:0.00397949;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00585711:0.0293909:0.328615;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.283526:-0.346554:-0.574583;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.405558:0.521782:1.29765;
		specparam tpw_XR_negedge = 0.335512:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.01944:0.00665868:0.00388529;
		specparam thold_XR_XS_posedge_posedge = 0.0400071:0.0576497:0.121024;
		specparam trecovery_XS_XC_adacond4_posedge_adacond4_negedge = -0.02542:-0.0750097:-0.341269;
		specparam tremoval_XS_XC_adacond4_posedge_adacond4_negedge = 0.106855:0.162217:0.534389;
		specparam tsetup_XS_XR_posedge_posedge = 0.0421581:0.0652049:0.191592;
		specparam thold_XS_XR_posedge_posedge = 0.0511317:0.0596125:0.043357;
		specparam tpw_XS_negedge = 0.191304:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.25908:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.25908:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$recovery (posedge XS &&& adacond4, negedge XC &&& adacond4, 
			 trecovery_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$hold (negedge XC &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSRQ 
`timescale 1ns/10ps
`celldefine
module SDFFNSRQX2 (Q, D, SIN, SMC, XR, XS, XC);
	output Q;
	input D, SIN, SMC, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.141716:0.276512:1.48874;
		specparam tpd_XR_Q_negedge_f = 0.133991:0.278857:1.22837;
		specparam tpd_XS_Q_negedge_r = 0.34545:0.515881:1.97299;
		specparam tpd_XS_Q_negedge_f = 0.34545:0.515881:1.97299;
		specparam tpd_XC_Q_negedge_r = 0.399271:0.571899:2.01956;
		specparam tpd_XC_Q_negedge_f = 0.335219:0.476913:1.37977;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.159023:0.119351:-0.119696;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0370873:-0.0111365:0.224263;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.159023:0.119351:-0.119696;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0370873:-0.0111365:0.224263;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.161498:0.126961:-0.0885788;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.040917:-0.0162706:0.195661;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.161498:0.126961:-0.0885788;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.040917:-0.0162706:0.195661;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.45196:0.413019:0.112551;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0188482:-0.00305833:0.231363;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.45196:0.413019:0.112551;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0188482:-0.00305833:0.231363;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.253404:-0.308858:-0.383388;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.381662:0.491827:1.20016;
		specparam tpw_XR_negedge = 0.333348:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.019024:0.00878685:0.0442402;
		specparam thold_XR_XS_posedge_posedge = 0.0269967:0.0359833:0.111576;
		specparam trecovery_XS_XC_adacond4_posedge_adacond4_negedge = -0.00300762:-0.0467969:-0.200579;
		specparam tremoval_XS_XC_adacond4_posedge_adacond4_negedge = 0.0800179:0.132922:0.424917;
		specparam tsetup_XS_XR_posedge_posedge = 0.0320321:0.0508196:0.18946;
		specparam thold_XS_XR_posedge_posedge = 0.0496903:0.0582862:0.0780376;
		specparam tpw_XS_negedge = 0.201205:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.282854:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.282854:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$recovery (posedge XS &&& adacond4, negedge XC &&& adacond4, 
			 trecovery_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$hold (negedge XC &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSRQ 
`timescale 1ns/10ps
`celldefine
module SDFFNSRQX4 (Q, D, SIN, SMC, XR, XS, XC);
	output Q;
	input D, SIN, SMC, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.143141:0.274543:1.43997;
		specparam tpd_XR_Q_negedge_f = 0.152143:0.301194:1.27869;
		specparam tpd_XS_Q_negedge_r = 0.391527:0.56145:2.0257;
		specparam tpd_XS_Q_negedge_f = 0.391527:0.56145:2.0257;
		specparam tpd_XC_Q_negedge_r = 0.44942:0.622527:2.06391;
		specparam tpd_XC_Q_negedge_f = 0.378541:0.51902:1.39782;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.13515:0.0970655:-0.173158;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0206351:0.00664156:0.272076;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.13515:0.0970655:-0.173158;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0206351:0.00664156:0.272076;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.149019:0.115105:-0.115905;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0323121:-0.00790384:0.216813;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.149019:0.115105:-0.115905;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0323121:-0.00790384:0.216813;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.455301:0.413471:0.0796783;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.00942158:0.00843849:0.258311;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.455301:0.413471:0.0796783;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.00942158:0.00843849:0.258311;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.272538:-0.347645:-0.489248;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.365769:0.480048:1.18746;
		specparam tpw_XR_negedge = 0.347218:0.433092:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0189482:0.0111938:0.0777004;
		specparam thold_XR_XS_posedge_posedge = 0.033421:0.0444951:0.137237;
		specparam trecovery_XS_XC_adacond4_posedge_adacond4_negedge = -0.0127272:-0.0559579:-0.20509;
		specparam tremoval_XS_XC_adacond4_posedge_adacond4_negedge = 0.0765305:0.129129:0.415254;
		specparam tsetup_XS_XR_posedge_posedge = 0.0175243:0.0224105:0.175708;
		specparam thold_XS_XR_posedge_posedge = 0.0531305:0.0622621:0.1056;
		specparam tpw_XS_negedge = 0.22326:0.354414:2.72095;
		specparam tpw_XC_posedge = 0.280245:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.280245:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$recovery (posedge XS &&& adacond4, negedge XC &&& adacond4, 
			 trecovery_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$hold (negedge XC &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSRQ 
`timescale 1ns/10ps
`celldefine
module SDFFNSRQXL (Q, D, SIN, SMC, XR, XS, XC);
	output Q;
	input D, SIN, SMC, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.123995:0.245389:1.41267;
		specparam tpd_XR_Q_negedge_f = 0.113869:0.248362:1.22471;
		specparam tpd_XS_Q_negedge_r = 0.322064:0.482533:1.91813;
		specparam tpd_XS_Q_negedge_f = 0.322064:0.482533:1.91813;
		specparam tpd_XC_Q_negedge_r = 0.406799:0.574426:2.07269;
		specparam tpd_XC_Q_negedge_f = 0.346879:0.486346:1.54893;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.130986:0.0885722:-0.233516;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0141435:0.0184703:0.332157;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.130986:0.0885722:-0.233516;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0141435:0.0184703:0.332157;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.164779:0.123438:-0.141225;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0356987:-0.00710232:0.246358;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.164779:0.123438:-0.141225;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0356987:-0.00710232:0.246358;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.424237:0.376503:-0.00571453;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0106495:0.00744825:0.271004;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.424237:0.376503:-0.00571453;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0106495:0.00744825:0.271004;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.284561:-0.347778:-0.591457;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.407912:0.524661:1.30486;
		specparam tpw_XR_negedge = 0.337323:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.017734:0.00874101:-0.00455945;
		specparam thold_XR_XS_posedge_posedge = 0.045951:0.0641407:0.126937;
		specparam trecovery_XS_XC_adacond4_posedge_adacond4_negedge = -0.0272195:-0.0764539:-0.349111;
		specparam tremoval_XS_XC_adacond4_posedge_adacond4_negedge = 0.11028:0.16607:0.538979;
		specparam tsetup_XS_XR_posedge_posedge = 0.0448832:0.0713222:0.188338;
		specparam thold_XS_XR_posedge_posedge = 0.0533898:0.0613222:0.0424261;
		specparam tpw_XS_negedge = 0.189454:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.259371:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.259371:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$recovery (posedge XS &&& adacond4, negedge XC &&& adacond4, 
			 trecovery_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$hold (negedge XC &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSRQX 
`timescale 1ns/10ps
`celldefine
module SDFFNSRQXX1 (Q, XQ, D, SIN, SMC, XR, XS, XC);
	output Q, XQ;
	input D, SIN, SMC, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_r, int_fwire_s;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.128148:0.254319:1.4381;
		specparam tpd_XR_Q_negedge_f = 0.120685:0.257699:1.19371;
		specparam tpd_XS_Q_negedge_r = 0.355226:0.517997:1.9766;
		specparam tpd_XS_Q_negedge_f = 0.355226:0.517997:1.9766;
		specparam tpd_XC_Q_negedge_r = 0.41441:0.585071:2.0985;
		specparam tpd_XC_Q_negedge_f = 0.358937:0.499309:1.49301;
		specparam tpd_XR_XQ_negedge_r = 0.268615:0.448376:1.89503;
		specparam tpd_XR_XQ_negedge_f = 0.268615:0.448376:1.89503;
		specparam tpd_XS_XQ_negedge_r = 0.1442:0.29599:1.55247;
		specparam tpd_XS_XQ_negedge_f = 0.139531:0.295811:1.43388;
		specparam tpd_XC_XQ_negedge_r = 0.468508:0.629297:2.14962;
		specparam tpd_XC_XQ_negedge_f = 0.509137:0.654323:1.78987;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.131932:0.0924397:-0.229577;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0142598:0.0201479:0.327175;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.131932:0.0924397:-0.229577;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0142598:0.0201479:0.327175;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.136925:0.0946691:-0.198639;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0153304:0.0153013:0.298682;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.136925:0.0946691:-0.198639;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0153304:0.0153013:0.298682;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.428451:0.38199:0.0040618;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00603443:0.0269141:0.331246;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.428451:0.38199:0.0040618;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00603443:0.0269141:0.331246;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.284975:-0.349612:-0.57663;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.403428:0.521782:1.29765;
		specparam tpw_XR_negedge = 0.337541:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0157636:0.00606375:0.0039804;
		specparam thold_XR_XS_posedge_posedge = 0.0545913:0.0745493:0.134709;
		specparam trecovery_XS_XC_adacond4_posedge_adacond4_negedge = -0.0285263:-0.0768878:-0.339789;
		specparam tremoval_XS_XC_adacond4_posedge_adacond4_negedge = 0.106818:0.163053:0.533399;
		specparam tsetup_XS_XR_posedge_posedge = 0.0544632:0.0849135:0.229108;
		specparam thold_XS_XR_posedge_posedge = 0.0157636:0.00606375:-0.0677645;
		specparam tpw_XS_negedge = 0.217642:0.341301:2.72095;
		specparam tpw_XC_posedge = 0.256761:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.256761:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$recovery (posedge XS &&& adacond4, negedge XC &&& adacond4, 
			 trecovery_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$hold (negedge XC &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSRQX 
`timescale 1ns/10ps
`celldefine
module SDFFNSRQXX2 (Q, XQ, D, SIN, SMC, XR, XS, XC);
	output Q, XQ;
	input D, SIN, SMC, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_r, int_fwire_s;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.144446:0.279463:1.48709;
		specparam tpd_XR_Q_negedge_f = 0.137134:0.281935:1.23275;
		specparam tpd_XS_Q_negedge_r = 0.409322:0.578416:2.06365;
		specparam tpd_XS_Q_negedge_f = 0.409322:0.578416:2.06365;
		specparam tpd_XC_Q_negedge_r = 0.407945:0.579866:2.02468;
		specparam tpd_XC_Q_negedge_f = 0.347506:0.490268:1.3937;
		specparam tpd_XR_XQ_negedge_r = 0.318628:0.502957:1.98849;
		specparam tpd_XR_XQ_negedge_f = 0.318628:0.502957:1.98849;
		specparam tpd_XS_XQ_negedge_r = 0.15774:0.315245:1.59565;
		specparam tpd_XS_XQ_negedge_f = 0.1534:0.313995:1.44714;
		specparam tpd_XC_XQ_negedge_r = 0.488328:0.649668:2.09845;
		specparam tpd_XC_XQ_negedge_f = 0.536976:0.677936:1.71117;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.157044:0.118147:-0.1242;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0373464:-0.0113283:0.227131;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.157044:0.118147:-0.1242;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0373464:-0.0113283:0.227131;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.157914:0.125944:-0.0883839;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0397872:-0.0156094:0.198148;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.157914:0.125944:-0.0883839;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0397872:-0.0156094:0.198148;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.449:0.411551:0.110585;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0161198:-0.00255007:0.233614;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.449:0.411551:0.110585;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0161198:-0.00255007:0.233614;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.256942:-0.313437:-0.386394;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.380263:0.492311:1.19668;
		specparam tpw_XR_negedge = 0.335166:0.427847:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0177213:0.00698327:0.0225248;
		specparam thold_XR_XS_posedge_posedge = 0.056425:0.0721995:0.122699;
		specparam trecovery_XS_XC_adacond4_posedge_adacond4_negedge = -0.00501365:-0.0491844:-0.202131;
		specparam tremoval_XS_XC_adacond4_posedge_adacond4_negedge = 0.0785456:0.129129:0.425768;
		specparam tsetup_XS_XR_posedge_posedge = 0.0592663:0.0891861:0.233421;
		specparam thold_XS_XR_posedge_posedge = 0.0177321:0.00698327:-0.0575309;
		specparam tpw_XS_negedge = 0.259298:0.383263:2.72095;
		specparam tpw_XC_posedge = 0.282551:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.282551:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$recovery (posedge XS &&& adacond4, negedge XC &&& adacond4, 
			 trecovery_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$hold (negedge XC &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSRQX 
`timescale 1ns/10ps
`celldefine
module SDFFNSRQXX4 (Q, XQ, D, SIN, SMC, XR, XS, XC);
	output Q, XQ;
	input D, SIN, SMC, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_r, int_fwire_s;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.144521:0.276077:1.43793;
		specparam tpd_XR_Q_negedge_f = 0.151989:0.300354:1.27389;
		specparam tpd_XS_Q_negedge_r = 0.436524:0.605437:2.086;
		specparam tpd_XS_Q_negedge_f = 0.436524:0.605437:2.086;
		specparam tpd_XC_Q_negedge_r = 0.460302:0.631893:2.0713;
		specparam tpd_XC_Q_negedge_f = 0.390954:0.531784:1.41122;
		specparam tpd_XR_XQ_negedge_r = 0.321477:0.497664:2.019;
		specparam tpd_XR_XQ_negedge_f = 0.321477:0.497664:2.019;
		specparam tpd_XS_XQ_negedge_r = 0.137683:0.283956:1.51173;
		specparam tpd_XS_XQ_negedge_f = 0.145169:0.302954:1.41786;
		specparam tpd_XC_XQ_negedge_r = 0.529479:0.68821:2.12986;
		specparam tpd_XC_XQ_negedge_f = 0.577442:0.713617:1.72958;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.134392:0.0951895:-0.176749;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0224246:0.00828647:0.273429;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.134392:0.0951895:-0.176749;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0224246:0.00828647:0.273429;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.166835:0.132059:-0.0747949;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0454076:-0.0197388:0.176738;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.166835:0.132059:-0.0747949;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0454076:-0.0197388:0.176738;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.448373:0.404305:0.0745707;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = -0.0191333:-0.00418132:0.213966;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.448373:0.404305:0.0745707;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = -0.0191333:-0.00418132:0.213966;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.27349:-0.353485:-0.489653;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.363904:0.480048:1.18554;
		specparam tpw_XR_negedge = 0.351379:0.435715:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0160341:0.00553392:0.0268162;
		specparam thold_XR_XS_posedge_posedge = 0.0546232:0.0689859:0.144192;
		specparam trecovery_XS_XC_adacond4_posedge_adacond4_negedge = -0.0128899:-0.0584187:-0.203772;
		specparam tremoval_XS_XC_adacond4_posedge_adacond4_negedge = 0.0763266:0.125335:0.412308;
		specparam tsetup_XS_XR_posedge_posedge = 0.0525706:0.0720198:0.224424;
		specparam thold_XS_XR_posedge_posedge = 0.0192698:0.00617576:-0.0760674;
		specparam tpw_XS_negedge = 0.276401:0.39113:2.72095;
		specparam tpw_XC_posedge = 0.280245:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.280245:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$recovery (posedge XS &&& adacond4, negedge XC &&& adacond4, 
			 trecovery_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$hold (negedge XC &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFNSRQX 
`timescale 1ns/10ps
`celldefine
module SDFFNSRQXXL (Q, XQ, D, SIN, SMC, XR, XS, XC);
	output Q, XQ;
	input D, SIN, SMC, XR, XS, XC;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_XC;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_clk, int_fwire_d, int_fwire_IQ;
	wire int_fwire_IXQ, int_fwire_r, int_fwire_s;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_clk, delayed_XC);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, int_fwire_clk, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.124738:0.247918:1.42892;
		specparam tpd_XR_Q_negedge_f = 0.115084:0.250448:1.23506;
		specparam tpd_XS_Q_negedge_r = 0.340472:0.50081:1.94663;
		specparam tpd_XS_Q_negedge_f = 0.340472:0.50081:1.94663;
		specparam tpd_XC_Q_negedge_r = 0.411231:0.579578:2.09192;
		specparam tpd_XC_Q_negedge_f = 0.353454:0.494301:1.56428;
		specparam tpd_XR_XQ_negedge_r = 0.259895:0.436779:1.87547;
		specparam tpd_XR_XQ_negedge_f = 0.259895:0.436779:1.87547;
		specparam tpd_XS_XQ_negedge_r = 0.152525:0.302018:1.57295;
		specparam tpd_XS_XQ_negedge_f = 0.13528:0.280215:1.32557;
		specparam tpd_XC_XQ_negedge_r = 0.457482:0.617126:2.15497;
		specparam tpd_XC_XQ_negedge_f = 0.491792:0.628938:1.68958;
		specparam tsetup_D_XC_adacond0_posedge_adacond0_negedge = 0.131224:0.0919969:-0.228581;
		specparam thold_D_XC_adacond0_posedge_adacond0_negedge = -0.0136954:0.0171797:0.326156;
		specparam tsetup_D_XC_adacond0_negedge_adacond0_negedge = 0.131224:0.0919969:-0.228581;
		specparam thold_D_XC_adacond0_negedge_adacond0_negedge = -0.0136954:0.0171797:0.326156;
		specparam tsetup_SIN_XC_adacond1_posedge_adacond1_negedge = 0.135245:0.093912:-0.204281;
		specparam thold_SIN_XC_adacond1_posedge_adacond1_negedge = -0.0177513:0.0123699:0.3002;
		specparam tsetup_SIN_XC_adacond1_negedge_adacond1_negedge = 0.135245:0.093912:-0.204281;
		specparam thold_SIN_XC_adacond1_negedge_adacond1_negedge = -0.0177513:0.0123699:0.3002;
		specparam tsetup_SMC_XC_adacond2_posedge_adacond2_negedge = 0.430316:0.382936:0.00121587;
		specparam thold_SMC_XC_adacond2_posedge_adacond2_negedge = 0.00490599:0.0274222:0.33493;
		specparam tsetup_SMC_XC_adacond2_negedge_adacond2_negedge = 0.430316:0.382936:0.00121587;
		specparam thold_SMC_XC_adacond2_negedge_adacond2_negedge = 0.00490599:0.0274222:0.33493;
		specparam trecovery_XR_XC_adacond3_posedge_adacond3_negedge = -0.287416:-0.350188:-0.593326;
		specparam tremoval_XR_XC_adacond3_posedge_adacond3_negedge = 0.406309:0.522266:1.30326;
		specparam tpw_XR_negedge = 0.339738:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.018753:0.00732426:-0.005393;
		specparam thold_XR_XS_posedge_posedge = 0.052432:0.0746485:0.138555;
		specparam trecovery_XS_XC_adacond4_posedge_adacond4_negedge = -0.0274509:-0.0779958:-0.34741;
		specparam tremoval_XS_XC_adacond4_posedge_adacond4_negedge = 0.106919:0.16607:0.538979;
		specparam tsetup_XS_XR_posedge_posedge = 0.0561484:0.0872597:0.219652;
		specparam thold_XS_XR_posedge_posedge = 0.018753:0.00732426:-0.0750148;
		specparam tpw_XS_negedge = 0.201974:0.330811:2.72095;
		specparam tpw_XC_posedge = 0.25908:0.330811:2.72095;
		specparam tpw_XC_negedge = 0.25908:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(negedge XC => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_Q_negedge_r , tpd_XC_Q_negedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(negedge XC => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_XC_XQ_negedge_r , tpd_XC_XQ_negedge_f );
		$setuphold (negedge XC &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_posedge_adacond0_negedge, 
			 thold_D_XC_adacond0_posedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_XC_adacond0_negedge_adacond0_negedge, 
			 thold_D_XC_adacond0_negedge_adacond0_negedge, notifier,,, delayed_XC, delayed_D);
		$setuphold (negedge XC &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_posedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_posedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_XC_adacond1_negedge_adacond1_negedge, 
			 thold_SIN_XC_adacond1_negedge_adacond1_negedge, notifier,,, delayed_XC, delayed_SIN);
		$setuphold (negedge XC &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_posedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_posedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (negedge XC &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_XC_adacond2_negedge_adacond2_negedge, 
			 thold_SMC_XC_adacond2_negedge_adacond2_negedge, notifier,,, delayed_XC, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, negedge XC &&& adacond3, 
			 trecovery_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$hold (negedge XC &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_XC_adacond3_posedge_adacond3_negedge, notifier);
		$recovery (posedge XS &&& adacond4, negedge XC &&& adacond4, 
			 trecovery_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$hold (negedge XC &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_XC_adacond4_posedge_adacond4_negedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge XC, tpw_XC_posedge, 0, notifier);
		$width (negedge XC, tpw_XC_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFQ 
`timescale 1ns/10ps
`celldefine
module SDFFQX1 (Q, D, SIN, SMC, C);
	output Q;
	input D, SIN, SMC, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	wire int_fwire_s =0;
	wire int_fwire_r =0;
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_C_Q_posedge_r = 0.357492:0.498602:1.64933;
		specparam tpd_C_Q_posedge_f = 0.31046:0.424252:1.03023;
		specparam tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge = 0.233727:0.22964:0.383949;
		specparam thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge = -0.135253:-0.165056:-0.332526;
		specparam tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge = 0.233727:0.22964:0.383949;
		specparam thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge = -0.135253:-0.165056:-0.332526;
		specparam tsetup_SIN_C_SMC_posedge_SMC_posedge = 0.232412:0.227466:0.384098;
		specparam thold_SIN_C_SMC_posedge_SMC_posedge = -0.134975:-0.16483:-0.330662;
		specparam tsetup_SIN_C_SMC_negedge_SMC_posedge = 0.232412:0.227466:0.384098;
		specparam thold_SIN_C_SMC_negedge_SMC_posedge = -0.134975:-0.16483:-0.330662;
		specparam tsetup_SMC_C_adacond0_posedge_adacond0_posedge = 0.368261:0.35721:0.390765;
		specparam thold_SMC_C_adacond0_posedge_adacond0_posedge = -0.113669:-0.154255:-0.246464;
		specparam tsetup_SMC_C_adacond0_negedge_adacond0_posedge = 0.368261:0.35721:0.390765;
		specparam thold_SMC_C_adacond0_negedge_adacond0_posedge = -0.113669:-0.154255:-0.246464;
		specparam tpw_C_posedge = 0.210936:0.330811:2.72095;
		specparam tpw_C_negedge = 0.210936:0.330811:2.72095;

		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_posedge_SMC_posedge, 
			 thold_SIN_C_SMC_posedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_negedge_SMC_posedge, 
			 thold_SIN_C_SMC_negedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_posedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_negedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFQ 
`timescale 1ns/10ps
`celldefine
module SDFFQX2 (Q, D, SIN, SMC, C);
	output Q;
	input D, SIN, SMC, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	wire int_fwire_s =0;
	wire int_fwire_r =0;
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_C_Q_posedge_r = 0.342188:0.48529:1.64383;
		specparam tpd_C_Q_posedge_f = 0.323971:0.444691:1.04645;
		specparam tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge = 0.218611:0.21998:0.38263;
		specparam thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge = -0.139086:-0.170828:-0.337346;
		specparam tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge = 0.218611:0.21998:0.38263;
		specparam thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge = -0.139086:-0.170828:-0.337346;
		specparam tsetup_SIN_C_SMC_posedge_SMC_posedge = 0.214604:0.218304:0.385259;
		specparam thold_SIN_C_SMC_posedge_SMC_posedge = -0.138229:-0.168828:-0.337633;
		specparam tsetup_SIN_C_SMC_negedge_SMC_posedge = 0.214604:0.218304:0.385259;
		specparam thold_SIN_C_SMC_negedge_SMC_posedge = -0.138229:-0.168828:-0.337633;
		specparam tsetup_SMC_C_adacond0_posedge_adacond0_posedge = 0.365521:0.356605:0.39185;
		specparam thold_SMC_C_adacond0_posedge_adacond0_posedge = -0.118365:-0.160345:-0.252249;
		specparam tsetup_SMC_C_adacond0_negedge_adacond0_posedge = 0.365521:0.356605:0.39185;
		specparam thold_SMC_C_adacond0_negedge_adacond0_posedge = -0.118365:-0.160345:-0.252249;
		specparam tpw_C_posedge = 0.200157:0.330811:2.72095;
		specparam tpw_C_negedge = 0.200157:0.330811:2.72095;

		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_posedge_SMC_posedge, 
			 thold_SIN_C_SMC_posedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_negedge_SMC_posedge, 
			 thold_SIN_C_SMC_negedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_posedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_negedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFQ 
`timescale 1ns/10ps
`celldefine
module SDFFQX4 (Q, D, SIN, SMC, C);
	output Q;
	input D, SIN, SMC, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	wire int_fwire_s =0;
	wire int_fwire_r =0;
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_C_Q_posedge_r = 0.369057:0.509079:1.64543;
		specparam tpd_C_Q_posedge_f = 0.33146:0.447367:1.03714;
		specparam tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge = 0.189272:0.194827:0.343955;
		specparam thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge = -0.125529:-0.153317:-0.303083;
		specparam tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge = 0.189272:0.194827:0.343955;
		specparam thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge = -0.125529:-0.153317:-0.303083;
		specparam tsetup_SIN_C_SMC_posedge_SMC_posedge = 0.185239:0.193358:0.342935;
		specparam thold_SIN_C_SMC_posedge_SMC_posedge = -0.121601:-0.151382:-0.299058;
		specparam tsetup_SIN_C_SMC_negedge_SMC_posedge = 0.185239:0.193358:0.342935;
		specparam thold_SIN_C_SMC_negedge_SMC_posedge = -0.121601:-0.151382:-0.299058;
		specparam tsetup_SMC_C_adacond0_posedge_adacond0_posedge = 0.331953:0.319279:0.345445;
		specparam thold_SMC_C_adacond0_posedge_adacond0_posedge = -0.100333:-0.141782:-0.216396;
		specparam tsetup_SMC_C_adacond0_negedge_adacond0_posedge = 0.331953:0.319279:0.345445;
		specparam thold_SMC_C_adacond0_negedge_adacond0_posedge = -0.100333:-0.141782:-0.216396;
		specparam tpw_C_posedge = 0.231514:0.330811:2.72095;
		specparam tpw_C_negedge = 0.231514:0.330811:2.72095;

		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_posedge_SMC_posedge, 
			 thold_SIN_C_SMC_posedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_negedge_SMC_posedge, 
			 thold_SIN_C_SMC_negedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_posedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_negedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFQ 
`timescale 1ns/10ps
`celldefine
module SDFFQXL (Q, D, SIN, SMC, C);
	output Q;
	input D, SIN, SMC, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	wire int_fwire_s =0;
	wire int_fwire_r =0;
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_C_Q_posedge_r = 0.340197:0.481196:1.63508;
		specparam tpd_C_Q_posedge_f = 0.310155:0.443994:1.41182;
		specparam tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge = 0.242185:0.233177:0.387842;
		specparam thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge = -0.135251:-0.167368:-0.332307;
		specparam tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge = 0.242185:0.233177:0.387842;
		specparam thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge = -0.135251:-0.167368:-0.332307;
		specparam tsetup_SIN_C_SMC_posedge_SMC_posedge = 0.23863:0.231902:0.388647;
		specparam thold_SIN_C_SMC_posedge_SMC_posedge = -0.134121:-0.164144:-0.330533;
		specparam tsetup_SIN_C_SMC_negedge_SMC_posedge = 0.23863:0.231902:0.388647;
		specparam thold_SIN_C_SMC_negedge_SMC_posedge = -0.134121:-0.164144:-0.330533;
		specparam tsetup_SMC_C_adacond0_posedge_adacond0_posedge = 0.369619:0.359091:0.394638;
		specparam thold_SMC_C_adacond0_posedge_adacond0_posedge = -0.112757:-0.156069:-0.253989;
		specparam tsetup_SMC_C_adacond0_negedge_adacond0_posedge = 0.369619:0.359091:0.394638;
		specparam thold_SMC_C_adacond0_negedge_adacond0_posedge = -0.112757:-0.156069:-0.253989;
		specparam tpw_C_posedge = 0.200157:0.330811:2.72095;
		specparam tpw_C_negedge = 0.200157:0.330811:2.72095;

		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_posedge_SMC_posedge, 
			 thold_SIN_C_SMC_posedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_negedge_SMC_posedge, 
			 thold_SIN_C_SMC_negedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_posedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_negedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFQX 
`timescale 1ns/10ps
`celldefine
module SDFFQXX1 (Q, XQ, D, SIN, SMC, C);
	output Q, XQ;
	input D, SIN, SMC, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	altos_dff_err (xcr_0, delayed_C, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, delayed_C, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_C_Q_posedge_r = 0.380013:0.525565:1.66857;
		specparam tpd_C_Q_posedge_f = 0.330868:0.450031:1.05716;
		specparam tpd_C_XQ_posedge_r = 0.416994:0.54472:1.67784;
		specparam tpd_C_XQ_posedge_f = 0.439208:0.538409:1.13867;
		specparam tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge = 0.231561:0.22764:0.384919;
		specparam thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge = -0.137829:-0.165423:-0.332247;
		specparam tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge = 0.231561:0.22764:0.384919;
		specparam thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge = -0.137829:-0.165423:-0.332247;
		specparam tsetup_SIN_C_SMC_posedge_SMC_posedge = 0.226441:0.225047:0.384018;
		specparam thold_SIN_C_SMC_posedge_SMC_posedge = -0.13199:-0.164295:-0.331281;
		specparam tsetup_SIN_C_SMC_negedge_SMC_posedge = 0.226441:0.225047:0.384018;
		specparam thold_SIN_C_SMC_negedge_SMC_posedge = -0.13199:-0.164295:-0.331281;
		specparam tsetup_SMC_C_adacond0_posedge_adacond0_posedge = 0.366513:0.35655:0.3895;
		specparam thold_SMC_C_adacond0_posedge_adacond0_posedge = -0.113574:-0.153161:-0.25073;
		specparam tsetup_SMC_C_adacond0_negedge_adacond0_posedge = 0.366513:0.35655:0.3895;
		specparam thold_SMC_C_adacond0_negedge_adacond0_posedge = -0.113574:-0.153161:-0.25073;
		specparam tpw_C_posedge = 0.223675:0.330811:2.72095;
		specparam tpw_C_negedge = 0.223675:0.330811:2.72095;

		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_posedge_SMC_posedge, 
			 thold_SIN_C_SMC_posedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_negedge_SMC_posedge, 
			 thold_SIN_C_SMC_negedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_posedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_negedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFQX 
`timescale 1ns/10ps
`celldefine
module SDFFQXX2 (Q, XQ, D, SIN, SMC, C);
	output Q, XQ;
	input D, SIN, SMC, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	altos_dff_err (xcr_0, delayed_C, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, delayed_C, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_C_Q_posedge_r = 0.363571:0.511555:1.66914;
		specparam tpd_C_Q_posedge_f = 0.347793:0.476728:1.08678;
		specparam tpd_C_XQ_posedge_r = 0.428429:0.552579:1.69211;
		specparam tpd_C_XQ_posedge_f = 0.444198:0.544664:1.13622;
		specparam tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge = 0.214512:0.218735:0.38505;
		specparam thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge = -0.139293:-0.170539:-0.337943;
		specparam tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge = 0.214512:0.218735:0.38505;
		specparam thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge = -0.139293:-0.170539:-0.337943;
		specparam tsetup_SIN_C_SMC_posedge_SMC_posedge = 0.212229:0.216832:0.385081;
		specparam thold_SIN_C_SMC_posedge_SMC_posedge = -0.136929:-0.168539:-0.338875;
		specparam tsetup_SIN_C_SMC_negedge_SMC_posedge = 0.212229:0.216832:0.385081;
		specparam thold_SIN_C_SMC_negedge_SMC_posedge = -0.136929:-0.168539:-0.338875;
		specparam tsetup_SMC_C_adacond0_posedge_adacond0_posedge = 0.361813:0.354495:0.38926;
		specparam thold_SMC_C_adacond0_posedge_adacond0_posedge = -0.11607:-0.160421:-0.251155;
		specparam tsetup_SMC_C_adacond0_negedge_adacond0_posedge = 0.361813:0.354495:0.38926;
		specparam thold_SMC_C_adacond0_negedge_adacond0_posedge = -0.11607:-0.160421:-0.251155;
		specparam tpw_C_posedge = 0.213507:0.330811:2.72095;
		specparam tpw_C_negedge = 0.213507:0.330811:2.72095;

		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_posedge_SMC_posedge, 
			 thold_SIN_C_SMC_posedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_negedge_SMC_posedge, 
			 thold_SIN_C_SMC_negedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_posedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_negedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFQX 
`timescale 1ns/10ps
`celldefine
module SDFFQXX4 (Q, XQ, D, SIN, SMC, C);
	output Q, XQ;
	input D, SIN, SMC, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	wire int_fwire_s =0;
	wire int_fwire_r =0;
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
//	altos_dff_err (xcr_0, delayed_C, int_fwire_d);
//	altos_dff (int_fwire_IQ, notifier, delayed_C, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_C_Q_posedge_r = 0.381585:0.525081:1.67831;
		specparam tpd_C_Q_posedge_f = 0.344179:0.465002:1.06717;
		specparam tpd_C_XQ_posedge_r = 0.450674:0.576608:1.72348;
		specparam tpd_C_XQ_posedge_f = 0.503598:0.609394:1.21092;
		specparam tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge = 0.189291:0.194827:0.347631;
		specparam thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge = -0.123736:-0.152353:-0.300867;
		specparam tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge = 0.189291:0.194827:0.347631;
		specparam thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge = -0.123736:-0.152353:-0.300867;
		specparam tsetup_SIN_C_SMC_posedge_SMC_posedge = 0.184567:0.193358:0.345344;
		specparam thold_SIN_C_SMC_posedge_SMC_posedge = -0.123776:-0.152458:-0.30292;
		specparam tsetup_SIN_C_SMC_negedge_SMC_posedge = 0.184567:0.193358:0.345344;
		specparam thold_SIN_C_SMC_negedge_SMC_posedge = -0.123776:-0.152458:-0.30292;
		specparam tsetup_SMC_C_adacond0_posedge_adacond0_posedge = 0.330735:0.319185:0.345146;
		specparam thold_SMC_C_adacond0_posedge_adacond0_posedge = -0.102522:-0.142718:-0.215751;
		specparam tsetup_SMC_C_adacond0_negedge_adacond0_posedge = 0.330735:0.319185:0.345146;
		specparam thold_SMC_C_adacond0_negedge_adacond0_posedge = -0.102522:-0.142718:-0.215751;
		specparam tpw_C_posedge = 0.239353:0.330811:2.72095;
		specparam tpw_C_negedge = 0.239353:0.330811:2.72095;

		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_posedge_SMC_posedge, 
			 thold_SIN_C_SMC_posedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_negedge_SMC_posedge, 
			 thold_SIN_C_SMC_negedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_posedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_negedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFQX 
`timescale 1ns/10ps
`celldefine
module SDFFQXXL (Q, XQ, D, SIN, SMC, C);
	output Q, XQ;
	input D, SIN, SMC, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	altos_dff_err (xcr_0, delayed_C, int_fwire_d);
	altos_dff (int_fwire_IQ, notifier, delayed_C, int_fwire_d, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, D__bar, int_twire_0;
	wire int_twire_1, SIN__bar;


	// Additional timing gates
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar);
	or (adacond0, int_twire_1, int_twire_0);

	specify
		specparam tpd_C_Q_posedge_r = 0.359921:0.50505:1.66272;
		specparam tpd_C_Q_posedge_f = 0.32906:0.468436:1.44123;
		specparam tpd_C_XQ_posedge_r = 0.380064:0.510008:1.64942;
		specparam tpd_C_XQ_posedge_f = 0.437123:0.561932:1.54549;
		specparam tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge = 0.238652:0.232168:0.387611;
		specparam thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge = -0.137866:-0.166156:-0.333881;
		specparam tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge = 0.238652:0.232168:0.387611;
		specparam thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge = -0.137866:-0.166156:-0.333881;
		specparam tsetup_SIN_C_SMC_posedge_SMC_posedge = 0.234591:0.23066:0.387908;
		specparam thold_SIN_C_SMC_posedge_SMC_posedge = -0.135845:-0.164881:-0.330362;
		specparam tsetup_SIN_C_SMC_negedge_SMC_posedge = 0.234591:0.23066:0.387908;
		specparam thold_SIN_C_SMC_negedge_SMC_posedge = -0.135845:-0.164881:-0.330362;
		specparam tsetup_SMC_C_adacond0_posedge_adacond0_posedge = 0.3692:0.358724:0.394548;
		specparam thold_SMC_C_adacond0_posedge_adacond0_posedge = -0.11374:-0.156513:-0.252848;
		specparam tsetup_SMC_C_adacond0_negedge_adacond0_posedge = 0.3692:0.358724:0.394548;
		specparam thold_SMC_C_adacond0_negedge_adacond0_posedge = -0.11374:-0.156513:-0.252848;
		specparam tpw_C_posedge = 0.210609:0.330811:2.72095;
		specparam tpw_C_negedge = 0.210609:0.330811:2.72095;

		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& ~SMC, posedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_posedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_posedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& ~SMC, negedge D &&& ~SMC, 
			 tsetup_D_C_NTB_SMC_negedge_NTB_SMC_posedge, 
			 thold_D_C_NTB_SMC_negedge_NTB_SMC_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& SMC, posedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_posedge_SMC_posedge, 
			 thold_SIN_C_SMC_posedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& SMC, negedge SIN &&& SMC, 
			 tsetup_SIN_C_SMC_negedge_SMC_posedge, 
			 thold_SIN_C_SMC_negedge_SMC_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond0, posedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_posedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond0, negedge SMC &&& adacond0, 
			 tsetup_SMC_C_adacond0_negedge_adacond0_posedge, 
			 thold_SMC_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_SMC);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFRQ 
`timescale 1ns/10ps
`celldefine
module SDFFRQX1 (Q, D, SIN, SMC, XR, C);
	output Q;
	input D, SIN, SMC, XR, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_r;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, XR);
	wire int_fwire_s =0;
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.121454:0.259894:1.19483;
		specparam tpd_XR_Q_negedge_f = 0.121454:0.259894:1.19483;
		specparam tpd_C_Q_posedge_r = 0.347465:0.487921:1.5948;
		specparam tpd_C_Q_posedge_f = 0.330528:0.443747:1.01713;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.227225:0.230416:0.456049;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.150259:-0.181342:-0.390821;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.227225:0.230416:0.456049;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.150259:-0.181342:-0.390821;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.22594:0.237977:0.484457;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.149526:-0.184458:-0.417853;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.22594:0.237977:0.484457;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.149526:-0.184458:-0.417853;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.354857:0.344185:0.456984;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.128206:-0.170664:-0.230066;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.354857:0.344185:0.456984;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.128206:-0.170664:-0.230066;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.184925:-0.230426:0.234895;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.248704:0.342846:0.709403;
		specparam tpw_XR_negedge = 0.297484:0.396376:2.72095;
		specparam tpw_C_posedge = 0.178738:0.330811:2.72095;
		specparam tpw_C_negedge = 0.178738:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFRQ 
`timescale 1ns/10ps
`celldefine
module SDFFRQX2 (Q, D, SIN, SMC, XR, C);
	output Q;
	input D, SIN, SMC, XR, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_r;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.133424:0.278408:1.22067;
		specparam tpd_XR_Q_negedge_f = 0.133424:0.278408:1.22067;
		specparam tpd_C_Q_posedge_r = 0.361129:0.509625:1.66223;
		specparam tpd_C_Q_posedge_f = 0.323557:0.443559:1.04055;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.210214:0.218744:0.381752;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.143924:-0.171028:-0.334549;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.210214:0.218744:0.381752;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.143924:-0.171028:-0.334549;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.215019:0.225907:0.414139;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.146579:-0.178566:-0.36597;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.215019:0.225907:0.414139;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.146579:-0.178566:-0.36597;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.363631:0.35235:0.388199;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.122288:-0.165107:-0.221111;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.363631:0.35235:0.388199;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.122288:-0.165107:-0.221111;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.183892:-0.235135:0.184329;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.250857:0.345753:0.765094;
		specparam tpw_XR_negedge = 0.297484:0.396376:2.72095;
		specparam tpw_C_posedge = 0.205376:0.330811:2.72095;
		specparam tpw_C_negedge = 0.205376:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFRQ 
`timescale 1ns/10ps
`celldefine
module SDFFRQX4 (Q, D, SIN, SMC, XR, C);
	output Q;
	input D, SIN, SMC, XR, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_r;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.15057:0.30109:1.27788;
		specparam tpd_XR_Q_negedge_f = 0.15057:0.30109:1.27788;
		specparam tpd_C_Q_posedge_r = 0.419345:0.569975:1.72559;
		specparam tpd_C_Q_posedge_f = 0.351011:0.469715:1.04804;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.183732:0.194296:0.327919;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.125037:-0.152346:-0.281476;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.183732:0.194296:0.327919;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.125037:-0.152346:-0.281476;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.189155:0.204702:0.37433;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.133328:-0.164074:-0.326081;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.189155:0.204702:0.37433;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.133328:-0.164074:-0.326081;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.373374:0.356056:0.34102;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.111962:-0.14892:-0.208467;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.373374:0.356056:0.34102;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.111962:-0.14892:-0.208467;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.184607:-0.262141:0.0762013;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.235809:0.334282:0.752971;
		specparam tpw_XR_negedge = 0.30786:0.404243:2.72095;
		specparam tpw_C_posedge = 0.262871:0.330811:2.72095;
		specparam tpw_C_negedge = 0.262871:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFRQ 
`timescale 1ns/10ps
`celldefine
module SDFFRQXL (Q, D, SIN, SMC, XR, C);
	output Q;
	input D, SIN, SMC, XR, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_r;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.113786:0.250103:1.23372;
		specparam tpd_XR_Q_negedge_f = 0.113786:0.250103:1.23372;
		specparam tpd_C_Q_posedge_r = 0.34101:0.478401:1.57866;
		specparam tpd_C_Q_posedge_f = 0.323591:0.436332:1.08485;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.227242:0.234612:0.459139;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.149277:-0.181931:-0.394111;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.227242:0.234612:0.459139;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.149277:-0.181931:-0.394111;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.229331:0.238751:0.49064;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.153043:-0.187394:-0.422384;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.229331:0.238751:0.49064;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.153043:-0.187394:-0.422384;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.352331:0.346091:0.466784;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.127609:-0.173451:-0.226953;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.352331:0.346091:0.466784;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.127609:-0.173451:-0.226953;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.185016:-0.228897:0.219659;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.248704:0.342846:0.710658;
		specparam tpw_XR_negedge = 0.299393:0.396376:2.72095;
		specparam tpw_C_posedge = 0.173675:0.330811:2.72095;
		specparam tpw_C_negedge = 0.173675:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFRQX 
`timescale 1ns/10ps
`celldefine
module SDFFRQXX1 (Q, XQ, D, SIN, SMC, XR, C);
	output Q, XQ;
	input D, SIN, SMC, XR, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.121538:0.259198:1.19188;
		specparam tpd_XR_Q_negedge_f = 0.121538:0.259198:1.19188;
		specparam tpd_C_Q_posedge_r = 0.353863:0.493173:1.59348;
		specparam tpd_C_Q_posedge_f = 0.332861:0.445411:1.01839;
		specparam tpd_XR_XQ_negedge_r = 0.218398:0.384154:1.82491;
		specparam tpd_XR_XQ_negedge_f = 0.218398:0.384154:1.82491;
		specparam tpd_C_XQ_posedge_r = 0.403851:0.530763:1.63745;
		specparam tpd_C_XQ_posedge_f = 0.435678:0.547385:1.28312;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.22229:0.230677:0.454529;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.148283:-0.179552:-0.389848;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.22229:0.230677:0.454529;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.148283:-0.179552:-0.389848;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.223893:0.236482:0.483777;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.149352:-0.184981:-0.420752;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.223893:0.236482:0.483777;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.149352:-0.184981:-0.420752;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.35538:0.348185:0.455436;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.128616:-0.170993:-0.22863;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.35538:0.348185:0.455436;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.128616:-0.170993:-0.22863;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.185818:-0.234044:0.224136;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.247522:0.340705:0.711544;
		specparam tpw_XR_negedge = 0.299393:0.396376:2.72095;
		specparam tpw_C_posedge = 0.187092:0.330811:2.72095;
		specparam tpw_C_negedge = 0.187092:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFRQX 
`timescale 1ns/10ps
`celldefine
module SDFFRQXX2 (Q, XQ, D, SIN, SMC, XR, C);
	output Q, XQ;
	input D, SIN, SMC, XR, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.137552:0.283247:1.23541;
		specparam tpd_XR_Q_negedge_f = 0.137552:0.283247:1.23541;
		specparam tpd_C_Q_posedge_r = 0.372169:0.520922:1.68264;
		specparam tpd_C_Q_posedge_f = 0.331534:0.452235:1.05542;
		specparam tpd_XR_XQ_negedge_r = 0.26349:0.42924:1.88189;
		specparam tpd_XR_XQ_negedge_f = 0.26349:0.42924:1.88189;
		specparam tpd_C_XQ_posedge_r = 0.430071:0.557168:1.68202;
		specparam tpd_C_XQ_posedge_f = 0.489472:0.601767:1.31213;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.211117:0.217748:0.382293;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.142307:-0.170823:-0.332331;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.211117:0.217748:0.382293;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.142307:-0.170823:-0.332331;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.214486:0.225003:0.413525;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.143986:-0.178075:-0.365907;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.214486:0.225003:0.413525;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.143986:-0.178075:-0.365907;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.363356:0.352863:0.383922;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.121002:-0.163808:-0.225279;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.363356:0.352863:0.383922;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.121002:-0.163808:-0.225279;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.186606:-0.237153:0.183859;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.25088:0.345753:0.765094;
		specparam tpw_XR_negedge = 0.299153:0.398998:2.72095;
		specparam tpw_C_posedge = 0.228619:0.330811:2.72095;
		specparam tpw_C_negedge = 0.228619:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFRQX 
`timescale 1ns/10ps
`celldefine
module SDFFRQXX4 (Q, XQ, D, SIN, SMC, XR, C);
	output Q, XQ;
	input D, SIN, SMC, XR, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.153784:0.303583:1.27995;
		specparam tpd_XR_Q_negedge_f = 0.153784:0.303583:1.27995;
		specparam tpd_C_Q_posedge_r = 0.433172:0.581984:1.72785;
		specparam tpd_C_Q_posedge_f = 0.362443:0.481085:1.05731;
		specparam tpd_XR_XQ_negedge_r = 0.274477:0.436877:1.95638;
		specparam tpd_XR_XQ_negedge_f = 0.274477:0.436877:1.95638;
		specparam tpd_C_XQ_posedge_r = 0.459901:0.587613:1.73071;
		specparam tpd_C_XQ_posedge_f = 0.541899:0.652553:1.36831;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.184439:0.194296:0.328996;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.124353:-0.154217:-0.28396;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.184439:0.194296:0.328996;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.124353:-0.154217:-0.28396;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.189337:0.205006:0.374526;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.133682:-0.163661:-0.326036;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.189337:0.205006:0.374526;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.133682:-0.163661:-0.326036;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.373711:0.356711:0.337887;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.108917:-0.150805:-0.207769;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.373711:0.356711:0.337887;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.108917:-0.150805:-0.207769;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.184868:-0.264846:0.0746209;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.236484:0.334282:0.754226;
		specparam tpw_XR_negedge = 0.311591:0.406866:2.72095;
		specparam tpw_C_posedge = 0.28869:0.330811:2.72095;
		specparam tpw_C_negedge = 0.28869:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFRQX 
`timescale 1ns/10ps
`celldefine
module SDFFRQXXL (Q, XQ, D, SIN, SMC, XR, C);
	output Q, XQ;
	input D, SIN, SMC, XR, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_r, XR);
	altos_dff_r_err (xcr_0, delayed_C, int_fwire_d, int_fwire_r);
	altos_dff_r (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR);
	and (adacond1, SMC, XR);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN, SMC);
	and (int_twire_3, D, SIN__bar, SMC__bar);
	and (int_twire_4, D, SIN);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XR_Q_negedge_r = 0.114704:0.251339:1.23955;
		specparam tpd_XR_Q_negedge_f = 0.114704:0.251339:1.23955;
		specparam tpd_C_Q_posedge_r = 0.34848:0.486458:1.59584;
		specparam tpd_C_Q_posedge_f = 0.327554:0.44097:1.09498;
		specparam tpd_XR_XQ_negedge_r = 0.206373:0.371302:1.7956;
		specparam tpd_XR_XQ_negedge_f = 0.206373:0.371302:1.7956;
		specparam tpd_C_XQ_posedge_r = 0.392821:0.520172:1.63147;
		specparam tpd_C_XQ_posedge_f = 0.414738:0.517726:1.16432;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.224552:0.233358:0.459691;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.149483:-0.182018:-0.39511;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.224552:0.233358:0.459691;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.149483:-0.182018:-0.39511;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.230733:0.237728:0.490152;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.149983:-0.185488:-0.425459;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.230733:0.237728:0.490152;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.149983:-0.185488:-0.425459;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.35177:0.346091:0.463183;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.129617:-0.171235:-0.226828;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.35177:0.346091:0.463183;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.129617:-0.171235:-0.226828;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.187922:-0.233972:0.221087;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.247522:0.340705:0.708801;
		specparam tpw_XR_negedge = 0.301517:0.396376:2.72095;
		specparam tpw_C_posedge = 0.18127:0.330811:2.72095;
		specparam tpw_C_negedge = 0.18127:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSQ 
`timescale 1ns/10ps
`celldefine
module SDFFSQX1 (Q, D, SIN, SMC, XS, C);
	output Q;
	input D, SIN, SMC, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_s;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, XS);
	wire int_fwire_r =0;
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.280292:0.437397:1.88119;
		specparam tpd_XS_Q_negedge_f = 0.280292:0.437397:1.88119;
		specparam tpd_C_Q_posedge_r = 0.303991:0.436726:1.54523;
		specparam tpd_C_Q_posedge_f = 0.333417:0.444705:1.04455;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.237188:0.238918:0.456815;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.142981:-0.175882:-0.381294;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.237188:0.238918:0.456815;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.142981:-0.175882:-0.381294;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.242944:0.246327:0.486487;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.14448:-0.180842:-0.408055;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.242944:0.246327:0.486487;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.14448:-0.180842:-0.408055;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.403575:0.387231:0.460294;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.122614:-0.165801:-0.240688;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.403575:0.387231:0.460294;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.122614:-0.165801:-0.240688;
		specparam trecovery_XS_C_adacond3_posedge_adacond3_posedge = -0.0362598:-0.0550443:0.172789;
		specparam tremoval_XS_C_adacond3_posedge_adacond3_posedge = 0.106758:0.126923:0.0335127;
		specparam tpw_XS_negedge = 0.166101:0.330811:2.72095;
		specparam tpw_C_posedge = 0.160643:0.330811:2.72095;
		specparam tpw_C_negedge = 0.160643:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XS &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSQ 
`timescale 1ns/10ps
`celldefine
module SDFFSQX2 (Q, D, SIN, SMC, XS, C);
	output Q;
	input D, SIN, SMC, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_s;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.296421:0.457133:1.90435;
		specparam tpd_XS_Q_negedge_f = 0.296421:0.457133:1.90435;
		specparam tpd_C_Q_posedge_r = 0.317235:0.456428:1.61442;
		specparam tpd_C_Q_posedge_f = 0.330086:0.447224:1.05838;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.219907:0.221108:0.380582;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.138602:-0.167835:-0.324936;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.219907:0.221108:0.380582;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.138602:-0.167835:-0.324936;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.223718:0.229295:0.415176;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.142813:-0.174717:-0.35385;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.223718:0.229295:0.415176;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.142813:-0.174717:-0.35385;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.414511:0.393509:0.385615;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.117931:-0.157965:-0.232017;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.414511:0.393509:0.385615;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.117931:-0.157965:-0.232017;
		specparam trecovery_XS_C_adacond3_posedge_adacond3_posedge = -0.0213946:-0.0428599:0.141027;
		specparam tremoval_XS_C_adacond3_posedge_adacond3_posedge = 0.0851825:0.105092:0.0596502;
		specparam tpw_XS_negedge = 0.176647:0.330811:2.72095;
		specparam tpw_C_posedge = 0.181559:0.330811:2.72095;
		specparam tpw_C_negedge = 0.181559:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XS &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSQ 
`timescale 1ns/10ps
`celldefine
module SDFFSQX4 (Q, D, SIN, SMC, XS, C);
	output Q;
	input D, SIN, SMC, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_s;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.338155:0.499079:1.94816;
		specparam tpd_XS_Q_negedge_f = 0.338155:0.499079:1.94816;
		specparam tpd_C_Q_posedge_r = 0.367409:0.507614:1.64636;
		specparam tpd_C_Q_posedge_f = 0.366897:0.483014:1.05462;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.191465:0.195765:0.33008;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.119585:-0.149369:-0.274906;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.191465:0.195765:0.33008;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.119585:-0.149369:-0.274906;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.197048:0.209286:0.373726;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.127327:-0.157906:-0.318194;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.197048:0.209286:0.373726;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.127327:-0.157906:-0.318194;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.423755:0.401615:0.333655;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.104284:-0.144754:-0.22423;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.423755:0.401615:0.333655;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.104284:-0.144754:-0.22423;
		specparam trecovery_XS_C_adacond3_posedge_adacond3_posedge = -0.0225217:-0.043226:0.16524;
		specparam tremoval_XS_C_adacond3_posedge_adacond3_posedge = 0.0838653:0.101728:0.0473518;
		specparam tpw_XS_negedge = 0.191731:0.333433:2.72095;
		specparam tpw_C_posedge = 0.231504:0.330811:2.72095;
		specparam tpw_C_negedge = 0.231504:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XS &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSQ 
`timescale 1ns/10ps
`celldefine
module SDFFSQXL (Q, D, SIN, SMC, XS, C);
	output Q;
	input D, SIN, SMC, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_s;
	wire xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.287087:0.444438:1.89814;
		specparam tpd_XS_Q_negedge_f = 0.287087:0.444438:1.89814;
		specparam tpd_C_Q_posedge_r = 0.308328:0.440706:1.5535;
		specparam tpd_C_Q_posedge_f = 0.325852:0.438363:1.13095;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.241581:0.240974:0.46452;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.146078:-0.177092:-0.384501;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.241581:0.240974:0.46452;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.146078:-0.177092:-0.384501;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.243431:0.249527:0.494412;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.14744:-0.181027:-0.41323;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.243431:0.249527:0.494412;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.14744:-0.181027:-0.41323;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.40293:0.387096:0.467434;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.122595:-0.1665:-0.238835;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.40293:0.387096:0.467434;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.122595:-0.1665:-0.238835;
		specparam trecovery_XS_C_adacond3_posedge_adacond3_posedge = -0.0344304:-0.051519:0.176732;
		specparam tremoval_XS_C_adacond3_posedge_adacond3_posedge = 0.107103:0.125:0.0299135;
		specparam tpw_XS_negedge = 0.165833:0.330811:2.72095;
		specparam tpw_C_posedge = 0.160643:0.330811:2.72095;
		specparam tpw_C_negedge = 0.160643:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XS &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSQX 
`timescale 1ns/10ps
`celldefine
module SDFFSQXX1 (Q, XQ, D, SIN, SMC, XS, C);
	output Q, XQ;
	input D, SIN, SMC, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.310802:0.466121:1.92389;
		specparam tpd_XS_Q_negedge_f = 0.310802:0.466121:1.92389;
		specparam tpd_C_Q_posedge_r = 0.307958:0.440487:1.55023;
		specparam tpd_C_Q_posedge_f = 0.338386:0.450357:1.05103;
		specparam tpd_XS_XQ_negedge_r = 0.139643:0.297561:1.4245;
		specparam tpd_XS_XQ_negedge_f = 0.139643:0.297561:1.4245;
		specparam tpd_C_XQ_posedge_r = 0.444638:0.578023:1.68181;
		specparam tpd_C_XQ_posedge_f = 0.396672:0.512016:1.25002;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.237843:0.239249:0.455067;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.143976:-0.175858:-0.382572;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.237843:0.239249:0.455067;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.143976:-0.175858:-0.382572;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.239042:0.241481:0.485535;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.143772:-0.180779:-0.410864;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.239042:0.241481:0.485535;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.143772:-0.180779:-0.410864;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.404945:0.387412:0.460176;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.122027:-0.166344:-0.241048;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.404945:0.387412:0.460176;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.122027:-0.166344:-0.241048;
		specparam trecovery_XS_C_adacond3_posedge_adacond3_posedge = -0.0362202:-0.0565572:0.168965;
		specparam tremoval_XS_C_adacond3_posedge_adacond3_posedge = 0.106758:0.126923:0.0306532;
		specparam tpw_XS_negedge = 0.195289:0.330811:2.72095;
		specparam tpw_C_posedge = 0.165812:0.330811:2.72095;
		specparam tpw_C_negedge = 0.165812:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XS &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSQX 
`timescale 1ns/10ps
`celldefine
module SDFFSQXX2 (Q, XQ, D, SIN, SMC, XS, C);
	output Q, XQ;
	input D, SIN, SMC, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.360314:0.519863:2.0121;
		specparam tpd_XS_Q_negedge_f = 0.360314:0.519863:2.0121;
		specparam tpd_C_Q_posedge_r = 0.325221:0.46447:1.62862;
		specparam tpd_C_Q_posedge_f = 0.341455:0.459984:1.07332;
		specparam tpd_XS_XQ_negedge_r = 0.152379:0.313897:1.43302;
		specparam tpd_XS_XQ_negedge_f = 0.152379:0.313897:1.43302;
		specparam tpd_C_XQ_posedge_r = 0.476019:0.614833:1.75841;
		specparam tpd_C_XQ_posedge_f = 0.439825:0.559784:1.30601;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.216485:0.220377:0.37947;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.137796:-0.167777:-0.32872;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.216485:0.220377:0.37947;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.137796:-0.167777:-0.32872;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.222283:0.226875:0.413738;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.138985:-0.174938:-0.355458;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.222283:0.226875:0.413738;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.138985:-0.174938:-0.355458;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.414218:0.393595:0.385597;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.116587:-0.159977:-0.235925;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.414218:0.393595:0.385597;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.116587:-0.159977:-0.235925;
		specparam trecovery_XS_C_adacond3_posedge_adacond3_posedge = -0.021775:-0.0438981:0.141871;
		specparam tremoval_XS_C_adacond3_posedge_adacond3_posedge = 0.0851825:0.105092:0.0540729;
		specparam tpw_XS_negedge = 0.232157:0.37015:2.72095;
		specparam tpw_C_posedge = 0.197659:0.330811:2.72095;
		specparam tpw_C_negedge = 0.197659:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XS &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSQX 
`timescale 1ns/10ps
`celldefine
module SDFFSQXX4 (Q, XQ, D, SIN, SMC, XS, C);
	output Q, XQ;
	input D, SIN, SMC, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.383796:0.544737:2.03864;
		specparam tpd_XS_Q_negedge_f = 0.383796:0.544737:2.03864;
		specparam tpd_C_Q_posedge_r = 0.375996:0.516601:1.67387;
		specparam tpd_C_Q_posedge_f = 0.378321:0.495787:1.07561;
		specparam tpd_XS_XQ_negedge_r = 0.144343:0.303181:1.4057;
		specparam tpd_XS_XQ_negedge_f = 0.144343:0.303181:1.4057;
		specparam tpd_C_XQ_posedge_r = 0.512448:0.648902:1.78401;
		specparam tpd_C_XQ_posedge_f = 0.481191:0.59574:1.31211;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.186715:0.195765:0.326245;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.122718:-0.146171:-0.271818;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.186715:0.195765:0.326245;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.122718:-0.146171:-0.271818;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.19711:0.208738:0.374079;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.126622:-0.159324:-0.31565;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.19711:0.208738:0.374079;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.126622:-0.159324:-0.31565;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.422538:0.401731:0.333728;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.104666:-0.143817:-0.225133;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.422538:0.401731:0.333728;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.104666:-0.143817:-0.225133;
		specparam trecovery_XS_C_adacond3_posedge_adacond3_posedge = -0.0250733:-0.0419187:0.170554;
		specparam tremoval_XS_C_adacond3_posedge_adacond3_posedge = 0.0838653:0.101728:0.0445168;
		specparam tpw_XS_negedge = 0.245991:0.375395:2.72095;
		specparam tpw_C_posedge = 0.249513:0.330811:2.72095;
		specparam tpw_C_negedge = 0.249513:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XS &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSQX 
`timescale 1ns/10ps
`celldefine
module SDFFSQXXL (Q, XQ, D, SIN, SMC, XS, C);
	output Q, XQ;
	input D, SIN, SMC, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, XS);
	altos_dff_s_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s);
	altos_dff_s (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, xcr_0);
	buf (Q, int_fwire_IQ);
	not (int_fwire_IXQ, int_fwire_IQ);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, D__bar, int_twire_0;
	wire int_twire_1, int_twire_2, int_twire_3;
	wire int_twire_4, SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XS);
	and (adacond1, SMC, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, D__bar, SIN__bar);
	and (int_twire_3, D__bar, SIN, SMC__bar);
	and (int_twire_4, D, SIN__bar, SMC);
	or (adacond3, int_twire_4, int_twire_3, int_twire_2);

	specify
		specparam tpd_XS_Q_negedge_r = 0.303636:0.458686:1.90472;
		specparam tpd_XS_Q_negedge_f = 0.303636:0.458686:1.90472;
		specparam tpd_C_Q_posedge_r = 0.312705:0.444267:1.54937;
		specparam tpd_C_Q_posedge_f = 0.331836:0.444607:1.13092;
		specparam tpd_XS_XQ_negedge_r = 0.132113:0.277714:1.30377;
		specparam tpd_XS_XQ_negedge_f = 0.132113:0.277714:1.30377;
		specparam tpd_C_XQ_posedge_r = 0.430824:0.56232:1.67289;
		specparam tpd_C_XQ_posedge_f = 0.388899:0.494515:1.14681;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.24269:0.241278:0.461071;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.144444:-0.177029:-0.386204;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.24269:0.241278:0.461071;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.144444:-0.177029:-0.386204;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.244185:0.248279:0.492512;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.14725:-0.181554:-0.411348;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.244185:0.248279:0.492512;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.14725:-0.181554:-0.411348;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.403115:0.387096:0.4636;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.122258:-0.167469:-0.237015;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.403115:0.387096:0.4636;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.122258:-0.167469:-0.237015;
		specparam trecovery_XS_C_adacond3_posedge_adacond3_posedge = -0.0349433:-0.0513397:0.17771;
		specparam tremoval_XS_C_adacond3_posedge_adacond3_posedge = 0.107103:0.125:0.025916;
		specparam tpw_XS_negedge = 0.18568:0.330811:2.72095;
		specparam tpw_C_posedge = 0.165812:0.330811:2.72095;
		specparam tpw_C_negedge = 0.165812:0.330811:2.72095;

		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$recovery (posedge XS &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XS &&& adacond3, 
			 tremoval_XS_C_adacond3_posedge_adacond3_posedge, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSRQ 
`timescale 1ns/10ps
`celldefine
module SDFFSRQX1 (Q, D, SIN, SMC, XR, XS, C);
	output Q;
	input D, SIN, SMC, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.123755:0.247715:1.41372;
		specparam tpd_XR_Q_negedge_f = 0.116677:0.25199:1.17506;
		specparam tpd_XS_Q_negedge_r = 0.324373:0.486878:1.92562;
		specparam tpd_XS_Q_negedge_f = 0.324373:0.486878:1.92562;
		specparam tpd_C_Q_posedge_r = 0.343447:0.482205:1.57352;
		specparam tpd_C_Q_posedge_f = 0.342771:0.453834:1.02373;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.248783:0.248663:0.463958;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.149181:-0.179853:-0.386866;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.248783:0.248663:0.463958;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.149181:-0.179853:-0.386866;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.250714:0.253072:0.497046;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.150169:-0.183765:-0.412313;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.250714:0.253072:0.497046;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.150169:-0.183765:-0.412313;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.407447:0.392502:0.469353;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.125965:-0.170286:-0.231624;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.407447:0.392502:0.469353;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.125965:-0.170286:-0.231624;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.19143:-0.231981:0.226518;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.273632:0.363343:0.736732;
		specparam tpw_XR_negedge = 0.337912:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0203264:0.00665868:0.00452136;
		specparam thold_XR_XS_posedge_posedge = 0.0414123:0.0577229:0.12472;
		specparam trecovery_XS_C_adacond4_posedge_adacond4_posedge = -0.0313879:-0.0535521:0.172943;
		specparam tremoval_XS_C_adacond4_posedge_adacond4_posedge = 0.125819:0.149845:0.0660077;
		specparam tsetup_XS_XR_posedge_posedge = 0.0418878:0.0670319:0.187811;
		specparam thold_XS_XR_posedge_posedge = 0.0522923:0.0607994:0.0412665;
		specparam tpw_XS_negedge = 0.191304:0.330811:2.72095;
		specparam tpw_C_posedge = 0.178738:0.330811:2.72095;
		specparam tpw_C_negedge = 0.178738:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$recovery (posedge XS &&& adacond4, posedge C &&& adacond4, 
			 trecovery_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$hold (posedge C &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSRQ 
`timescale 1ns/10ps
`celldefine
module SDFFSRQX2 (Q, D, SIN, SMC, XR, XS, C);
	output Q;
	input D, SIN, SMC, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.141629:0.274581:1.46144;
		specparam tpd_XR_Q_negedge_f = 0.134504:0.278175:1.21523;
		specparam tpd_XS_Q_negedge_r = 0.345684:0.514001:1.94578;
		specparam tpd_XS_Q_negedge_f = 0.345684:0.514001:1.94578;
		specparam tpd_C_Q_posedge_r = 0.364474:0.511774:1.64316;
		specparam tpd_C_Q_posedge_f = 0.344629:0.463537:1.05269;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.224937:0.226577:0.390482;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.142633:-0.170907:-0.331498;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.224937:0.226577:0.390482;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.142633:-0.170907:-0.331498;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.230926:0.235919:0.42288;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.145476:-0.178476:-0.360402;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.230926:0.235919:0.42288;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.145476:-0.178476:-0.360402;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.416703:0.3954:0.39454;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.122383:-0.162027:-0.22691;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.416703:0.3954:0.39454;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.122383:-0.162027:-0.22691;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.189555:-0.236356:0.188192;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.275915:0.368314:0.794319;
		specparam tpw_XR_negedge = 0.333348:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0188554:0.00865447:0.0441122;
		specparam thold_XR_XS_posedge_posedge = 0.0269967:0.0359833:0.111576;
		specparam trecovery_XS_C_adacond4_posedge_adacond4_posedge = -0.021648:-0.0446427:0.138316;
		specparam tremoval_XS_C_adacond4_posedge_adacond4_posedge = 0.103884:0.129129:0.0888732;
		specparam tsetup_XS_XR_posedge_posedge = 0.035635:0.0509407:0.188099;
		specparam thold_XS_XR_posedge_posedge = 0.0496903:0.0582862:0.0780327;
		specparam tpw_XS_negedge = 0.203195:0.330811:2.72095;
		specparam tpw_C_posedge = 0.210936:0.330811:2.72095;
		specparam tpw_C_negedge = 0.210936:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$recovery (posedge XS &&& adacond4, posedge C &&& adacond4, 
			 trecovery_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$hold (posedge C &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSRQ 
`timescale 1ns/10ps
`celldefine
module SDFFSRQX4 (Q, D, SIN, SMC, XR, XS, C);
	output Q;
	input D, SIN, SMC, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.143225:0.274532:1.43925;
		specparam tpd_XR_Q_negedge_f = 0.152634:0.302101:1.28025;
		specparam tpd_XS_Q_negedge_r = 0.391599:0.56148:2.02564;
		specparam tpd_XS_Q_negedge_f = 0.391599:0.56148:2.02564;
		specparam tpd_C_Q_posedge_r = 0.421567:0.571443:1.71537;
		specparam tpd_C_Q_posedge_f = 0.380062:0.498692:1.0719;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.196129:0.201233:0.334147;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.123788:-0.151335:-0.275311;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.196129:0.201233:0.334147;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.123788:-0.151335:-0.275311;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.205191:0.215478:0.378033;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.128726:-0.161994:-0.325879;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.205191:0.215478:0.378033;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.128726:-0.161994:-0.325879;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.425802:0.404269:0.346786;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.108078:-0.147546:-0.212966;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.425802:0.404269:0.346786;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.108078:-0.147546:-0.212966;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.191982:-0.265579:0.0718523;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.258333:0.352248:0.778164;
		specparam tpw_XR_negedge = 0.347218:0.433092:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0187123:0.0114331:0.0770791;
		specparam thold_XR_XS_posedge_posedge = 0.0320748:0.0444951:0.137237;
		specparam trecovery_XS_C_adacond4_posedge_adacond4_posedge = -0.0223429:-0.0450837:0.164682;
		specparam tremoval_XS_C_adacond4_posedge_adacond4_posedge = 0.10214:0.121541:0.0703786;
		specparam tsetup_XS_XR_posedge_posedge = 0.0163812:0.0235633:0.175637;
		specparam thold_XS_XR_posedge_posedge = 0.0540763:0.0622621:0.106637;
		specparam tpw_XS_negedge = 0.22326:0.354414:2.72095;
		specparam tpw_C_posedge = 0.265484:0.330811:2.72095;
		specparam tpw_C_negedge = 0.265484:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$recovery (posedge XS &&& adacond4, posedge C &&& adacond4, 
			 trecovery_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$hold (posedge C &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSRQ 
`timescale 1ns/10ps
`celldefine
module SDFFSRQXL (Q, D, SIN, SMC, XR, XS, C);
	output Q;
	input D, SIN, SMC, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_r;
	wire int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.123343:0.245487:1.42014;
		specparam tpd_XR_Q_negedge_f = 0.114092:0.249266:1.23133;
		specparam tpd_XS_Q_negedge_r = 0.321985:0.483088:1.9278;
		specparam tpd_XS_Q_negedge_f = 0.321985:0.483088:1.9278;
		specparam tpd_C_Q_posedge_r = 0.342143:0.479241:1.57376;
		specparam tpd_C_Q_posedge_f = 0.342982:0.455732:1.10305;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.251607:0.24741:0.471137;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.149846:-0.178338:-0.390238;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.251607:0.24741:0.471137;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.149846:-0.178338:-0.390238;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.251836:0.255813:0.498665;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.149925:-0.184717:-0.414419;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.251836:0.255813:0.498665;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.149925:-0.184717:-0.414419;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.405976:0.387346:0.474063;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.127471:-0.168855:-0.228739;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.405976:0.387346:0.474063;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.127471:-0.168855:-0.228739;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.193348:-0.229981:0.21978;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.271853:0.361124:0.733467;
		specparam tpw_XR_negedge = 0.339738:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0171954:0.00743541:-0.00394227;
		specparam thold_XR_XS_posedge_posedge = 0.0447904:0.0630319:0.129747;
		specparam trecovery_XS_C_adacond4_posedge_adacond4_posedge = -0.0362988:-0.0551914:0.172193;
		specparam tremoval_XS_C_adacond4_posedge_adacond4_posedge = 0.125526:0.150661:0.0649588;
		specparam tsetup_XS_XR_posedge_posedge = 0.0465529:0.0723054:0.192234;
		specparam thold_XS_XR_posedge_posedge = 0.0520275:0.0607994:0.0430453;
		specparam tpw_XS_negedge = 0.189036:0.330811:2.72095;
		specparam tpw_C_posedge = 0.176207:0.330811:2.72095;
		specparam tpw_C_negedge = 0.176207:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$recovery (posedge XS &&& adacond4, posedge C &&& adacond4, 
			 trecovery_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$hold (posedge C &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSRQX 
`timescale 1ns/10ps
`celldefine
module SDFFSRQXX1 (Q, XQ, D, SIN, SMC, XR, XS, C);
	output Q, XQ;
	input D, SIN, SMC, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.128154:0.254352:1.43858;
		specparam tpd_XR_Q_negedge_f = 0.120684:0.257681:1.19396;
		specparam tpd_XS_Q_negedge_r = 0.355194:0.517985:1.97677;
		specparam tpd_XS_Q_negedge_f = 0.355194:0.517985:1.97677;
		specparam tpd_C_Q_posedge_r = 0.352569:0.492735:1.59984;
		specparam tpd_C_Q_posedge_f = 0.352166:0.465243:1.04376;
		specparam tpd_XR_XQ_negedge_r = 0.268656:0.447658:1.88571;
		specparam tpd_XR_XQ_negedge_f = 0.268656:0.447658:1.88571;
		specparam tpd_XS_XQ_negedge_r = 0.144258:0.295276:1.54297;
		specparam tpd_XS_XQ_negedge_f = 0.139496:0.295292:1.4272;
		specparam tpd_C_XQ_posedge_r = 0.461681:0.59476:1.6899;
		specparam tpd_C_XQ_posedge_f = 0.447237:0.561571:1.28491;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.245383:0.246374:0.461622;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.147997:-0.178875:-0.385458;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.245383:0.246374:0.461622;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.147997:-0.178875:-0.385458;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.247163:0.250982:0.492613;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.150858:-0.182749:-0.415676;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.247163:0.250982:0.492613;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.150858:-0.182749:-0.415676;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.406539:0.39248:0.465109;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.127211:-0.168957:-0.233358;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.406539:0.39248:0.465109;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.127211:-0.168957:-0.233358;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.193593:-0.233908:0.22191;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.271853:0.361124:0.736209;
		specparam tpw_XR_negedge = 0.337541:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0197611:0.00606375:0.00307415;
		specparam thold_XR_XS_posedge_posedge = 0.0545913:0.0745493:0.134709;
		specparam trecovery_XS_C_adacond4_posedge_adacond4_posedge = -0.0323615:-0.0546672:0.171645;
		specparam tremoval_XS_C_adacond4_posedge_adacond4_posedge = 0.125819:0.149845:0.0630555;
		specparam tsetup_XS_XR_posedge_posedge = 0.0519166:0.0849135:0.229127;
		specparam thold_XS_XR_posedge_posedge = 0.0197611:0.00606375:-0.0677645;
		specparam tpw_XS_negedge = 0.217642:0.341301:2.72095;
		specparam tpw_C_posedge = 0.18737:0.330811:2.72095;
		specparam tpw_C_negedge = 0.18737:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$recovery (posedge XS &&& adacond4, posedge C &&& adacond4, 
			 trecovery_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$hold (posedge C &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSRQX 
`timescale 1ns/10ps
`celldefine
module SDFFSRQXX2 (Q, XQ, D, SIN, SMC, XR, XS, C);
	output Q, XQ;
	input D, SIN, SMC, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.144441:0.278621:1.47576;
		specparam tpd_XR_Q_negedge_f = 0.137135:0.281448:1.22756;
		specparam tpd_XS_Q_negedge_r = 0.408959:0.576949:2.05185;
		specparam tpd_XS_Q_negedge_f = 0.408959:0.576949:2.05185;
		specparam tpd_C_Q_posedge_r = 0.373832:0.521645:1.66514;
		specparam tpd_C_Q_posedge_f = 0.353871:0.474015:1.07132;
		specparam tpd_XR_XQ_negedge_r = 0.318646:0.502947:1.98823;
		specparam tpd_XR_XQ_negedge_f = 0.318646:0.502947:1.98823;
		specparam tpd_XS_XQ_negedge_r = 0.157751:0.315217:1.59538;
		specparam tpd_XS_XQ_negedge_f = 0.153397:0.313993:1.44699;
		specparam tpd_C_XQ_posedge_r = 0.494617:0.633843:1.78151;
		specparam tpd_C_XQ_posedge_f = 0.502787:0.620696:1.36217;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.226039:0.226577:0.388693;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.140226:-0.168725:-0.330064;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.226039:0.226577:0.388693;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.140226:-0.168725:-0.330064;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.229046:0.233813:0.419442;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.14319:-0.176335:-0.360171;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.229046:0.233813:0.419442;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.14319:-0.176335:-0.360171;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.418548:0.397159:0.392254;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.122783:-0.163481:-0.229133;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.418548:0.397159:0.392254;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.122783:-0.163481:-0.229133;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.193578:-0.238518:0.179996;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.27664:0.366085:0.793806;
		specparam tpw_XR_negedge = 0.335166:0.427847:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0185844:0.00821074:0.0213908;
		specparam thold_XR_XS_posedge_posedge = 0.056425:0.0721995:0.122699;
		specparam trecovery_XS_C_adacond4_posedge_adacond4_posedge = -0.025516:-0.045211:0.140892;
		specparam tremoval_XS_C_adacond4_posedge_adacond4_posedge = 0.103884:0.129129:0.0859307;
		specparam tsetup_XS_XR_posedge_posedge = 0.0629586:0.0883097:0.23238;
		specparam thold_XS_XR_posedge_posedge = 0.0185952:0.00821074:-0.0586669;
		specparam tpw_XS_negedge = 0.259298:0.383263:2.72095;
		specparam tpw_C_posedge = 0.231514:0.330811:2.72095;
		specparam tpw_C_negedge = 0.231514:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$recovery (posedge XS &&& adacond4, posedge C &&& adacond4, 
			 trecovery_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$hold (posedge C &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSRQX 
`timescale 1ns/10ps
`celldefine
module SDFFSRQXX4 (Q, XQ, D, SIN, SMC, XR, XS, C);
	output Q, XQ;
	input D, SIN, SMC, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.144465:0.276047:1.4379;
		specparam tpd_XR_Q_negedge_f = 0.151952:0.300337:1.27391;
		specparam tpd_XS_Q_negedge_r = 0.436834:0.606088:2.08568;
		specparam tpd_XS_Q_negedge_f = 0.436834:0.606088:2.08568;
		specparam tpd_C_Q_posedge_r = 0.432958:0.581577:1.72302;
		specparam tpd_C_Q_posedge_f = 0.390642:0.50936:1.08218;
		specparam tpd_XR_XQ_negedge_r = 0.321481:0.497477:2.0164;
		specparam tpd_XR_XQ_negedge_f = 0.321481:0.497477:2.0164;
		specparam tpd_XS_XQ_negedge_r = 0.137695:0.283757:1.50923;
		specparam tpd_XS_XQ_negedge_f = 0.145161:0.302818:1.41629;
		specparam tpd_C_XQ_posedge_r = 0.529115:0.665759:1.79836;
		specparam tpd_C_XQ_posedge_f = 0.550221:0.66322:1.37954;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.194313:0.201233:0.335634;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.12254:-0.1517:-0.276469;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.194313:0.201233:0.335634;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.12254:-0.1517:-0.276469;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.201891:0.212512:0.380157;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.131634:-0.161554:-0.324955;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.201891:0.212512:0.380157;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.131634:-0.161554:-0.324955;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.425949:0.404675:0.346838;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.107777:-0.147734:-0.214201;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.425949:0.404675:0.346838;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.107777:-0.147734:-0.214201;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.193822:-0.267909:0.0698085;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.256725:0.350029:0.778534;
		specparam tpw_XR_negedge = 0.351001:0.435715:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0162607:0.00551711:0.0268028;
		specparam thold_XR_XS_posedge_posedge = 0.0552996:0.0689859:0.144192;
		specparam trecovery_XS_C_adacond4_posedge_adacond4_posedge = -0.0258043:-0.0452946:0.169904;
		specparam tremoval_XS_C_adacond4_posedge_adacond4_posedge = 0.0981422:0.121541:0.0674361;
		specparam tsetup_XS_XR_posedge_posedge = 0.0525702:0.0720198:0.224423;
		specparam thold_XS_XR_posedge_posedge = 0.0192698:0.00617576:-0.0760674;
		specparam tpw_XS_negedge = 0.276401:0.39113:2.72095;
		specparam tpw_C_posedge = 0.291302:0.330811:2.72095;
		specparam tpw_C_negedge = 0.291302:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$recovery (posedge XS &&& adacond4, posedge C &&& adacond4, 
			 trecovery_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$hold (posedge C &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: SDFFSRQX 
`timescale 1ns/10ps
`celldefine
module SDFFSRQXXL (Q, XQ, D, SIN, SMC, XR, XS, C);
	output Q, XQ;
	input D, SIN, SMC, XR, XS, C;
	reg notifier;
	wire delayed_D, delayed_SIN, delayed_SMC, delayed_XR, delayed_XS, delayed_C;

	// Function
	wire delayed_SMC__bar, int_fwire_0, int_fwire_1;
	wire int_fwire_d, int_fwire_IQ, int_fwire_IXQ;
	wire int_fwire_r, int_fwire_s, xcr_0;

	and (int_fwire_0, delayed_SIN, delayed_SMC);
	not (delayed_SMC__bar, delayed_SMC);
	and (int_fwire_1, delayed_D, delayed_SMC__bar);
	or (int_fwire_d, int_fwire_1, int_fwire_0);
	not (int_fwire_s, delayed_XS);
	not (int_fwire_r, delayed_XR);
	altos_dff_sr_err (xcr_0, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r);
	altos_dff_sr_0 (int_fwire_IQ, notifier, delayed_C, int_fwire_d, int_fwire_s, int_fwire_r, xcr_0);
	buf (Q, int_fwire_IQ);
	nor (int_fwire_IXQ, int_fwire_IQ, int_fwire_s);
	buf (XQ, int_fwire_IXQ);

	// Timing

	// Additional timing wires
	wire adacond0, adacond1, adacond2;
	wire adacond3, adacond4, D__bar;
	wire int_twire_0, int_twire_1, int_twire_2;
	wire int_twire_3, int_twire_4, int_twire_5;
	wire SIN__bar, SMC__bar;


	// Additional timing gates
	not (SMC__bar, SMC);
	and (adacond0, SMC__bar, XR, XS);
	and (adacond1, SMC, XR, XS);
	not (D__bar, D);
	and (int_twire_0, D__bar, SIN, XR, XS);
	not (SIN__bar, SIN);
	and (int_twire_1, D, SIN__bar, XR, XS);
	or (adacond2, int_twire_1, int_twire_0);
	and (int_twire_2, SMC__bar, D, XS);
	and (int_twire_3, SMC, SIN, XS);
	or (adacond3, int_twire_3, int_twire_2);
	and (int_twire_4, SMC__bar, D__bar, XR);
	and (int_twire_5, SMC, SIN__bar, XR);
	or (adacond4, int_twire_5, int_twire_4);

	specify
		specparam tpd_XR_Q_negedge_r = 0.125006:0.248393:1.43698;
		specparam tpd_XR_Q_negedge_f = 0.115034:0.250858:1.24009;
		specparam tpd_XS_Q_negedge_r = 0.340401:0.501276:1.95496;
		specparam tpd_XS_Q_negedge_f = 0.340401:0.501276:1.95496;
		specparam tpd_C_Q_posedge_r = 0.348156:0.486057:1.59466;
		specparam tpd_C_Q_posedge_f = 0.347251:0.460877:1.11549;
		specparam tpd_XR_XQ_negedge_r = 0.259967:0.435369:1.85638;
		specparam tpd_XR_XQ_negedge_f = 0.259967:0.435369:1.85638;
		specparam tpd_XS_XQ_negedge_r = 0.152662:0.300556:1.55367;
		specparam tpd_XS_XQ_negedge_f = 0.135239:0.279251:1.3142;
		specparam tpd_C_XQ_posedge_r = 0.451355:0.582121:1.68066;
		specparam tpd_C_XQ_posedge_f = 0.428681:0.533934:1.17328;
		specparam tsetup_D_C_adacond0_posedge_adacond0_posedge = 0.249846:0.245889:0.4691;
		specparam thold_D_C_adacond0_posedge_adacond0_posedge = -0.146662:-0.1784:-0.389691;
		specparam tsetup_D_C_adacond0_negedge_adacond0_posedge = 0.249846:0.245889:0.4691;
		specparam thold_D_C_adacond0_negedge_adacond0_posedge = -0.146662:-0.1784:-0.389691;
		specparam tsetup_SIN_C_adacond1_posedge_adacond1_posedge = 0.250324:0.254615:0.497995;
		specparam thold_SIN_C_adacond1_posedge_adacond1_posedge = -0.150169:-0.183765:-0.417152;
		specparam tsetup_SIN_C_adacond1_negedge_adacond1_posedge = 0.250324:0.254615:0.497995;
		specparam thold_SIN_C_adacond1_negedge_adacond1_posedge = -0.150169:-0.183765:-0.417152;
		specparam tsetup_SMC_C_adacond2_posedge_adacond2_posedge = 0.406091:0.391346:0.47377;
		specparam thold_SMC_C_adacond2_posedge_adacond2_posedge = -0.127034:-0.170697:-0.231271;
		specparam tsetup_SMC_C_adacond2_negedge_adacond2_posedge = 0.406091:0.391346:0.47377;
		specparam thold_SMC_C_adacond2_negedge_adacond2_posedge = -0.127034:-0.170697:-0.231271;
		specparam trecovery_XR_C_adacond3_posedge_adacond3_posedge = -0.193319:-0.235239:0.225342;
		specparam tremoval_XR_C_adacond3_posedge_adacond3_posedge = 0.271853:0.361124:0.734361;
		specparam tpw_XR_negedge = 0.339738:0.425224:2.72095;
		specparam tsetup_XR_XS_posedge_posedge = 0.0197138:0.0084736:-0.00682191;
		specparam thold_XR_XS_posedge_posedge = 0.052432:0.0746485:0.137461;
		specparam trecovery_XS_C_adacond4_posedge_adacond4_posedge = -0.035112:-0.053727:0.17358;
		specparam tremoval_XS_C_adacond4_posedge_adacond4_posedge = 0.126739:0.150661:0.0609613;
		specparam tsetup_XS_XR_posedge_posedge = 0.0561484:0.0872597:0.222765;
		specparam thold_XS_XR_posedge_posedge = 0.018753:0.00732426:-0.0750148;
		specparam tpw_XS_negedge = 0.204715:0.330811:2.72095;
		specparam tpw_C_posedge = 0.182226:0.330811:2.72095;
		specparam tpw_C_negedge = 0.182226:0.330811:2.72095;

		(negedge XR => (Q+:1'b0)) = ( tpd_XR_Q_negedge_r , tpd_XR_Q_negedge_f );
		(negedge XS => (Q+:1'b1)) = ( tpd_XS_Q_negedge_r , tpd_XS_Q_negedge_f );
		(posedge C => (Q+:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_Q_posedge_r , tpd_C_Q_posedge_f );
		(negedge XR => (XQ-:1'b0)) = ( tpd_XR_XQ_negedge_r , tpd_XR_XQ_negedge_f );
		(negedge XS => (XQ-:1'b1)) = ( tpd_XS_XQ_negedge_r , tpd_XS_XQ_negedge_f );
		(posedge C => (XQ-:((D && SIN) || (D && !SIN && !SMC) || (!D && SIN && SMC)))) = ( tpd_C_XQ_posedge_r , tpd_C_XQ_posedge_f );
		$setuphold (posedge C &&& adacond0, posedge D &&& adacond0, 
			 tsetup_D_C_adacond0_posedge_adacond0_posedge, 
			 thold_D_C_adacond0_posedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond0, negedge D &&& adacond0, 
			 tsetup_D_C_adacond0_negedge_adacond0_posedge, 
			 thold_D_C_adacond0_negedge_adacond0_posedge, notifier,,, delayed_C, delayed_D);
		$setuphold (posedge C &&& adacond1, posedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_posedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_posedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond1, negedge SIN &&& adacond1, 
			 tsetup_SIN_C_adacond1_negedge_adacond1_posedge, 
			 thold_SIN_C_adacond1_negedge_adacond1_posedge, notifier,,, delayed_C, delayed_SIN);
		$setuphold (posedge C &&& adacond2, posedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_posedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_posedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge C &&& adacond2, negedge SMC &&& adacond2, 
			 tsetup_SMC_C_adacond2_negedge_adacond2_posedge, 
			 thold_SMC_C_adacond2_negedge_adacond2_posedge, notifier,,, delayed_C, delayed_SMC);
		$setuphold (posedge XS, posedge XR, 
			 tsetup_XR_XS_posedge_posedge, 
			 thold_XR_XS_posedge_posedge, notifier,,, delayed_XS, delayed_XR);
		$setuphold (posedge XR, posedge XS, 
			 tsetup_XS_XR_posedge_posedge, 
			 thold_XS_XR_posedge_posedge, notifier,,, delayed_XR, delayed_XS);
		$recovery (posedge XR &&& adacond3, posedge C &&& adacond3, 
			 trecovery_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$hold (posedge C &&& adacond3, posedge XR &&& adacond3, 
			 tremoval_XR_C_adacond3_posedge_adacond3_posedge, notifier);
		$recovery (posedge XS &&& adacond4, posedge C &&& adacond4, 
			 trecovery_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$hold (posedge C &&& adacond4, posedge XS &&& adacond4, 
			 tremoval_XS_C_adacond4_posedge_adacond4_posedge, notifier);
		$width (negedge XR, tpw_XR_negedge, 0, notifier);
		$width (negedge XS, tpw_XS_negedge, 0, notifier);
		$width (posedge C, tpw_C_posedge, 0, notifier);
		$width (negedge C, tpw_C_negedge, 0, notifier);
	endspecify
endmodule
`endcelldefine

// type: TBUF 
`timescale 1ns/10ps
`celldefine
module TBUFX1 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	bufif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.111744:0.213586:1.08195;
		specparam tpd_A_Y_f = 0.111713:0.214117:1.00576;
		specparam tpd_EN_Y_r = 0.0499162:0.126111:1.03899;
		specparam tpd_EN_Y_f = 0.0584156:0.126116:1.03899;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TBUF 
`timescale 1ns/10ps
`celldefine
module TBUFX12 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	bufif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.098575:0.244736:1.42347;
		specparam tpd_A_Y_f = 0.127243:0.292763:1.71715;
		specparam tpd_EN_Y_r = 0.169084:0.233645:0.448088;
		specparam tpd_EN_Y_f = 0.190076:0.271317:0.714094;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TBUF 
`timescale 1ns/10ps
`celldefine
module TBUFX2 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	bufif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0741837:0.200253:1.34469;
		specparam tpd_A_Y_f = 0.0950206:0.253478:1.66222;
		specparam tpd_EN_Y_r = 0.1303:0.184449:0.349381;
		specparam tpd_EN_Y_f = 0.113557:0.192554:0.546781;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TBUF 
`timescale 1ns/10ps
`celldefine
module TBUFX4 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	bufif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.091254:0.232141:1.41318;
		specparam tpd_A_Y_f = 0.110429:0.272806:1.67869;
		specparam tpd_EN_Y_r = 0.14101:0.196316:0.362256;
		specparam tpd_EN_Y_f = 0.152589:0.233101:0.628946;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TBUF 
`timescale 1ns/10ps
`celldefine
module TBUFX8 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	bufif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0838202:0.21876:1.36931;
		specparam tpd_A_Y_f = 0.107682:0.27017:1.68546;
		specparam tpd_EN_Y_r = 0.157662:0.221418:0.434055;
		specparam tpd_EN_Y_f = 0.149063:0.230104:0.634422;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TBUF 
`timescale 1ns/10ps
`celldefine
module TBUFXL (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	bufif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.140311:0.22568:0.892237;
		specparam tpd_A_Y_f = 0.159727:0.274193:1.14494;
		specparam tpd_EN_Y_r = 0.0681574:0.136737:1.03896;
		specparam tpd_EN_Y_f = 0.0795204:0.152575:1.03895;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TIEH 
`timescale 1ns/10ps
`celldefine
module TIEH (HI);
	output HI;

	// Function
	buf (HI, 1'b1);

	// Timing
	specify

	endspecify
endmodule
`endcelldefine

// type: TIEL 
`timescale 1ns/10ps
`celldefine
module TIEL (LO);
	output LO;

	// Function
	buf (LO, 1'b0);

	// Timing
	specify

	endspecify
endmodule
`endcelldefine

// type: TINV 
`timescale 1ns/10ps
`celldefine
module TINVX1 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	notif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0698518:0.192424:1.47381;
		specparam tpd_A_Y_f = 0.0738098:0.18506:1.34784;
		specparam tpd_EN_Y_r = 0.0527733:0.1261:1.03899;
		specparam tpd_EN_Y_f = 0.062198:0.1261:1.03898;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TINV 
`timescale 1ns/10ps
`celldefine
module TINVX12 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	notif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.221186:0.391384:1.7541;
		specparam tpd_A_Y_f = 0.232659:0.388947:1.62737;
		specparam tpd_EN_Y_r = 0.175746:0.240198:0.453946;
		specparam tpd_EN_Y_f = 0.190621:0.271395:0.707564;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TINV 
`timescale 1ns/10ps
`celldefine
module TINVX2 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	notif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.146927:0.294954:1.57266;
		specparam tpd_A_Y_f = 0.170326:0.330089:1.62835;
		specparam tpd_EN_Y_r = 0.132779:0.187582:0.352366;
		specparam tpd_EN_Y_f = 0.112834:0.191669:0.542884;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TINV 
`timescale 1ns/10ps
`celldefine
module TINVX4 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	notif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.165109:0.320105:1.60161;
		specparam tpd_A_Y_f = 0.186453:0.343531:1.60337;
		specparam tpd_EN_Y_r = 0.144235:0.198374:0.365417;
		specparam tpd_EN_Y_f = 0.152651:0.233034:0.630381;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TINV 
`timescale 1ns/10ps
`celldefine
module TINVX8 (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	notif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.203595:0.367595:1.72768;
		specparam tpd_A_Y_f = 0.213795:0.371318:1.62274;
		specparam tpd_EN_Y_r = 0.163847:0.22827:0.44006;
		specparam tpd_EN_Y_f = 0.151311:0.230517:0.628853;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: TINV 
`timescale 1ns/10ps
`celldefine
module TINVXL (Y, A, EN);
	output Y;
	input A, EN;

	// Function
	notif1 (Y, A, EN);

	// Timing
	specify
		specparam tpd_A_Y_r = 0.0843509:0.214261:1.53487;
		specparam tpd_A_Y_f = 0.0696099:0.15695:1.04061;
		specparam tpd_EN_Y_r = 0.0719439:0.142461:1.03896;
		specparam tpd_EN_Y_f = 0.0841645:0.158992:1.03896;

		(A => Y) = ( tpd_A_Y_r , tpd_A_Y_f );
		(EN => Y) = ( tpd_EN_Y_r , tpd_EN_Y_f );
	endspecify
endmodule
`endcelldefine

// type: XNOR2 
`timescale 1ns/10ps
`celldefine
module XNOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.102241:0.181796:0.692644;
		specparam tpd_A_Y_posedge_f = 0.136114:0.242077:1.03125;
		specparam tpd_A_Y_negedge_r = 0.097558:0.232457:1.77441;
		specparam tpd_A_Y_negedge_f = 0.0546693:0.123806:0.895759;
		specparam tpd_B_Y_posedge_r = 0.110429:0.18358:0.675613;
		specparam tpd_B_Y_posedge_f = 0.136671:0.250281:1.06076;
		specparam tpd_B_Y_negedge_r = 0.122557:0.239684:1.60201;
		specparam tpd_B_Y_negedge_f = 0.0689522:0.146957:0.953125;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XNOR2 
`timescale 1ns/10ps
`celldefine
module XNOR2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.172604:0.330865:1.65085;
		specparam tpd_A_Y_posedge_f = 0.211714:0.381118:1.7941;
		specparam tpd_A_Y_negedge_r = 0.198782:0.348317:1.68715;
		specparam tpd_A_Y_negedge_f = 0.258194:0.421133:1.65867;
		specparam tpd_B_Y_posedge_r = 0.182877:0.327659:1.59368;
		specparam tpd_B_Y_posedge_f = 0.226958:0.401176:1.84033;
		specparam tpd_B_Y_negedge_r = 0.222175:0.357229:1.61924;
		specparam tpd_B_Y_negedge_f = 0.272123:0.442946:1.76367;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XNOR2 
`timescale 1ns/10ps
`celldefine
module XNOR2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.239656:0.406194:1.79254;
		specparam tpd_A_Y_posedge_f = 0.280767:0.436454:1.52663;
		specparam tpd_A_Y_negedge_r = 0.253126:0.413941:1.80494;
		specparam tpd_A_Y_negedge_f = 0.300337:0.44602:1.24843;
		specparam tpd_B_Y_posedge_r = 0.249643:0.403172:1.71832;
		specparam tpd_B_Y_posedge_f = 0.296545:0.456462:1.57189;
		specparam tpd_B_Y_negedge_r = 0.277099:0.4204:1.74229;
		specparam tpd_B_Y_negedge_f = 0.30277:0.456307:1.33003;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XNOR2 
`timescale 1ns/10ps
`celldefine
module XNOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar);
	and (int_fwire_1, A, B);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.12872:0.206588:0.684138;
		specparam tpd_A_Y_posedge_f = 0.185146:0.302069:1.24633;
		specparam tpd_A_Y_negedge_r = 0.114011:0.250519:1.82875;
		specparam tpd_A_Y_negedge_f = 0.0795691:0.151941:1.01863;
		specparam tpd_B_Y_posedge_r = 0.136745:0.203161:0.638015;
		specparam tpd_B_Y_posedge_f = 0.186386:0.313161:1.35662;
		specparam tpd_B_Y_negedge_r = 0.144145:0.266752:1.67927;
		specparam tpd_B_Y_negedge_f = 0.0921865:0.159736:0.923737;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XNOR3 
`timescale 1ns/10ps
`celldefine
module XNOR3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C__bar);
	and (int_fwire_1, A__bar, B, C);
	and (int_fwire_2, A, B__bar, C);
	and (int_fwire_3, A, B, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.122337:0.273554:1.44985;
		specparam tpd_A_Y_posedge_f = 0.169384:0.3702:1.87842;
		specparam tpd_A_Y_negedge_r = 0.162603:0.332596:1.63971;
		specparam tpd_A_Y_negedge_f = 0.23603:0.391016:1.54759;
		specparam tpd_B_Y_posedge_r = 0.254138:0.416868:1.74273;
		specparam tpd_B_Y_posedge_f = 0.387877:0.583231:2.06172;
		specparam tpd_B_Y_negedge_r = 0.364339:0.512441:1.87934;
		specparam tpd_B_Y_negedge_f = 0.398142:0.578962:1.72531;
		specparam tpd_C_Y_posedge_r = 0.385224:0.535657:1.75776;
		specparam tpd_C_Y_posedge_f = 0.398691:0.595518:2.08267;
		specparam tpd_C_Y_negedge_r = 0.377447:0.527462:1.91445;
		specparam tpd_C_Y_negedge_f = 0.409187:0.605402:1.85726;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
		(posedge C => (Y:C)) = ( tpd_C_Y_posedge_r , tpd_C_Y_posedge_f );
		(negedge C => (Y:C)) = ( tpd_C_Y_negedge_r , tpd_C_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XNOR3 
`timescale 1ns/10ps
`celldefine
module XNOR3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C__bar);
	and (int_fwire_1, A__bar, B, C);
	and (int_fwire_2, A, B__bar, C);
	and (int_fwire_3, A, B, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.1746:0.34342:1.6478;
		specparam tpd_A_Y_posedge_f = 0.199982:0.395827:1.72716;
		specparam tpd_A_Y_negedge_r = 0.203224:0.388492:1.73716;
		specparam tpd_A_Y_negedge_f = 0.229512:0.373734:1.32316;
		specparam tpd_B_Y_posedge_r = 0.324532:0.499204:1.91662;
		specparam tpd_B_Y_posedge_f = 0.423204:0.613037:1.90614;
		specparam tpd_B_Y_negedge_r = 0.430915:0.593642:1.97248;
		specparam tpd_B_Y_negedge_f = 0.42994:0.604834:1.56455;
		specparam tpd_C_Y_posedge_r = 0.332068:0.494015:1.83952;
		specparam tpd_C_Y_posedge_f = 0.430809:0.621155:1.92039;
		specparam tpd_C_Y_negedge_r = 0.441164:0.605311:2.0031;
		specparam tpd_C_Y_negedge_f = 0.441558:0.6296:1.67885;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
		(posedge C => (Y:C)) = ( tpd_C_Y_posedge_r , tpd_C_Y_posedge_f );
		(negedge C => (Y:C)) = ( tpd_C_Y_negedge_r , tpd_C_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XNOR3 
`timescale 1ns/10ps
`celldefine
module XNOR3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C__bar);
	and (int_fwire_1, A__bar, B, C);
	and (int_fwire_2, A, B__bar, C);
	and (int_fwire_3, A, B, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.175794:0.34899:1.64613;
		specparam tpd_A_Y_posedge_f = 0.275753:0.490455:1.95597;
		specparam tpd_A_Y_negedge_r = 0.236609:0.43295:1.79453;
		specparam tpd_A_Y_negedge_f = 0.282255:0.444015:1.48971;
		specparam tpd_B_Y_posedge_r = 0.362346:0.547515:1.99447;
		specparam tpd_B_Y_posedge_f = 0.504478:0.713136:2.13058;
		specparam tpd_B_Y_negedge_r = 0.427811:0.594392:1.97268;
		specparam tpd_B_Y_negedge_f = 0.509796:0.702694:1.76925;
		specparam tpd_C_Y_posedge_r = 0.369887:0.542378:1.91082;
		specparam tpd_C_Y_posedge_f = 0.511556:0.720655:2.14285;
		specparam tpd_C_Y_negedge_r = 0.438281:0.606249:2.00416;
		specparam tpd_C_Y_negedge_f = 0.519236:0.723952:1.86308;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
		(posedge C => (Y:C)) = ( tpd_C_Y_posedge_r , tpd_C_Y_posedge_f );
		(negedge C => (Y:C)) = ( tpd_C_Y_negedge_r , tpd_C_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XNOR3 
`timescale 1ns/10ps
`celldefine
module XNOR3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (C__bar, C);
	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C__bar);
	and (int_fwire_1, A__bar, B, C);
	and (int_fwire_2, A, B__bar, C);
	and (int_fwire_3, A, B, C__bar);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.162477:0.313897:1.47814;
		specparam tpd_A_Y_posedge_f = 0.184069:0.408047:2.12292;
		specparam tpd_A_Y_negedge_r = 0.176337:0.360174:1.69956;
		specparam tpd_A_Y_negedge_f = 0.312223:0.481447:1.76543;
		specparam tpd_B_Y_posedge_r = 0.350653:0.516292:1.85163;
		specparam tpd_B_Y_posedge_f = 0.515657:0.739076:2.45174;
		specparam tpd_B_Y_negedge_r = 0.459666:0.61943:2.04367;
		specparam tpd_B_Y_negedge_f = 0.537283:0.737246:2.06981;
		specparam tpd_C_Y_posedge_r = 0.508968:0.657965:1.89987;
		specparam tpd_C_Y_posedge_f = 0.525977:0.751918:2.47669;
		specparam tpd_C_Y_negedge_r = 0.473322:0.635358:2.08433;
		specparam tpd_C_Y_negedge_f = 0.565574:0.776507:2.2207;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
		(posedge C => (Y:C)) = ( tpd_C_Y_posedge_r , tpd_C_Y_posedge_f );
		(negedge C => (Y:C)) = ( tpd_C_Y_negedge_r , tpd_C_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XOR2 
`timescale 1ns/10ps
`celldefine
module XOR2X1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, B);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.105101:0.217903:1.26522;
		specparam tpd_A_Y_posedge_f = 0.128615:0.246231:1.15662;
		specparam tpd_A_Y_negedge_r = 0.0840643:0.207142:1.61407;
		specparam tpd_A_Y_negedge_f = 0.0920741:0.220949:1.70514;
		specparam tpd_B_Y_posedge_r = 0.112652:0.23916:1.37299;
		specparam tpd_B_Y_posedge_f = 0.150611:0.252163:1.10254;
		specparam tpd_B_Y_negedge_r = 0.092001:0.21445:1.60036;
		specparam tpd_B_Y_negedge_f = 0.101106:0.218077:1.60466;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XOR2 
`timescale 1ns/10ps
`celldefine
module XOR2X2 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, B);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.144023:0.278867:1.46272;
		specparam tpd_A_Y_posedge_f = 0.208249:0.38617:1.81844;
		specparam tpd_A_Y_negedge_r = 0.227756:0.394882:1.76115;
		specparam tpd_A_Y_negedge_f = 0.189805:0.324637:1.40682;
		specparam tpd_B_Y_posedge_r = 0.170965:0.313414:1.55855;
		specparam tpd_B_Y_posedge_f = 0.233266:0.395805:1.71916;
		specparam tpd_B_Y_negedge_r = 0.220756:0.389215:1.79437;
		specparam tpd_B_Y_negedge_f = 0.198826:0.324325:1.37262;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XOR2 
`timescale 1ns/10ps
`celldefine
module XOR2X4 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, B);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.183199:0.329772:1.55588;
		specparam tpd_A_Y_posedge_f = 0.27046:0.450096:1.82031;
		specparam tpd_A_Y_negedge_r = 0.266906:0.443938:1.81617;
		specparam tpd_A_Y_negedge_f = 0.220569:0.357138:1.32117;
		specparam tpd_B_Y_posedge_r = 0.211391:0.363792:1.64664;
		specparam tpd_B_Y_posedge_f = 0.295347:0.460698:1.70079;
		specparam tpd_B_Y_negedge_r = 0.260776:0.438087:1.848;
		specparam tpd_B_Y_negedge_f = 0.229875:0.357037:1.28898;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XOR2 
`timescale 1ns/10ps
`celldefine
module XOR2XL (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire A__bar, B__bar, int_fwire_0;
	wire int_fwire_1;

	not (A__bar, A);
	and (int_fwire_0, A__bar, B);
	not (B__bar, B);
	and (int_fwire_1, A, B__bar);
	or (Y, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.169205:0.275861:1.35813;
		specparam tpd_A_Y_posedge_f = 0.123851:0.220312:0.911603;
		specparam tpd_A_Y_negedge_r = 0.128776:0.260063:1.74236;
		specparam tpd_A_Y_negedge_f = 0.0779022:0.167997:1.113;
		specparam tpd_B_Y_posedge_r = 0.174399:0.291937:1.44442;
		specparam tpd_B_Y_posedge_f = 0.147354:0.229952:0.861748;
		specparam tpd_B_Y_negedge_r = 0.145764:0.277145:1.74701;
		specparam tpd_B_Y_negedge_f = 0.0873134:0.15881:0.966507;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XOR3 
`timescale 1ns/10ps
`celldefine
module XOR3X1 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C);
	not (C__bar, C);
	and (int_fwire_1, A__bar, B, C__bar);
	and (int_fwire_2, A, B__bar, C__bar);
	and (int_fwire_3, A, B, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.122606:0.282184:1.53562;
		specparam tpd_A_Y_posedge_f = 0.16467:0.339491:1.76622;
		specparam tpd_A_Y_negedge_r = 0.186923:0.340038:1.64835;
		specparam tpd_A_Y_negedge_f = 0.170709:0.368055:1.55949;
		specparam tpd_B_Y_posedge_r = 0.277523:0.442469:1.80939;
		specparam tpd_B_Y_posedge_f = 0.369035:0.561811:2.00053;
		specparam tpd_B_Y_negedge_r = 0.352234:0.49952:1.84297;
		specparam tpd_B_Y_negedge_f = 0.343379:0.505351:1.71005;
		specparam tpd_C_Y_posedge_r = 0.28648:0.438543:1.73949;
		specparam tpd_C_Y_posedge_f = 0.379505:0.573342:2.02179;
		specparam tpd_C_Y_negedge_r = 0.364564:0.513393:1.87945;
		specparam tpd_C_Y_negedge_f = 0.388955:0.580955:1.80014;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
		(posedge C => (Y:C)) = ( tpd_C_Y_posedge_r , tpd_C_Y_posedge_f );
		(negedge C => (Y:C)) = ( tpd_C_Y_negedge_r , tpd_C_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XOR3 
`timescale 1ns/10ps
`celldefine
module XOR3X2 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C);
	not (C__bar, C);
	and (int_fwire_1, A__bar, B, C__bar);
	and (int_fwire_2, A, B__bar, C__bar);
	and (int_fwire_3, A, B, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.142235:0.311571:1.59569;
		specparam tpd_A_Y_posedge_f = 0.19839:0.382495:1.85462;
		specparam tpd_A_Y_negedge_r = 0.202666:0.362638:1.66619;
		specparam tpd_A_Y_negedge_f = 0.203572:0.412479:1.63688;
		specparam tpd_B_Y_posedge_r = 0.2983:0.469892:1.85033;
		specparam tpd_B_Y_posedge_f = 0.411159:0.612804:2.08236;
		specparam tpd_B_Y_negedge_r = 0.37014:0.52393:1.86325;
		specparam tpd_B_Y_negedge_f = 0.37718:0.548449:1.76751;
		specparam tpd_C_Y_posedge_r = 0.307256:0.466097:1.77628;
		specparam tpd_C_Y_posedge_f = 0.421158:0.623645:2.10142;
		specparam tpd_C_Y_negedge_r = 0.382614:0.537869:1.89925;
		specparam tpd_C_Y_negedge_f = 0.429651:0.630142:1.86696;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
		(posedge C => (Y:C)) = ( tpd_C_Y_posedge_r , tpd_C_Y_posedge_f );
		(negedge C => (Y:C)) = ( tpd_C_Y_negedge_r , tpd_C_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XOR3 
`timescale 1ns/10ps
`celldefine
module XOR3X4 (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C);
	not (C__bar, C);
	and (int_fwire_1, A__bar, B, C__bar);
	and (int_fwire_2, A, B__bar, C__bar);
	and (int_fwire_3, A, B, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.191465:0.369873:1.72246;
		specparam tpd_A_Y_posedge_f = 0.258724:0.440175:1.78006;
		specparam tpd_A_Y_negedge_r = 0.241922:0.412427:1.7326;
		specparam tpd_A_Y_negedge_f = 0.264883:0.469604:1.55667;
		specparam tpd_B_Y_posedge_r = 0.347554:0.527692:1.95436;
		specparam tpd_B_Y_posedge_f = 0.479509:0.678702:2.00559;
		specparam tpd_B_Y_negedge_r = 0.412794:0.576123:1.93469;
		specparam tpd_B_Y_negedge_f = 0.486911:0.669479:1.64734;
		specparam tpd_C_Y_posedge_r = 0.356552:0.523825:1.87298;
		specparam tpd_C_Y_posedge_f = 0.488912:0.688413:2.02087;
		specparam tpd_C_Y_negedge_r = 0.425539:0.590305:1.97016;
		specparam tpd_C_Y_negedge_f = 0.493976:0.688339:1.73859;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
		(posedge C => (Y:C)) = ( tpd_C_Y_posedge_r , tpd_C_Y_posedge_f );
		(negedge C => (Y:C)) = ( tpd_C_Y_negedge_r , tpd_C_Y_negedge_f );
	endspecify
endmodule
`endcelldefine

// type: XOR3 
`timescale 1ns/10ps
`celldefine
module XOR3XL (Y, A, B, C);
	output Y;
	input A, B, C;

	// Function
	wire A__bar, B__bar, C__bar;
	wire int_fwire_0, int_fwire_1, int_fwire_2;
	wire int_fwire_3;

	not (B__bar, B);
	not (A__bar, A);
	and (int_fwire_0, A__bar, B__bar, C);
	not (C__bar, C);
	and (int_fwire_1, A__bar, B, C__bar);
	and (int_fwire_2, A, B__bar, C__bar);
	and (int_fwire_3, A, B, C);
	or (Y, int_fwire_3, int_fwire_2, int_fwire_1, int_fwire_0);

	// Timing
	specify
		specparam tpd_A_Y_posedge_r = 0.1374:0.30513:1.51344;
		specparam tpd_A_Y_posedge_f = 0.249269:0.44973:2.18015;
		specparam tpd_A_Y_negedge_r = 0.232917:0.395459:1.72783;
		specparam tpd_A_Y_negedge_f = 0.203154:0.429605:1.81765;
		specparam tpd_B_Y_posedge_r = 0.348615:0.515109:1.85852;
		specparam tpd_B_Y_posedge_f = 0.515176:0.739369:2.45977;
		specparam tpd_B_Y_negedge_r = 0.459046:0.619377:2.05144;
		specparam tpd_B_Y_negedge_f = 0.536957:0.737698:2.07831;
		specparam tpd_C_Y_posedge_r = 0.508338:0.657908:1.908;
		specparam tpd_C_Y_posedge_f = 0.525658:0.75242:2.48433;
		specparam tpd_C_Y_negedge_r = 0.472701:0.635307:2.09249;
		specparam tpd_C_Y_negedge_f = 0.565101:0.776768:2.22921;

		(posedge A => (Y:A)) = ( tpd_A_Y_posedge_r , tpd_A_Y_posedge_f );
		(negedge A => (Y:A)) = ( tpd_A_Y_negedge_r , tpd_A_Y_negedge_f );
		(posedge B => (Y:B)) = ( tpd_B_Y_posedge_r , tpd_B_Y_posedge_f );
		(negedge B => (Y:B)) = ( tpd_B_Y_negedge_r , tpd_B_Y_negedge_f );
		(posedge C => (Y:C)) = ( tpd_C_Y_posedge_r , tpd_C_Y_posedge_f );
		(negedge C => (Y:C)) = ( tpd_C_Y_negedge_r , tpd_C_Y_negedge_f );
	endspecify
endmodule
`endcelldefine


`ifdef _udp_def_altos_latch_
`else
`define _udp_def_altos_latch_
primitive altos_latch (q, v, clk, d);
	output q;
	reg q;
	input v, clk, d;

	table
		* ? ? : ? : x;
		? 1 0 : ? : 0;
		? 1 1 : ? : 1;
		? x 0 : 0 : -;
		? x 1 : 1 : -;
		? 0 ? : ? : -;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_err_
`else
`define _udp_def_altos_dff_err_
primitive altos_dff_err (q, clk, d);
	output q;
	reg q;
	input clk, d;

	table
		(0x) ? : ? : 0;
		(1x) ? : ? : 1;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_
`else
`define _udp_def_altos_dff_
primitive altos_dff (q, v, clk, d, xcr);
	output q;
	reg q;
	input v, clk, d, xcr;

	table
		*  ?   ? ? : ? : x;
		? (x1) 0 0 : ? : 0;
		? (x1) 1 0 : ? : 1;
		? (x1) 0 1 : 0 : 0;
		? (x1) 1 1 : 1 : 1;
		? (x1) ? x : ? : -;
		? (bx) 0 ? : 0 : -;
		? (bx) 1 ? : 1 : -;
		? (x0) b ? : ? : -;
		? (x0) ? x : ? : -;
		? (01) 0 ? : ? : 0;
		? (01) 1 ? : ? : 1;
		? (10) ? ? : ? : -;
		?  b   * ? : ? : -;
		?  ?   ? * : ? : -;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_r_err_
`else
`define _udp_def_altos_dff_r_err_
primitive altos_dff_r_err (q, clk, d, r);
	output q;
	reg q;
	input clk, d, r;

	table
		 ?   0 (0x) : ? : -;
		 ?   0 (x0) : ? : -;
		(0x) ?  0   : ? : 0;
		(0x) 0  x   : ? : 0;
		(1x) ?  0   : ? : 1;
		(1x) 0  x   : ? : 1;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_r_
`else
`define _udp_def_altos_dff_r_
primitive altos_dff_r (q, v, clk, d, r, xcr);
	output q;
	reg q;
	input v, clk, d, r, xcr;

	table
		*  ?   ?  ?   ? : ? : x;
		?  ?   ?  1   ? : ? : 0;
		?  b   ? (1?) ? : 0 : -;
		?  x   0 (1?) ? : 0 : -;
		?  ?   ? (10) ? : ? : -;
		?  ?   ? (x0) ? : ? : -;
		?  ?   ? (0x) ? : 0 : -;
		? (x1) 0  ?   0 : ? : 0;
		? (x1) 1  0   0 : ? : 1;
		? (x1) 0  ?   1 : 0 : 0;
		? (x1) 1  0   1 : 1 : 1;
		? (x1) ?  ?   x : ? : -;
		? (bx) 0  ?   ? : 0 : -;
		? (bx) 1  0   ? : 1 : -;
		? (x0) 0  ?   ? : ? : -;
		? (x0) 1  0   ? : ? : -;
		? (x0) ?  0   x : ? : -;
		? (01) 0  ?   ? : ? : 0;
		? (01) 1  0   ? : ? : 1;
		? (10) ?  ?   ? : ? : -;
		?  b   *  ?   ? : ? : -;
		?  ?   ?  ?   * : ? : -;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_s_err_
`else
`define _udp_def_altos_dff_s_err_
primitive altos_dff_s_err (q, clk, d, s);
	output q;
	reg q;
	input clk, d, s;

	table
		 ?   1 (0x) : ? : -;
		 ?   1 (x0) : ? : -;
		(0x) ?  0   : ? : 0;
		(0x) 1  x   : ? : 0;
		(1x) ?  0   : ? : 1;
		(1x) 1  x   : ? : 1;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_s_
`else
`define _udp_def_altos_dff_s_
primitive altos_dff_s (q, v, clk, d, s, xcr);
	output q;
	reg q;
	input v, clk, d, s, xcr;

	table
		*  ?   ?  ?   ? : ? : x;
		?  ?   ?  1   ? : ? : 1;
		?  b   ? (1?) ? : 1 : -;
		?  x   1 (1?) ? : 1 : -;
		?  ?   ? (10) ? : ? : -;
		?  ?   ? (x0) ? : ? : -;
		?  ?   ? (0x) ? : 1 : -;
		? (x1) 0  0   0 : ? : 0;
		? (x1) 1  ?   0 : ? : 1;
		? (x1) 1  ?   1 : 1 : 1;
		? (x1) 0  0   1 : 0 : 0;
		? (x1) ?  ?   x : ? : -;
		? (bx) 1  ?   ? : 1 : -;
		? (bx) 0  0   ? : 0 : -;
		? (x0) 1  ?   ? : ? : -;
		? (x0) 0  0   ? : ? : -;
		? (x0) ?  0   x : ? : -;
		? (01) 1  ?   ? : ? : 1;
		? (01) 0  0   ? : ? : 0;
		? (10) ?  ?   ? : ? : -;
		?  b   *  ?   ? : ? : -;
		?  ?   ?  ?   * : ? : -;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_sr_err_
`else
`define _udp_def_altos_dff_sr_err_
primitive altos_dff_sr_err (q, clk, d, s, r);
	output q;
	reg q;
	input clk, d, s, r;

	table
		 ?   1 (0x)  ?   : ? : -;
		 ?   0  ?   (0x) : ? : -;
		 ?   0  ?   (x0) : ? : -;
		(0x) ?  0    0   : ? : 0;
		(0x) 1  x    0   : ? : 0;
		(0x) 0  0    x   : ? : 0;
		(1x) ?  0    0   : ? : 1;
		(1x) 1  x    0   : ? : 1;
		(1x) 0  0    x   : ? : 1;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_sr_0
`else
`define _udp_def_altos_dff_sr_0
primitive altos_dff_sr_0 (q, v, clk, d, s, r, xcr);
	output q;
	reg q;
	input v, clk, d, s, r, xcr;

	table
	//	v,  clk, d, s, r : q' : q;

		*  ?   ?   ?   ?   ? : ? : x;
		?  ?   ?   ?   1   ? : ? : 0;
		?  ?   ?   1   0   ? : ? : 1;
		?  b   ? (1?)  0   ? : 1 : -;
		?  x   1 (1?)  0   ? : 1 : -;
		?  ?   ? (10)  0   ? : ? : -;
		?  ?   ? (x0)  0   ? : ? : -;
		?  ?   ? (0x)  0   ? : 1 : -;
		?  b   ?  0   (1?) ? : 0 : -;
		?  x   0  0   (1?) ? : 0 : -;
		?  ?   ?  0   (10) ? : ? : -;
		?  ?   ?  0   (x0) ? : ? : -;
		?  ?   ?  0   (0x) ? : 0 : -;
		? (x1) 0  0    ?   0 : ? : 0;
		? (x1) 1  ?    0   0 : ? : 1;
		? (x1) 0  0    ?   1 : 0 : 0;
		? (x1) 1  ?    0   1 : 1 : 1;
		? (x1) ?  ?    0   x : ? : -;
		? (x1) ?  0    ?   x : ? : -;
		? (1x) 0  0    ?   ? : 0 : -;
		? (1x) 1  ?    0   ? : 1 : -;
		? (x0) 0  0    ?   ? : ? : -;
		? (x0) 1  ?    0   ? : ? : -;
		? (x0) ?  0    0   x : ? : -;
		? (0x) 0  0    ?   ? : 0 : -;
		? (0x) 1  ?    0   ? : 1 : -;
		? (01) 0  0    ?   ? : ? : 0;
		? (01) 1  ?    0   ? : ? : 1;
		? (10) ?  0    ?   ? : ? : -;
		? (10) ?  ?    0   ? : ? : -;
		?  b   *  0    ?   ? : ? : -;
		?  b   *  ?    0   ? : ? : -;
		?  ?   ?  ?    ?   * : ? : -;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_dff_sr_1
`else
`define _udp_def_altos_dff_sr_1
primitive altos_dff_sr_1 (q, v, clk, d, s, r, xcr);
	output q;
	reg q;
	input v, clk, d, s, r, xcr;

	table
	//	v,  clk, d, s, r : q' : q;

		*  ?   ?   ?   ?   ? : ? : x;
		?  ?   ?   0   1   ? : ? : 0;
		?  ?   ?   1   ?   ? : ? : 1;
		?  b   ? (1?)  0   ? : 1 : -;
		?  x   1 (1?)  0   ? : 1 : -;
		?  ?   ? (10)  0   ? : ? : -;
		?  ?   ? (x0)  0   ? : ? : -;
		?  ?   ? (0x)  0   ? : 1 : -;
		?  b   ?  0   (1?) ? : 0 : -;
		?  x   0  0   (1?) ? : 0 : -;
		?  ?   ?  0   (10) ? : ? : -;
		?  ?   ?  0   (x0) ? : ? : -;
		?  ?   ?  0   (0x) ? : 0 : -;
		? (x1) 0  0    ?   0 : ? : 0;
		? (x1) 1  ?    0   0 : ? : 1;
		? (x1) 0  0    ?   1 : 0 : 0;
		? (x1) 1  ?    0   1 : 1 : 1;
		? (x1) ?  ?    0   x : ? : -;
		? (x1) ?  0    ?   x : ? : -;
		? (1x) 0  0    ?   ? : 0 : -;
		? (1x) 1  ?    0   ? : 1 : -;
		? (x0) 0  0    ?   ? : ? : -;
		? (x0) 1  ?    0   ? : ? : -;
		? (x0) ?  0    0   x : ? : -;
		? (0x) 0  0    ?   ? : 0 : -;
		? (0x) 1  ?    0   ? : 1 : -;
		? (01) 0  0    ?   ? : ? : 0;
		? (01) 1  ?    0   ? : ? : 1;
		? (10) ?  0    ?   ? : ? : -;
		? (10) ?  ?    0   ? : ? : -;
		?  b   *  0    ?   ? : ? : -;
		?  b   *  ?    0   ? : ? : -;
		?  ?   ?  ?    ?   * : ? : -;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_latch_r_
`else
`define _udp_def_altos_latch_r_
primitive altos_latch_r (q, v, clk, d, r);
	output q;
	reg q;
	input v, clk, d, r;

	table
		* ? ? ? : ? : x;
		? ? ? 1 : ? : 0;
		? 0 ? 0 : ? : -;
		? 0 ? x : 0 : -;
		? 1 0 0 : ? : 0;
		? 1 0 x : ? : 0;
		? 1 1 0 : ? : 1;
		? x 0 0 : 0 : -;
		? x 0 x : 0 : -;
		? x 1 0 : 1 : -;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_latch_s_
`else
`define _udp_def_altos_latch_s_
primitive altos_latch_s (q, v, clk, d, s);
	output q;
	reg q;
	input v, clk, d, s;

	table
		* ? ? ? : ? : x;
		? ? ? 1 : ? : 1;
		? 0 ? 0 : ? : -;
		? 0 ? x : 1 : -;
		? 1 1 0 : ? : 1;
		? 1 1 x : ? : 1;
		? 1 0 0 : ? : 0;
		? x 1 0 : 1 : -;
		? x 1 x : 1 : -;
		? x 0 0 : 0 : -;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_latch_sr_0
`else
`define _udp_def_altos_latch_sr_0
primitive altos_latch_sr_0 (q, v, clk, d, s, r);
	output q;
	reg q;
	input v, clk, d, s, r;

	table
		* ? ? ? ? : ? : x;
		? 1 1 ? 0 : ? : 1;
		? 1 0 0 ? : ? : 0;
		? ? ? 1 0 : ? : 1;
		? ? ? ? 1 : ? : 0;
		? 0 * ? ? : ? : -;
		? 0 ? * 0 : 1 : 1;
		? 0 ? 0 * : 0 : 0;
		? * 1 ? 0 : 1 : 1;
		? * 0 0 ? : 0 : 0;
		? ? 1 * 0 : 1 : 1;
		? ? 0 0 * : 0 : 0;
	endtable
endprimitive
`endif

`ifdef _udp_def_altos_latch_sr_1
`else
`define _udp_def_altos_latch_sr_1
primitive altos_latch_sr_1 (q, v, clk, d, s, r);
	output q;
	reg q;
	input v, clk, d, s, r;

	table
		* ? ? ? ? : ? : x;
		? 1 1 ? 0 : ? : 1;
		? 1 0 0 ? : ? : 0;
		? ? ? 1 ? : ? : 1;
		? ? ? 0 1 : ? : 0;
		? 0 * ? ? : ? : -;
		? 0 ? * 0 : 1 : 1;
		? 0 ? 0 * : 0 : 0;
		? * 1 ? 0 : 1 : 1;
		? * 0 0 ? : 0 : 0;
		? ? 1 * 0 : 1 : 1;
		? ? 0 0 * : 0 : 0;
	endtable
endprimitive
`endif
