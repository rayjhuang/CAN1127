
module chiptop_1127a0 ( CSP, CSN, VFB, COMP, SW, BST, VDRV, LG, HG, GATE, DP, 
        DN, CC1, CC2, TST, GPIO_TS, SCL, SDA, GPIO1, GPIO2, GPIO3, GPIO4, 
        GPIO5 );
  input TST;
  output LG, HG, GATE;
  inout CSP,  CSN,  VFB,  COMP,  SW,  BST,  VDRV,  DP,  DN,  CC1,  CC2, 
     GPIO_TS,  SCL,  SDA,  GPIO1,  GPIO2,  GPIO3,  GPIO4,  GPIO5;
  wire   SRAM_WEB, SRAM_CEB, SRAM_OEB, PWREN_HOLD, RD_ENB, STB_RP, DRP_OSC,
         IMP_OSC, TX_EN, TX_DAT, RX_DAT, RX_SQL, DAC1_EN, AD_RST, AD_HOLD,
         COMP_O, CCI2C_EN, RSTB, SLEEP, OSC_LOW, OSC_STOP, PWRDN, VPP_0V,
         VPP_SEL, LDO3P9V, OSC_O, RD_DET, OCP_SEL, CC1_DOB, CC2_DOB, CC1_DI,
         CC2_DI, DP_COMP, DN_COMP, DN_FAULT, LFOSC_ENB, VPP_OTP, IO_RSTB5,
         V1P1, ANAP_TS, TS_ANA_R, ANAP_GP1, GP1_ANA_R, ANAP_GP2, GP2_ANA_R,
         ANAP_GP3, GP3_ANA_R, ANAP_GP4, GP4_ANA_R, ANAP_GP5, GP5_ANA_R, DI_TST,
         DI_TS, SRAM_CLK, PMEM_RE, PMEM_PGM, PMEM_CSB, do_ccctl_0_,
         do_srcctl_0, tm_atpg, n1, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17;
  wire   [10:0] SRAM_A;
  wire   [7:0] SRAM_D;
  wire   [7:0] ANAOPT;
  wire   [1:0] FSW;
  wire   [1:0] RP_EN;
  wire   [1:0] VCONN_EN;
  wire   [17:0] SAMPL_SEL;
  wire   [4:0] DUMMY_IN;
  wire   [55:0] REGTRM;
  wire   [7:0] PWR_I;
  wire   [1:0] OVP_SEL;
  wire   [1:0] CC_SLOPE;
  wire   [5:0] DAC3_V;
  wire   [10:0] DAC0;
  wire   [3:0] ANA_TM;
  wire   [9:0] DAC1;
  wire   [1:0] RP_SEL;
  wire   [1:0] IE_GPIO;
  wire   [6:0] DI_GPIO;
  wire   [6:0] OE_GPIO;
  wire   [6:0] DO_GPIO;
  wire   [6:0] PU_GPIO;
  wire   [6:0] PD_GPIO;
  wire   [3:0] DO_TS;
  wire   [1:0] PMEM_CLK;
  wire   [7:0] PMEM_Q1;
  wire   [7:0] PMEM_Q0;
  wire   [1:0] PMEM_SAP;
  wire   [1:0] PMEM_TWLB;
  wire   [15:0] PMEM_A;
  wire   [7:0] bck_regx0;
  wire   [7:2] bck_regx1;
  wire   [7:2] do_xana1;
  wire   [7:0] do_xana0;
  wire   [3:0] do_regx_xtm;
  wire   [5:2] do_cvctl;
  wire   [3:0] do_vooc;
  wire   [5:0] do_dpdm;
  wire   [5:4] do_srcctl;
  wire   [7:0] do_cctrx;
  wire   [5:0] di_xanav;
  wire   [5:0] srci;
  tri   CSP;
  tri   CSN;
  tri   VFB;
  tri   COMP;
  tri   SW;
  tri   BST;
  tri   VDRV;
  tri   DP;
  tri   DN;
  tri   CC1;
  tri   CC2;
  tri   TST;
  tri   GPIO_TS;
  tri   SCL;
  tri   SDA;
  tri   GPIO1;
  tri   GPIO2;
  tri   GPIO3;
  tri   GPIO4;
  tri   GPIO5;
  tri   [7:0] xdat_o;

  anatop_1127a0 U0_ANALOG_TOP ( .CC1(CC1), .CC2(CC2), .DP(DP), .DN(DN), .VFB(
        VFB), .CSP(CSP), .CSN(CSN), .COMP(COMP), .SW(SW), .BST(BST), .VDRV(
        VDRV), .LG(LG), .HG(HG), .GATE(GATE), .BST_SET(bck_regx0[0]), 
        .DCM_SEL(bck_regx0[1]), .HGOFF(bck_regx0[2]), .HGON(bck_regx0[4]), 
        .LGOFF(bck_regx0[3]), .LGON(bck_regx0[5]), .EN_DRV(bck_regx0[6]), 
        .FSW(FSW), .EN_OSC(bck_regx1[2]), .MAXDS(bck_regx1[3]), .EN_GM(
        bck_regx1[4]), .EN_ODLDO(bck_regx1[5]), .EN_IBUK(bck_regx1[6]), 
        .EN_CP(do_srcctl_0), .EXT_CP(bck_regx1[7]), .INT_CP(bck_regx0[7]), 
        .ANTI_INRUSH(do_cvctl[5]), .PWREN_HOLD(PWREN_HOLD), .RP_SEL(RP_SEL), 
        .RP1_EN(RP_EN[0]), .RP2_EN(RP_EN[1]), .VCONN1_EN(VCONN_EN[0]), 
        .VCONN2_EN(VCONN_EN[1]), .SGP({do_cctrx[0], do_regx_xtm}), .S20U(
        do_cctrx[1]), .S100U(do_cctrx[2]), .TX_EN(TX_EN), .TX_DAT(TX_DAT), 
        .CC_SEL(do_ccctl_0_), .TRA(do_cctrx[4]), .TFA(do_cctrx[5]), .LSR(
        do_cctrx[6]), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .SEL_RX_TH(do_cctrx[7]), .DAC1_EN(DAC1_EN), .DPDN_SHORT(do_dpdm[0]), .DP_2V7_EN(do_dpdm[4]), 
        .DN_2V7_EN(do_dpdm[3]), .DP_0P6V_EN(do_xana1[3]), .DN_0P6V_EN(
        do_xana1[2]), .DP_DWN_EN(do_dpdm[2]), .DN_DWN_EN(do_dpdm[1]), 
        .CC_SLOPE(CC_SLOPE), .DAC2(PWR_I), .DAC3(DAC3_V), .DAC1(DAC1), .CV2(
        do_xana0[0]), .LFOSC_ENB(LFOSC_ENB), .VO_DISCHG(do_srcctl[4]), 
        .DISCHG_SEL(do_srcctl[5]), .CMP_SEL_VO10(SAMPL_SEL[1]), .CMP_SEL_VO20(
        SAMPL_SEL[10]), .CMP_SEL_GP1(SAMPL_SEL[17]), .CMP_SEL_GP2(
        SAMPL_SEL[16]), .CMP_SEL_GP3(SAMPL_SEL[15]), .CMP_SEL_GP4(
        SAMPL_SEL[14]), .CMP_SEL_GP5(SAMPL_SEL[13]), .CMP_SEL_VIN20(
        SAMPL_SEL[0]), .CMP_SEL_TS(SAMPL_SEL[3]), .CMP_SEL_IS(SAMPL_SEL[2]), 
        .CMP_SEL_CC2(SAMPL_SEL[7]), .CMP_SEL_CC1(SAMPL_SEL[6]), 
        .CMP_SEL_CC2_4(SAMPL_SEL[12]), .CMP_SEL_CC1_4(SAMPL_SEL[11]), 
        .CMP_SEL_DP(SAMPL_SEL[4]), .CMP_SEL_DP_3(SAMPL_SEL[8]), .CMP_SEL_DN(
        SAMPL_SEL[5]), .CMP_SEL_DN_3(SAMPL_SEL[9]), .OCP_EN(do_cvctl[2]), 
        .COMP_O(COMP_O), .CCI2C_EN(CCI2C_EN), .UVP_SEL(do_xana0[7]), .TM(
        ANA_TM), .V5OCP(srci[4]), .RSTB(RSTB), .DAC0(DAC0), .SLEEP(SLEEP), 
        .OSC_LOW(OSC_LOW), .OSC_STOP(OSC_STOP), .PWRDN(PWRDN), .VPP_ZERO(
        VPP_0V), .OSC_O(OSC_O), .RD_DET(RD_DET), .IMP_OSC(IMP_OSC), .DRP_OSC(
        DRP_OSC), .STB_RP(STB_RP), .RD_ENB(RD_ENB), .OCP(srci[1]), .SCP(
        srci[3]), .UVP(srci[0]), .LDO3P9V(LDO3P9V), .VPP_SEL(VPP_SEL), 
        .CC1_DOB(CC1_DOB), .CC2_DOB(CC2_DOB), .CC1_DI(CC1_DI), .CC2_DI(CC2_DI), 
        .OTPI(srci[5]), .OVP_SEL(OVP_SEL), .OVP(srci[2]), .DN_COMP(DN_COMP), 
        .DP_COMP(DP_COMP), .DPDN_VTH(do_xana0[5]), .DPDEN(do_vooc[3]), .DPDO(
        do_vooc[2]), .DPIE(do_dpdm[5]), .DNDEN(do_vooc[1]), .DNDO(do_vooc[0]), 
        .DNIE(do_dpdm[5]), .CP_CLKX2(ANAOPT[7]), .SEL_CONST_OVP(ANAOPT[6]), 
        .LP_EN(ANAOPT[5]), .DNCHK_EN(ANAOPT[3]), .IRP_EN(ANAOPT[2]), .CCFBEN(
        ANAOPT[0]), .REGTRM(REGTRM), .AD_RST(AD_RST), .AD_HOLD(AD_HOLD), 
        .DN_FAULT(DN_FAULT), .SEL_CCGAIN(do_xana0[3]), .VFB_SWB(do_xana0[1]), 
        .CPVSEL(do_xana1[6]), .CLAMPV_EN(do_xana1[5]), .HVNG_CPEN(do_xana1[7]), 
        .OCP_SEL(OCP_SEL), .OCP_80M(di_xanav[1]), .OCP_160M(di_xanav[0]), 
        .DMY_OUT(di_xanav[5:2]), .DMY_IN(DUMMY_IN), .VPP_OTP(VPP_OTP), 
        .RSTB_5(IO_RSTB5), .V1P1(V1P1), .TS_ANA_R(TS_ANA_R), .GP5_ANA_R(
        GP5_ANA_R), .GP4_ANA_R(GP4_ANA_R), .GP3_ANA_R(GP3_ANA_R), .GP2_ANA_R(
        GP2_ANA_R), .GP1_ANA_R(GP1_ANA_R), .TS_ANA_P(ANAP_TS), .GP5_ANA_P(
        ANAP_GP5), .GP4_ANA_P(ANAP_GP4), .GP3_ANA_P(ANAP_GP3), .GP2_ANA_P(
        ANAP_GP2), .GP1_ANA_P(ANAP_GP1) );
  IODMURUDA_A0 PAD_SCL ( .DO(DO_GPIO[0]), .IE(IE_GPIO[1]), .OE(OE_GPIO[0]), 
        .PD(PD_GPIO[0]), .PU(PU_GPIO[0]), .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(
        SCL), .ANA_R(), .DI(DI_GPIO[0]) );
  IODMURUDA_A0 PAD_SDA ( .DO(DO_GPIO[1]), .IE(IE_GPIO[1]), .OE(OE_GPIO[1]), 
        .PD(PD_GPIO[1]), .PU(PU_GPIO[1]), .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(
        SDA), .ANA_R(), .DI(DI_GPIO[1]) );
  IOBMURUDA_A0 PAD_TST ( .DO(1'b0), .IE(1'b1), .OE(1'b0), .PD(1'b1), .PU(1'b0), 
        .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(TST), .ANA_R(), .DI(DI_TST) );
  IOBMURUDA_A1 PAD_GPIO1 ( .ANA_P(ANAP_GP1), .DO(DO_GPIO[2]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[2]), .PD(PD_GPIO[2]), .PU(PU_GPIO[2]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO1), .ANA_R(GP1_ANA_R), .DI(DI_GPIO[2]) );
  IOBMURUDA_A1 PAD_GPIO2 ( .ANA_P(ANAP_GP2), .DO(DO_GPIO[3]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[3]), .PD(PD_GPIO[3]), .PU(PU_GPIO[3]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO2), .ANA_R(GP2_ANA_R), .DI(DI_GPIO[3]) );
  IOBMURUDA_A1 PAD_GPIO3 ( .ANA_P(ANAP_GP3), .DO(DO_GPIO[4]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[4]), .PD(PD_GPIO[4]), .PU(PU_GPIO[4]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO3), .ANA_R(GP3_ANA_R), .DI(DI_GPIO[4]) );
  IOBMURUDA_A1 PAD_GPIO4 ( .ANA_P(ANAP_GP4), .DO(DO_GPIO[5]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[5]), .PD(PD_GPIO[5]), .PU(PU_GPIO[5]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO4), .ANA_R(GP4_ANA_R), .DI(DI_GPIO[5]) );
  IOBMURUDA_A1 PAD_GPIO5 ( .ANA_P(ANAP_GP5), .DO(DO_GPIO[6]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[6]), .PD(PD_GPIO[6]), .PU(PU_GPIO[6]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO5), .ANA_R(GP5_ANA_R), .DI(DI_GPIO[6]) );
  IOBMURUDA_A1 PAD_GPIO_TS ( .ANA_P(ANAP_TS), .DO(DO_TS[3]), .IE(IE_GPIO[0]), 
        .OE(DO_TS[2]), .PD(DO_TS[0]), .PU(DO_TS[1]), .RSTB_5(IO_RSTB5), .VB(
        V1P1), .PAD(GPIO_TS), .ANA_R(TS_ANA_R), .DI(DI_TS) );
  MSL18B_1536X8_RW10TM4_16_20221107 U0_SRAM ( .A(SRAM_A), .DI(SRAM_D), .DO(
        xdat_o), .CK(SRAM_CLK), .WEB(SRAM_WEB), .CSB(SRAM_CEB), .OEB(SRAM_OEB)
         );
  ATO0008KX8MX180LBX4DA U0_CODE_0_ ( .A(PMEM_A), .TWLB(PMEM_TWLB), .Q(PMEM_Q0), 
        .SAP(PMEM_SAP), .CSB(PMEM_CSB), .CLK(PMEM_CLK[0]), .PGM(n1), .RE(
        PMEM_RE), .VDDP(VPP_OTP), .VDD(), .VSS() );
  ATO0008KX8MX180LBX4DA U0_CODE_1_ ( .A(PMEM_A), .TWLB(PMEM_TWLB), .Q(PMEM_Q1), 
        .SAP(PMEM_SAP), .CSB(PMEM_CSB), .CLK(PMEM_CLK[1]), .PGM(PMEM_PGM), 
        .RE(PMEM_RE), .VDDP(VPP_OTP), .VDD(), .VSS() );
  core_a0 U0_CORE ( .SRCI(srci), .XANAV(di_xanav), .BCK_REGX({bck_regx1, FSW, 
        bck_regx0}), .ANA_REGX({do_xana1[7:5], SYNOPSYS_UNCONNECTED_1, 
        do_xana1[3:2], SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        do_xana0[7], SYNOPSYS_UNCONNECTED_4, do_xana0[5], 
        SYNOPSYS_UNCONNECTED_5, do_xana0[3], SYNOPSYS_UNCONNECTED_6, 
        do_xana0[1:0]}), .LFOSC_ENB(LFOSC_ENB), .STB_RP(STB_RP), .RD_ENB(
        RD_ENB), .OCP_SEL(OCP_SEL), .PWREN_HOLD(PWREN_HOLD), .CC1_DI(CC1_DI), 
        .CC2_DI(CC2_DI), .DRP_OSC(DRP_OSC), .IMP_OSC(IMP_OSC), .CC1_DOB(
        CC1_DOB), .CC2_DOB(CC2_DOB), .DAC1_EN(DAC1_EN), .SH_RST(AD_RST), 
        .SH_HOLD(AD_HOLD), .LDO3P9V(LDO3P9V), .XTM(do_regx_xtm), .DO_CVCTL({
        OVP_SEL, do_cvctl[5], SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        do_cvctl[2], SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10}), 
        .DO_CCTRX({do_cctrx[7:4], SYNOPSYS_UNCONNECTED_11, do_cctrx[2:0]}), 
        .DO_SRCCTL({CC_SLOPE, do_srcctl, VCONN_EN, SYNOPSYS_UNCONNECTED_12, 
        do_srcctl_0}), .DO_CCCTL({RP_EN, RP_SEL, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, do_ccctl_0_}), 
        .DO_DAC0(DAC0), .DO_DPDN(do_dpdm), .DO_VOOC(do_vooc), .DO_PWR_I(PWR_I), 
        .PMEM_A(PMEM_A), .PMEM_Q0(PMEM_Q0), .PMEM_Q1(PMEM_Q1), .PMEM_TWLB(
        PMEM_TWLB), .PMEM_SAP(PMEM_SAP), .PMEM_CLK(PMEM_CLK), .PMEM_CSB(
        PMEM_CSB), .PMEM_RE(PMEM_RE), .PMEM_PGM(PMEM_PGM), .VPP_SEL(VPP_SEL), 
        .VPP_0V(VPP_0V), .SRAM_WEB(SRAM_WEB), .SRAM_CEB(SRAM_CEB), .SRAM_OEB(
        SRAM_OEB), .SRAM_CLK(SRAM_CLK), .SRAM_A(SRAM_A), .SRAM_D(SRAM_D), 
        .SRAM_RDAT(xdat_o), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .RD_DET(RD_DET), 
        .TX_DAT(TX_DAT), .TX_EN(TX_EN), .OSC_STOP(OSC_STOP), .OSC_LOW(OSC_LOW), 
        .SLEEP(SLEEP), .PWRDN(PWRDN), .OCDRV_ENZ(), .DAC1_V(DAC1), .SAMPL_SEL(
        SAMPL_SEL), .DAC1_COMP(COMP_O), .CCI2C_EN(CCI2C_EN), .ANA_TM(ANA_TM), 
        .DM_FAULT(DN_FAULT), .DM_COMP(DN_COMP), .DP_COMP(DP_COMP), .DI_GPIO(
        DI_GPIO), .DO_GPIO(DO_GPIO), .OE_GPIO(OE_GPIO), .GPIO_PU(PU_GPIO), 
        .GPIO_PD(PD_GPIO), .GPIO_IE(IE_GPIO), .DO_TS(DO_TS), .DI_TS(DI_TS), 
        .REGTRM(REGTRM), .ANAOPT({ANAOPT[7:5], SYNOPSYS_UNCONNECTED_16, 
        ANAOPT[3:2], SYNOPSYS_UNCONNECTED_17, ANAOPT[0]}), .DUMMY_IN(DUMMY_IN), 
        .DAC3_V(DAC3_V), .i_clk(OSC_O), .i_rstz(RSTB), .atpg_en(tm_atpg), 
        .di_tst(DI_TST), .tm_atpg(tm_atpg) );
  BUFX12 U3 ( .A(PMEM_PGM), .Y(n1) );
endmodule


module core_a0 ( SRCI, XANAV, BCK_REGX, ANA_REGX, LFOSC_ENB, STB_RP, RD_ENB, 
        OCP_SEL, PWREN_HOLD, CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, CC1_DOB, 
        CC2_DOB, DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, XTM, DO_CVCTL, DO_CCTRX, 
        DO_SRCCTL, DO_CCCTL, DO_DAC0, DO_DPDN, DO_VOOC, DO_PWR_I, PMEM_A, 
        PMEM_Q0, PMEM_Q1, PMEM_TWLB, PMEM_SAP, PMEM_CLK, PMEM_CSB, PMEM_RE, 
        PMEM_PGM, VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, 
        SRAM_A, SRAM_D, SRAM_RDAT, RX_DAT, RX_SQL, RD_DET, TX_DAT, TX_EN, 
        OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, DAC1_V, SAMPL_SEL, 
        DAC1_COMP, CCI2C_EN, ANA_TM, DM_FAULT, DM_COMP, DP_COMP, DI_GPIO, 
        DO_GPIO, OE_GPIO, GPIO_PU, GPIO_PD, GPIO_IE, DO_TS, DI_TS, REGTRM, 
        ANAOPT, DUMMY_IN, DAC3_V, i_clk, i_rstz, atpg_en, di_tst, tm_atpg );
  input [5:0] SRCI;
  input [5:0] XANAV;
  output [15:0] BCK_REGX;
  output [15:0] ANA_REGX;
  output [3:0] XTM;
  output [7:0] DO_CVCTL;
  output [7:0] DO_CCTRX;
  output [7:0] DO_SRCCTL;
  output [7:0] DO_CCCTL;
  output [10:0] DO_DAC0;
  output [5:0] DO_DPDN;
  output [3:0] DO_VOOC;
  output [7:0] DO_PWR_I;
  output [15:0] PMEM_A;
  input [7:0] PMEM_Q0;
  input [7:0] PMEM_Q1;
  output [1:0] PMEM_TWLB;
  output [1:0] PMEM_SAP;
  output [1:0] PMEM_CLK;
  output [10:0] SRAM_A;
  output [7:0] SRAM_D;
  input [7:0] SRAM_RDAT;
  output [9:0] DAC1_V;
  output [17:0] SAMPL_SEL;
  output [3:0] ANA_TM;
  input [6:0] DI_GPIO;
  output [6:0] DO_GPIO;
  output [6:0] OE_GPIO;
  output [6:0] GPIO_PU;
  output [6:0] GPIO_PD;
  output [1:0] GPIO_IE;
  output [3:0] DO_TS;
  output [55:0] REGTRM;
  output [7:0] ANAOPT;
  output [4:0] DUMMY_IN;
  output [5:0] DAC3_V;
  input CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, RX_DAT, RX_SQL, RD_DET, DAC1_COMP,
         DM_FAULT, DM_COMP, DP_COMP, DI_TS, i_clk, i_rstz, atpg_en, di_tst;
  output LFOSC_ENB, STB_RP, RD_ENB, OCP_SEL, PWREN_HOLD, CC1_DOB, CC2_DOB,
         DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, PMEM_CSB, PMEM_RE, PMEM_PGM,
         VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, TX_DAT,
         TX_EN, OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, CCI2C_EN, tm_atpg;
  wire   N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N268, n687, n688, aswclk, detclk, tclk_sel, s_clk, aswkup, x_clk,
         t_di_gpio4, t_pmem_clk, pmem_csb, t_pmem_csb, r_osc_gate, t_osc_gate,
         g_clk, xram_ce, iram_ce, r_i2c_attr, esfrm_oe, esfrm_we, sfrack,
         ictlr_psrack, esfrm_rrdy, memwr, memrd, memrd_c, memack, o_cpurst,
         hit_xd, hit_xr, hit_ps, hit_ps_c, mcu_ram_r, mcu_ram_w, regx_re,
         iram_we, xram_we, regx_we, bist_en, bist_wr, srstz, prl_cany0w,
         prl_cany0r, mempsrd, r_bclk_sel, r_hold_mcu, t0_intr, fcp_intr,
         dpdm_urx, s0_rxdoe, mcuo_scl, mcuo_sda, mempsack, mempswr, mempsrd_c,
         sfr_w, sfr_r, ictlr_psack, ictlr_inc, set_hold, bkpt_hold, bkpt_ena,
         r_psrd, r_pswr, prl_cany0, prl_c0set, pmem_pgm, pmem_re, we_twlb,
         r_otp_wpls, pwrdn_rst, r_otp_pwdn_en, ramacc, frc_lg_on, gating_pwr,
         cc1_di, cc2_di, r_sleep, ps_pwrdn, r_pwrdn, r_ocdrv_enz, r_osc_stop,
         r_pwrv_upd, r_otpi_gate, r_fcpre, r_fortxdat, r_fortxrdy, r_fortxen,
         r_gpio_tm, pid_goidle, pid_gobusy, bus_idle, sse_idle, r_exist1st,
         r_ordrs4, r_fifopsh, r_fifopop, r_unlock, r_first, r_last, r_fiforst,
         r_set_cpmsgid, r_txendk, r_txshrt, r_auto_discard, r_dat_portrole,
         r_dat_datarole, r_pshords, r_discard, r_strtch, r_i2c_ninc,
         r_i2c_fwnak, r_i2c_fwack, hwi2c_stretch, i2c_ev_6_, i2c_ev_3,
         i2c_ev_2, prl_discard, prl_GCTxDone, pff_obsd, pff_empty, pff_full,
         ptx_ack, clk_1p0m, clk_500, prstz, sse_rdrdy, upd_rdrdy, sse_prefetch,
         slvo_sda, slvo_re, slvo_early, dm_comp, dp_comp, di_sqlch, ptx_cc,
         ptx_oe, sh_rst, sh_hold, fcp_oe, fcp_do, sdischg_duty, clk_100k,
         r_bck2_2_, r_imp_osc, clk_500k, r_vpp_en, r_vpp0v_en, di_ts,
         di_aswk_0, r_xana_23, r_xana_19, r_xana_18, divff_o1, clk_50k, N448,
         o_dodat0_15_, N568, N569, N570, N571, N572, N575, N576, N577, N578,
         N579, N580, N581, N582, N583, N584, N1478, N1483, net8853, n123, n126,
         n128, n129, n131, n133, n135, n137, n138, n140, n508, n509, n510,
         n511, n4, n300, n297, n296, n299, n298, n58, n82, n83, n84, n531,
         n532, n557, n558, n559, n560, n561, n562, n563, n564, n10, n43, n50,
         n51, n142, n145, n680, n681, n682, n683, n684, n685, n686, n722, n723,
         n724, n762, n812, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n941, n942, n943, n952, n953, n954, n955, n956, n957, n959, n960,
         n961, n962, n964, n965, n966, n973, n975, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1133, n1134,
         n1135, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1152, n1153, n1154, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1, n2, n3, n5, n6, n7, n8,
         n9, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n29, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n44, n45, n46, n47, n48, n49, n52, n53, n54, n55, n56, n57, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n124, n125, n127, n130,
         n132, n134, n136, n139, n141, n143, n144, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108;
  wire   [9:0] aswclk_ps;
  wire   [9:0] detclk_ps;
  wire   [1:0] pmem_clk;
  wire   [7:0] sse_wdat;
  wire   [7:0] prx_fifowdat;
  wire   [7:0] sse_adr;
  wire   [7:0] prl_cany0adr;
  wire   [7:0] esfrm_wdat;
  wire   [6:0] esfrm_adr;
  wire   [7:0] mcu_esfrrdat;
  wire   [7:0] delay_inst;
  wire   [7:0] esfrm_rdat;
  wire   [3:0] r_pg0_sel;
  wire   [15:0] memaddr;
  wire   [15:0] memaddr_c;
  wire   [7:0] memdatao;
  wire   [7:0] idat_adr;
  wire   [7:0] idat_wdat;
  wire   [10:0] iram_a;
  wire   [10:0] xram_a;
  wire   [7:0] iram_d;
  wire   [7:0] xram_d;
  wire   [1:0] sram_rdat;
  wire   [7:0] regx_rdat;
  wire   [10:0] bist_adr;
  wire   [7:0] bist_wdat;
  wire   [7:0] memdatai;
  wire   [7:0] ictlr_inst;
  wire   [15:0] mcu_pc;
  wire   [22:16] mcu_dbgpo;
  wire   [3:2] sfr_intr;
  wire   [7:0] exint;
  wire   [7:0] ff_p0;
  wire   [6:0] do_p0;
  wire   [7:0] sfr_rdat;
  wire   [7:0] sfr_wdat;
  wire   [6:0] sfr_adr;
  wire   [14:0] bkpt_pc;
  wire   [14:0] r_inst_ofs;
  wire   [7:0] pmem_q0;
  wire   [7:0] pmem_q1;
  wire   [1:0] pmem_twlb;
  wire   [1:0] wd_twlb;
  wire   [1:0] r_sqlch;
  wire   [3:2] r_ccrx;
  wire   [1:0] r_rxdb_opt;
  wire   [7:4] r_pwrctl;
  wire   [5:2] di_pro;
  wire   [1:0] lg_pulse_len;
  wire   [7:0] r_srcctl;
  wire   [7:0] r_dpdmctl;
  wire   [11:0] r_fw_pwrv;
  wire   [5:0] r_cvcwr;
  wire   [15:0] r_cvofs;
  wire   [7:0] r_cctrx;
  wire   [7:0] r_ccctl;
  wire   [6:0] r_fcpwr;
  wire   [7:0] fcp_r_dat;
  wire   [7:0] fcp_r_sta;
  wire   [7:0] fcp_r_msk;
  wire   [7:0] fcp_r_ctl;
  wire   [7:0] fcp_r_crc;
  wire   [7:0] fcp_r_acc;
  wire   [7:0] fcp_r_tui;
  wire   [7:0] r_accctl;
  wire   [7:5] r_comp_opt;
  wire   [14:0] sfr_dacwr;
  wire   [17:0] r_dac_en;
  wire   [17:0] r_sar_en;
  wire   [7:0] r_isofs;
  wire   [7:0] r_adofs;
  wire   [7:0] dac_r_ctl;
  wire   [7:0] dac_r_cmpsta;
  wire   [17:0] dac_r_comp;
  wire   [143:0] dac_r_vs;
  wire   [5:0] x_daclsb;
  wire   [6:0] REVID;
  wire   [6:0] r_pu_gpio;
  wire   [6:0] r_pd_gpio;
  wire   [6:0] r_gpio_oe;
  wire   [1:0] r_gpio_ie;
  wire   [55:0] r_regtrm;
  wire   [3:0] r_ana_tm;
  wire   [7:0] i2c_ltbuf;
  wire   [7:0] i2c_lt_ofs;
  wire   [4:0] r_txnumk;
  wire   [1:0] r_auto_gdcrc;
  wire   [1:0] r_spec;
  wire   [1:0] r_dat_spec;
  wire   [6:0] r_txauto;
  wire   [6:0] r_rxords_ena;
  wire   [7:1] r_i2c_deva;
  wire   [2:0] prl_cpmsgid;
  wire   [1:0] pff_ack;
  wire   [7:0] pff_rdat;
  wire   [15:0] pff_rxpart;
  wire   [5:0] pff_ptr;
  wire   [6:0] prx_setsta;
  wire   [1:0] prx_rst;
  wire   [4:0] prx_rcvinf;
  wire   [5:0] prx_adpn;
  wire   [3:0] prx_fsm;
  wire   [2:0] ptx_fsm;
  wire   [3:0] prl_fsm;
  wire   [3:0] slvo_ev;
  wire   [1:0] r_i2cslv_route;
  wire   [5:4] r_i2crout;
  wire   [1:0] r_i2cmcu_route;
  wire   [18:17] upd_dbgpo;
  wire   [7:0] r_dacwdat;
  wire   [17:8] wr_dacv;
  wire   [10:7] r_dacwr;
  wire   [17:0] dacmux_sel;
  wire   [3:0] comp_smpl;
  wire   [7:0] r_cvcwdat;
  wire   [7:0] r_sdischg;
  wire   [7:0] r_vcomp;
  wire   [7:0] r_idacsh;
  wire   [7:0] r_cvofsx;
  wire   [7:0] r_xtm;
  wire   [6:0] bist_r_ctl;
  wire   [1:0] regx_hitbst;
  wire   [7:0] bist_r_dat;
  wire   [1:0] regx_wrpwm;
  wire   [15:0] r_pwm;
  wire   [1:0] r_sap;
  wire   [3:0] lt_gpi;
  wire   [6:0] r_do_ts;
  wire   [3:0] r_dpdo_sel;
  wire   [3:0] r_dndo_sel;
  wire   [4:2] di_aswk;
  wire   [7:0] r_bck0;
  wire   [7:0] r_bck1;
  wire   [15:0] r_xana;
  wire   [5:0] di_xanav;
  wire   [7:0] r_aopt;
  wire   [6:0] di_gpio;
  wire   [7:6] do_opt;
  wire   [1:0] pwm_o;
  wire   [15:0] d_dodat;
  wire   [3:0] r_lt_gpi;
  tri   [7:0] SRAM_RDAT;

  CKBUFX1 U0_ASWCLK_BUF_0_ ( .A(aswclk_ps[0]), .Y(aswclk_ps[1]) );
  CKBUFX1 U0_ASWCLK_BUF_1_ ( .A(aswclk_ps[1]), .Y(aswclk_ps[2]) );
  CKBUFX1 U0_ASWCLK_BUF_2_ ( .A(aswclk_ps[2]), .Y(aswclk_ps[3]) );
  CKBUFX1 U0_ASWCLK_BUF_3_ ( .A(aswclk_ps[3]), .Y(aswclk_ps[4]) );
  CKBUFX1 U0_ASWCLK_BUF_4_ ( .A(aswclk_ps[4]), .Y(aswclk_ps[5]) );
  CKBUFX1 U0_ASWCLK_BUF_5_ ( .A(aswclk_ps[5]), .Y(aswclk_ps[6]) );
  CKBUFX1 U0_ASWCLK_BUF_6_ ( .A(aswclk_ps[6]), .Y(aswclk_ps[7]) );
  CKBUFX1 U0_ASWCLK_BUF_7_ ( .A(aswclk_ps[7]), .Y(aswclk_ps[8]) );
  CKBUFX1 U0_ASWCLK_BUF_8_ ( .A(aswclk_ps[8]), .Y(aswclk_ps[9]) );
  CKBUFX1 U0_ASWCLK_BUF_9_ ( .A(aswclk_ps[9]), .Y(aswclk) );
  CKBUFX1 U0_DETCLK_BUF_0_ ( .A(detclk_ps[0]), .Y(detclk_ps[1]) );
  CKBUFX1 U0_DETCLK_BUF_1_ ( .A(detclk_ps[1]), .Y(detclk_ps[2]) );
  CKBUFX1 U0_DETCLK_BUF_2_ ( .A(detclk_ps[2]), .Y(detclk_ps[3]) );
  CKBUFX1 U0_DETCLK_BUF_3_ ( .A(detclk_ps[3]), .Y(detclk_ps[4]) );
  CKBUFX1 U0_DETCLK_BUF_4_ ( .A(detclk_ps[4]), .Y(detclk_ps[5]) );
  CKBUFX1 U0_DETCLK_BUF_5_ ( .A(detclk_ps[5]), .Y(detclk_ps[6]) );
  CKBUFX1 U0_DETCLK_BUF_6_ ( .A(detclk_ps[6]), .Y(detclk_ps[7]) );
  CKBUFX1 U0_DETCLK_BUF_7_ ( .A(detclk_ps[7]), .Y(detclk_ps[8]) );
  CKBUFX1 U0_DETCLK_BUF_8_ ( .A(detclk_ps[8]), .Y(detclk_ps[9]) );
  CKBUFX1 U0_DETCLK_BUF_9_ ( .A(detclk_ps[9]), .Y(detclk) );
  AND2X1 U0_SCAN_EN ( .A(DI_GPIO[2]), .B(n95), .Y(n10) );
  CKMUX2X1 U0_CLK_MUX ( .D0(i_clk), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(s_clk)
         );
  CKMUX2X1 U0_DCLKMUX ( .D0(RD_DET), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        detclk_ps[0]) );
  CKMUX2X1 U0_ACLKMUX ( .D0(aswkup), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        aswclk_ps[0]) );
  CKBUFX1 U0_MCK_BUF ( .A(i_clk), .Y(x_clk) );
  CKBUFX1 U0_TCK_BUF ( .A(DI_GPIO[4]), .Y(t_di_gpio4) );
  CKBUFX1 U0_BUF_NEG0 ( .A(pmem_clk[0]), .Y(t_pmem_clk) );
  CKBUFX1 U0_BUF_NEG1 ( .A(pmem_csb), .Y(t_pmem_csb) );
  CKBUFX1 U0_BUF_NEG2 ( .A(r_osc_gate), .Y(t_osc_gate) );
  CLKDLX1 U0_MCLK_ICG ( .CK(s_clk), .E(n289), .SE(n113), .ECK(g_clk) );
  CLKDLX1 U0_SRAM_ICG ( .CK(g_clk), .E(n208), .SE(n112), .ECK(SRAM_CLK) );
  INVX1 U0_REVIDZ_0_ ( .A(1'b0), .Y(REVID[0]) );
  INVX1 U0_REVIDZ_1_ ( .A(1'b1), .Y(REVID[1]) );
  INVX1 U0_REVIDZ_2_ ( .A(1'b1), .Y(REVID[2]) );
  INVX1 U0_REVIDZ_3_ ( .A(1'b1), .Y(REVID[3]) );
  INVX1 U0_REVIDZ_4_ ( .A(1'b0), .Y(REVID[4]) );
  INVX1 U0_REVIDZ_5_ ( .A(1'b0), .Y(REVID[5]) );
  INVX1 U0_REVIDZ_6_ ( .A(1'b1), .Y(REVID[6]) );
  INVX1 U147 ( .A(n84), .Y(n82) );
  INVX1 U162 ( .A(n84), .Y(n83) );
  INVX1 U198 ( .A(srstz), .Y(n84) );
  MUX2X1 U1044 ( .D0(n687), .D1(DUMMY_IN[4]), .S(n10), .Y(DO_GPIO[6]) );
  MUX2X1 U1045 ( .D0(n688), .D1(PMEM_A[15]), .S(n10), .Y(DO_GPIO[5]) );
  mpb_a0 u0_mpb ( .i_rd({prl_cany0r, n762}), .i_wr({prl_cany0w, i2c_ev_3}), 
        .wdat0(sse_wdat), .wdat1(prx_fifowdat), .addr0(sse_adr), .addr1(
        prl_cany0adr), .r_i2c_attr(r_i2c_attr), .esfrm_oe(esfrm_oe), 
        .esfrm_we(esfrm_we), .sfrack(sfrack), .esfrm_wdat(esfrm_wdat), 
        .esfrm_adr(esfrm_adr), .mcu_esfr_rdat(mcu_esfrrdat), .delay_rdat(
        delay_inst), .delay_rrdy(ictlr_psrack), .esfrm_rrdy(esfrm_rrdy), 
        .esfrm_rdat(esfrm_rdat), .channel_sel(1'b0), .r_pg0_sel(r_pg0_sel), 
        .dma_w(1'b0), .dma_r(1'b0), .dma_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_wdat({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_ack(), .memaddr(memaddr), 
        .memaddr_c({memaddr_c[15:7], n44, memaddr_c[5], n42, memaddr_c[3:0]}), 
        .memwr(memwr), .memrd(memrd), .memrd_c(memrd_c), .cpurst(o_cpurst), 
        .memdatao(memdatao), .memack(memack), .hit_xd(hit_xd), .hit_xr(hit_xr), 
        .hit_ps(hit_ps), .hit_ps_c(hit_ps_c), .idat_r(mcu_ram_r), .idat_w(
        mcu_ram_w), .idat_adr(idat_adr), .idat_wdat(idat_wdat), .iram_ce(
        iram_ce), .xram_ce(xram_ce), .regx_re(regx_re), .iram_we(iram_we), 
        .xram_we(xram_we), .regx_we(regx_we), .iram_a(iram_a), .xram_a(xram_a), 
        .iram_d(iram_d), .xram_d(xram_d), .iram_rdat({n129, n131, n133, n135, 
        n138, n140, sram_rdat}), .xram_rdat({n129, n131, n133, n135, n138, 
        n140, sram_rdat}), .regx_rdat({regx_rdat[7], n6, regx_rdat[5:1], n5}), 
        .bist_en(bist_en), .bist_wr(bist_wr), .bist_adr(bist_adr), .bist_wdat(
        bist_wdat), .bist_xram(1'b0), .mclk(g_clk), .srstz(srstz), .test_si(
        n145), .test_so(n142), .test_se(n10) );
  mcu51_a0 u0_mcu ( .bclki2c(r_bclk_sel), .pc_ini({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .slp2wakeup(1'b0), .r_hold_mcu(r_hold_mcu), .wdt_slow(1'b0), .wdtov({n145, 
        SYNOPSYS_UNCONNECTED_1}), .mdubsy(), .cs_run(), .t0_intr(t0_intr), 
        .clki2c(g_clk), .clkmdu(g_clk), .clkur0(g_clk), .clktm0(g_clk), 
        .clktm1(g_clk), .clkwdt(g_clk), .i2c_autoack(1'b0), .i2c_con_ens1(), 
        .clkcpu(g_clk), .clkper(g_clk), .reset(n84), .ro(o_cpurst), .port0i({
        n4, di_gpio[6:4], n137, di_gpio[2:0]}), .exint_9(fcp_intr), .exint({
        exint[7:4], n724, n723, exint[1:0]}), .clkcpuen(), .clkperen(), 
        .port0o({SYNOPSYS_UNCONNECTED_2, do_p0}), .port0ff(ff_p0), .rxd0o(
        do_opt[7]), .txd0(do_opt[6]), .rxd0i(dpdm_urx), .rxd0oe(s0_rxdoe), 
        .scli(n509), .sdai(n511), .sclo(mcuo_scl), .sdao(mcuo_sda), 
        .waitstaten(), .mempsack(mempsack), .memack(memack), .memdatai(
        memdatai), .memdatao(memdatao), .memaddr(memaddr), .mempswr(mempswr), 
        .mempsrd(mempsrd), .memwr(memwr), .memrd(memrd), .memdatao_comb({
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10}), .memaddr_comb(
        memaddr_c), .mempswr_comb(), .mempsrd_comb(mempsrd_c), .memwr_comb(), 
        .memrd_comb(memrd_c), .ramdatai({n129, n131, n133, n135, n138, n140, 
        sram_rdat}), .ramdatao(idat_wdat), .ramaddr(idat_adr), .ramwe(
        mcu_ram_w), .ramoe(mcu_ram_r), .dbgpo({SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, mcu_dbgpo, mcu_pc}), 
        .sfrack(sfrack), .sfrdatai(sfr_rdat), .sfrdatao(sfr_wdat), .sfraddr(
        sfr_adr), .sfrwe(sfr_w), .sfroe(sfr_r), .esfrm_wrdata(esfrm_wdat), 
        .esfrm_addr(esfrm_adr), .esfrm_we(esfrm_we), .esfrm_oe(esfrm_oe), 
        .esfrm_rddata(mcu_esfrrdat), .test_si2(DI_GPIO[1]), .test_si1(n681), 
        .test_so1(n680), .test_se(n10) );
  ictlr_a0 u0_ictlr ( .bkpt_ena(bkpt_ena), .bkpt_pc(bkpt_pc), .memaddr_c({
        memaddr_c[14:7], n44, n12, n11, n19, n45, n21, n20}), .memaddr(
        memaddr[14:0]), .mcu_psr_c(mempsrd_c), .mcu_psw(mempswr), .hit_ps_c(
        hit_ps_c), .hit_ps(hit_ps), .mempsack(ictlr_psack), .memdatao(memdatao), .o_set_hold(set_hold), .o_bkp_hold(bkpt_hold), .o_ofs_inc(ictlr_inc), 
        .o_inst(ictlr_inst), .d_inst(delay_inst), .sfr_psrack(ictlr_psrack), 
        .sfr_psofs(r_inst_ofs), .sfr_psr(r_psrd), .sfr_psw(r_pswr), .dw_rst(
        prl_c0set), .dw_ena(prl_cany0), .sfr_wdat({n66, n64, n62, n60, n57, 
        n55, n53, n48}), .pmem_pgm(pmem_pgm), .pmem_re(pmem_re), .pmem_csb(
        pmem_csb), .pmem_clk(pmem_clk), .pmem_a(PMEM_A), .pmem_q0(pmem_q0), 
        .pmem_q1(pmem_q1), .pmem_twlb(pmem_twlb), .wd_twlb(wd_twlb), .we_twlb(
        we_twlb), .pwrdn_rst(pwrdn_rst), .r_pwdn_en(r_otp_pwdn_en), .r_multi(
        r_otp_wpls), .r_hold_mcu(r_hold_mcu), .clk(g_clk), .srst(o_cpurst), 
        .test_si3(n680), .test_si2(slvo_sda), .test_si1(n686), .test_so2(n681), 
        .test_so1(n685), .test_se(n10) );
  regbank_a0 u0_regbank ( .srci({di_pro[5], n531, n532, di_pro[2], n126, n128}), .lg_pulse_len(lg_pulse_len), .dm_fault(n1171), .cc1_di(cc1_di), .cc2_di(
        cc2_di), .di_rd_det(di_aswk[2]), .i_tmrf(t0_intr), .i_vcbyval(r_xtm[4]), .dnchk_en(n1170), .r_pwrv_upd(r_pwrv_upd), .aswkup(aswkup), .lg_dischg(
        frc_lg_on), .gating_pwr(gating_pwr), .ps_pwrdn(ps_pwrdn), .r_sleep(
        r_sleep), .r_pwrdn(r_pwrdn), .r_ocdrv_enz(r_ocdrv_enz), .r_osc_stop(
        r_osc_stop), .r_osc_lo(o_dodat0_15_), .r_osc_gate(r_osc_gate), 
        .r_fw_pwrv(r_fw_pwrv), .r_cvcwr(r_cvcwr[1:0]), .r_cvofs(r_cvofs), 
        .r_otpi_gate(r_otpi_gate), .r_pwrctl(r_pwrctl), .r_pwr_i(DO_PWR_I), 
        .r_cvctl(DO_CVCTL), .r_srcctl(r_srcctl), .r_dpdmctl(r_dpdmctl), 
        .r_ccrx({r_sqlch, SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        r_ccrx, r_rxdb_opt}), .r_cctrx(r_cctrx), .r_ccctl(r_ccctl), .r_fcpwr(
        r_fcpwr), .r_fcpre(r_fcpre), .fcp_r_dat(fcp_r_dat), .fcp_r_sta(
        fcp_r_sta), .fcp_r_msk(fcp_r_msk), .fcp_r_ctl(fcp_r_ctl), .fcp_r_crc(
        fcp_r_crc), .fcp_r_acc(fcp_r_acc), .fcp_r_tui(fcp_r_tui), .r_accctl(
        r_accctl), .r_bclk_sel(r_bclk_sel), .r_dacwr(sfr_dacwr), .r_dac_en(
        r_dac_en[7:0]), .r_sar_en(r_sar_en[7:0]), .r_adofs(r_adofs), .r_isofs(
        r_isofs), .x_daclsb(x_daclsb), .r_comp_opt({r_comp_opt, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}), .dac_r_ctl(dac_r_ctl), .dac_r_comp(
        dac_r_comp[7:0]), .dac_r_cmpsta(dac_r_cmpsta), .dac_r_vs(
        dac_r_vs[63:0]), .REVID(REVID), .atpg_en(n91), .sfr_r(sfr_r), .sfr_w(
        sfr_w), .set_hold(set_hold), .bkpt_hold(bkpt_hold), .cpurst(o_cpurst), 
        .sfr_addr({1'b1, sfr_adr}), .sfr_wdat({n66, n64, n62, n60, n57, n55, 
        n53, n48}), .sfr_rdat(sfr_rdat), .ff_p0(ff_p0), .di_p0({n4, 
        di_gpio[6:4], n137, di_gpio[2:0]}), .ictlr_idle(pmem_csb), .ictlr_inc(
        ictlr_inc), .r_inst_ofs(r_inst_ofs), .r_psrd(r_psrd), .r_pswr(r_pswr), 
        .r_fortxdat(r_fortxdat), .r_fortxrdy(r_fortxrdy), .r_fortxen(r_fortxen), .r_ana_tm(r_ana_tm), .r_gpio_tm(r_gpio_tm), .r_gpio_ie(r_gpio_ie), 
        .r_gpio_oe(r_gpio_oe), .r_gpio_pu(r_pu_gpio), .r_gpio_pd(r_pd_gpio), 
        .r_gpio_s0({N268, N267, N266}), .r_gpio_s1({N265, N264, N263}), 
        .r_gpio_s2({N262, N261, N260}), .r_gpio_s3({N259, N258, N257}), 
        .r_regtrm(r_regtrm), .i_pc(mcu_pc), .i_goidle(pid_goidle), .i_gobusy(
        pid_gobusy), .i_i2c_idle(sse_idle), .bus_idle(bus_idle), .i2c_stretch(
        hwi2c_stretch), .i_i2c_rwbuf(sse_wdat), .i_i2c_ltbuf(i2c_ltbuf), 
        .i_i2c_ofs(i2c_lt_ofs), .o_intr({exint[6], sfr_intr, exint[5:4]}), 
        .r_auto_gdcrc(r_auto_gdcrc), .r_exist1st(r_exist1st), .r_ordrs4(
        r_ordrs4), .r_fifopsh(r_fifopsh), .r_fifopop(r_fifopop), .r_unlock(
        r_unlock), .r_first(r_first), .r_last(r_last), .r_fiforst(r_fiforst), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_txendk(r_txendk), .r_txnumk(r_txnumk), .r_txshrt(r_txshrt), .r_auto_discard(r_auto_discard), .r_hold_mcu(r_hold_mcu), .r_txauto(r_txauto), .r_rxords_ena(r_rxords_ena), .r_spec(r_spec), 
        .r_dat_spec(r_dat_spec), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_discard(r_discard), .r_pshords(
        r_pshords), .r_pg0_sel(r_pg0_sel), .r_strtch(r_strtch), .r_i2c_attr(
        r_i2c_attr), .r_i2c_ninc(r_i2c_ninc), .r_hwi2c_en(), .r_i2c_fwnak(
        r_i2c_fwnak), .r_i2c_fwack(r_i2c_fwack), .r_i2c_deva(r_i2c_deva), 
        .i2c_ev({n762, i2c_ev_6_, slvo_ev[3:2], i2c_ev_3, i2c_ev_2, 
        slvo_ev[1:0]}), .prl_c0set(prl_c0set), .prl_cany0(prl_cany0), 
        .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_cpmsgid(
        prl_cpmsgid), .pff_ack(pff_ack), .prx_rst(prx_rst), .pff_obsd(pff_obsd), .pff_full(pff_full), .pff_empty(pff_empty), .ptx_ack(ptx_ack), .pff_ptr(
        pff_ptr), .prx_adpn(prx_adpn), .pff_rdat(pff_rdat), .pff_rxpart(
        pff_rxpart), .prx_rcvinf(prx_rcvinf), .ptx_fsm(ptx_fsm), .prx_fsm(
        prx_fsm), .prl_fsm(prl_fsm), .prx_setsta(prx_setsta), .clk_1p0m(
        clk_1p0m), .clk_500(clk_500), .clk(g_clk), .xrstz(i_rstz), .xclk(s_clk), .dbgpo({SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58}), .srstz(srstz), 
        .prstz(prstz), .test_si2(r_pwm[15]), .test_si1(n685), .test_so2(n51), 
        .test_so1(n684), .test_se(n10) );
  i2cslv_a0 u0_i2cslv ( .i_sda(n510), .i_scl(n508), .o_sda(slvo_sda), .i_deva(
        r_i2c_deva), .i_inc(n722), .i_fwnak(r_i2c_fwnak), .i_fwack(r_i2c_fwack), .o_we(i2c_ev_3), .o_re(slvo_re), .o_r_early(slvo_early), .o_idle(sse_idle), 
        .o_dec(), .o_busev(slvo_ev), .o_ofs(sse_adr), .o_lt_ofs(i2c_lt_ofs), 
        .o_wdat(sse_wdat), .o_lt_buf(i2c_ltbuf), .o_dbgpo({
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66}), .i_rdat(esfrm_rdat), .i_rd_mem(sse_rdrdy), .i_clk(g_clk), .i_rstz(n83), .i_prefetch(sse_prefetch), 
        .test_si(n682), .test_se(n10) );
  updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 u0_updphy ( .i_cc(n58), .i_cc_49(n123), 
        .i_sqlch(di_sqlch), .r_sqlch(r_sqlch), .r_adprx_en(r_ccrx[3]), 
        .r_adp2nd(r_ccrx[2]), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), 
        .r_fifopsh(r_fifopsh), .r_fifopop(r_fifopop), .r_fiforst(r_fiforst), 
        .r_unlock(r_unlock), .r_first(r_first), .r_last(r_last), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_rdy(upd_rdrdy), .r_wdat({n66, n64, 
        n62, n60, n57, n55, n52, sfr_wdat[0]}), .r_rdat(esfrm_rdat), 
        .r_txnumk(r_txnumk), .r_txendk(r_txendk), .r_txshrt(r_txshrt), 
        .r_auto_discard(r_auto_discard), .r_txauto(r_txauto), .r_rxords_ena(
        r_rxords_ena), .r_spec(r_spec), .r_dat_spec(r_dat_spec), 
        .r_auto_gdcrc(r_auto_gdcrc), .r_rxdb_opt(r_rxdb_opt), .r_pshords(
        r_pshords), .r_dat_portrole(r_dat_portrole), .r_dat_datarole(
        r_dat_datarole), .r_discard(r_discard), .pid_goidle(pid_goidle), 
        .pid_gobusy(pid_gobusy), .pff_ack(pff_ack), .pff_rdat(pff_rdat), 
        .pff_rxpart(pff_rxpart), .prx_rcvinf(prx_rcvinf), .pff_obsd(pff_obsd), 
        .pff_ptr(pff_ptr), .pff_empty(pff_empty), .pff_full(pff_full), 
        .ptx_ack(ptx_ack), .ptx_cc(ptx_cc), .ptx_oe(ptx_oe), .prx_setsta(
        prx_setsta), .prx_rst(prx_rst), .prl_c0set(prl_c0set), .prl_cany0(
        prl_cany0), .prl_cany0r(prl_cany0r), .prl_cany0w(prl_cany0w), 
        .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_cany0adr(
        prl_cany0adr), .prl_cpmsgid(prl_cpmsgid), .prx_fifowdat(prx_fifowdat), 
        .ptx_fsm(ptx_fsm), .prl_fsm(prl_fsm), .prx_fsm(prx_fsm), .prx_adpn(
        prx_adpn), .dbgpo({SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, upd_dbgpo, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .clk(g_clk), 
        .srstz(prstz), .test_si(bist_r_ctl[3]), .test_so(n43), .test_se(n10)
         );
  dacmux_a0 u0_dacmux ( .clk(g_clk), .srstz(n82), .i_comp(n4), .r_comp_opt(
        r_comp_opt), .r_wdat(r_dacwdat), .r_adofs(r_adofs), .r_isofs(r_isofs), 
        .r_wr({n23, r_dacwr[9:7], sfr_dacwr[14:8]}), .dacv_wr({wr_dacv[17:16], 
        n18, n15, wr_dacv[13], n14, n13, n17, n22, n16, sfr_dacwr[7:0]}), 
        .o_dacv(dac_r_vs), .o_shrst(sh_rst), .o_hold(sh_hold), .o_dac1(DAC1_V), 
        .o_daci_sel(dacmux_sel), .o_dat(dac_r_comp), .r_dac_en(r_dac_en), 
        .r_sar_en(r_sar_en), .o_dactl(dac_r_ctl), .o_cmpsta(dac_r_cmpsta), 
        .x_daclsb(x_daclsb), .o_intr(exint[7]), .o_smpl({
        SYNOPSYS_UNCONNECTED_97, comp_smpl}), .test_si2(r_vcomp[7]), 
        .test_si1(DI_GPIO[0]), .test_so1(n686), .test_se(n10) );
  fcp_a0 u0_fcp ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(1'b0), .intr(
        fcp_intr), .tx_en(fcp_oe), .tx_dat(fcp_do), .r_dat(fcp_r_dat), .r_sta(
        fcp_r_sta), .r_ctl(fcp_r_ctl), .r_msk(fcp_r_msk), .r_crc(fcp_r_crc), 
        .r_acc(fcp_r_acc), .r_dpdmsta(r_accctl), .r_wdat({n66, n64, n62, n60, 
        n57, n55, n52, n48}), .r_wr(r_fcpwr), .r_re(r_fcpre), .clk(g_clk), 
        .srstz(n83), .r_tui(fcp_r_tui), .test_si(n683), .test_so(n682), 
        .test_se(n10) );
  cvctl_a0 u0_cvctl ( .r_cvcwr(r_cvcwr), .wdat(r_cvcwdat), .r_sdischg(
        r_sdischg), .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), .r_cvofsx(r_cvofsx), .r_cvofs(r_cvofs), .sdischg_duty(sdischg_duty), .r_hlsb_en(r_pwrctl[4]), 
        .r_hlsb_sel(r_pwrctl[5]), .r_hlsb_freq(r_xtm[5]), .r_hlsb_duty(
        r_xtm[6]), .r_fw_pwrv(r_fw_pwrv), .r_dac0(DO_DAC0), .r_dac3(DAC3_V), 
        .clk_100k(clk_100k), .clk(g_clk), .srstz(n83), .test_si(d_dodat[15]), 
        .test_se(n10) );
  regx_a0 u0_regx ( .regx_r(regx_re), .regx_w(regx_we), .di_drposc(di_aswk_0), 
        .di_imposc(di_aswk[4]), .di_rd_det(di_aswk[2]), .clk_500k(clk_500k), 
        .r_imp_osc(r_imp_osc), .regx_addr({n1, xram_a[5:0]}), .regx_wdat({
        xram_d[7:2], n70, n68}), .regx_rdat(regx_rdat), .regx_hitbst(
        regx_hitbst), .regx_wrpwm(regx_wrpwm), .regx_wrcvc({r_cvcwr[2], 
        r_cvcwr[5:3]}), .r_sdischg(r_sdischg), .r_bistctl(bist_r_ctl), 
        .r_bistdat(bist_r_dat), .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), 
        .r_cvofsx(r_cvofsx), .r_pwm(r_pwm), .regx_wrdac({wr_dacv[17:16], 
        r_dacwr[10:9], wr_dacv[15:8], r_dacwr[8:7]}), .dac_r_vs(
        dac_r_vs[143:64]), .dac_comp(dac_r_comp[17:8]), .r_dac_en(
        r_dac_en[17:8]), .r_sar_en(r_sar_en[17:8]), .r_aopt(r_aopt), .r_xtm(
        r_xtm), .r_adummyi({SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, DUMMY_IN}), .r_bck0(r_bck0), .r_bck1(r_bck1), 
        .r_bck2({SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, r_bck2_2_, lg_pulse_len}), .r_i2crout({
        r_i2crout, r_i2cmcu_route, r_i2cslv_route}), .r_xana({r_xana_23, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, r_xana_19, r_xana_18, OCP_SEL, PWREN_HOLD, 
        r_xana}), .di_xanav(di_xanav), .lt_gpi(lt_gpi), .di_tst(di_tst), 
        .bkpt_pc(bkpt_pc), .bkpt_ena(bkpt_ena), .we_twlb(we_twlb), .r_vpp_en(
        r_vpp_en), .r_vpp0v_en(r_vpp0v_en), .r_otp_pwdn_en(r_otp_pwdn_en), 
        .r_otp_wpls(r_otp_wpls), .wd_twlb(wd_twlb), .r_sap(r_sap), .r_twlb(
        pmem_twlb), .upd_pwrv(r_pwrv_upd), .ramacc(ramacc), .sse_idle(sse_idle), .bus_idle(bus_idle), .r_do_ts(r_do_ts), .r_dpdo_sel(r_dpdo_sel), 
        .r_dndo_sel(r_dndo_sel), .di_ts(di_ts), .detclk(detclk), .aswclk(
        aswclk), .atpg_en(n95), .di_aswk({di_aswk[4], n1171, di_aswk[2], 1'b0, 
        di_aswk_0}), .clk(g_clk), .rrstz(n82), .test_si2(n43), .test_si1(n51), 
        .test_so1(n50), .test_se(n10) );
  srambist_a0 u0_srambist ( .clk(g_clk), .srstz(n83), .reg_hit(regx_hitbst), 
        .reg_w(regx_we), .reg_r(regx_re), .reg_wdat({xram_d[7:2], n70, n68}), 
        .iram_rdat({n129, n131, n133, n135, n138, n140, sram_rdat}), 
        .xram_rdat({n129, n131, n133, n135, n138, n140, sram_rdat}), .bist_en(
        bist_en), .bist_xram(), .bist_wr(bist_wr), .bist_adr(bist_adr), 
        .bist_wdat(bist_wdat), .o_bistctl(bist_r_ctl), .o_bistdat(bist_r_dat), 
        .test_si(n50), .test_se(n10) );
  divclk_a0 u0_divclk ( .mclk(g_clk), .srstz(n83), .atpg_en(n72), .clk_1p0m(
        clk_1p0m), .clk_500k(clk_500k), .clk_100k(clk_100k), .clk_50k(clk_50k), 
        .clk_500(clk_500), .divff_o1(divff_o1), .divff_o2(), .test_si(
        r_sar_en[17]), .test_so(n683), .test_se(n10) );
  glpwm_a0_0 u0_pwm_0_ ( .clk(g_clk), .rstz(n83), .clk_base(clk_50k), .we(
        regx_wrpwm[0]), .wdat({xram_d[7:2], n70, n68}), .r_pwm(r_pwm[7:0]), 
        .pwm_o(pwm_o[0]), .test_si(n142), .test_se(n10) );
  glpwm_a0_1 u0_pwm_1_ ( .clk(g_clk), .rstz(n82), .clk_base(clk_50k), .we(
        regx_wrpwm[1]), .wdat({xram_d[7:2], n70, n68}), .r_pwm(r_pwm[15:8]), 
        .pwm_o(pwm_o[1]), .test_si(r_pwm[7]), .test_se(n10) );
  SNPS_CLOCK_GATE_HIGH_core_a0 clk_gate_d_dodat_reg ( .CLK(g_clk), .EN(N568), 
        .ENCLK(net8853), .TE(n10) );
  DLNQX1 r_lt_gpi_reg_2_ ( .D(DI_GPIO[1]), .XG(i_rstz), .Q(r_lt_gpi[2]) );
  DLNQX1 r_lt_gpi_reg_0_ ( .D(DI_GPIO[3]), .XG(i_rstz), .Q(r_lt_gpi[0]) );
  DLNQX1 r_lt_gpi_reg_3_ ( .D(DI_GPIO[0]), .XG(i_rstz), .Q(r_lt_gpi[3]) );
  DLNQX1 r_lt_gpi_reg_1_ ( .D(DI_GPIO[2]), .XG(i_rstz), .Q(r_lt_gpi[1]) );
  SDFFQX1 d_dodat_reg_10_ ( .D(N1483), .SIN(d_dodat[9]), .SMC(n10), .C(net8853), .Q(d_dodat[10]) );
  SDFFQX1 d_dodat_reg_11_ ( .D(N1478), .SIN(d_dodat[10]), .SMC(n10), .C(
        net8853), .Q(d_dodat[11]) );
  SDFFQX1 d_dodat_reg_12_ ( .D(N572), .SIN(d_dodat[11]), .SMC(n10), .C(net8853), .Q(d_dodat[12]) );
  SDFFQX1 d_dodat_reg_15_ ( .D(N569), .SIN(d_dodat[14]), .SMC(n10), .C(net8853), .Q(d_dodat[15]) );
  SDFFQX1 d_dodat_reg_9_ ( .D(N575), .SIN(d_dodat[8]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[9]) );
  SDFFQX1 d_dodat_reg_14_ ( .D(N570), .SIN(d_dodat[13]), .SMC(n10), .C(net8853), .Q(d_dodat[14]) );
  SDFFQX1 d_dodat_reg_8_ ( .D(N576), .SIN(d_dodat[7]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[8]) );
  SDFFQX1 d_dodat_reg_13_ ( .D(N571), .SIN(d_dodat[12]), .SMC(n10), .C(net8853), .Q(d_dodat[13]) );
  SDFFQX1 d_dodat_reg_2_ ( .D(N582), .SIN(d_dodat[1]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[2]) );
  SDFFQX1 d_dodat_reg_1_ ( .D(N583), .SIN(d_dodat[0]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[1]) );
  SDFFQX1 d_dodat_reg_3_ ( .D(N581), .SIN(d_dodat[2]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[3]) );
  SDFFQX1 d_dodat_reg_0_ ( .D(N584), .SIN(n684), .SMC(n10), .C(net8853), .Q(
        d_dodat[0]) );
  SDFFQX1 d_dodat_reg_5_ ( .D(N579), .SIN(d_dodat[4]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[5]) );
  SDFFQX1 d_dodat_reg_6_ ( .D(N578), .SIN(d_dodat[5]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[6]) );
  SDFFQX1 d_dodat_reg_4_ ( .D(N580), .SIN(d_dodat[3]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[4]) );
  SDFFQX1 d_dodat_reg_7_ ( .D(N577), .SIN(d_dodat[6]), .SMC(n10), .C(net8853), 
        .Q(d_dodat[7]) );
  MUX4X1 U728 ( .D0(n226), .D1(n240), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N263), 
        .S1(N264), .Y(n562) );
  MUX4X1 U727 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N263), .S1(N264), .Y(n561) );
  MUX2X1 U726 ( .D0(n562), .D1(n561), .S(N265), .Y(DO_GPIO[1]) );
  MUX4X1 U725 ( .D0(n226), .D1(n240), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N266), 
        .S1(N267), .Y(n564) );
  MUX4X1 U724 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N266), .S1(N267), .Y(n563) );
  MUX2X1 U723 ( .D0(n564), .D1(n563), .S(N268), .Y(DO_GPIO[0]) );
  MUX4X1 U713 ( .D0(n226), .D1(n240), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N260), 
        .S1(N261), .Y(n560) );
  MUX4X1 U712 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N260), .S1(N261), .Y(n559) );
  MUX2X1 U711 ( .D0(n560), .D1(n559), .S(N262), .Y(N448) );
  MUX4X1 U710 ( .D0(n226), .D1(n240), .D2(do_p0[0]), .D3(do_p0[1]), .S0(N257), 
        .S1(N258), .Y(n558) );
  MUX4X1 U709 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N257), .S1(N258), .Y(n557) );
  INVX2 U3 ( .A(regx_rdat[1]), .Y(n182) );
  INVXL U4 ( .A(n34), .Y(memdatai[7]) );
  INVX2 U5 ( .A(regx_rdat[0]), .Y(n180) );
  INVX2 U6 ( .A(regx_rdat[4]), .Y(n188) );
  BUFX3 U7 ( .A(xram_a[6]), .Y(n1) );
  OR2X2 U8 ( .A(wr_dacv[14]), .B(wr_dacv[15]), .Y(n8) );
  MUX2IX2 U9 ( .D0(n69), .D1(n49), .S(n175), .Y(r_dacwdat[0]) );
  MUX2IX4 U10 ( .D0(n199), .D1(n61), .S(n9), .Y(r_dacwdat[4]) );
  NOR8X2 U11 ( .A(n169), .B(n173), .C(n8), .D(n172), .E(n171), .F(r_dacwr[7]), 
        .G(n170), .H(wr_dacv[13]), .Y(n9) );
  OR2X1 U12 ( .A(slvo_early), .B(slvo_re), .Y(n762) );
  NAND21X1 U13 ( .B(r_dacwr[10]), .A(n165), .Y(n172) );
  AND2X1 U14 ( .A(n176), .B(n177), .Y(sse_prefetch) );
  BUFX3 U15 ( .A(memaddr_c[6]), .Y(n44) );
  OAI211X1 U16 ( .C(n198), .D(n180), .A(n194), .B(n179), .Y(memdatai[0]) );
  INVX1 U17 ( .A(regx_rdat[2]), .Y(n184) );
  INVX1 U18 ( .A(regx_rdat[6]), .Y(n193) );
  INVX1 U19 ( .A(wr_dacv[9]), .Y(n168) );
  INVX1 U20 ( .A(r_dacwr[8]), .Y(n166) );
  AO21X1 U21 ( .B(SRAM_RDAT[6]), .C(n114), .A(n162), .Y(n131) );
  AO21X1 U22 ( .B(SRAM_RDAT[4]), .C(n110), .A(n122), .Y(n135) );
  AO21X1 U23 ( .B(SRAM_RDAT[5]), .C(n100), .A(n161), .Y(n133) );
  AO21X1 U24 ( .B(SRAM_RDAT[3]), .C(n110), .A(n143), .Y(n138) );
  AO21X1 U25 ( .B(SRAM_RDAT[7]), .C(n96), .A(n163), .Y(n129) );
  AOI21X1 U26 ( .B(n41), .C(n139), .A(n202), .Y(n2) );
  BUFXL U27 ( .A(xram_ce), .Y(n3) );
  INVX8 U28 ( .A(n29), .Y(PMEM_PGM) );
  BUFXL U29 ( .A(regx_rdat[0]), .Y(n5) );
  BUFXL U30 ( .A(regx_rdat[6]), .Y(n6) );
  NAND21X1 U31 ( .B(wr_dacv[17]), .A(n164), .Y(n173) );
  BUFXL U32 ( .A(xram_a[1]), .Y(n7) );
  INVX3 U33 ( .A(r_dacwr[9]), .Y(n165) );
  BUFXL U34 ( .A(n42), .Y(n11) );
  BUFX1 U35 ( .A(memaddr_c[4]), .Y(n42) );
  BUFXL U36 ( .A(memaddr_c[5]), .Y(n12) );
  INVXL U37 ( .A(n167), .Y(n13) );
  INVX2 U38 ( .A(wr_dacv[11]), .Y(n167) );
  NAND21X1 U39 ( .B(wr_dacv[8]), .A(n166), .Y(n171) );
  BUFXL U40 ( .A(wr_dacv[12]), .Y(n14) );
  BUFXL U41 ( .A(memaddr_c[2]), .Y(n45) );
  BUFXL U42 ( .A(wr_dacv[14]), .Y(n15) );
  BUFXL U43 ( .A(wr_dacv[8]), .Y(n16) );
  INVXL U44 ( .A(n9), .Y(n46) );
  BUFXL U45 ( .A(wr_dacv[10]), .Y(n17) );
  BUFXL U46 ( .A(wr_dacv[15]), .Y(n18) );
  BUFXL U47 ( .A(memaddr_c[3]), .Y(n19) );
  BUFXL U48 ( .A(memaddr_c[0]), .Y(n20) );
  BUFXL U49 ( .A(memaddr_c[1]), .Y(n21) );
  INVXL U50 ( .A(n168), .Y(n22) );
  BUFXL U51 ( .A(r_dacwr[10]), .Y(n23) );
  NAND21X2 U52 ( .B(wr_dacv[12]), .A(n167), .Y(n170) );
  OR2X2 U53 ( .A(wr_dacv[15]), .B(wr_dacv[14]), .Y(n174) );
  BUFX3 U54 ( .A(iram_ce), .Y(n24) );
  BUFX3 U55 ( .A(n297), .Y(PMEM_TWLB[0]) );
  NOR21XL U56 ( .B(pmem_twlb[0]), .A(atpg_en), .Y(n297) );
  BUFX3 U57 ( .A(n296), .Y(PMEM_TWLB[1]) );
  NOR21XL U58 ( .B(pmem_twlb[1]), .A(n113), .Y(n296) );
  BUFX4 U59 ( .A(n299), .Y(PMEM_SAP[0]) );
  NOR21XL U60 ( .B(r_sap[0]), .A(atpg_en), .Y(n299) );
  BUFX4 U61 ( .A(n298), .Y(PMEM_SAP[1]) );
  NOR21XL U62 ( .B(r_sap[1]), .A(n111), .Y(n298) );
  INVX1 U63 ( .A(n300), .Y(n29) );
  NOR21XL U64 ( .B(pmem_pgm), .A(n112), .Y(n300) );
  AOI221XL U65 ( .A(t_pmem_csb), .B(n962), .C(comp_smpl[1]), .D(n960), .E(
        n1131), .Y(n1130) );
  INVX2 U66 ( .A(regx_rdat[3]), .Y(n186) );
  XOR3XL U67 ( .A(SRAM_A[6]), .B(n687), .C(n31), .Y(N578) );
  NOR4XL U68 ( .A(r_cvcwr[3]), .B(r_cvcwr[2]), .C(r_cvcwr[5]), .D(r_cvcwr[4]), 
        .Y(n820) );
  INVX1 U69 ( .A(n198), .Y(n35) );
  XNOR2XL U70 ( .A(SRAM_D[2]), .B(n964), .Y(n31) );
  XOR3X1 U71 ( .A(SRAM_D[1]), .B(n688), .C(n32), .Y(N579) );
  XNOR2XL U72 ( .A(SRAM_A[5]), .B(n941), .Y(n32) );
  AO22AXL U73 ( .A(iram_d[4]), .B(iram_we), .C(xram_d[4]), .D(n217), .Y(
        SRAM_D[4]) );
  INVX1 U74 ( .A(xram_d[0]), .Y(n69) );
  OR4X1 U75 ( .A(n160), .B(n159), .C(n158), .D(n33), .Y(n688) );
  AO222XL U76 ( .A(n978), .B(TX_DAT), .C(upd_dbgpo[17]), .D(n285), .E(n953), 
        .F(n205), .Y(n33) );
  NOR21XL U77 ( .B(r_ccctl[1]), .A(n88), .Y(DO_CCCTL[1]) );
  NOR21XL U78 ( .B(r_ccctl[2]), .A(n88), .Y(DO_CCCTL[2]) );
  NOR21XL U79 ( .B(r_ccctl[3]), .A(n88), .Y(DO_CCCTL[3]) );
  NOR21XL U80 ( .B(r_aopt[1]), .A(n81), .Y(ANAOPT[1]) );
  NOR21XL U81 ( .B(r_aopt[4]), .A(n81), .Y(ANAOPT[4]) );
  NOR21XL U82 ( .B(r_xana[12]), .A(n85), .Y(ANA_REGX[12]) );
  NOR21XL U83 ( .B(r_xana[2]), .A(n85), .Y(ANA_REGX[2]) );
  NOR21XL U84 ( .B(r_xana[4]), .A(n85), .Y(ANA_REGX[4]) );
  NOR21XL U85 ( .B(r_xana[6]), .A(n86), .Y(ANA_REGX[6]) );
  NOR21XL U86 ( .B(r_xana[8]), .A(n86), .Y(ANA_REGX[8]) );
  NOR21XL U87 ( .B(r_xana[9]), .A(n86), .Y(ANA_REGX[9]) );
  NOR21XL U88 ( .B(r_cctrx[3]), .A(n89), .Y(DO_CCTRX[3]) );
  INVX1 U89 ( .A(n820), .Y(n207) );
  INVX1 U90 ( .A(n99), .Y(n79) );
  INVX1 U91 ( .A(n99), .Y(n78) );
  INVX1 U92 ( .A(n97), .Y(n77) );
  INVX1 U93 ( .A(n99), .Y(n76) );
  INVX1 U94 ( .A(n98), .Y(n75) );
  INVX1 U95 ( .A(n108), .Y(n74) );
  INVX1 U96 ( .A(n99), .Y(n80) );
  INVX1 U97 ( .A(n100), .Y(n73) );
  INVX1 U98 ( .A(n97), .Y(n87) );
  INVX1 U99 ( .A(n98), .Y(n81) );
  INVX1 U100 ( .A(n99), .Y(n85) );
  INVX1 U101 ( .A(n98), .Y(n86) );
  INVX1 U102 ( .A(n98), .Y(n88) );
  INVX1 U103 ( .A(n98), .Y(n89) );
  INVX1 U104 ( .A(n97), .Y(n90) );
  INVX1 U105 ( .A(n98), .Y(n91) );
  INVX1 U106 ( .A(n97), .Y(n92) );
  INVX1 U107 ( .A(n109), .Y(n72) );
  INVX1 U108 ( .A(n99), .Y(n94) );
  INVX1 U109 ( .A(n97), .Y(n93) );
  INVX1 U110 ( .A(n97), .Y(n95) );
  INVX1 U111 ( .A(wr_dacv[16]), .Y(n164) );
  INVX1 U112 ( .A(n197), .Y(n191) );
  INVX1 U113 ( .A(n61), .Y(n60) );
  INVX1 U114 ( .A(n59), .Y(n57) );
  NAND2X1 U115 ( .A(n287), .B(n1144), .Y(n1150) );
  INVX1 U116 ( .A(n285), .Y(n1144) );
  NAND2X1 U117 ( .A(n96), .B(n208), .Y(SRAM_CEB) );
  INVX1 U118 ( .A(n67), .Y(n66) );
  INVX1 U119 ( .A(n63), .Y(n62) );
  INVX1 U120 ( .A(n54), .Y(n53) );
  INVX1 U121 ( .A(n65), .Y(n64) );
  INVX1 U122 ( .A(n56), .Y(n55) );
  INVX1 U123 ( .A(n54), .Y(n52) );
  NOR2X1 U124 ( .A(n93), .B(n209), .Y(OSC_LOW) );
  INVX1 U125 ( .A(n49), .Y(n48) );
  INVX1 U126 ( .A(n112), .Y(n101) );
  INVX1 U127 ( .A(n113), .Y(n110) );
  INVX1 U128 ( .A(n112), .Y(n102) );
  INVX1 U129 ( .A(n111), .Y(n109) );
  INVX1 U130 ( .A(atpg_en), .Y(n108) );
  INVX1 U131 ( .A(n111), .Y(n106) );
  INVX1 U132 ( .A(n111), .Y(n107) );
  INVX1 U133 ( .A(n112), .Y(n104) );
  INVX1 U134 ( .A(atpg_en), .Y(n103) );
  INVX1 U135 ( .A(n111), .Y(n105) );
  INVX1 U136 ( .A(n112), .Y(n96) );
  INVX1 U137 ( .A(n113), .Y(n99) );
  INVX1 U138 ( .A(n113), .Y(n97) );
  INVX1 U139 ( .A(n113), .Y(n98) );
  INVX1 U140 ( .A(n112), .Y(n100) );
  NAND21X1 U141 ( .B(hit_xr), .A(n178), .Y(n197) );
  OAI22X1 U142 ( .A(n291), .B(n259), .C(n292), .D(n258), .Y(n1075) );
  INVX1 U143 ( .A(sfr_wdat[4]), .Y(n61) );
  AOI21X1 U144 ( .B(n287), .C(n37), .A(n293), .Y(n1135) );
  INVX1 U145 ( .A(sfr_wdat[0]), .Y(n49) );
  INVX1 U146 ( .A(sfr_wdat[3]), .Y(n59) );
  MUX2IX1 U148 ( .D0(n216), .D1(n56), .S(n47), .Y(r_dacwdat[2]) );
  MUX2AXL U149 ( .D0(n215), .D1(n57), .S(n47), .Y(r_dacwdat[3]) );
  MUX2AXL U150 ( .D0(n214), .D1(n62), .S(n47), .Y(r_dacwdat[5]) );
  MUX2AXL U151 ( .D0(n212), .D1(n66), .S(n47), .Y(r_dacwdat[7]) );
  MUX2AXL U152 ( .D0(n213), .D1(n64), .S(n47), .Y(r_dacwdat[6]) );
  NAND21X1 U153 ( .B(n979), .A(n148), .Y(n286) );
  NAND21X1 U154 ( .B(n973), .A(n37), .Y(n285) );
  OR4X1 U155 ( .A(n954), .B(n959), .C(n978), .D(n956), .Y(n1145) );
  NAND2X1 U156 ( .A(n200), .B(n2), .Y(n1042) );
  INVX1 U157 ( .A(n955), .Y(n287) );
  INVX1 U158 ( .A(n977), .Y(n148) );
  NAND43X1 U159 ( .B(n286), .C(n962), .D(n960), .A(n1154), .Y(n200) );
  NOR4XL U160 ( .A(n1150), .B(n1145), .C(n975), .D(n953), .Y(n1154) );
  INVX1 U161 ( .A(n1032), .Y(n226) );
  INVX1 U163 ( .A(n141), .Y(n201) );
  NAND21X1 U164 ( .B(n200), .A(n2), .Y(n141) );
  OR3XL U165 ( .A(n957), .B(n977), .C(n1145), .Y(n1163) );
  OR2X1 U166 ( .A(n959), .B(n975), .Y(n1134) );
  INVX1 U167 ( .A(n979), .Y(n151) );
  INVX1 U168 ( .A(s0_rxdoe), .Y(n288) );
  INVX1 U169 ( .A(n897), .Y(SRAM_D[7]) );
  INVX1 U170 ( .A(n899), .Y(n208) );
  OAI22X1 U171 ( .A(n67), .B(n207), .C(n820), .D(n212), .Y(r_cvcwdat[7]) );
  OAI22X1 U172 ( .A(n59), .B(n207), .C(n820), .D(n215), .Y(r_cvcwdat[3]) );
  OAI22X1 U173 ( .A(n63), .B(n207), .C(n820), .D(n214), .Y(r_cvcwdat[5]) );
  OAI22X1 U174 ( .A(n65), .B(n207), .C(n820), .D(n213), .Y(r_cvcwdat[6]) );
  OAI22X1 U175 ( .A(n56), .B(n207), .C(n820), .D(n216), .Y(r_cvcwdat[2]) );
  INVX1 U176 ( .A(sfr_wdat[7]), .Y(n67) );
  INVX1 U177 ( .A(sfr_wdat[6]), .Y(n65) );
  INVX1 U178 ( .A(sfr_wdat[1]), .Y(n54) );
  INVX1 U179 ( .A(sfr_wdat[5]), .Y(n63) );
  INVX1 U180 ( .A(sfr_wdat[2]), .Y(n56) );
  INVX1 U181 ( .A(n898), .Y(SRAM_D[0]) );
  INVX1 U182 ( .A(fcp_oe), .Y(n265) );
  XNOR2XL U183 ( .A(DO_DAC0[0]), .B(DAC3_V[5]), .Y(n942) );
  INVX1 U184 ( .A(xram_we), .Y(n217) );
  NOR2X1 U185 ( .A(n243), .B(n236), .Y(n1047) );
  INVX1 U186 ( .A(o_dodat0_15_), .Y(n209) );
  NOR2X1 U187 ( .A(n94), .B(n229), .Y(STB_RP) );
  NOR2X1 U188 ( .A(n94), .B(n230), .Y(ANAOPT[3]) );
  AOI21X1 U189 ( .B(n242), .C(n238), .A(atpg_en), .Y(CCI2C_EN) );
  NOR2X1 U190 ( .A(n93), .B(n221), .Y(DO_SRCCTL[3]) );
  NOR2X1 U191 ( .A(n92), .B(n220), .Y(DO_SRCCTL[2]) );
  NOR2X1 U192 ( .A(n92), .B(n218), .Y(BCK_REGX[2]) );
  NOR2X1 U193 ( .A(n93), .B(n219), .Y(DO_SRCCTL[0]) );
  NOR2X1 U194 ( .A(n93), .B(n211), .Y(OSC_STOP) );
  OR2X1 U195 ( .A(sh_hold), .B(n95), .Y(SH_HOLD) );
  OR2X1 U196 ( .A(n202), .B(n111), .Y(tclk_sel) );
  INVX1 U197 ( .A(n115), .Y(n112) );
  INVX1 U199 ( .A(n114), .Y(n113) );
  INVX1 U200 ( .A(n115), .Y(n111) );
  AOI221X1 U201 ( .A(regx_rdat[7]), .B(n35), .C(n129), .D(n191), .E(n36), .Y(
        n34) );
  AO21X1 U202 ( .B(ictlr_inst[7]), .C(n196), .A(n195), .Y(n36) );
  OAI211X1 U203 ( .C(n198), .D(n193), .A(n194), .B(n192), .Y(memdatai[6]) );
  AOI22X1 U204 ( .A(n191), .B(n131), .C(ictlr_inst[6]), .D(n196), .Y(n192) );
  OAI211X1 U205 ( .C(n198), .D(n188), .A(n194), .B(n187), .Y(memdatai[4]) );
  AOI22X1 U206 ( .A(n191), .B(n135), .C(ictlr_inst[4]), .D(n196), .Y(n187) );
  OAI211X1 U207 ( .C(n198), .D(n186), .A(n194), .B(n185), .Y(memdatai[3]) );
  AOI22X1 U208 ( .A(n191), .B(n138), .C(ictlr_inst[3]), .D(n196), .Y(n185) );
  OAI211X1 U209 ( .C(n198), .D(n190), .A(n194), .B(n189), .Y(memdatai[5]) );
  AOI22X1 U210 ( .A(n191), .B(n133), .C(ictlr_inst[5]), .D(n196), .Y(n189) );
  INVX2 U211 ( .A(regx_rdat[5]), .Y(n190) );
  OAI211X1 U212 ( .C(n198), .D(n184), .A(n194), .B(n183), .Y(memdatai[2]) );
  AOI22X1 U213 ( .A(n191), .B(n140), .C(ictlr_inst[2]), .D(n196), .Y(n183) );
  OAI211X1 U214 ( .C(n198), .D(n182), .A(n194), .B(n181), .Y(memdatai[1]) );
  AOI22X1 U215 ( .A(n191), .B(sram_rdat[1]), .C(ictlr_inst[1]), .D(n196), .Y(
        n181) );
  AOI22X1 U216 ( .A(n191), .B(sram_rdat[0]), .C(ictlr_inst[0]), .D(n196), .Y(
        n179) );
  INVX1 U217 ( .A(n69), .Y(n68) );
  NAND21X1 U218 ( .B(n196), .A(hit_xr), .Y(n198) );
  XNOR2XL U219 ( .A(n1012), .B(n1013), .Y(N570) );
  XNOR2XL U220 ( .A(n1014), .B(n1015), .Y(n1013) );
  XNOR2XL U221 ( .A(n1017), .B(n1018), .Y(n1012) );
  XNOR2XL U222 ( .A(DAC1_V[8]), .B(TX_EN), .Y(n1014) );
  INVX1 U223 ( .A(n194), .Y(n195) );
  INVX1 U224 ( .A(n196), .Y(n178) );
  OAI22X1 U225 ( .A(n218), .B(n1061), .C(n1062), .D(n228), .Y(n1063) );
  OAI22X1 U226 ( .A(n931), .B(n259), .C(n229), .D(n258), .Y(n1066) );
  INVX1 U227 ( .A(r_xana_19), .Y(n229) );
  XNOR2XL U228 ( .A(n999), .B(n1000), .Y(N572) );
  XNOR2XL U229 ( .A(n1001), .B(n1002), .Y(n1000) );
  XNOR2XL U230 ( .A(n210), .B(n1003), .Y(n999) );
  XNOR2XL U231 ( .A(dacmux_sel[12]), .B(DO_DAC0[7]), .Y(n1001) );
  INVX1 U232 ( .A(n137), .Y(n225) );
  AOI221XL U233 ( .A(n1095), .B(di_pro[5]), .C(n253), .D(n4), .E(n1096), .Y(
        n1093) );
  OAI22X1 U234 ( .A(n220), .B(n1097), .C(n291), .D(n254), .Y(n1096) );
  INVX1 U235 ( .A(n126), .Y(n291) );
  INVX1 U236 ( .A(n1171), .Y(n290) );
  INVX1 U237 ( .A(n128), .Y(n292) );
  OR2X1 U238 ( .A(n881), .B(di_gpio[2]), .Y(n877) );
  XNOR2XL U239 ( .A(DO_GPIO[3]), .B(SRAM_A[3]), .Y(n932) );
  XNOR2XL U240 ( .A(n926), .B(DO_GPIO[2]), .Y(n925) );
  XNOR2XL U241 ( .A(DO_GPIO[4]), .B(SRAM_A[4]), .Y(n938) );
  XNOR2XL U242 ( .A(n980), .B(n981), .Y(N577) );
  XNOR2XL U243 ( .A(n982), .B(n983), .Y(n981) );
  XOR2X1 U244 ( .A(n984), .B(n985), .Y(n980) );
  XNOR2XL U245 ( .A(DO_DAC0[2]), .B(DAC1_V[1]), .Y(n982) );
  XNOR2XL U246 ( .A(n934), .B(n935), .Y(N580) );
  XNOR2XL U247 ( .A(n936), .B(n937), .Y(n935) );
  XNOR2XL U248 ( .A(n938), .B(n939), .Y(n934) );
  XNOR2XL U249 ( .A(DAC3_V[4]), .B(n898), .Y(n936) );
  XNOR2XL U250 ( .A(n927), .B(n928), .Y(N581) );
  XNOR2XL U251 ( .A(n929), .B(n930), .Y(n928) );
  XNOR2XL U252 ( .A(n932), .B(n933), .Y(n927) );
  XNOR2XL U253 ( .A(DAC3_V[3]), .B(n931), .Y(n929) );
  XNOR2XL U254 ( .A(n921), .B(n922), .Y(N582) );
  XNOR2XL U255 ( .A(n923), .B(n924), .Y(n922) );
  XNOR2XL U256 ( .A(n925), .B(n230), .Y(n921) );
  XNOR2XL U257 ( .A(dacmux_sel[2]), .B(DO_PWR_I[2]), .Y(n924) );
  AO22X1 U258 ( .A(n979), .B(di_pro[5]), .C(n961), .D(r_osc_stop), .Y(n1149)
         );
  AOI222XL U259 ( .A(n838), .B(n839), .C(n840), .D(n841), .E(n236), .F(n842), 
        .Y(n511) );
  ENOX1 U260 ( .A(n855), .B(n856), .C(n223), .D(n855), .Y(n852) );
  AOI22AXL U261 ( .A(n857), .B(n224), .D(n857), .C(n858), .Y(n856) );
  OAI21X1 U262 ( .B(di_gpio[2]), .C(n276), .A(n859), .Y(n858) );
  NAND4X1 U263 ( .A(n850), .B(n276), .C(n225), .D(n274), .Y(n859) );
  AOI222XL U264 ( .A(n251), .B(di_sqlch), .C(n1095), .D(n205), .E(n253), .F(
        cc1_di), .Y(n1106) );
  AOI222XL U265 ( .A(n251), .B(n123), .C(n1095), .D(TX_DAT), .E(n253), .F(
        cc2_di), .Y(n1094) );
  AOI222XL U266 ( .A(n843), .B(n839), .C(n844), .D(n841), .E(n243), .F(n842), 
        .Y(n510) );
  AOI222XL U267 ( .A(n843), .B(n852), .C(n844), .D(n853), .E(n243), .F(n854), 
        .Y(n508) );
  AOI221XL U268 ( .A(n1086), .B(n128), .C(n251), .D(di_pro[2]), .E(n1107), .Y(
        n1105) );
  OAI22X1 U269 ( .A(n1101), .B(n231), .C(n221), .D(n250), .Y(n1107) );
  INVX1 U270 ( .A(n123), .Y(n293) );
  AOI222XL U271 ( .A(n838), .B(n852), .C(n840), .D(n853), .E(n236), .F(n854), 
        .Y(n509) );
  XNOR2XL U272 ( .A(n965), .B(n966), .Y(n964) );
  XNOR2XL U273 ( .A(n942), .B(n943), .Y(n941) );
  XNOR2XL U274 ( .A(r_xana_19), .B(r_srcctl[0]), .Y(n1002) );
  XNOR2XL U275 ( .A(n228), .B(dacmux_sel[11]), .Y(n1036) );
  XNOR2XL U276 ( .A(n1034), .B(n1035), .Y(N1478) );
  XNOR2XL U277 ( .A(n1037), .B(n907), .Y(n1034) );
  XNOR2XL U278 ( .A(DO_DAC0[6]), .B(n1036), .Y(n1035) );
  XNOR2XL U279 ( .A(DAC1_V[5]), .B(n897), .Y(n1037) );
  OA21X1 U280 ( .B(n233), .C(dm_comp), .A(n1119), .Y(n1118) );
  INVX1 U281 ( .A(n1170), .Y(n230) );
  NOR3XL U282 ( .A(n840), .B(n844), .C(n293), .Y(n58) );
  INVX1 U283 ( .A(n822), .Y(n162) );
  INVX1 U284 ( .A(n825), .Y(n143) );
  INVX1 U285 ( .A(n824), .Y(n122) );
  INVX1 U286 ( .A(n823), .Y(n161) );
  INVX1 U287 ( .A(n821), .Y(n163) );
  INVX1 U288 ( .A(n532), .Y(n150) );
  INVX1 U289 ( .A(n531), .Y(n147) );
  INVX1 U290 ( .A(n826), .Y(n127) );
  INVX1 U291 ( .A(n4), .Y(n149) );
  AO21X1 U292 ( .B(n124), .C(n40), .A(n161), .Y(n955) );
  AO21X1 U293 ( .B(n124), .C(n39), .A(n162), .Y(n977) );
  AO21X1 U294 ( .B(n124), .C(n146), .A(n163), .Y(n979) );
  AO21X1 U295 ( .B(n124), .C(n125), .A(n122), .Y(n953) );
  OAI21BBX1 U296 ( .A(n132), .B(n40), .C(n831), .Y(n956) );
  OAI22X1 U297 ( .A(n244), .B(n1041), .C(mcuo_scl), .D(n241), .Y(n1032) );
  OAI21BBX1 U298 ( .A(n130), .B(n40), .C(n835), .Y(n954) );
  OAI21BBX1 U299 ( .A(n125), .B(n130), .C(n836), .Y(n978) );
  OAI21BBX1 U300 ( .A(n132), .B(n146), .C(n829), .Y(n959) );
  OAI21BBX1 U301 ( .A(n132), .B(n39), .C(n830), .Y(n957) );
  OR2X1 U302 ( .A(n957), .B(n961), .Y(n975) );
  AO21X1 U303 ( .B(n144), .C(n39), .A(n127), .Y(n973) );
  NOR21XL U304 ( .B(dacmux_sel[9]), .A(n73), .Y(SAMPL_SEL[9]) );
  NOR21XL U305 ( .B(dacmux_sel[5]), .A(n73), .Y(SAMPL_SEL[5]) );
  NOR21XL U306 ( .B(dacmux_sel[8]), .A(n73), .Y(SAMPL_SEL[8]) );
  NOR21XL U307 ( .B(dacmux_sel[4]), .A(n73), .Y(SAMPL_SEL[4]) );
  NOR21XL U308 ( .B(dacmux_sel[12]), .A(n74), .Y(SAMPL_SEL[12]) );
  NOR21XL U309 ( .B(dacmux_sel[6]), .A(n73), .Y(SAMPL_SEL[6]) );
  NOR21XL U310 ( .B(dacmux_sel[7]), .A(n73), .Y(SAMPL_SEL[7]) );
  NOR21XL U311 ( .B(dacmux_sel[2]), .A(n74), .Y(SAMPL_SEL[2]) );
  NOR21XL U312 ( .B(dacmux_sel[3]), .A(n73), .Y(SAMPL_SEL[3]) );
  NOR21XL U313 ( .B(dacmux_sel[0]), .A(n74), .Y(SAMPL_SEL[0]) );
  NOR21XL U314 ( .B(dacmux_sel[13]), .A(n74), .Y(SAMPL_SEL[13]) );
  NOR21XL U315 ( .B(dacmux_sel[14]), .A(n74), .Y(SAMPL_SEL[14]) );
  NOR21XL U316 ( .B(dacmux_sel[15]), .A(n74), .Y(SAMPL_SEL[15]) );
  NOR21XL U317 ( .B(dacmux_sel[16]), .A(n74), .Y(SAMPL_SEL[16]) );
  NOR21XL U318 ( .B(dacmux_sel[17]), .A(n74), .Y(SAMPL_SEL[17]) );
  NOR21XL U319 ( .B(dacmux_sel[1]), .A(n74), .Y(SAMPL_SEL[1]) );
  AOI21X1 U320 ( .B(n146), .C(n144), .A(n143), .Y(n37) );
  NOR2X1 U321 ( .A(n1042), .B(n295), .Y(n1004) );
  INVX1 U322 ( .A(n1165), .Y(n206) );
  NOR2X1 U323 ( .A(n93), .B(n984), .Y(DO_TS[3]) );
  NOR2X1 U324 ( .A(n94), .B(n907), .Y(OE_GPIO[3]) );
  NOR2X1 U325 ( .A(n94), .B(n908), .Y(OE_GPIO[2]) );
  AND2X1 U326 ( .A(dacmux_sel[11]), .B(n100), .Y(SAMPL_SEL[11]) );
  OR2X1 U327 ( .A(n904), .B(n95), .Y(OE_GPIO[6]) );
  OR2X1 U328 ( .A(n905), .B(n95), .Y(OE_GPIO[5]) );
  INVX1 U329 ( .A(pwm_o[0]), .Y(n227) );
  NOR2X1 U330 ( .A(n93), .B(n266), .Y(SAMPL_SEL[10]) );
  OAI21BBX1 U331 ( .A(n132), .B(n125), .C(n832), .Y(n962) );
  AO21X1 U332 ( .B(n130), .C(n146), .A(n156), .Y(n960) );
  INVX1 U333 ( .A(xram_d[7]), .Y(n212) );
  INVX1 U334 ( .A(n71), .Y(n70) );
  INVX1 U335 ( .A(n1033), .Y(n240) );
  NOR2X1 U336 ( .A(n93), .B(n906), .Y(OE_GPIO[4]) );
  NOR2X1 U337 ( .A(n94), .B(n267), .Y(SH_RST) );
  INVX1 U338 ( .A(n843), .Y(n244) );
  INVX1 U339 ( .A(n838), .Y(n241) );
  XNOR2XL U340 ( .A(DAC3_V[2]), .B(n900), .Y(n923) );
  XNOR2XL U341 ( .A(DAC3_V[1]), .B(n901), .Y(n919) );
  INVX1 U342 ( .A(xram_d[2]), .Y(n216) );
  INVX1 U343 ( .A(xram_d[6]), .Y(n213) );
  INVX1 U344 ( .A(xram_d[5]), .Y(n214) );
  INVX1 U345 ( .A(xram_d[3]), .Y(n215) );
  XNOR2XL U346 ( .A(n915), .B(n916), .Y(N583) );
  XNOR2XL U347 ( .A(n917), .B(n918), .Y(n916) );
  XNOR2XL U348 ( .A(n919), .B(n920), .Y(n915) );
  XNOR2XL U349 ( .A(DO_PWR_I[1]), .B(DO_GPIO[1]), .Y(n917) );
  NOR2X1 U350 ( .A(n94), .B(n909), .Y(OE_GPIO[1]) );
  NOR2X1 U351 ( .A(n94), .B(n910), .Y(OE_GPIO[0]) );
  INVX1 U352 ( .A(n833), .Y(n156) );
  INVX1 U353 ( .A(n1016), .Y(n205) );
  XNOR2XL U354 ( .A(n902), .B(SRAM_D[6]), .Y(n1029) );
  XNOR2XL U355 ( .A(n1026), .B(n1027), .Y(N1483) );
  XNOR2XL U356 ( .A(DAC1_V[4]), .B(n1028), .Y(n1027) );
  XNOR2XL U357 ( .A(n1029), .B(n908), .Y(n1026) );
  XNOR2XL U358 ( .A(DO_DAC0[5]), .B(n266), .Y(n1028) );
  INVX1 U359 ( .A(n952), .Y(TX_DAT) );
  NOR2X1 U360 ( .A(n273), .B(n274), .Y(n880) );
  INVX1 U361 ( .A(n900), .Y(SRAM_A[2]) );
  INVX1 U362 ( .A(n901), .Y(SRAM_A[1]) );
  AO22XL U363 ( .A(xram_a[4]), .B(xram_ce), .C(iram_a[4]), .D(iram_ce), .Y(
        SRAM_A[4]) );
  XNOR2XL U364 ( .A(n899), .B(n904), .Y(n1017) );
  XNOR2XL U365 ( .A(SRAM_A[7]), .B(SRAM_D[3]), .Y(n985) );
  XNOR2XL U366 ( .A(SRAM_D[5]), .B(SRAM_A[9]), .Y(n996) );
  XNOR2XL U367 ( .A(SRAM_A[8]), .B(SRAM_D[4]), .Y(n990) );
  XNOR2XL U368 ( .A(n911), .B(n912), .Y(N584) );
  XNOR2XL U369 ( .A(DO_PWR_I[0]), .B(n914), .Y(n911) );
  XNOR2XL U370 ( .A(n903), .B(n913), .Y(n912) );
  XNOR2XL U371 ( .A(dacmux_sel[16]), .B(dacmux_sel[0]), .Y(n914) );
  XNOR2XL U372 ( .A(n986), .B(n987), .Y(N576) );
  XNOR2XL U373 ( .A(n988), .B(n989), .Y(n987) );
  XOR2X1 U374 ( .A(n910), .B(n990), .Y(n986) );
  XNOR2XL U375 ( .A(DO_DAC0[3]), .B(DAC1_V[2]), .Y(n988) );
  XNOR2XL U376 ( .A(n992), .B(n993), .Y(N575) );
  XNOR2XL U377 ( .A(n994), .B(n995), .Y(n993) );
  XOR2X1 U378 ( .A(n909), .B(n996), .Y(n992) );
  XNOR2XL U379 ( .A(DO_DAC0[4]), .B(DAC1_V[3]), .Y(n994) );
  AOI22X1 U380 ( .A(xram_d[7]), .B(xram_we), .C(iram_we), .D(iram_d[7]), .Y(
        n897) );
  ENOX1 U381 ( .A(n213), .B(n217), .C(iram_d[6]), .D(iram_we), .Y(SRAM_D[6])
         );
  NOR2X1 U382 ( .A(xram_ce), .B(n24), .Y(n899) );
  INVX1 U383 ( .A(n902), .Y(SRAM_A[10]) );
  INVX1 U384 ( .A(n903), .Y(SRAM_A[0]) );
  OAI22X1 U385 ( .A(n54), .B(n207), .C(n820), .D(n71), .Y(r_cvcwdat[1]) );
  ENOX1 U386 ( .A(n214), .B(n217), .C(iram_d[5]), .D(iram_we), .Y(SRAM_D[5])
         );
  XNOR2XL U387 ( .A(dacmux_sel[6]), .B(DO_PWR_I[6]), .Y(n966) );
  XNOR2XL U388 ( .A(dacmux_sel[5]), .B(DO_PWR_I[5]), .Y(n943) );
  OAI22X1 U389 ( .A(n207), .B(n49), .C(n820), .D(n69), .Y(r_cvcwdat[0]) );
  OAI22X1 U390 ( .A(n207), .B(n61), .C(n820), .D(n199), .Y(r_cvcwdat[4]) );
  INVXL U391 ( .A(xram_d[4]), .Y(n199) );
  ENOX1 U392 ( .A(n215), .B(n217), .C(iram_d[3]), .D(iram_we), .Y(SRAM_D[3])
         );
  XNOR2XL U393 ( .A(dacmux_sel[7]), .B(DO_PWR_I[7]), .Y(n983) );
  XNOR2XL U394 ( .A(dacmux_sel[4]), .B(DO_PWR_I[4]), .Y(n937) );
  XNOR2XL U395 ( .A(dacmux_sel[3]), .B(DO_PWR_I[3]), .Y(n930) );
  XNOR2XL U396 ( .A(n1005), .B(n1006), .Y(N571) );
  XNOR2XL U397 ( .A(n1009), .B(n1010), .Y(n1005) );
  XNOR2XL U398 ( .A(n1007), .B(n1008), .Y(n1006) );
  XNOR2XL U399 ( .A(n235), .B(n905), .Y(n1009) );
  XNOR2XL U400 ( .A(n1019), .B(n1020), .Y(N569) );
  XNOR2XL U401 ( .A(n1023), .B(n1024), .Y(n1019) );
  XNOR2XL U402 ( .A(n1021), .B(n1022), .Y(n1020) );
  XNOR2XL U403 ( .A(n1025), .B(n952), .Y(n1023) );
  XNOR2XL U404 ( .A(dacmux_sel[1]), .B(dacmux_sel[17]), .Y(n918) );
  XNOR2XL U405 ( .A(r_srcctl[1]), .B(dacmux_sel[13]), .Y(n1008) );
  XNOR2XL U406 ( .A(o_dodat0_15_), .B(dacmux_sel[15]), .Y(n1022) );
  XNOR2XL U407 ( .A(r_srcctl[3]), .B(dacmux_sel[8]), .Y(n989) );
  XNOR2XL U408 ( .A(dacmux_sel[14]), .B(DO_DAC0[9]), .Y(n1015) );
  XNOR2XL U409 ( .A(r_srcctl[2]), .B(dacmux_sel[9]), .Y(n995) );
  AOI22XL U410 ( .A(n68), .B(xram_we), .C(iram_d[0]), .D(iram_we), .Y(n898) );
  ENOX1 U411 ( .A(n216), .B(n217), .C(iram_d[2]), .D(iram_we), .Y(SRAM_D[2])
         );
  ENOX1 U412 ( .A(n71), .B(n217), .C(iram_d[1]), .D(iram_we), .Y(SRAM_D[1]) );
  NOR2X1 U413 ( .A(n93), .B(n210), .Y(DO_VOOC[0]) );
  NOR21XL U414 ( .B(n1018), .A(n90), .Y(DO_VOOC[2]) );
  OAI22X1 U415 ( .A(n1041), .B(n242), .C(mcuo_scl), .D(n238), .Y(n1166) );
  INVX1 U416 ( .A(n933), .Y(CC1_DOB) );
  INVX1 U417 ( .A(r_osc_gate), .Y(n289) );
  NOR2X1 U418 ( .A(sh_hold), .B(n267), .Y(N568) );
  INVX1 U419 ( .A(di_gpio[0]), .Y(n223) );
  INVX1 U420 ( .A(r_srcctl[2]), .Y(n220) );
  INVX1 U421 ( .A(r_srcctl[3]), .Y(n221) );
  INVX1 U422 ( .A(di_gpio[1]), .Y(n224) );
  INVX1 U423 ( .A(n840), .Y(n238) );
  INVX1 U424 ( .A(n844), .Y(n242) );
  NOR21XL U425 ( .B(n1010), .A(n91), .Y(DO_VOOC[1]) );
  INVX1 U426 ( .A(r_osc_stop), .Y(n211) );
  INVX1 U427 ( .A(r_srcctl[0]), .Y(n219) );
  OAI32X1 U428 ( .A(n254), .B(n263), .C(n284), .D(n250), .E(n264), .Y(n1111)
         );
  OAI22X1 U429 ( .A(n1041), .B(n1080), .C(mcuo_scl), .D(n1081), .Y(n1046) );
  OAI22X1 U430 ( .A(n219), .B(n1101), .C(n250), .D(n272), .Y(n1100) );
  INVX1 U431 ( .A(n926), .Y(n218) );
  AND2X1 U432 ( .A(n1025), .B(n100), .Y(DO_VOOC[3]) );
  INVX1 U433 ( .A(n1097), .Y(n251) );
  INVX1 U434 ( .A(n1112), .Y(n235) );
  INVX1 U435 ( .A(n1101), .Y(n253) );
  INVX1 U436 ( .A(n1095), .Y(n250) );
  INVX1 U437 ( .A(n1058), .Y(n258) );
  INVX1 U438 ( .A(n1059), .Y(n259) );
  INVX1 U439 ( .A(n1081), .Y(n236) );
  INVX1 U440 ( .A(n1080), .Y(n243) );
  INVX1 U441 ( .A(n1086), .Y(n254) );
  OAI21X1 U442 ( .B(xram_we), .C(iram_we), .A(n102), .Y(SRAM_WEB) );
  OR2X1 U443 ( .A(iram_we), .B(xram_we), .Y(n1024) );
  INVX1 U444 ( .A(n1062), .Y(n261) );
  INVX1 U445 ( .A(n1061), .Y(n260) );
  INVX1 U446 ( .A(n939), .Y(CC2_DOB) );
  NOR2X1 U447 ( .A(n1016), .B(n92), .Y(TX_EN) );
  NAND2X1 U448 ( .A(n228), .B(n96), .Y(RD_ENB) );
  NOR21XL U449 ( .B(PWRDN), .A(n263), .Y(VPP_0V) );
  XNOR2XL U450 ( .A(DO_GPIO[0]), .B(DAC3_V[0]), .Y(n913) );
  NOR2X1 U451 ( .A(n284), .B(n92), .Y(PWRDN) );
  NOR2X1 U452 ( .A(n93), .B(n931), .Y(BCK_REGX[5]) );
  NOR2X1 U453 ( .A(n94), .B(n1112), .Y(ANAOPT[5]) );
  NOR2X1 U454 ( .A(n92), .B(n920), .Y(DO_SRCCTL[4]) );
  XNOR2XL U455 ( .A(DO_DAC0[1]), .B(DAC1_V[0]), .Y(n965) );
  NAND2X1 U456 ( .A(n272), .B(n96), .Y(SLEEP) );
  NOR2X1 U457 ( .A(n92), .B(n264), .Y(BCK_REGX[4]) );
  XNOR2XL U458 ( .A(DO_DAC0[8]), .B(DAC1_V[7]), .Y(n1007) );
  XNOR2XL U459 ( .A(DO_DAC0[10]), .B(DAC1_V[9]), .Y(n1021) );
  XNOR2XL U460 ( .A(DAC1_V[6]), .B(n906), .Y(n1003) );
  AND2XL U461 ( .A(n762), .B(n177), .Y(i2c_ev_6_) );
  INVX1 U462 ( .A(n851), .Y(n275) );
  INVX1 U463 ( .A(n860), .Y(n276) );
  NOR21XL U464 ( .B(r_srcctl[1]), .A(n90), .Y(DO_SRCCTL[1]) );
  OR2X2 U465 ( .A(pmem_csb), .B(n95), .Y(PMEM_CSB) );
  INVX1 U466 ( .A(n812), .Y(n139) );
  NAND2X1 U467 ( .A(n1152), .B(n204), .Y(n812) );
  INVX1 U468 ( .A(n136), .Y(n202) );
  NAND32X1 U469 ( .B(n204), .C(n134), .A(n41), .Y(n136) );
  INVX1 U470 ( .A(n1152), .Y(n134) );
  INVX1 U471 ( .A(n1153), .Y(n144) );
  INVX1 U472 ( .A(atpg_en), .Y(n114) );
  INVX1 U473 ( .A(atpg_en), .Y(n115) );
  NOR2X1 U474 ( .A(n94), .B(n203), .Y(lt_gpi[3]) );
  NOR2X1 U475 ( .A(n94), .B(n204), .Y(lt_gpi[0]) );
  NAND2X1 U476 ( .A(n283), .B(n115), .Y(OCDRV_ENZ) );
  INVX1 U477 ( .A(n998), .Y(n294) );
  NAND43X1 U478 ( .B(n155), .C(n154), .D(n153), .A(n152), .Y(n687) );
  AO2222XL U479 ( .A(do_p0[6]), .B(n201), .C(mcu_dbgpo[17]), .D(n975), .E(
        fcp_oe), .F(n956), .G(r_accctl[4]), .H(n954), .Y(n154) );
  OA2222XL U480 ( .A(n151), .B(n150), .C(n287), .D(n149), .E(n293), .F(n37), 
        .G(n148), .H(n147), .Y(n152) );
  AO2222XL U481 ( .A(n978), .B(r_ccctl[0]), .C(n953), .D(TX_DAT), .E(
        mcu_dbgpo[16]), .F(n959), .G(n58), .H(n973), .Y(n153) );
  AO222X1 U482 ( .A(comp_smpl[3]), .B(n960), .C(pmem_pgm), .D(n962), .E(x_clk), 
        .F(n202), .Y(n155) );
  AO2222XL U483 ( .A(r_dpdmctl[6]), .B(n954), .C(mcu_dbgpo[22]), .D(n959), .E(
        di_pro[2]), .F(n286), .G(fcp_do), .H(n956), .Y(n159) );
  AO2222XL U484 ( .A(mcu_dbgpo[19]), .B(n957), .C(n201), .D(n157), .E(n955), 
        .F(dp_comp), .G(o_dodat0_15_), .H(n961), .Y(n158) );
  AO222X1 U485 ( .A(comp_smpl[2]), .B(n960), .C(pmem_re), .D(n962), .E(i_rstz), 
        .F(n202), .Y(n160) );
  NAND42X1 U486 ( .C(r_pg0_sel[1]), .D(r_pg0_sel[0]), .A(r_pg0_sel[3]), .B(
        r_pg0_sel[2]), .Y(n176) );
  INVX1 U487 ( .A(sse_adr[7]), .Y(n177) );
  NAND3X1 U488 ( .A(n1128), .B(n1129), .C(n1130), .Y(DO_GPIO[4]) );
  AOI222XL U489 ( .A(slvo_sda), .B(n953), .C(n205), .D(n978), .E(upd_dbgpo[18]), .F(n973), .Y(n1128) );
  AOI221XL U490 ( .A(n201), .B(n1133), .C(mcu_dbgpo[18]), .D(n1134), .E(n1135), 
        .Y(n1129) );
  OAI21BBX1 U491 ( .A(SRAM_RDAT[0]), .B(n114), .C(n828), .Y(sram_rdat[0]) );
  OAI21BBX1 U492 ( .A(SRAM_RDAT[1]), .B(n96), .C(n827), .Y(sram_rdat[1]) );
  AO21X1 U493 ( .B(SRAM_RDAT[2]), .C(n110), .A(n127), .Y(n140) );
  AND2X1 U494 ( .A(r_vpp0v_en), .B(ps_pwrdn), .Y(pwrdn_rst) );
  NAND3X1 U495 ( .A(n1138), .B(n1139), .C(n1140), .Y(DO_GPIO[3]) );
  AOI22X1 U496 ( .A(cc2_di), .B(n953), .C(mcu_dbgpo[21]), .D(n1145), .Y(n1138)
         );
  AOI221XL U497 ( .A(n123), .B(n955), .C(prx_rcvinf[4]), .D(n285), .E(n1142), 
        .Y(n1139) );
  AOI221XL U498 ( .A(r_vpp_en), .B(n962), .C(comp_smpl[0]), .D(n960), .E(n1141), .Y(n1140) );
  AO21X1 U499 ( .B(mempsrd), .C(hit_ps), .A(n178), .Y(n194) );
  OAI21X1 U500 ( .B(hit_xd), .C(hit_xr), .A(memrd), .Y(n196) );
  OAI21BBX1 U501 ( .A(DI_GPIO[3]), .B(n106), .C(n825), .Y(n137) );
  OAI21BBX1 U502 ( .A(DRP_OSC), .B(n105), .C(n829), .Y(di_aswk_0) );
  OAI221X1 U503 ( .A(r_dpdo_sel[3]), .B(n1048), .C(n1049), .D(n262), .E(n1050), 
        .Y(n1018) );
  NAND4X1 U504 ( .A(n255), .B(n262), .C(n257), .D(n1051), .Y(n1050) );
  AOI22X1 U505 ( .A(r_dpdo_sel[2]), .B(n1068), .C(n1069), .D(n255), .Y(n1048)
         );
  AOI22X1 U506 ( .A(r_dpdo_sel[2]), .B(n1054), .C(n1055), .D(n255), .Y(n1049)
         );
  OAI22AX1 U507 ( .D(n882), .C(n883), .A(n223), .B(n882), .Y(exint[0]) );
  NAND3X1 U508 ( .A(n282), .B(n281), .C(N268), .Y(n882) );
  AOI22AXL U509 ( .A(n884), .B(n885), .D(n885), .C(di_gpio[1]), .Y(n883) );
  NAND3X1 U510 ( .A(n280), .B(n279), .C(N265), .Y(n885) );
  INVX1 U511 ( .A(r_xana_18), .Y(n228) );
  OAI22X1 U512 ( .A(n1056), .B(n257), .C(r_dpdo_sel[1]), .D(n1057), .Y(n1055)
         );
  AOI221XL U513 ( .A(n1058), .B(pwm_o[0]), .C(n1059), .D(pwm_o[1]), .E(n1060), 
        .Y(n1057) );
  AOI221XL U514 ( .A(n1058), .B(di_aswk[2]), .C(r_bck0[3]), .D(n1059), .E(
        n1063), .Y(n1056) );
  OAI22X1 U515 ( .A(n211), .B(n1061), .C(n209), .D(n1062), .Y(n1060) );
  OAI22X1 U516 ( .A(n1064), .B(n257), .C(r_dpdo_sel[1]), .D(n1065), .Y(n1054)
         );
  AOI221XL U517 ( .A(n261), .B(n1170), .C(r_srcctl[5]), .D(n260), .E(n1067), 
        .Y(n1064) );
  AOI221XL U518 ( .A(n261), .B(di_aswk[4]), .C(n260), .D(di_aswk_0), .E(n1066), 
        .Y(n1065) );
  OAI22X1 U519 ( .A(n920), .B(n259), .C(n264), .D(n258), .Y(n1067) );
  ENOX1 U520 ( .A(n886), .B(n887), .C(di_gpio[2]), .D(n886), .Y(n884) );
  NOR32XL U521 ( .B(n277), .C(N262), .A(N261), .Y(n886) );
  NOR4XL U522 ( .A(N258), .B(N257), .C(n137), .D(n273), .Y(n887) );
  OAI21BBX1 U523 ( .A(SRCI[1]), .B(n104), .C(n836), .Y(n126) );
  OAI21BBX1 U524 ( .A(DM_FAULT), .B(n103), .C(n832), .Y(n1171) );
  NOR21XL U525 ( .B(bist_r_ctl[5]), .A(n73), .Y(SRAM_OEB) );
  OAI21BBX1 U526 ( .A(SRCI[0]), .B(n104), .C(n821), .Y(n128) );
  NAND42X1 U527 ( .C(N258), .D(n137), .A(n880), .B(n881), .Y(n878) );
  OAI21BBX1 U528 ( .A(DI_GPIO[2]), .B(n106), .C(n826), .Y(di_gpio[2]) );
  OAI21BBX1 U529 ( .A(IMP_OSC), .B(n107), .C(n822), .Y(di_aswk[4]) );
  OAI22X1 U530 ( .A(n888), .B(n248), .C(r_i2crout[5]), .D(n889), .Y(dpdm_urx)
         );
  AOI22AXL U531 ( .A(r_pwrctl[7]), .B(n247), .D(r_pwrctl[7]), .C(n890), .Y(
        n888) );
  AOI22X1 U532 ( .A(r_pwrctl[6]), .B(n247), .C(n890), .D(n269), .Y(n889) );
  INVX1 U533 ( .A(n854), .Y(n247) );
  OAI22AX1 U534 ( .D(n875), .C(n876), .A(n223), .B(n875), .Y(exint[1]) );
  NAND3X1 U535 ( .A(N266), .B(n281), .C(N268), .Y(n875) );
  AOI32X1 U536 ( .A(n877), .B(n878), .C(n879), .D(n278), .E(di_gpio[1]), .Y(
        n876) );
  INVX1 U537 ( .A(n879), .Y(n278) );
  OAI31XL U538 ( .A(n861), .B(o_cpurst), .C(hit_ps), .D(n862), .Y(mempsack) );
  NOR2X1 U539 ( .A(mempsrd), .B(mempswr), .Y(n861) );
  NAND2X1 U540 ( .A(ictlr_psack), .B(hit_ps), .Y(n862) );
  AOI22BXL U541 ( .B(n891), .A(n223), .D(n892), .C(n891), .Y(n890) );
  AOI22AXL U542 ( .A(n893), .B(n894), .D(n894), .C(n224), .Y(n892) );
  OAI21X1 U543 ( .B(di_gpio[2]), .C(n895), .A(n896), .Y(n893) );
  NAND4X1 U544 ( .A(N258), .B(n880), .C(n895), .D(n225), .Y(n896) );
  OAI22X1 U545 ( .A(n1073), .B(n257), .C(r_dpdo_sel[1]), .D(n1074), .Y(n1068)
         );
  AOI221XL U546 ( .A(n1058), .B(n531), .C(n1059), .D(di_pro[5]), .E(n1076), 
        .Y(n1073) );
  AOI221XL U547 ( .A(n261), .B(n532), .C(n260), .D(di_pro[2]), .E(n1075), .Y(
        n1074) );
  OAI22X1 U548 ( .A(n231), .B(n1061), .C(n290), .D(n1062), .Y(n1076) );
  AOI22X1 U549 ( .A(r_dndo_sel[3]), .B(n1091), .C(n1092), .D(n256), .Y(n1084)
         );
  OAI22X1 U550 ( .A(n1098), .B(n249), .C(r_dndo_sel[2]), .D(n1099), .Y(n1091)
         );
  OAI22X1 U551 ( .A(n1093), .B(n249), .C(r_dndo_sel[2]), .D(n1094), .Y(n1092)
         );
  AOI221XL U552 ( .A(n1086), .B(pwm_o[1]), .C(n251), .D(o_dodat0_15_), .E(
        n1100), .Y(n1099) );
  INVX1 U553 ( .A(n1082), .Y(n210) );
  OAI221X1 U554 ( .A(r_dpdmctl[0]), .B(n1083), .C(n1084), .D(n270), .E(n1085), 
        .Y(n1082) );
  INVX1 U555 ( .A(r_dpdmctl[0]), .Y(n270) );
  OAI211X1 U556 ( .C(fcp_do), .D(n265), .A(n1086), .B(n1087), .Y(n1085) );
  XNOR2XL U557 ( .A(n1169), .B(r_aopt[3]), .Y(n1170) );
  NAND2X1 U558 ( .A(r_imp_osc), .B(di_aswk[4]), .Y(n1169) );
  GEN2XL U559 ( .D(n1113), .E(n1114), .C(n1115), .B(r_do_ts[6]), .A(n1116), 
        .Y(n984) );
  AOI21X1 U560 ( .B(n1119), .C(di_pro[5]), .A(n233), .Y(n1113) );
  AOI211X1 U561 ( .C(r_do_ts[4]), .D(n1117), .A(n232), .B(n1118), .Y(n1116) );
  AOI22X1 U562 ( .A(r_do_ts[4]), .B(n1126), .C(n1121), .D(n531), .Y(n1114) );
  OAI21BBX1 U563 ( .A(SRCI[3]), .B(n110), .C(n834), .Y(n532) );
  AO21X1 U564 ( .B(SRCI[4]), .C(n110), .A(n156), .Y(n531) );
  OAI21BBX1 U565 ( .A(DAC1_COMP), .B(n104), .C(n836), .Y(n4) );
  OAI21BBX1 U566 ( .A(RX_DAT), .B(n103), .C(n835), .Y(n123) );
  AO222X1 U567 ( .A(n954), .B(r_dpdmctl[4]), .C(n956), .D(dm_comp), .E(n286), 
        .F(n126), .Y(n1131) );
  OAI21BBX1 U568 ( .A(CC2_DI), .B(n103), .C(n830), .Y(cc2_di) );
  OAI21BBX1 U569 ( .A(CC1_DI), .B(n102), .C(n831), .Y(cc1_di) );
  OAI21BBX1 U570 ( .A(SRCI[5]), .B(n102), .C(n832), .Y(di_pro[5]) );
  OAI21BBX1 U571 ( .A(SRCI[2]), .B(n105), .C(n835), .Y(di_pro[2]) );
  OAI21BBX1 U572 ( .A(DM_COMP), .B(n103), .C(n829), .Y(dm_comp) );
  OAI21BBX1 U573 ( .A(RD_DET), .B(n105), .C(n830), .Y(di_aswk[2]) );
  OAI21BBX1 U574 ( .A(RX_SQL), .B(n103), .C(n834), .Y(di_sqlch) );
  ENOX1 U575 ( .A(n845), .B(n846), .C(n223), .D(n845), .Y(n839) );
  AOI22AXL U576 ( .A(n847), .B(n224), .D(n847), .C(n848), .Y(n846) );
  OAI21X1 U577 ( .B(di_gpio[2]), .C(n275), .A(n849), .Y(n848) );
  NAND4X1 U578 ( .A(N257), .B(n850), .C(n275), .D(n225), .Y(n849) );
  NAND3X1 U579 ( .A(n1146), .B(n1147), .C(n1148), .Y(DO_GPIO[2]) );
  AOI22X1 U580 ( .A(di_sqlch), .B(n1150), .C(N448), .D(n1042), .Y(n1147) );
  AOI22X1 U581 ( .A(mcu_dbgpo[20]), .B(n1163), .C(cc1_di), .D(n953), .Y(n1146)
         );
  AOI221XL U582 ( .A(t_pmem_clk), .B(n962), .C(n4), .D(n960), .E(n1149), .Y(
        n1148) );
  OAI22X1 U583 ( .A(n1070), .B(n257), .C(r_dpdo_sel[1]), .D(n1071), .Y(n1069)
         );
  AOI22X1 U584 ( .A(n261), .B(n123), .C(n260), .D(di_sqlch), .Y(n1071) );
  AOI221XL U585 ( .A(n261), .B(cc2_di), .C(n260), .D(cc1_di), .E(n1072), .Y(
        n1070) );
  OAI22X1 U586 ( .A(n952), .B(n259), .C(n1016), .D(n258), .Y(n1072) );
  AOI221XL U587 ( .A(n1086), .B(r_vpp_en), .C(n251), .D(di_aswk[4]), .E(n1102), 
        .Y(n1098) );
  OAI22X1 U588 ( .A(n939), .B(n1101), .C(n920), .D(n250), .Y(n1102) );
  AOI221XL U589 ( .A(n1121), .B(di_xanav[0]), .C(n1119), .D(di_xanav[1]), .E(
        n1124), .Y(n1115) );
  OAI21BX1 U590 ( .C(r_do_ts[4]), .B(n1125), .A(n233), .Y(n1124) );
  AOI22X1 U591 ( .A(n126), .B(n234), .C(r_do_ts[3]), .D(n532), .Y(n1125) );
  AOI22X1 U592 ( .A(r_dndo_sel[3]), .B(n1103), .C(n1104), .D(n256), .Y(n1083)
         );
  OAI22X1 U593 ( .A(n1108), .B(n249), .C(r_dndo_sel[2]), .D(n1109), .Y(n1103)
         );
  OAI22X1 U594 ( .A(n1105), .B(n249), .C(r_dndo_sel[2]), .D(n1106), .Y(n1104)
         );
  AOI221XL U595 ( .A(n253), .B(CC1_DOB), .C(n235), .D(n251), .E(n1111), .Y(
        n1108) );
  AO22AXL U596 ( .A(n975), .B(mcu_dbgpo[16]), .C(n286), .D(n292), .Y(n1141) );
  ENOX1 U597 ( .A(n290), .B(n234), .C(n234), .D(t_pmem_clk), .Y(n1126) );
  NAND21X1 U598 ( .B(n101), .A(d_dodat[0]), .Y(n828) );
  NAND21X1 U599 ( .B(n115), .A(d_dodat[4]), .Y(n824) );
  NAND21X1 U600 ( .B(n101), .A(d_dodat[1]), .Y(n827) );
  NAND21X1 U601 ( .B(n114), .A(d_dodat[5]), .Y(n823) );
  NAND21X1 U602 ( .B(n101), .A(d_dodat[3]), .Y(n825) );
  NAND21X1 U603 ( .B(n101), .A(d_dodat[6]), .Y(n822) );
  NAND21X1 U604 ( .B(n102), .A(d_dodat[7]), .Y(n821) );
  AO21X1 U605 ( .B(DP_COMP), .C(n110), .A(n156), .Y(dp_comp) );
  OAI21BBX1 U606 ( .A(XANAV[0]), .B(n104), .C(n828), .Y(di_xanav[0]) );
  OAI21BBX1 U607 ( .A(XANAV[1]), .B(n104), .C(n827), .Y(di_xanav[1]) );
  INVX1 U608 ( .A(n1120), .Y(n232) );
  AOI31X1 U609 ( .A(r_do_ts[5]), .B(dp_comp), .C(n1121), .D(r_do_ts[6]), .Y(
        n1120) );
  NAND21X1 U610 ( .B(n101), .A(d_dodat[2]), .Y(n826) );
  OAI22X1 U611 ( .A(dp_comp), .B(n248), .C(r_i2crout[5]), .D(dm_comp), .Y(n854) );
  OAI22X1 U612 ( .A(r_i2crout[5]), .B(dp_comp), .C(dm_comp), .D(n248), .Y(n842) );
  OAI22X1 U613 ( .A(r_i2crout[4]), .B(cc2_di), .C(cc1_di), .D(n246), .Y(n853)
         );
  OAI22X1 U614 ( .A(cc2_di), .B(n246), .C(r_i2crout[4]), .D(cc1_di), .Y(n841)
         );
  XOR2X1 U615 ( .A(do_p0[5]), .B(pwm_o[1]), .Y(n157) );
  OAI21BBX1 U616 ( .A(DI_GPIO[5]), .B(n106), .C(n823), .Y(di_gpio[5]) );
  OAI21BBX1 U617 ( .A(DI_GPIO[6]), .B(n106), .C(n822), .Y(di_gpio[6]) );
  OAI21BBX1 U618 ( .A(DI_TS), .B(n106), .C(n831), .Y(di_ts) );
  INVX1 U619 ( .A(dacmux_sel[10]), .Y(n266) );
  INVX1 U620 ( .A(n118), .Y(n146) );
  NAND32X1 U621 ( .B(n204), .C(n117), .A(n206), .Y(n118) );
  INVX1 U622 ( .A(r_lt_gpi[1]), .Y(n117) );
  OAI211X1 U623 ( .C(r_gpio_tm), .D(di_tst), .A(n102), .B(i_rstz), .Y(n1165)
         );
  NOR21XL U624 ( .B(n1042), .A(n1143), .Y(n1142) );
  AOI22X1 U625 ( .A(n558), .B(n273), .C(n557), .D(N259), .Y(n1143) );
  NAND32X1 U626 ( .B(r_gpio_oe[5]), .C(n1004), .A(n2), .Y(n905) );
  NAND32X1 U627 ( .B(r_gpio_oe[6]), .C(n1004), .A(n2), .Y(n904) );
  XNOR2XL U628 ( .A(do_p0[4]), .B(n227), .Y(n1133) );
  NAND2X1 U629 ( .A(n38), .B(n834), .Y(n961) );
  NAND4X1 U630 ( .A(r_lt_gpi[1]), .B(n204), .C(n130), .D(n206), .Y(n38) );
  OAI21X1 U631 ( .B(n1004), .C(n1038), .A(n998), .Y(n907) );
  AND2X1 U632 ( .A(n1039), .B(r_gpio_oe[3]), .Y(n1038) );
  AOI32X1 U633 ( .A(n880), .B(n288), .C(N258), .D(n850), .E(n1040), .Y(n1039)
         );
  OAI22X1 U634 ( .A(N257), .B(n1032), .C(n274), .D(n1033), .Y(n1040) );
  OAI21X1 U635 ( .B(n1004), .C(n1030), .A(n998), .Y(n908) );
  AOI221XL U636 ( .A(n240), .B(n851), .C(n226), .D(n860), .E(n1031), .Y(n1030)
         );
  OAI21X1 U637 ( .B(s0_rxdoe), .C(n895), .A(r_gpio_oe[2]), .Y(n1031) );
  NOR2X1 U638 ( .A(n1165), .B(r_lt_gpi[1]), .Y(n1164) );
  OAI22X1 U639 ( .A(n1122), .B(n233), .C(r_do_ts[5]), .D(n1123), .Y(n1117) );
  AOI22X1 U640 ( .A(divff_o1), .B(n234), .C(r_do_ts[3]), .D(x_clk), .Y(n1123)
         );
  AOI22X1 U641 ( .A(pwm_o[0]), .B(n234), .C(r_do_ts[3]), .D(pwm_o[1]), .Y(
        n1122) );
  INVX1 U642 ( .A(n120), .Y(n125) );
  NAND21X1 U643 ( .B(r_lt_gpi[0]), .A(n1164), .Y(n120) );
  OAI21BBX1 U644 ( .A(XANAV[2]), .B(n107), .C(n826), .Y(di_xanav[2]) );
  OAI21BBX1 U645 ( .A(XANAV[3]), .B(n107), .C(n825), .Y(di_xanav[3]) );
  OAI21BBX1 U646 ( .A(XANAV[4]), .B(n107), .C(n824), .Y(di_xanav[4]) );
  OAI21BBX1 U647 ( .A(XANAV[5]), .B(n107), .C(n823), .Y(di_xanav[5]) );
  OAI21X1 U648 ( .B(pmem_pgm), .C(hwi2c_stretch), .A(r_strtch), .Y(n1041) );
  AND3X1 U649 ( .A(r_lt_gpi[1]), .B(n204), .C(n206), .Y(n39) );
  AND2X1 U650 ( .A(n1164), .B(r_lt_gpi[0]), .Y(n40) );
  OAI22X1 U651 ( .A(slvo_sda), .B(n244), .C(mcuo_sda), .D(n241), .Y(n1033) );
  NOR2X1 U652 ( .A(r_i2cmcu_route[0]), .B(r_i2cmcu_route[1]), .Y(n838) );
  NOR2X1 U653 ( .A(r_i2cslv_route[0]), .B(r_i2cslv_route[1]), .Y(n843) );
  NAND2X1 U654 ( .A(d_dodat[14]), .B(n91), .Y(n830) );
  NAND2X1 U655 ( .A(d_dodat[15]), .B(n92), .Y(n829) );
  NAND2X1 U656 ( .A(d_dodat[13]), .B(n92), .Y(n831) );
  NAND2X1 U657 ( .A(d_dodat[9]), .B(n92), .Y(n835) );
  NAND2X1 U658 ( .A(d_dodat[8]), .B(n92), .Y(n836) );
  NOR2X1 U659 ( .A(n1004), .B(r_gpio_oe[4]), .Y(n906) );
  INVX1 U660 ( .A(xram_d[1]), .Y(n71) );
  INVX1 U661 ( .A(sh_rst), .Y(n267) );
  NAND21X1 U662 ( .B(n115), .A(d_dodat[10]), .Y(n834) );
  NAND21X1 U663 ( .B(n101), .A(d_dodat[12]), .Y(n832) );
  NAND21X1 U664 ( .B(n110), .A(d_dodat[11]), .Y(n833) );
  NOR2XL U665 ( .A(ptx_oe), .B(r_fortxen), .Y(n1016) );
  NOR2X1 U666 ( .A(n239), .B(r_i2cmcu_route[1]), .Y(n840) );
  NOR2X1 U667 ( .A(n245), .B(r_i2cslv_route[1]), .Y(n844) );
  OAI211X1 U668 ( .C(s0_rxdoe), .D(n891), .A(r_gpio_oe[0]), .B(n991), .Y(n910)
         );
  AOI221XL U669 ( .A(n226), .B(n855), .C(n240), .D(n845), .E(n294), .Y(n991)
         );
  OAI211X1 U670 ( .C(s0_rxdoe), .D(n894), .A(r_gpio_oe[1]), .B(n997), .Y(n909)
         );
  AOI221XL U671 ( .A(n226), .B(n857), .C(n240), .D(n847), .E(n294), .Y(n997)
         );
  INVX1 U672 ( .A(r_i2cmcu_route[0]), .Y(n239) );
  INVX1 U673 ( .A(r_i2cslv_route[0]), .Y(n245) );
  MUX2IX1 U674 ( .D0(ptx_cc), .D1(r_fortxdat), .S(r_fortxrdy), .Y(n952) );
  AOI22X1 U675 ( .A(xram_a[10]), .B(n3), .C(iram_a[10]), .D(iram_ce), .Y(n902)
         );
  NOR3XL U676 ( .A(N261), .B(N262), .C(N260), .Y(n860) );
  NOR3XL U677 ( .A(N261), .B(N262), .C(n277), .Y(n851) );
  INVX1 U678 ( .A(N257), .Y(n274) );
  INVX1 U679 ( .A(r_do_ts[3]), .Y(n234) );
  INVX1 U680 ( .A(N260), .Y(n277) );
  NOR3XL U681 ( .A(N267), .B(N268), .C(n282), .Y(n845) );
  INVX1 U682 ( .A(N259), .Y(n273) );
  INVX1 U683 ( .A(N266), .Y(n282) );
  NAND3X1 U684 ( .A(N262), .B(N260), .C(N261), .Y(n895) );
  INVX1 U685 ( .A(r_do_ts[5]), .Y(n233) );
  NOR2X1 U686 ( .A(r_do_ts[3]), .B(r_do_ts[4]), .Y(n1121) );
  NOR2X1 U687 ( .A(n234), .B(r_do_ts[4]), .Y(n1119) );
  AOI22XL U688 ( .A(xram_a[0]), .B(n3), .C(iram_a[0]), .D(n24), .Y(n903) );
  AO22X1 U689 ( .A(xram_a[7]), .B(xram_ce), .C(iram_a[7]), .D(iram_ce), .Y(
        SRAM_A[7]) );
  AO22X1 U690 ( .A(xram_ce), .B(xram_a[9]), .C(iram_ce), .D(iram_a[9]), .Y(
        SRAM_A[9]) );
  AO22X1 U691 ( .A(xram_a[8]), .B(xram_ce), .C(iram_a[8]), .D(iram_ce), .Y(
        SRAM_A[8]) );
  NOR2X1 U692 ( .A(N258), .B(N259), .Y(n850) );
  NOR3XL U693 ( .A(N264), .B(N265), .C(n280), .Y(n847) );
  NOR3XL U694 ( .A(N264), .B(N265), .C(N263), .Y(n857) );
  NOR3XL U695 ( .A(N267), .B(N268), .C(N266), .Y(n855) );
  INVX1 U696 ( .A(N263), .Y(n280) );
  NAND3X1 U697 ( .A(N268), .B(N266), .C(N267), .Y(n891) );
  NAND3X1 U698 ( .A(N265), .B(N263), .C(N264), .Y(n894) );
  NOR21XL U699 ( .B(r_do_ts[2]), .A(n90), .Y(DO_TS[2]) );
  OR2X1 U700 ( .A(r_gpio_ie[1]), .B(n95), .Y(GPIO_IE[1]) );
  AOI221XL U701 ( .A(t_osc_gate), .B(n1095), .C(n253), .D(n926), .E(n1110), 
        .Y(n1109) );
  OAI22X1 U702 ( .A(n211), .B(n1097), .C(n227), .D(n254), .Y(n1110) );
  OAI22X1 U703 ( .A(n246), .B(n1166), .C(r_i2crout[4]), .D(n1167), .Y(n933) );
  OAI21BBX1 U704 ( .A(DI_GPIO[1]), .B(n105), .C(n827), .Y(di_gpio[1]) );
  OAI22X1 U705 ( .A(r_i2crout[4]), .B(n1166), .C(n246), .D(n1167), .Y(n939) );
  NOR21XL U706 ( .B(esfrm_rrdy), .A(prl_cany0), .Y(sse_rdrdy) );
  OAI21BBX1 U707 ( .A(DI_GPIO[0]), .B(n105), .C(n828), .Y(di_gpio[0]) );
  OAI22X1 U708 ( .A(slvo_sda), .B(n242), .C(mcuo_sda), .D(n238), .Y(n1167) );
  INVX1 U714 ( .A(r_pwrdn), .Y(n284) );
  NAND31X1 U715 ( .C(r_otpi_gate), .A(n1127), .B(r_srcctl[4]), .Y(n920) );
  NAND21X1 U716 ( .B(sdischg_duty), .A(r_sdischg[6]), .Y(n1127) );
  NAND21X1 U717 ( .B(r_bck0[2]), .A(n1168), .Y(n926) );
  NAND21X1 U718 ( .B(r_bck2_2_), .A(gating_pwr), .Y(n1168) );
  OAI21BBX1 U719 ( .A(r_xtm[7]), .B(n283), .C(r_aopt[5]), .Y(n1112) );
  NOR2X1 U720 ( .A(r_dndo_sel[0]), .B(r_dndo_sel[1]), .Y(n1086) );
  NOR2X1 U721 ( .A(n252), .B(r_dndo_sel[0]), .Y(n1095) );
  NOR2X1 U722 ( .A(r_dpdo_sel[0]), .B(r_dpdmctl[2]), .Y(n1058) );
  NOR2X1 U729 ( .A(n271), .B(r_dpdo_sel[0]), .Y(n1059) );
  OAI221X1 U730 ( .A(r_pwrctl[7]), .B(n1043), .C(r_i2crout[5]), .D(n237), .E(
        n1044), .Y(n1025) );
  INVX1 U731 ( .A(n1045), .Y(n237) );
  OAI21X1 U732 ( .B(s0_rxdoe), .C(n248), .A(r_pwrctl[7]), .Y(n1044) );
  AOI22X1 U733 ( .A(r_i2crout[5]), .B(n1046), .C(r_dpdmctl[3]), .D(n1047), .Y(
        n1043) );
  NAND2X1 U734 ( .A(r_dndo_sel[0]), .B(r_dndo_sel[1]), .Y(n1101) );
  NAND2X1 U735 ( .A(r_dpdo_sel[0]), .B(r_dpdmctl[2]), .Y(n1062) );
  NAND2X1 U736 ( .A(r_dpdo_sel[0]), .B(n271), .Y(n1061) );
  NAND2X1 U737 ( .A(r_i2cmcu_route[1]), .B(n239), .Y(n1081) );
  NAND2X1 U738 ( .A(r_dndo_sel[0]), .B(n252), .Y(n1097) );
  NAND2X1 U739 ( .A(r_i2cslv_route[1]), .B(n245), .Y(n1080) );
  INVX1 U740 ( .A(r_ocdrv_enz), .Y(n283) );
  OAI211X1 U741 ( .C(r_pwrctl[6]), .D(n1077), .A(n265), .B(n1078), .Y(n1010)
         );
  AOI22X1 U742 ( .A(r_pwrctl[6]), .B(n1079), .C(r_i2crout[5]), .D(n1045), .Y(
        n1078) );
  AOI22X1 U743 ( .A(n1046), .B(n248), .C(r_dpdmctl[1]), .D(n1047), .Y(n1077)
         );
  NAND2X1 U744 ( .A(n288), .B(n248), .Y(n1079) );
  INVX1 U745 ( .A(r_dpdmctl[2]), .Y(n271) );
  NOR2X1 U746 ( .A(r_bck0[5]), .B(frc_lg_on), .Y(n931) );
  INVX1 U747 ( .A(r_i2crout[4]), .Y(n246) );
  INVX1 U748 ( .A(r_dndo_sel[1]), .Y(n252) );
  AOI211X1 U749 ( .C(n1088), .D(n265), .A(r_dndo_sel[3]), .B(r_dndo_sel[2]), 
        .Y(n1087) );
  OAI21BBX1 U750 ( .A(n1089), .B(r_pwrctl[6]), .C(n1090), .Y(n1088) );
  OAI22X1 U751 ( .A(n248), .B(do_opt[6]), .C(do_opt[7]), .D(r_i2crout[5]), .Y(
        n1089) );
  OAI21BBX1 U752 ( .A(n1047), .B(r_dpdmctl[0]), .C(n269), .Y(n1090) );
  INVX1 U753 ( .A(r_bck0[4]), .Y(n264) );
  INVX1 U754 ( .A(r_sleep), .Y(n272) );
  OAI22X1 U755 ( .A(slvo_sda), .B(n1080), .C(mcuo_sda), .D(n1081), .Y(n1045)
         );
  INVX1 U756 ( .A(r_i2crout[5]), .Y(n248) );
  AOI211X1 U757 ( .C(r_pwrctl[7]), .D(n1052), .A(r_dpdo_sel[0]), .B(n1053), 
        .Y(n1051) );
  OAI22X1 U758 ( .A(do_opt[7]), .B(n248), .C(r_i2crout[5]), .D(do_opt[6]), .Y(
        n1052) );
  AOI21X1 U759 ( .B(r_dpdmctl[2]), .C(n1047), .A(r_pwrctl[7]), .Y(n1053) );
  INVX1 U760 ( .A(r_vpp0v_en), .Y(n263) );
  INVX1 U761 ( .A(r_pwrctl[6]), .Y(n269) );
  INVX1 U762 ( .A(PWREN_HOLD), .Y(n231) );
  AND2X1 U763 ( .A(esfrm_rrdy), .B(prl_cany0), .Y(upd_rdrdy) );
  INVX1 U764 ( .A(r_dpdo_sel[1]), .Y(n257) );
  INVX1 U765 ( .A(r_dndo_sel[2]), .Y(n249) );
  INVX1 U766 ( .A(r_dpdo_sel[2]), .Y(n255) );
  INVX1 U767 ( .A(r_dndo_sel[3]), .Y(n256) );
  INVX1 U768 ( .A(r_dpdo_sel[3]), .Y(n262) );
  NOR21XL U769 ( .B(r_vpp_en), .A(n73), .Y(VPP_SEL) );
  NOR21XL U770 ( .B(r_srcctl[5]), .A(n90), .Y(DO_SRCCTL[5]) );
  NOR21XL U771 ( .B(r_dpdmctl[6]), .A(n89), .Y(DO_DPDN[3]) );
  NOR21XL U772 ( .B(r_regtrm[0]), .A(n111), .Y(REGTRM[0]) );
  NOR21XL U773 ( .B(r_regtrm[1]), .A(n79), .Y(REGTRM[1]) );
  NOR21XL U774 ( .B(r_regtrm[2]), .A(n78), .Y(REGTRM[2]) );
  NOR21XL U775 ( .B(r_regtrm[3]), .A(n77), .Y(REGTRM[3]) );
  NOR21XL U776 ( .B(r_regtrm[4]), .A(n76), .Y(REGTRM[4]) );
  NOR21XL U777 ( .B(r_regtrm[5]), .A(n75), .Y(REGTRM[5]) );
  NOR21XL U778 ( .B(r_regtrm[6]), .A(n75), .Y(REGTRM[6]) );
  NOR21XL U779 ( .B(r_regtrm[7]), .A(n75), .Y(REGTRM[7]) );
  NOR21XL U780 ( .B(r_regtrm[8]), .A(n75), .Y(REGTRM[8]) );
  NOR21XL U781 ( .B(r_regtrm[9]), .A(n74), .Y(REGTRM[9]) );
  NOR21XL U782 ( .B(r_regtrm[10]), .A(n111), .Y(REGTRM[10]) );
  NOR21XL U783 ( .B(r_regtrm[11]), .A(atpg_en), .Y(REGTRM[11]) );
  NOR21XL U784 ( .B(r_regtrm[12]), .A(n111), .Y(REGTRM[12]) );
  NOR21XL U785 ( .B(r_regtrm[13]), .A(n79), .Y(REGTRM[13]) );
  NOR21XL U786 ( .B(r_regtrm[14]), .A(n79), .Y(REGTRM[14]) );
  NOR21XL U787 ( .B(r_regtrm[15]), .A(n79), .Y(REGTRM[15]) );
  NOR21XL U788 ( .B(r_regtrm[16]), .A(n79), .Y(REGTRM[16]) );
  NOR21XL U789 ( .B(r_regtrm[17]), .A(n79), .Y(REGTRM[17]) );
  NOR21XL U790 ( .B(r_regtrm[18]), .A(n79), .Y(REGTRM[18]) );
  NOR21XL U791 ( .B(r_regtrm[19]), .A(n79), .Y(REGTRM[19]) );
  NOR21XL U792 ( .B(r_regtrm[20]), .A(n79), .Y(REGTRM[20]) );
  NOR21XL U793 ( .B(r_regtrm[21]), .A(n79), .Y(REGTRM[21]) );
  NOR21XL U794 ( .B(r_regtrm[22]), .A(n78), .Y(REGTRM[22]) );
  NOR21XL U795 ( .B(r_regtrm[23]), .A(n78), .Y(REGTRM[23]) );
  NOR21XL U796 ( .B(r_regtrm[40]), .A(n76), .Y(REGTRM[40]) );
  NOR21XL U797 ( .B(r_regtrm[41]), .A(n89), .Y(REGTRM[41]) );
  NOR21XL U798 ( .B(r_regtrm[42]), .A(n76), .Y(REGTRM[42]) );
  NOR21XL U799 ( .B(r_regtrm[43]), .A(n76), .Y(REGTRM[43]) );
  NOR21XL U800 ( .B(r_regtrm[44]), .A(n76), .Y(REGTRM[44]) );
  NOR21XL U801 ( .B(r_regtrm[45]), .A(n76), .Y(REGTRM[45]) );
  NOR21XL U802 ( .B(r_regtrm[46]), .A(n76), .Y(REGTRM[46]) );
  NOR21XL U803 ( .B(r_regtrm[47]), .A(n76), .Y(REGTRM[47]) );
  NOR21XL U804 ( .B(r_regtrm[48]), .A(n76), .Y(REGTRM[48]) );
  NOR21XL U805 ( .B(r_regtrm[49]), .A(n76), .Y(REGTRM[49]) );
  NOR21XL U806 ( .B(r_regtrm[50]), .A(n75), .Y(REGTRM[50]) );
  NOR21XL U807 ( .B(r_regtrm[51]), .A(n75), .Y(REGTRM[51]) );
  NOR21XL U808 ( .B(r_regtrm[52]), .A(n75), .Y(REGTRM[52]) );
  NOR21XL U809 ( .B(r_regtrm[53]), .A(n75), .Y(REGTRM[53]) );
  NOR21XL U810 ( .B(r_regtrm[54]), .A(n75), .Y(REGTRM[54]) );
  NOR21XL U811 ( .B(r_regtrm[55]), .A(n75), .Y(REGTRM[55]) );
  NOR21XL U812 ( .B(r_sdischg[7]), .A(n80), .Y(LDO3P9V) );
  NOR21XL U813 ( .B(r_srcctl[6]), .A(n90), .Y(DO_SRCCTL[6]) );
  NOR21XL U814 ( .B(r_srcctl[7]), .A(n91), .Y(DO_SRCCTL[7]) );
  NOR21XL U815 ( .B(r_dpdmctl[5]), .A(n89), .Y(DO_DPDN[2]) );
  NOR21XL U816 ( .B(r_dpdmctl[7]), .A(n89), .Y(DO_DPDN[4]) );
  NOR21XL U817 ( .B(r_xtm[0]), .A(n73), .Y(XTM[0]) );
  NOR21XL U818 ( .B(r_xtm[1]), .A(n72), .Y(XTM[1]) );
  NOR21XL U819 ( .B(r_ccctl[7]), .A(n88), .Y(DO_CCCTL[7]) );
  NOR21XL U820 ( .B(r_ccctl[6]), .A(n88), .Y(DO_CCCTL[6]) );
  NOR21XL U821 ( .B(r_ccctl[4]), .A(n88), .Y(DO_CCCTL[4]) );
  NOR21XL U822 ( .B(r_ccctl[5]), .A(n88), .Y(DO_CCCTL[5]) );
  NOR21XL U823 ( .B(r_xana[0]), .A(n81), .Y(ANA_REGX[0]) );
  NOR21XL U824 ( .B(r_accctl[4]), .A(n89), .Y(DO_DPDN[0]) );
  NOR21XL U825 ( .B(r_bck0[3]), .A(n87), .Y(BCK_REGX[3]) );
  NOR21XL U826 ( .B(r_xana[15]), .A(n85), .Y(ANA_REGX[15]) );
  NOR21XL U827 ( .B(r_xana[13]), .A(n85), .Y(ANA_REGX[13]) );
  NOR21XL U828 ( .B(r_xana[14]), .A(n85), .Y(ANA_REGX[14]) );
  NOR21XL U829 ( .B(r_xana[1]), .A(n85), .Y(ANA_REGX[1]) );
  NOR21XL U830 ( .B(r_xana[3]), .A(n85), .Y(ANA_REGX[3]) );
  NOR21XL U831 ( .B(r_regtrm[24]), .A(n78), .Y(REGTRM[24]) );
  NOR21XL U832 ( .B(r_regtrm[25]), .A(n78), .Y(REGTRM[25]) );
  NOR21XL U833 ( .B(r_regtrm[26]), .A(n78), .Y(REGTRM[26]) );
  NOR21XL U834 ( .B(r_regtrm[27]), .A(n78), .Y(REGTRM[27]) );
  NOR21XL U835 ( .B(r_regtrm[28]), .A(n78), .Y(REGTRM[28]) );
  NOR21XL U836 ( .B(r_regtrm[29]), .A(n78), .Y(REGTRM[29]) );
  NOR21XL U837 ( .B(r_regtrm[30]), .A(n78), .Y(REGTRM[30]) );
  NOR21XL U838 ( .B(r_regtrm[31]), .A(n77), .Y(REGTRM[31]) );
  NOR21XL U839 ( .B(r_regtrm[32]), .A(n77), .Y(REGTRM[32]) );
  NOR21XL U840 ( .B(r_regtrm[33]), .A(n77), .Y(REGTRM[33]) );
  NOR21XL U841 ( .B(r_regtrm[34]), .A(n77), .Y(REGTRM[34]) );
  NOR21XL U842 ( .B(r_regtrm[35]), .A(n77), .Y(REGTRM[35]) );
  NOR21XL U843 ( .B(r_regtrm[36]), .A(n77), .Y(REGTRM[36]) );
  NOR21XL U844 ( .B(r_regtrm[37]), .A(n77), .Y(REGTRM[37]) );
  NOR21XL U845 ( .B(r_regtrm[38]), .A(n77), .Y(REGTRM[38]) );
  NOR21XL U846 ( .B(r_regtrm[39]), .A(n77), .Y(REGTRM[39]) );
  NOR21XL U847 ( .B(r_aopt[0]), .A(n81), .Y(ANAOPT[0]) );
  NOR21XL U848 ( .B(r_aopt[2]), .A(n81), .Y(ANAOPT[2]) );
  NOR21XL U849 ( .B(r_aopt[6]), .A(n81), .Y(ANAOPT[6]) );
  NOR21XL U850 ( .B(r_aopt[7]), .A(n81), .Y(ANAOPT[7]) );
  NOR21XL U851 ( .B(r_accctl[3]), .A(n90), .Y(DO_DPDN[5]) );
  NOR21XL U852 ( .B(r_xana[5]), .A(n85), .Y(ANA_REGX[5]) );
  NOR21XL U853 ( .B(r_ana_tm[0]), .A(n86), .Y(ANA_TM[0]) );
  NOR21XL U854 ( .B(r_ana_tm[1]), .A(n86), .Y(ANA_TM[1]) );
  NOR21XL U855 ( .B(r_ana_tm[2]), .A(n86), .Y(ANA_TM[2]) );
  NOR21XL U856 ( .B(r_ana_tm[3]), .A(n86), .Y(ANA_TM[3]) );
  NOR21XL U859 ( .B(r_xana[7]), .A(n86), .Y(ANA_REGX[7]) );
  NOR21XL U860 ( .B(r_xana_23), .A(n80), .Y(LFOSC_ENB) );
  NOR21XL U861 ( .B(r_xana[10]), .A(n81), .Y(ANA_REGX[10]) );
  NOR21XL U862 ( .B(r_xana[11]), .A(n85), .Y(ANA_REGX[11]) );
  NOR21XL U863 ( .B(x_daclsb[2]), .A(n88), .Y(DAC1_EN) );
  NOR21XL U864 ( .B(r_cctrx[7]), .A(n89), .Y(DO_CCTRX[7]) );
  NOR21XL U865 ( .B(r_cctrx[6]), .A(n89), .Y(DO_CCTRX[6]) );
  NOR21XL U866 ( .B(r_cctrx[5]), .A(n89), .Y(DO_CCTRX[5]) );
  NOR21XL U867 ( .B(r_cctrx[4]), .A(n89), .Y(DO_CCTRX[4]) );
  NOR21XL U868 ( .B(r_xtm[2]), .A(n72), .Y(XTM[2]) );
  NOR21XL U869 ( .B(r_xtm[3]), .A(n72), .Y(XTM[3]) );
  NOR21XL U870 ( .B(r_cctrx[0]), .A(n88), .Y(DO_CCTRX[0]) );
  NOR21XL U871 ( .B(r_bck0[7]), .A(n87), .Y(BCK_REGX[7]) );
  NOR21XL U872 ( .B(r_bck1[7]), .A(n87), .Y(BCK_REGX[15]) );
  NOR21XL U873 ( .B(r_bck1[6]), .A(n87), .Y(BCK_REGX[14]) );
  NOR21XL U874 ( .B(r_bck1[5]), .A(n87), .Y(BCK_REGX[13]) );
  NOR21XL U875 ( .B(r_bck1[4]), .A(n87), .Y(BCK_REGX[12]) );
  NOR21XL U876 ( .B(r_bck1[3]), .A(n87), .Y(BCK_REGX[11]) );
  NOR21XL U877 ( .B(r_bck1[2]), .A(n86), .Y(BCK_REGX[10]) );
  NOR21XL U878 ( .B(r_bck1[0]), .A(n87), .Y(BCK_REGX[8]) );
  NOR21XL U879 ( .B(r_bck1[1]), .A(n88), .Y(BCK_REGX[9]) );
  NOR21XL U880 ( .B(r_bck0[6]), .A(n87), .Y(BCK_REGX[6]) );
  NOR21XL U881 ( .B(r_bck0[1]), .A(n87), .Y(BCK_REGX[1]) );
  NOR21XL U882 ( .B(r_bck0[0]), .A(n86), .Y(BCK_REGX[0]) );
  AND2X1 U883 ( .A(r_dpdmctl[4]), .B(n100), .Y(DO_DPDN[1]) );
  OR2XL U884 ( .A(mcu_ram_r), .B(mcu_ram_w), .Y(ramacc) );
  NOR2X1 U885 ( .A(n93), .B(n268), .Y(DO_CCCTL[0]) );
  INVX1 U886 ( .A(r_ccctl[0]), .Y(n268) );
  OR2X1 U887 ( .A(r_cctrx[2]), .B(n95), .Y(DO_CCTRX[2]) );
  OR2X1 U888 ( .A(r_cctrx[1]), .B(n95), .Y(DO_CCTRX[1]) );
  OR2X1 U889 ( .A(r_gpio_ie[0]), .B(n95), .Y(GPIO_IE[0]) );
  INVX1 U890 ( .A(sfr_intr[2]), .Y(n723) );
  NOR21XL U891 ( .B(i2c_ev_3), .A(sse_adr[7]), .Y(i2c_ev_2) );
  NAND32X1 U892 ( .B(N261), .C(n277), .A(N262), .Y(n881) );
  NAND3X1 U893 ( .A(N263), .B(n279), .C(N265), .Y(n879) );
  INVX1 U894 ( .A(N264), .Y(n279) );
  INVX1 U895 ( .A(N267), .Y(n281) );
  OAI21BBX1 U896 ( .A(PMEM_Q1[7]), .B(n114), .C(n821), .Y(pmem_q1[7]) );
  OAI21BBX1 U897 ( .A(PMEM_Q0[7]), .B(n108), .C(n829), .Y(pmem_q0[7]) );
  OAI21BBX1 U898 ( .A(PMEM_Q1[1]), .B(n109), .C(n827), .Y(pmem_q1[1]) );
  OAI21BBX1 U899 ( .A(PMEM_Q0[1]), .B(n107), .C(n835), .Y(pmem_q0[1]) );
  OAI21BBX1 U900 ( .A(PMEM_Q1[5]), .B(n109), .C(n823), .Y(pmem_q1[5]) );
  OAI21BBX1 U901 ( .A(PMEM_Q0[5]), .B(n108), .C(n831), .Y(pmem_q0[5]) );
  OAI21BBX1 U902 ( .A(PMEM_Q0[3]), .B(n105), .C(n833), .Y(pmem_q0[3]) );
  OAI21BBX1 U903 ( .A(PMEM_Q1[3]), .B(n109), .C(n825), .Y(pmem_q1[3]) );
  OAI21BBX1 U904 ( .A(PMEM_Q1[6]), .B(n115), .C(n822), .Y(pmem_q1[6]) );
  OAI21BBX1 U905 ( .A(PMEM_Q0[6]), .B(n108), .C(n830), .Y(pmem_q0[6]) );
  OAI21BBX1 U906 ( .A(PMEM_Q1[2]), .B(n109), .C(n826), .Y(pmem_q1[2]) );
  OAI21BBX1 U907 ( .A(PMEM_Q0[2]), .B(n104), .C(n834), .Y(pmem_q0[2]) );
  OAI21BBX1 U908 ( .A(PMEM_Q1[0]), .B(n108), .C(n828), .Y(pmem_q1[0]) );
  OAI21BBX1 U909 ( .A(PMEM_Q0[0]), .B(n103), .C(n836), .Y(pmem_q0[0]) );
  OAI21BBX1 U910 ( .A(PMEM_Q1[4]), .B(n109), .C(n824), .Y(pmem_q1[4]) );
  OAI21BBX1 U911 ( .A(PMEM_Q0[4]), .B(n108), .C(n832), .Y(pmem_q0[4]) );
  INVX1 U912 ( .A(r_i2c_ninc), .Y(n722) );
  INVX1 U913 ( .A(sfr_intr[3]), .Y(n724) );
  OAI21BBX1 U914 ( .A(t_di_gpio4), .B(n106), .C(n824), .Y(di_gpio[4]) );
  NOR21X2 U915 ( .B(pmem_re), .A(n113), .Y(PMEM_RE) );
  NOR21X1 U916 ( .B(pmem_clk[0]), .A(n80), .Y(PMEM_CLK[0]) );
  NOR21X1 U917 ( .B(pmem_clk[1]), .A(n80), .Y(PMEM_CLK[1]) );
  NOR21XL U918 ( .B(di_tst), .A(n812), .Y(tm_atpg) );
  NOR21XL U919 ( .B(r_do_ts[1]), .A(n91), .Y(DO_TS[1]) );
  NOR21XL U920 ( .B(r_do_ts[0]), .A(n90), .Y(DO_TS[0]) );
  NOR21XL U921 ( .B(r_pu_gpio[6]), .A(n80), .Y(GPIO_PU[6]) );
  NOR21XL U922 ( .B(r_pu_gpio[5]), .A(n80), .Y(GPIO_PU[5]) );
  NOR21XL U923 ( .B(r_pu_gpio[4]), .A(n80), .Y(GPIO_PU[4]) );
  NOR21XL U924 ( .B(r_pd_gpio[3]), .A(n91), .Y(GPIO_PD[3]) );
  NOR21XL U925 ( .B(r_pd_gpio[2]), .A(n91), .Y(GPIO_PD[2]) );
  NOR21XL U926 ( .B(r_pd_gpio[1]), .A(n90), .Y(GPIO_PD[1]) );
  NOR21XL U927 ( .B(r_pd_gpio[0]), .A(n91), .Y(GPIO_PD[0]) );
  NOR21XL U928 ( .B(r_pd_gpio[6]), .A(n81), .Y(GPIO_PD[6]) );
  NOR21XL U929 ( .B(r_pd_gpio[5]), .A(n90), .Y(GPIO_PD[5]) );
  NOR21XL U930 ( .B(r_pd_gpio[4]), .A(n90), .Y(GPIO_PD[4]) );
  NOR21XL U931 ( .B(r_pu_gpio[3]), .A(n80), .Y(GPIO_PU[3]) );
  NOR21XL U932 ( .B(r_pu_gpio[2]), .A(n80), .Y(GPIO_PU[2]) );
  NOR21XL U933 ( .B(r_pu_gpio[1]), .A(n80), .Y(GPIO_PU[1]) );
  NOR21XL U934 ( .B(r_pu_gpio[0]), .A(n81), .Y(GPIO_PU[0]) );
  NAND21X1 U935 ( .B(r_lt_gpi[2]), .A(n203), .Y(n1153) );
  NOR21XL U936 ( .B(r_lt_gpi[1]), .A(n72), .Y(lt_gpi[1]) );
  NOR21XL U937 ( .B(r_lt_gpi[2]), .A(n72), .Y(lt_gpi[2]) );
  NOR2X1 U938 ( .A(n1153), .B(r_lt_gpi[1]), .Y(n1152) );
  NAND2X1 U939 ( .A(di_tst), .B(n295), .Y(n998) );
  INVX1 U940 ( .A(r_lt_gpi[0]), .Y(n204) );
  INVX1 U941 ( .A(r_lt_gpi[3]), .Y(n203) );
  INVX1 U942 ( .A(n116), .Y(n130) );
  NAND21X1 U943 ( .B(r_lt_gpi[2]), .A(r_lt_gpi[3]), .Y(n116) );
  INVX1 U944 ( .A(n121), .Y(n124) );
  NAND21X1 U945 ( .B(r_lt_gpi[3]), .A(r_lt_gpi[2]), .Y(n121) );
  INVX1 U946 ( .A(n119), .Y(n132) );
  NAND21X1 U947 ( .B(n203), .A(r_lt_gpi[2]), .Y(n119) );
  AND2X1 U948 ( .A(di_tst), .B(n114), .Y(n41) );
  INVX1 U949 ( .A(i_rstz), .Y(n295) );
  NAND21X1 U950 ( .B(wr_dacv[10]), .A(n168), .Y(n169) );
  NOR8X2 U951 ( .A(n169), .B(n173), .C(n174), .D(n172), .E(n171), .F(
        r_dacwr[7]), .G(n170), .H(wr_dacv[13]), .Y(n175) );
  AOI22XL U952 ( .A(xram_a[2]), .B(xram_ce), .C(iram_a[2]), .D(iram_ce), .Y(
        n900) );
  AO22XL U953 ( .A(xram_ce), .B(xram_a[5]), .C(iram_a[5]), .D(iram_ce), .Y(
        SRAM_A[5]) );
  AO22XL U954 ( .A(n1), .B(n3), .C(iram_a[6]), .D(n24), .Y(SRAM_A[6]) );
  INVXL U955 ( .A(n46), .Y(n47) );
  AO22XL U956 ( .A(xram_a[3]), .B(xram_ce), .C(iram_a[3]), .D(iram_ce), .Y(
        SRAM_A[3]) );
  AOI22XL U957 ( .A(n7), .B(xram_ce), .C(iram_a[1]), .D(iram_ce), .Y(n901) );
  MUX2XL U958 ( .D0(n70), .D1(n53), .S(n47), .Y(r_dacwdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_core_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_1 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o, test_si, 
        test_se );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we, test_si, test_se;
  output pwm_o;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, net8871, n1, n2, n3, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [6:0] pwmcnt;

  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  glreg_a0_1 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm), .test_si(pwmcnt[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8871), .TE(test_se) );
  SDFFSQX1 pwmcnt_reg_6_ ( .D(N20), .SIN(pwmcnt[5]), .SMC(test_se), .C(net8871), .XS(n2), .Q(pwmcnt[6]) );
  SDFFSQX1 pwmcnt_reg_4_ ( .D(N18), .SIN(pwmcnt[3]), .SMC(test_se), .C(net8871), .XS(n2), .Q(pwmcnt[4]) );
  SDFFSQX1 pwmcnt_reg_5_ ( .D(N19), .SIN(pwmcnt[4]), .SMC(test_se), .C(net8871), .XS(n2), .Q(pwmcnt[5]) );
  SDFFSQX1 pwmcnt_reg_2_ ( .D(N16), .SIN(pwmcnt[1]), .SMC(test_se), .C(net8871), .XS(n2), .Q(pwmcnt[2]) );
  SDFFSQX1 pwmcnt_reg_3_ ( .D(N17), .SIN(pwmcnt[2]), .SMC(test_se), .C(net8871), .XS(n2), .Q(pwmcnt[3]) );
  SDFFSQX1 pwmcnt_reg_1_ ( .D(N15), .SIN(pwmcnt[0]), .SMC(test_se), .C(net8871), .XS(n1), .Q(pwmcnt[1]) );
  SDFFSQX1 pwmcnt_reg_0_ ( .D(N14), .SIN(test_si), .SMC(test_se), .C(net8871), 
        .XS(n1), .Q(pwmcnt[0]) );
  INVX1 U6 ( .A(n33), .Y(n4) );
  INVX1 U7 ( .A(n36), .Y(n13) );
  INVX1 U8 ( .A(n27), .Y(n7) );
  NOR21XL U9 ( .B(we), .A(wdat[7]), .Y(n33) );
  NAND2X1 U10 ( .A(n8), .B(n4), .Y(N13) );
  INVX1 U11 ( .A(n35), .Y(n12) );
  INVX1 U12 ( .A(n34), .Y(n11) );
  OAI221X1 U13 ( .A(n19), .B(n20), .C(pwmcnt[6]), .D(n6), .E(n21), .Y(pwm_o)
         );
  AOI32X1 U14 ( .A(n22), .B(n14), .C(r_pwm[4]), .D(r_pwm[5]), .E(n15), .Y(n20)
         );
  OAI211X1 U15 ( .C(r_pwm[4]), .D(n14), .A(n22), .B(n23), .Y(n21) );
  INVX1 U16 ( .A(pwmcnt[4]), .Y(n14) );
  NOR2X1 U17 ( .A(pwmcnt[1]), .B(pwmcnt[0]), .Y(n36) );
  AOI21X1 U18 ( .B(n24), .C(n25), .A(n19), .Y(n23) );
  AOI32X1 U19 ( .A(n7), .B(n17), .C(r_pwm[2]), .D(r_pwm[3]), .E(n18), .Y(n24)
         );
  OAI221X1 U20 ( .A(n9), .B(n16), .C(r_pwm[2]), .D(n17), .E(n26), .Y(n25) );
  INVX1 U21 ( .A(pwmcnt[2]), .Y(n17) );
  AOI211X1 U22 ( .C(n13), .D(n5), .A(n27), .B(n28), .Y(n26) );
  INVX1 U23 ( .A(r_pwm[1]), .Y(n5) );
  AOI21X1 U24 ( .B(r_pwm[1]), .C(n16), .A(r_pwm[0]), .Y(n28) );
  INVX1 U25 ( .A(pwmcnt[1]), .Y(n16) );
  NOR2X1 U26 ( .A(n18), .B(r_pwm[3]), .Y(n27) );
  INVX1 U27 ( .A(pwmcnt[3]), .Y(n18) );
  NAND21X1 U28 ( .B(r_pwm[5]), .A(pwmcnt[5]), .Y(n22) );
  AND2X1 U29 ( .A(pwmcnt[6]), .B(n6), .Y(n19) );
  INVX1 U30 ( .A(r_pwm[6]), .Y(n6) );
  INVX1 U31 ( .A(pwmcnt[5]), .Y(n15) );
  INVX1 U32 ( .A(pwmcnt[0]), .Y(n9) );
  GEN2XL U33 ( .D(pwmcnt[1]), .E(pwmcnt[0]), .C(n36), .B(r_pwm[7]), .A(n33), 
        .Y(N15) );
  GEN2XL U34 ( .D(pwmcnt[2]), .E(n13), .C(n35), .B(r_pwm[7]), .A(n33), .Y(N16)
         );
  GEN2XL U35 ( .D(pwmcnt[4]), .E(n11), .C(n31), .B(r_pwm[7]), .A(n33), .Y(N18)
         );
  GEN2XL U36 ( .D(pwmcnt[3]), .E(n12), .C(n34), .B(r_pwm[7]), .A(n33), .Y(N17)
         );
  OAI21X1 U37 ( .B(n32), .C(n8), .A(n4), .Y(N19) );
  XNOR2XL U38 ( .A(n31), .B(pwmcnt[5]), .Y(n32) );
  OAI21X1 U39 ( .B(n29), .C(n8), .A(n4), .Y(N20) );
  XNOR2XL U40 ( .A(pwmcnt[6]), .B(n30), .Y(n29) );
  NOR2X1 U41 ( .A(pwmcnt[5]), .B(n10), .Y(n30) );
  INVX1 U42 ( .A(n31), .Y(n10) );
  OAI21X1 U43 ( .B(pwmcnt[0]), .C(n8), .A(n4), .Y(N14) );
  NOR2X1 U44 ( .A(n11), .B(pwmcnt[4]), .Y(n31) );
  NOR2X1 U45 ( .A(n13), .B(pwmcnt[2]), .Y(n35) );
  NOR2X1 U46 ( .A(n12), .B(pwmcnt[3]), .Y(n34) );
  INVX1 U47 ( .A(r_pwm[7]), .Y(n8) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8889;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8889), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8889), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8889), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8889), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8889), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8889), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8889), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8889), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8889), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_0 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o, test_si, 
        test_se );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we, test_si, test_se;
  output pwm_o;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, net8907, n1, n2, n3, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [6:0] pwmcnt;

  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  glreg_a0_0 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm), .test_si(pwmcnt[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8907), .TE(test_se) );
  SDFFSQX1 pwmcnt_reg_6_ ( .D(N20), .SIN(pwmcnt[5]), .SMC(test_se), .C(net8907), .XS(n2), .Q(pwmcnt[6]) );
  SDFFSQX1 pwmcnt_reg_4_ ( .D(N18), .SIN(pwmcnt[3]), .SMC(test_se), .C(net8907), .XS(n2), .Q(pwmcnt[4]) );
  SDFFSQX1 pwmcnt_reg_2_ ( .D(N16), .SIN(pwmcnt[1]), .SMC(test_se), .C(net8907), .XS(n2), .Q(pwmcnt[2]) );
  SDFFSQX1 pwmcnt_reg_5_ ( .D(N19), .SIN(pwmcnt[4]), .SMC(test_se), .C(net8907), .XS(n2), .Q(pwmcnt[5]) );
  SDFFSQX1 pwmcnt_reg_1_ ( .D(N15), .SIN(pwmcnt[0]), .SMC(test_se), .C(net8907), .XS(n1), .Q(pwmcnt[1]) );
  SDFFSQX1 pwmcnt_reg_3_ ( .D(N17), .SIN(pwmcnt[2]), .SMC(test_se), .C(net8907), .XS(n2), .Q(pwmcnt[3]) );
  SDFFSQX1 pwmcnt_reg_0_ ( .D(N14), .SIN(test_si), .SMC(test_se), .C(net8907), 
        .XS(n1), .Q(pwmcnt[0]) );
  INVX1 U6 ( .A(n33), .Y(n4) );
  INVX1 U7 ( .A(n36), .Y(n14) );
  INVX1 U8 ( .A(n27), .Y(n7) );
  NOR21XL U9 ( .B(we), .A(wdat[7]), .Y(n33) );
  NAND2X1 U10 ( .A(n8), .B(n4), .Y(N13) );
  INVX1 U11 ( .A(n35), .Y(n12) );
  INVX1 U12 ( .A(n34), .Y(n11) );
  OAI221X1 U13 ( .A(n19), .B(n20), .C(pwmcnt[6]), .D(n6), .E(n21), .Y(pwm_o)
         );
  AOI32X1 U14 ( .A(n22), .B(n15), .C(r_pwm[4]), .D(r_pwm[5]), .E(n16), .Y(n20)
         );
  OAI211X1 U15 ( .C(r_pwm[4]), .D(n15), .A(n22), .B(n23), .Y(n21) );
  INVX1 U16 ( .A(pwmcnt[4]), .Y(n15) );
  NOR2X1 U17 ( .A(n18), .B(r_pwm[3]), .Y(n27) );
  NOR2X1 U18 ( .A(pwmcnt[1]), .B(pwmcnt[0]), .Y(n36) );
  AOI211X1 U19 ( .C(n14), .D(n5), .A(n27), .B(n28), .Y(n26) );
  INVX1 U20 ( .A(r_pwm[1]), .Y(n5) );
  AOI21X1 U21 ( .B(r_pwm[1]), .C(n17), .A(r_pwm[0]), .Y(n28) );
  AOI21X1 U22 ( .B(n24), .C(n25), .A(n19), .Y(n23) );
  AOI32X1 U23 ( .A(n7), .B(n9), .C(r_pwm[2]), .D(r_pwm[3]), .E(n18), .Y(n24)
         );
  OAI221X1 U24 ( .A(n13), .B(n17), .C(r_pwm[2]), .D(n9), .E(n26), .Y(n25) );
  INVX1 U25 ( .A(pwmcnt[2]), .Y(n9) );
  INVX1 U26 ( .A(pwmcnt[3]), .Y(n18) );
  INVX1 U27 ( .A(pwmcnt[1]), .Y(n17) );
  AND2X1 U28 ( .A(pwmcnt[6]), .B(n6), .Y(n19) );
  INVX1 U29 ( .A(r_pwm[6]), .Y(n6) );
  INVX1 U30 ( .A(pwmcnt[5]), .Y(n16) );
  INVX1 U31 ( .A(pwmcnt[0]), .Y(n13) );
  NAND21X1 U32 ( .B(r_pwm[5]), .A(pwmcnt[5]), .Y(n22) );
  GEN2XL U33 ( .D(pwmcnt[1]), .E(pwmcnt[0]), .C(n36), .B(r_pwm[7]), .A(n33), 
        .Y(N15) );
  GEN2XL U34 ( .D(pwmcnt[2]), .E(n14), .C(n35), .B(r_pwm[7]), .A(n33), .Y(N16)
         );
  GEN2XL U35 ( .D(pwmcnt[4]), .E(n11), .C(n31), .B(r_pwm[7]), .A(n33), .Y(N18)
         );
  GEN2XL U36 ( .D(pwmcnt[3]), .E(n12), .C(n34), .B(r_pwm[7]), .A(n33), .Y(N17)
         );
  OAI21X1 U37 ( .B(n32), .C(n8), .A(n4), .Y(N19) );
  XNOR2XL U38 ( .A(n31), .B(pwmcnt[5]), .Y(n32) );
  OAI21X1 U39 ( .B(pwmcnt[0]), .C(n8), .A(n4), .Y(N14) );
  OAI21X1 U40 ( .B(n29), .C(n8), .A(n4), .Y(N20) );
  XNOR2XL U41 ( .A(pwmcnt[6]), .B(n30), .Y(n29) );
  NOR2X1 U42 ( .A(pwmcnt[5]), .B(n10), .Y(n30) );
  INVX1 U43 ( .A(n31), .Y(n10) );
  NOR2X1 U44 ( .A(n11), .B(pwmcnt[4]), .Y(n31) );
  NOR2X1 U45 ( .A(n14), .B(pwmcnt[2]), .Y(n35) );
  NOR2X1 U46 ( .A(n12), .B(pwmcnt[3]), .Y(n34) );
  INVX1 U47 ( .A(r_pwm[7]), .Y(n8) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8925;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8925), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8925), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8925), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8925), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8925), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8925), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8925), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8925), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8925), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module divclk_a0 ( mclk, srstz, atpg_en, clk_1p0m, clk_500k, clk_100k, clk_50k, 
        clk_500, divff_o1, divff_o2, test_si, test_so, test_se );
  input mclk, srstz, atpg_en, test_si, test_se;
  output clk_1p0m, clk_500k, clk_100k, clk_50k, clk_500, divff_o1, divff_o2,
         test_so;
  wire   div500k_5_0, div1p0m_2, div100k_2, N23, N24, N25, N26, N37, N38, N39,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         n22, n23, n24, n1, n2, n3, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n25, n26, n27, n4, n5, n6, n7, n8, n9, n10;
  wire   [2:0] div12;
  wire   [6:0] div50k_100;

  CLKDLX1 U0_D1P0M_ICG ( .CK(mclk), .E(n22), .SE(atpg_en), .ECK(clk_1p0m) );
  CLKDLX1 U0_D500K_ICG ( .CK(clk_1p0m), .E(div1p0m_2), .SE(atpg_en), .ECK(
        clk_500k) );
  CLKDLX1 U0_D100K_ICG ( .CK(clk_500k), .E(n23), .SE(atpg_en), .ECK(clk_100k)
         );
  CLKDLX1 U0_D50K_ICG ( .CK(clk_100k), .E(div100k_2), .SE(atpg_en), .ECK(
        clk_50k) );
  CLKDLX1 U0_D0P5K_ICG ( .CK(clk_50k), .E(n24), .SE(atpg_en), .ECK(clk_500) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(srstz), .Y(n3) );
  divclk_a0_DW01_inc_0 add_60 ( .A(div50k_100), .SUM({N52, N51, N50, N49, N48, 
        N47, N46}) );
  SDFFRQX1 div1p0m_2_reg ( .D(n4), .SIN(test_si), .SMC(test_se), .C(clk_1p0m), 
        .XR(n1), .Q(div1p0m_2) );
  SDFFRQX1 div100k_2_reg ( .D(n5), .SIN(div50k_100[6]), .SMC(test_se), .C(
        clk_100k), .XR(n1), .Q(div100k_2) );
  SDFFRQX1 div50k_100_reg_6_ ( .D(N59), .SIN(div50k_100[5]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[6]) );
  SDFFRQX1 div50k_100_reg_5_ ( .D(N58), .SIN(div50k_100[4]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[5]) );
  SDFFRQX1 div50k_100_reg_4_ ( .D(N57), .SIN(div50k_100[3]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[4]) );
  SDFFRQX1 div50k_100_reg_3_ ( .D(N56), .SIN(div50k_100[2]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[3]) );
  SDFFRQX1 div500k_5_reg_1_ ( .D(N38), .SIN(div500k_5_0), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(divff_o2) );
  SDFFRQX1 div500k_5_reg_0_ ( .D(N37), .SIN(div100k_2), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(div500k_5_0) );
  SDFFRQX1 div12_reg_0_ ( .D(N23), .SIN(div1p0m_2), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(div12[0]) );
  SDFFRQX1 div50k_100_reg_1_ ( .D(N54), .SIN(div50k_100[0]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[1]) );
  SDFFRQX1 div50k_100_reg_2_ ( .D(N55), .SIN(div50k_100[1]), .SMC(test_se), 
        .C(clk_50k), .XR(n2), .Q(div50k_100[2]) );
  SDFFRQX1 div500k_5_reg_2_ ( .D(N39), .SIN(divff_o2), .SMC(test_se), .C(
        clk_500k), .XR(n1), .Q(test_so) );
  SDFFRQX1 div50k_100_reg_0_ ( .D(N53), .SIN(divff_o1), .SMC(test_se), .C(
        clk_50k), .XR(n1), .Q(div50k_100[0]) );
  SDFFRQX1 div12_reg_1_ ( .D(N24), .SIN(div12[0]), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(div12[1]) );
  SDFFRQX1 div12_reg_2_ ( .D(N25), .SIN(div12[1]), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(div12[2]) );
  SDFFRQX1 div12_reg_3_ ( .D(N26), .SIN(div12[2]), .SMC(test_se), .C(mclk), 
        .XR(n1), .Q(divff_o1) );
  XNOR2XL U6 ( .A(n19), .B(n18), .Y(n16) );
  XNOR2XL U7 ( .A(n14), .B(n16), .Y(N25) );
  INVX1 U8 ( .A(n26), .Y(n9) );
  NOR2X1 U9 ( .A(n25), .B(n26), .Y(n18) );
  NOR2X1 U10 ( .A(n15), .B(n20), .Y(N24) );
  XOR2X1 U11 ( .A(n16), .B(n21), .Y(n20) );
  XNOR2XL U12 ( .A(n9), .B(n25), .Y(n21) );
  NOR21XL U13 ( .B(n14), .A(n15), .Y(N26) );
  NOR21XL U14 ( .B(N48), .A(n24), .Y(N55) );
  NOR21XL U15 ( .B(N49), .A(n24), .Y(N56) );
  NOR21XL U16 ( .B(N47), .A(n24), .Y(N54) );
  NOR21XL U17 ( .B(N50), .A(n24), .Y(N57) );
  NOR21XL U18 ( .B(N51), .A(n24), .Y(N58) );
  NOR2X1 U19 ( .A(n11), .B(n10), .Y(n15) );
  NOR2X1 U20 ( .A(N23), .B(n11), .Y(n22) );
  XNOR2XL U21 ( .A(n19), .B(div12[1]), .Y(n26) );
  XNOR2XL U22 ( .A(n10), .B(div12[2]), .Y(n19) );
  XNOR2XL U23 ( .A(n9), .B(div12[0]), .Y(n25) );
  XNOR2XL U24 ( .A(n17), .B(divff_o1), .Y(n14) );
  NAND2X1 U25 ( .A(n18), .B(n19), .Y(n17) );
  INVX1 U26 ( .A(divff_o1), .Y(n10) );
  AND4X1 U27 ( .A(div50k_100[5]), .B(div50k_100[1]), .C(div50k_100[6]), .D(n12), .Y(n24) );
  NOR41XL U28 ( .D(div50k_100[0]), .A(div50k_100[4]), .B(div50k_100[3]), .C(
        div50k_100[2]), .Y(n12) );
  NOR21XL U29 ( .B(N46), .A(n24), .Y(N53) );
  NOR21XL U30 ( .B(N52), .A(n24), .Y(N59) );
  OAI32X1 U31 ( .A(n7), .B(test_so), .C(n8), .D(n13), .E(n6), .Y(N39) );
  INVX1 U32 ( .A(div500k_5_0), .Y(n8) );
  AOI21BBXL U33 ( .B(n23), .C(divff_o2), .A(N37), .Y(n13) );
  NOR3XL U34 ( .A(div500k_5_0), .B(divff_o2), .C(n6), .Y(n23) );
  NOR2X1 U35 ( .A(n23), .B(div500k_5_0), .Y(N37) );
  INVX1 U36 ( .A(test_so), .Y(n6) );
  NAND31X1 U37 ( .C(div12[0]), .A(div12[1]), .B(div12[2]), .Y(n11) );
  XOR2X1 U38 ( .A(n27), .B(div12[1]), .Y(N23) );
  XNOR2XL U39 ( .A(divff_o1), .B(div12[2]), .Y(n27) );
  XNOR2XL U40 ( .A(n7), .B(div500k_5_0), .Y(N38) );
  INVX1 U41 ( .A(divff_o2), .Y(n7) );
  INVX1 U42 ( .A(div100k_2), .Y(n5) );
  INVX1 U43 ( .A(div1p0m_2), .Y(n4) );
endmodule


module divclk_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module srambist_a0 ( clk, srstz, reg_hit, reg_w, reg_r, reg_wdat, iram_rdat, 
        xram_rdat, bist_en, bist_xram, bist_wr, bist_adr, bist_wdat, o_bistctl, 
        o_bistdat, test_si, test_se );
  input [1:0] reg_hit;
  input [7:0] reg_wdat;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  output [10:0] bist_adr;
  output [7:0] bist_wdat;
  output [6:0] o_bistctl;
  output [7:0] o_bistdat;
  input clk, srstz, reg_w, reg_r, test_si, test_se;
  output bist_en, bist_xram, bist_wr;
  wire   we_1_, bistctl_re, N21, busy_dly, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, r_bistfault, upd_fault, wd_fault, net8943, n110, n111, n10,
         n11, n12, n24, n25, n29, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n84, n85, n89, n120, n121, n122,
         n3, n4, n5, n6, n7, n8, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n26, n27, n28, n30, n31, n32, n64, n65, n66, n80, n81, n82, n83,
         n86, n87, n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n112, n113,
         n114, n115, n116, n117, n118, n119, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133;
  wire   [1:0] rw_sta;

  INVX1 U17 ( .A(n12), .Y(n11) );
  INVX1 U18 ( .A(n12), .Y(n10) );
  INVX1 U19 ( .A(srstz), .Y(n12) );
  INVX8 U146 ( .A(n11), .Y(n24) );
  glreg_WIDTH1_0 u0_bistfault ( .clk(clk), .arstz(n11), .we(upd_fault), .wdat(
        wd_fault), .rdat(o_bistctl[3]), .test_si(o_bistdat[7]), .test_se(
        test_se) );
  glreg_WIDTH5_1 u0_bistctl ( .clk(clk), .arstz(n11), .we(n25), .wdat({
        reg_wdat[6:4], reg_wdat[2:1]}), .rdat({o_bistctl[6:4], o_bistctl[2:1]}), .test_si(rw_sta[1]), .test_se(test_se) );
  glreg_a0_6 u0_bistdat ( .clk(clk), .arstz(n10), .we(we_1_), .wdat(reg_wdat), 
        .rdat(o_bistdat), .test_si(o_bistctl[6]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_srambist_a0 clk_gate_adr_reg ( .CLK(clk), .EN(N86), 
        .ENCLK(net8943), .TE(test_se) );
  srambist_a0_DW01_inc_0 add_65 ( .A(bist_adr), .SUM({N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64}) );
  SDFFQX1 busy_dly_reg ( .D(o_bistctl[0]), .SIN(bistctl_re), .SMC(test_se), 
        .C(clk), .Q(busy_dly) );
  SDFFQX1 r_bistfault_reg ( .D(n110), .SIN(busy_dly), .SMC(test_se), .C(clk), 
        .Q(r_bistfault) );
  SDFFRQX1 bistctl_re_reg ( .D(N21), .SIN(bist_adr[10]), .SMC(test_se), .C(clk), .XR(n11), .Q(bistctl_re) );
  SDFFQX1 rw_sta_reg_1_ ( .D(n130), .SIN(rw_sta[0]), .SMC(test_se), .C(clk), 
        .Q(rw_sta[1]) );
  SDFFQX1 rw_sta_reg_0_ ( .D(n111), .SIN(r_bistfault), .SMC(test_se), .C(clk), 
        .Q(rw_sta[0]) );
  SDFFQX1 adr_reg_9_ ( .D(N96), .SIN(bist_adr[8]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[9]) );
  SDFFQX1 adr_reg_10_ ( .D(N97), .SIN(bist_adr[9]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[10]) );
  SDFFQX1 adr_reg_5_ ( .D(N92), .SIN(bist_adr[4]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[5]) );
  SDFFQX1 adr_reg_6_ ( .D(N93), .SIN(bist_adr[5]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[6]) );
  SDFFQX1 adr_reg_8_ ( .D(N95), .SIN(bist_adr[7]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[8]) );
  SDFFQX1 adr_reg_7_ ( .D(N94), .SIN(bist_adr[6]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[7]) );
  SDFFQX1 adr_reg_3_ ( .D(N90), .SIN(bist_adr[2]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[3]) );
  SDFFQX1 adr_reg_4_ ( .D(N91), .SIN(bist_adr[3]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[4]) );
  SDFFQX1 adr_reg_1_ ( .D(N88), .SIN(bist_adr[0]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[1]) );
  SDFFQX1 adr_reg_2_ ( .D(N89), .SIN(bist_adr[1]), .SMC(test_se), .C(net8943), 
        .Q(bist_adr[2]) );
  SDFFQX1 adr_reg_0_ ( .D(N87), .SIN(test_si), .SMC(test_se), .C(net8943), .Q(
        bist_adr[0]) );
  INVX1 U3 ( .A(1'b1), .Y(bist_xram) );
  NAND21X1 U5 ( .B(n105), .A(n104), .Y(n106) );
  AND2X1 U6 ( .A(bist_adr[6]), .B(bist_adr[3]), .Y(n103) );
  INVX1 U7 ( .A(n95), .Y(n3) );
  BUFXL U8 ( .A(o_bistctl[0]), .Y(bist_en) );
  AO21XL U9 ( .B(n101), .C(n92), .A(n91), .Y(n93) );
  INVXL U10 ( .A(iram_rdat[4]), .Y(n133) );
  XOR2XL U11 ( .A(bist_wdat[1]), .B(iram_rdat[1]), .Y(n70) );
  XOR2XL U12 ( .A(iram_rdat[1]), .B(n48), .Y(n42) );
  NAND21XL U13 ( .B(n90), .A(bist_adr[1]), .Y(n101) );
  OAI21BBX1 U14 ( .A(N64), .B(n89), .C(n4), .Y(N87) );
  AOI21XL U15 ( .B(n97), .C(n90), .A(n88), .Y(n4) );
  NAND32XL U16 ( .B(rw_sta[1]), .C(n131), .A(o_bistctl[0]), .Y(n115) );
  OAI21BBXL U20 ( .A(n8), .B(o_bistctl[0]), .C(n10), .Y(n113) );
  NAND21XL U21 ( .B(bist_adr[9]), .A(n105), .Y(n96) );
  INVX1 U22 ( .A(n121), .Y(n25) );
  NAND2X1 U23 ( .A(reg_hit[0]), .B(reg_w), .Y(n121) );
  INVX1 U24 ( .A(n91), .Y(n97) );
  AND2X1 U25 ( .A(reg_w), .B(reg_hit[1]), .Y(we_1_) );
  INVX1 U26 ( .A(n49), .Y(n123) );
  INVX1 U27 ( .A(n99), .Y(n105) );
  INVX1 U28 ( .A(n82), .Y(n86) );
  INVX1 U29 ( .A(n20), .Y(n22) );
  INVX1 U30 ( .A(n66), .Y(n81) );
  INVX1 U31 ( .A(n32), .Y(n65) );
  INVX1 U32 ( .A(n28), .Y(n31) );
  INVX1 U33 ( .A(n23), .Y(n27) );
  OAI22AX1 U34 ( .D(n75), .C(n72), .A(n127), .B(n75), .Y(bist_wdat[4]) );
  OAI21X1 U35 ( .B(n127), .C(n119), .A(n72), .Y(bist_wdat[0]) );
  NAND2X1 U36 ( .A(n74), .B(n117), .Y(n75) );
  NAND2X1 U37 ( .A(n127), .B(n119), .Y(n72) );
  INVX1 U38 ( .A(n73), .Y(n117) );
  INVX1 U39 ( .A(n77), .Y(n119) );
  OR2X1 U40 ( .A(n85), .B(n84), .Y(n19) );
  OR2X1 U41 ( .A(n84), .B(n120), .Y(n91) );
  NOR21XL U42 ( .B(n84), .A(n120), .Y(n89) );
  OAI2B11X1 U43 ( .D(N65), .C(n95), .A(n94), .B(n93), .Y(N88) );
  INVX1 U44 ( .A(n88), .Y(n94) );
  INVX1 U45 ( .A(n89), .Y(n95) );
  AND2X1 U46 ( .A(reg_r), .B(reg_hit[0]), .Y(N21) );
  XNOR2XL U47 ( .A(n127), .B(n79), .Y(bist_wdat[1]) );
  AOI21X1 U48 ( .B(n75), .C(n74), .A(n77), .Y(n79) );
  XNOR2XL U49 ( .A(n127), .B(n78), .Y(bist_wdat[2]) );
  AOI21X1 U50 ( .B(n75), .C(n117), .A(n77), .Y(n78) );
  OAI22X1 U51 ( .A(n72), .B(n75), .C(n76), .D(n127), .Y(bist_wdat[3]) );
  NOR2X1 U52 ( .A(n77), .B(n75), .Y(n76) );
  OAI22X1 U53 ( .A(n72), .B(n117), .C(n73), .D(n127), .Y(bist_wdat[6]) );
  XNOR2XL U54 ( .A(iram_rdat[2]), .B(n51), .Y(n44) );
  AOI21X1 U55 ( .B(n49), .C(n124), .A(n50), .Y(n51) );
  AOI31XL U56 ( .A(iram_rdat[7]), .B(n42), .C(n43), .D(n128), .Y(n38) );
  AOI21X1 U57 ( .B(n123), .C(n133), .A(n44), .Y(n43) );
  AOI21X1 U58 ( .B(n49), .C(n41), .A(n50), .Y(n48) );
  XOR2XL U59 ( .A(bist_wdat[3]), .B(iram_rdat[3]), .Y(n67) );
  XNOR2XL U60 ( .A(n127), .B(iram_rdat[7]), .Y(n69) );
  XNOR2XL U61 ( .A(iram_rdat[6]), .B(n60), .Y(n52) );
  OAI22X1 U62 ( .A(n126), .B(n124), .C(n61), .D(n128), .Y(n60) );
  XNOR2XL U63 ( .A(iram_rdat[0]), .B(n59), .Y(n53) );
  NAND2X1 U64 ( .A(n126), .B(n57), .Y(n59) );
  INVXL U65 ( .A(iram_rdat[5]), .Y(n132) );
  NOR43XL U66 ( .B(n5), .C(n6), .D(n7), .A(n67), .Y(n63) );
  XOR2X1 U67 ( .A(bist_wdat[5]), .B(n132), .Y(n5) );
  XNOR2XL U68 ( .A(bist_wdat[0]), .B(iram_rdat[0]), .Y(n6) );
  XNOR2XL U69 ( .A(bist_wdat[6]), .B(iram_rdat[6]), .Y(n7) );
  NOR4XL U70 ( .A(n68), .B(n69), .C(n70), .D(n71), .Y(n62) );
  XNOR2XL U71 ( .A(n133), .B(bist_wdat[4]), .Y(n68) );
  XOR2X1 U72 ( .A(bist_wdat[2]), .B(iram_rdat[2]), .Y(n71) );
  INVX1 U73 ( .A(n115), .Y(bist_wr) );
  NAND2X1 U74 ( .A(n41), .B(n124), .Y(n49) );
  INVX1 U75 ( .A(n61), .Y(n124) );
  INVX1 U76 ( .A(n58), .Y(n126) );
  NAND2X1 U77 ( .A(n131), .B(n116), .Y(n29) );
  NAND3X1 U78 ( .A(bist_adr[9]), .B(bist_adr[10]), .C(n106), .Y(o_bistctl[0])
         );
  NAND21X1 U79 ( .B(bist_adr[1]), .A(n90), .Y(n92) );
  NAND21X1 U80 ( .B(bist_adr[7]), .A(n27), .Y(n20) );
  NAND21X1 U81 ( .B(bist_adr[8]), .A(n22), .Y(n99) );
  NAND21X1 U82 ( .B(bist_adr[3]), .A(n86), .Y(n66) );
  NAND21X1 U83 ( .B(bist_adr[4]), .A(n81), .Y(n32) );
  NAND21X1 U84 ( .B(bist_adr[5]), .A(n65), .Y(n28) );
  NAND21X1 U85 ( .B(bist_adr[6]), .A(n31), .Y(n23) );
  INVX1 U86 ( .A(bist_adr[0]), .Y(n90) );
  OR2X1 U87 ( .A(bist_adr[2]), .B(n92), .Y(n82) );
  NOR43XL U88 ( .B(bist_adr[4]), .C(bist_adr[8]), .D(bist_adr[5]), .A(n101), 
        .Y(n102) );
  NAND4X1 U89 ( .A(bist_adr[2]), .B(bist_adr[7]), .C(n103), .D(n102), .Y(n104)
         );
  NOR2X1 U90 ( .A(o_bistdat[2]), .B(o_bistdat[3]), .Y(n77) );
  NOR2X1 U91 ( .A(n118), .B(o_bistdat[3]), .Y(n73) );
  INVX1 U92 ( .A(o_bistdat[5]), .Y(n127) );
  INVX1 U93 ( .A(o_bistdat[2]), .Y(n118) );
  NAND2X1 U94 ( .A(o_bistdat[3]), .B(n118), .Y(n74) );
  NAND21X1 U95 ( .B(n24), .A(n19), .Y(n88) );
  NAND42XL U96 ( .C(o_bistdat[6]), .D(n121), .A(reg_wdat[0]), .B(o_bistdat[7]), 
        .Y(n85) );
  OAI22AX1 U97 ( .D(n121), .C(o_bistctl[1]), .A(reg_wdat[1]), .B(n121), .Y(n84) );
  AO21X1 U98 ( .B(N66), .C(n89), .A(n87), .Y(N89) );
  GEN2XL U99 ( .D(bist_adr[2]), .E(n92), .C(n86), .B(n97), .A(n88), .Y(n87) );
  AO21X1 U100 ( .B(N71), .C(n89), .A(n26), .Y(N94) );
  GEN2XL U101 ( .D(bist_adr[7]), .E(n23), .C(n22), .B(n97), .A(n88), .Y(n26)
         );
  AO21X1 U102 ( .B(N70), .C(n89), .A(n30), .Y(N93) );
  GEN2XL U103 ( .D(bist_adr[6]), .E(n28), .C(n27), .B(n97), .A(n88), .Y(n30)
         );
  AO21X1 U104 ( .B(N67), .C(n89), .A(n83), .Y(N90) );
  GEN2XL U105 ( .D(bist_adr[3]), .E(n82), .C(n81), .B(n97), .A(n88), .Y(n83)
         );
  AO21X1 U106 ( .B(N68), .C(n89), .A(n80), .Y(N91) );
  GEN2XL U107 ( .D(bist_adr[4]), .E(n66), .C(n65), .B(n97), .A(n88), .Y(n80)
         );
  AO21X1 U108 ( .B(N69), .C(n89), .A(n64), .Y(N92) );
  GEN2XL U109 ( .D(bist_adr[5]), .E(n32), .C(n31), .B(n97), .A(n88), .Y(n64)
         );
  AO21X1 U110 ( .B(N72), .C(n89), .A(n21), .Y(N95) );
  GEN2XL U111 ( .D(bist_adr[8]), .E(n20), .C(n105), .B(n97), .A(n88), .Y(n21)
         );
  AO21X1 U112 ( .B(N73), .C(n89), .A(n100), .Y(N96) );
  GEN2XL U113 ( .D(bist_adr[9]), .E(n99), .C(n98), .B(n97), .A(n114), .Y(n100)
         );
  INVX1 U114 ( .A(n96), .Y(n98) );
  NAND3X1 U115 ( .A(n85), .B(n29), .C(n122), .Y(n120) );
  AOI22X1 U116 ( .A(rw_sta[1]), .B(n129), .C(o_bistctl[2]), .D(rw_sta[0]), .Y(
        n122) );
  NAND43X1 U117 ( .B(n18), .C(n17), .D(n16), .A(n15), .Y(N97) );
  INVX1 U118 ( .A(n19), .Y(n17) );
  NAND21X1 U119 ( .B(n91), .A(n14), .Y(n15) );
  AND2X1 U120 ( .A(N74), .B(n3), .Y(n18) );
  NAND3X1 U121 ( .A(n120), .B(n85), .C(n11), .Y(N86) );
  ENOX1 U122 ( .A(n72), .B(n74), .C(n74), .D(o_bistdat[5]), .Y(bist_wdat[5])
         );
  NOR42XL U123 ( .C(n116), .D(n10), .A(n131), .B(n35), .Y(n34) );
  NOR4XL U124 ( .A(n36), .B(n37), .C(n38), .D(n39), .Y(n35) );
  NAND3X1 U125 ( .A(n52), .B(n53), .C(n54), .Y(n36) );
  XNOR2XL U126 ( .A(n40), .B(n132), .Y(n39) );
  OAI22X1 U127 ( .A(bistctl_re), .B(n112), .C(n114), .D(n109), .Y(n110) );
  INVX1 U128 ( .A(wd_fault), .Y(n109) );
  AOI31X1 U129 ( .A(busy_dly), .B(n11), .C(n33), .D(n34), .Y(n112) );
  AOI211X1 U130 ( .C(n62), .D(n63), .A(n29), .B(n129), .Y(n33) );
  OAI22X1 U131 ( .A(o_bistdat[4]), .B(n45), .C(n123), .D(n46), .Y(n37) );
  XNOR2XL U132 ( .A(n126), .B(n133), .Y(n46) );
  NOR32XL U133 ( .B(n47), .C(n44), .A(n42), .Y(n45) );
  AOI21XL U134 ( .B(iram_rdat[4]), .C(n123), .A(iram_rdat[7]), .Y(n47) );
  XNOR2XL U135 ( .A(iram_rdat[3]), .B(n55), .Y(n54) );
  NAND2X1 U136 ( .A(n56), .B(n57), .Y(n55) );
  OAI22X1 U137 ( .A(o_bistdat[4]), .B(n123), .C(n58), .D(n49), .Y(n56) );
  NOR2X1 U138 ( .A(n125), .B(o_bistdat[1]), .Y(n61) );
  INVX1 U139 ( .A(o_bistdat[0]), .Y(n125) );
  NAND2X1 U140 ( .A(o_bistdat[1]), .B(n125), .Y(n41) );
  OR2X1 U141 ( .A(n131), .B(n116), .Y(n8) );
  NOR2X1 U142 ( .A(n50), .B(o_bistdat[4]), .Y(n58) );
  NOR2X1 U143 ( .A(o_bistdat[0]), .B(o_bistdat[1]), .Y(n50) );
  OAI32X1 U144 ( .A(n115), .B(n114), .C(n129), .D(n116), .E(n113), .Y(n130) );
  ENOX1 U145 ( .A(n126), .B(n41), .C(n41), .D(o_bistdat[4]), .Y(n40) );
  INVX1 U147 ( .A(rw_sta[0]), .Y(n131) );
  NAND2X1 U148 ( .A(n50), .B(o_bistdat[4]), .Y(n57) );
  MUX2IX1 U149 ( .D0(n131), .D1(n108), .S(n113), .Y(n111) );
  NAND21X1 U151 ( .B(n24), .A(n107), .Y(n108) );
  INVX1 U152 ( .A(n29), .Y(n107) );
  XNOR2XL U153 ( .A(n96), .B(bist_adr[10]), .Y(n14) );
  INVX1 U154 ( .A(o_bistdat[4]), .Y(n128) );
  INVX1 U155 ( .A(o_bistctl[2]), .Y(n129) );
  INVX1 U156 ( .A(rw_sta[1]), .Y(n116) );
  OR2X1 U157 ( .A(bistctl_re), .B(r_bistfault), .Y(upd_fault) );
  NOR21XL U158 ( .B(r_bistfault), .A(bistctl_re), .Y(wd_fault) );
  BUFX3 U159 ( .A(o_bistdat[5]), .Y(bist_wdat[7]) );
  INVX8 U160 ( .A(srstz), .Y(n16) );
  INVX8 U161 ( .A(srstz), .Y(n114) );
endmodule


module srambist_a0_DW01_inc_0 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1XL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_srambist_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_6 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8961;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8961), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8961), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8961), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net8961), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net8961), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8961), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net8961), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8961), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8961), 
        .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net8979;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8979), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net8979), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net8979), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net8979), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net8979), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net8979), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module regx_a0 ( regx_r, regx_w, di_drposc, di_imposc, di_rd_det, clk_500k, 
        r_imp_osc, regx_addr, regx_wdat, regx_rdat, regx_hitbst, regx_wrpwm, 
        regx_wrcvc, r_sdischg, r_bistctl, r_bistdat, r_vcomp, r_idacsh, 
        r_cvofsx, r_pwm, regx_wrdac, dac_r_vs, dac_comp, r_dac_en, r_sar_en, 
        r_aopt, r_xtm, r_adummyi, r_bck0, r_bck1, r_bck2, r_i2crout, r_xana, 
        di_xanav, lt_gpi, di_tst, bkpt_pc, bkpt_ena, we_twlb, r_vpp_en, 
        r_vpp0v_en, r_otp_pwdn_en, r_otp_wpls, wd_twlb, r_sap, r_twlb, 
        upd_pwrv, ramacc, sse_idle, bus_idle, r_do_ts, r_dpdo_sel, r_dndo_sel, 
        di_ts, detclk, aswclk, atpg_en, di_aswk, clk, rrstz, test_si2, 
        test_si1, test_so1, test_se );
  input [6:0] regx_addr;
  input [7:0] regx_wdat;
  output [7:0] regx_rdat;
  output [1:0] regx_hitbst;
  output [1:0] regx_wrpwm;
  output [3:0] regx_wrcvc;
  input [7:0] r_sdischg;
  input [6:0] r_bistctl;
  input [7:0] r_bistdat;
  input [7:0] r_vcomp;
  input [7:0] r_idacsh;
  input [7:0] r_cvofsx;
  input [15:0] r_pwm;
  output [13:0] regx_wrdac;
  input [79:0] dac_r_vs;
  input [9:0] dac_comp;
  input [9:0] r_dac_en;
  input [9:0] r_sar_en;
  output [7:0] r_aopt;
  output [7:0] r_xtm;
  output [7:0] r_adummyi;
  output [7:0] r_bck0;
  output [7:0] r_bck1;
  output [7:0] r_bck2;
  output [5:0] r_i2crout;
  output [23:0] r_xana;
  input [5:0] di_xanav;
  input [3:0] lt_gpi;
  output [14:0] bkpt_pc;
  output [1:0] wd_twlb;
  output [1:0] r_sap;
  input [1:0] r_twlb;
  output [6:0] r_do_ts;
  output [3:0] r_dpdo_sel;
  output [3:0] r_dndo_sel;
  input [4:0] di_aswk;
  input regx_r, regx_w, di_drposc, di_imposc, di_rd_det, clk_500k, di_tst,
         upd_pwrv, ramacc, sse_idle, bus_idle, di_ts, detclk, aswclk, atpg_en,
         clk, rrstz, test_si2, test_si1, test_se;
  output r_imp_osc, bkpt_ena, we_twlb, r_vpp_en, r_vpp0v_en, r_otp_pwdn_en,
         r_otp_wpls, test_so1;
  wire   we_19, we_7, we_6, we_5, we_4, reg1B_3_, reg10_7_, lt_drp,
         i2c_mode_upd, N8, d_we16, lt_reg1C_0, net8997, n148, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n24, n33, n35, n38, n39, n40, n41, n42,
         n43, n44, n46, n47, n49, n50, n1, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27,
         n28, n29, n30, n31, n32, n34, n36, n37, n45, n48, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n61, n62, n63, n64, n65, n66, n67, n68, n95,
         n96, n98, n99, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n141,
         n142, n143, n144, n145, n146, n147, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151,
         SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153,
         SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155,
         SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157,
         SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159,
         SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161,
         SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163,
         SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165,
         SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167,
         SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169,
         SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171,
         SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173,
         SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175,
         SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177,
         SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179,
         SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181,
         SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183,
         SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185,
         SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187,
         SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189,
         SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191,
         SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193,
         SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195,
         SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197,
         SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199,
         SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201,
         SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203,
         SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205,
         SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207,
         SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209,
         SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211,
         SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213,
         SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215,
         SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217,
         SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219,
         SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221,
         SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223,
         SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225,
         SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227,
         SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229,
         SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231,
         SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233,
         SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235,
         SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237,
         SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239,
         SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241,
         SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243,
         SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245,
         SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247,
         SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249,
         SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251,
         SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253,
         SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255,
         SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257,
         SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259,
         SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261,
         SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263,
         SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265,
         SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267,
         SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269,
         SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271,
         SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273,
         SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275,
         SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277,
         SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279,
         SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281,
         SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283,
         SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285,
         SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287,
         SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289,
         SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291,
         SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293,
         SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295,
         SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297,
         SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299,
         SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301,
         SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303,
         SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305,
         SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307,
         SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309,
         SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311,
         SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313,
         SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315,
         SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317,
         SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319,
         SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321,
         SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323,
         SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325,
         SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327,
         SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329,
         SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331,
         SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333,
         SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335,
         SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337,
         SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339,
         SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341,
         SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343,
         SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345,
         SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347,
         SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349,
         SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351,
         SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353,
         SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355,
         SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357,
         SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359,
         SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361,
         SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363,
         SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365,
         SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367,
         SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369,
         SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371,
         SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373,
         SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375,
         SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377,
         SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379,
         SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381,
         SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383,
         SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385,
         SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387,
         SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389,
         SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391,
         SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393,
         SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395,
         SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397,
         SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399,
         SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401,
         SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403,
         SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405,
         SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407,
         SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409,
         SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411,
         SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413,
         SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415,
         SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417,
         SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419,
         SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421,
         SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423,
         SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425,
         SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427,
         SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429,
         SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431,
         SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433,
         SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435,
         SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437,
         SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439,
         SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441,
         SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443,
         SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445,
         SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447,
         SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449,
         SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451,
         SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453,
         SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455,
         SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457,
         SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459,
         SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461,
         SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463,
         SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465,
         SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467,
         SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469,
         SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471,
         SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473,
         SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475,
         SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477,
         SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479,
         SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481,
         SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483,
         SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485,
         SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487,
         SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489,
         SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491,
         SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493,
         SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495,
         SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497,
         SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499,
         SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501,
         SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503,
         SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505,
         SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507,
         SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509,
         SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511,
         SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513,
         SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515,
         SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517,
         SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519,
         SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521,
         SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523,
         SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525,
         SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527,
         SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529,
         SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531,
         SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533,
         SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535,
         SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537,
         SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539,
         SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541,
         SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543,
         SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545,
         SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547,
         SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549,
         SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551,
         SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553,
         SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555,
         SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557,
         SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559,
         SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561,
         SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563,
         SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565,
         SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567,
         SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569,
         SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571,
         SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573,
         SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575,
         SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577,
         SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579,
         SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581,
         SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583,
         SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585,
         SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587,
         SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589,
         SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591,
         SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593,
         SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595,
         SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597,
         SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599,
         SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601,
         SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603,
         SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605,
         SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607,
         SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609,
         SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611,
         SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613,
         SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615,
         SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617,
         SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619,
         SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621,
         SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623,
         SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625,
         SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627,
         SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629,
         SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631,
         SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633,
         SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635,
         SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637,
         SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639,
         SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641,
         SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643,
         SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645,
         SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647,
         SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649,
         SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651,
         SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653,
         SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655,
         SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657,
         SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659,
         SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661,
         SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663,
         SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665,
         SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667,
         SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669,
         SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671,
         SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673,
         SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675,
         SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677,
         SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679,
         SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681,
         SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683,
         SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685,
         SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687,
         SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689,
         SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691,
         SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693,
         SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695,
         SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697,
         SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699,
         SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701,
         SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703,
         SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705,
         SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707,
         SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709,
         SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711,
         SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713,
         SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715,
         SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717,
         SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719,
         SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721,
         SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723,
         SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725,
         SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727,
         SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729,
         SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731,
         SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733,
         SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735,
         SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737,
         SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739,
         SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741,
         SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743,
         SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745,
         SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747,
         SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749,
         SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751,
         SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753,
         SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755,
         SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757,
         SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759,
         SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761,
         SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763,
         SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765,
         SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767,
         SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769,
         SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771,
         SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773,
         SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775,
         SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777,
         SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779,
         SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781,
         SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783,
         SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785,
         SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787,
         SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789,
         SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791,
         SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793,
         SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795,
         SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797,
         SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799,
         SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801,
         SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803,
         SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805,
         SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807,
         SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809,
         SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811,
         SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813,
         SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815,
         SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817,
         SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819,
         SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821,
         SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823,
         SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825,
         SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827,
         SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829,
         SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831,
         SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833,
         SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835,
         SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837,
         SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839,
         SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841,
         SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843,
         SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845,
         SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847,
         SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849,
         SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851,
         SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853,
         SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855,
         SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857,
         SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859,
         SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861,
         SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863,
         SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865,
         SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867,
         SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869,
         SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871,
         SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873,
         SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875,
         SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877,
         SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879,
         SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881,
         SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883,
         SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885,
         SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887,
         SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889,
         SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891,
         SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893,
         SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895,
         SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897,
         SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899,
         SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901,
         SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903,
         SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905,
         SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907,
         SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909,
         SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911,
         SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913,
         SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915,
         SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917,
         SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919,
         SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921,
         SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923,
         SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925,
         SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927,
         SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929,
         SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931,
         SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933,
         SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935,
         SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937,
         SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939,
         SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941,
         SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943,
         SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945,
         SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947,
         SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949,
         SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951,
         SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953,
         SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955,
         SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957,
         SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959,
         SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961,
         SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963,
         SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965,
         SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967,
         SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969,
         SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971,
         SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973,
         SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975,
         SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977,
         SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979,
         SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981,
         SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983,
         SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985,
         SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987,
         SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989,
         SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991,
         SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993,
         SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995,
         SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997,
         SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999,
         SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001,
         SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003,
         SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005,
         SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007,
         SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009,
         SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011,
         SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013,
         SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015,
         SYNOPSYS_UNCONNECTED_1016;
  wire   [30:23] we;
  wire   [6:0] d_regx_addr;
  wire   [7:0] reg1F;
  wire   [3:2] reg1E;
  wire   [3:0] reg14;
  wire   [3:0] d_lt_gpi;
  wire   [5:0] lt_reg15_5_0;
  wire   [5:0] i2c_mode_wdat;
  wire   [5:0] d_lt_aswk;
  wire   [5:0] lt_aswk;
  wire   [7:0] wd18;

  INVX1 U116 ( .A(n92), .Y(n91) );
  INVX1 U117 ( .A(n92), .Y(n88) );
  INVX1 U118 ( .A(n93), .Y(n90) );
  INVX1 U119 ( .A(n92), .Y(n89) );
  INVX1 U120 ( .A(n93), .Y(n80) );
  INVX1 U121 ( .A(n93), .Y(n81) );
  INVX1 U122 ( .A(n92), .Y(n82) );
  INVX1 U123 ( .A(n93), .Y(n79) );
  INVX1 U124 ( .A(n94), .Y(n78) );
  INVX1 U125 ( .A(n94), .Y(n77) );
  INVX1 U126 ( .A(n94), .Y(n76) );
  INVX1 U127 ( .A(n92), .Y(n75) );
  INVX1 U128 ( .A(n93), .Y(n74) );
  INVX1 U129 ( .A(n92), .Y(n73) );
  INVX1 U130 ( .A(n93), .Y(n72) );
  INVX1 U131 ( .A(n93), .Y(n71) );
  INVX1 U132 ( .A(n92), .Y(n70) );
  INVX1 U133 ( .A(n93), .Y(n83) );
  INVX1 U134 ( .A(n93), .Y(n84) );
  INVX1 U135 ( .A(n92), .Y(n87) );
  INVX1 U136 ( .A(n92), .Y(n85) );
  INVX1 U137 ( .A(n93), .Y(n86) );
  INVX1 U140 ( .A(rrstz), .Y(n94) );
  INVX1 U141 ( .A(rrstz), .Y(n92) );
  INVX1 U142 ( .A(rrstz), .Y(n93) );
  glreg_a0_19 u0_reg04 ( .clk(clk), .arstz(n70), .we(we_4), .wdat({
        regx_wdat[7], n14, n11, n19, n8, n22, wd_twlb}), .rdat(r_bck0), 
        .test_si(r_xana[23]), .test_se(test_se) );
  glreg_a0_18 u0_reg05 ( .clk(clk), .arstz(n71), .we(we_5), .wdat({n118, n13, 
        regx_wdat[5], n19, n8, regx_wdat[2], wd_twlb}), .rdat(r_bck1), 
        .test_si(r_bck0[7]), .test_se(test_se) );
  glreg_a0_17 u0_reg06 ( .clk(clk), .arstz(n72), .we(we_6), .wdat({n16, n14, 
        n11, n18, n8, n22, wd_twlb}), .rdat(r_bck2), .test_si(r_bck1[7]), 
        .test_se(test_se) );
  glreg_a0_16 u0_reg07 ( .clk(clk), .arstz(n73), .we(we_7), .wdat({n118, n13, 
        n10, n18, regx_wdat[3], n21, wd_twlb}), .rdat(r_adummyi), .test_si2(
        test_si2), .test_si1(r_bck2[7]), .test_se(test_se) );
  glreg_WIDTH1_2 u0_reg10 ( .clk(clk), .arstz(n91), .we(1'b1), .wdat(ramacc), 
        .rdat(reg10_7_), .test_si(r_adummyi[7]), .test_se(test_se) );
  glreg_6_00000002 u0_reg12 ( .clk(clk), .arstz(n84), .we(we_twlb), .wdat({
        regx_wdat[7], n14, n11, n18, n8, n22}), .rdat({r_vpp_en, r_vpp0v_en, 
        r_otp_pwdn_en, r_otp_wpls, r_sap}), .test_si(reg10_7_), .test_se(
        test_se) );
  glreg_a0_15 u0_reg13 ( .clk(clk), .arstz(n74), .we(we_19), .wdat({n118, n14, 
        n10, n19, n8, n21, wd_twlb}), .rdat({r_dpdo_sel, r_dndo_sel}), 
        .test_si(r_vpp_en), .test_se(test_se) );
  glreg_WIDTH6_1 u0_reg15 ( .clk(clk), .arstz(n86), .we(n49), .wdat({n11, n18, 
        regx_wdat[3], n22, wd_twlb}), .rdat(lt_reg15_5_0), .test_si(
        r_dpdo_sel[3]), .test_se(test_se) );
  glreg_WIDTH6_0 u1_reg15 ( .clk(clk), .arstz(n85), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat({n148, r_i2crout[4:0]}), .test_si(r_xana[0]), 
        .test_se(test_se) );
  glreg_a0_14 u0_reg17 ( .clk(clk), .arstz(n75), .we(we[23]), .wdat({n16, n14, 
        n10, n19, n8, n21, wd_twlb}), .rdat(r_aopt), .test_si(lt_reg15_5_0[5]), 
        .test_se(test_se) );
  glreg_a0_13 u0_tmp18 ( .clk(clk), .arstz(n76), .we(we[24]), .wdat({n118, n13, 
        n11, n19, regx_wdat[3], n22, wd_twlb[1], n98}), .rdat(wd18), .test_si(
        bkpt_ena), .test_se(test_se) );
  glreg_a0_12 u0_reg18 ( .clk(clk), .arstz(n77), .we(n50), .wdat(wd18), .rdat(
        bkpt_pc[7:0]), .test_si(r_aopt[7]), .test_se(test_se) );
  glreg_a0_11 u0_reg19 ( .clk(clk), .arstz(n78), .we(n50), .wdat({n118, n14, 
        n11, n19, n8, n22, n101, n98}), .rdat({bkpt_ena, bkpt_pc[14:8]}), 
        .test_si(bkpt_pc[7]), .test_se(test_se) );
  glreg_a0_10 u0_reg1A ( .clk(clk), .arstz(n79), .we(we[26]), .wdat({n118, n14, 
        n11, n18, regx_wdat[3], n22, n101, n98}), .rdat(r_xtm), .test_si(n138), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_8 u0_ts_db ( .o_dbc(reg1B_3_), .o_chg(), .i_org(di_ts), 
        .clk(clk), .rstz(n89), .test_si(wd18[7]), .test_so(n137), .test_se(
        test_se) );
  glreg_WIDTH7_0 u0_reg1B ( .clk(clk), .arstz(n83), .we(we[27]), .wdat({n16, 
        n14, n10, n19, n21, n101, n98}), .rdat(r_do_ts), .test_si(r_xtm[7]), 
        .test_se(test_se) );
  glreg_WIDTH1_1 u1_reg1C ( .clk(clk), .arstz(n91), .we(upd_pwrv), .wdat(
        lt_reg1C_0), .rdat(r_xana[0]), .test_si(n136), .test_se(test_se) );
  glreg_a0_9 u0_reg1C ( .clk(clk), .arstz(n82), .we(we[28]), .wdat({n118, n13, 
        n11, n18, n8, n22, n101, n98}), .rdat({r_xana[7:1], lt_reg1C_0}), 
        .test_si(r_do_ts[6]), .test_se(test_se) );
  glreg_a0_8 u0_reg1D ( .clk(clk), .arstz(n81), .we(we[29]), .wdat({n118, n14, 
        n11, n19, regx_wdat[3], n22, n101, n98}), .rdat(r_xana[15:8]), 
        .test_si(r_xana[7]), .test_se(test_se) );
  glreg_a0_7 u0_reg1E ( .clk(clk), .arstz(n80), .we(we[30]), .wdat({n118, n14, 
        n11, n18, n8, n22, wd_twlb}), .rdat({r_xana[23], r_imp_osc, 
        r_xana[21:20], reg1E, r_xana[17:16]}), .test_si(r_xana[15]), .test_se(
        test_se) );
  dbnc_WIDTH2_TIMEOUT2_7 u0_dosc_db ( .o_dbc(reg14[1]), .o_chg(), .i_org(
        di_imposc), .clk(clk), .rstz(n91), .test_si(lt_drp), .test_so(n140), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_6 u0_iosc_db ( .o_dbc(reg14[2]), .o_chg(), .i_org(
        di_drposc), .clk(clk), .rstz(n91), .test_si(n140), .test_so(n139), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_5 u0_xana_db ( .o_dbc(reg1F[0]), .o_chg(), .i_org(
        di_xanav[0]), .clk(clk), .rstz(n90), .test_si(n137), .test_so(n136), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_4 u1_xana_db ( .o_dbc(reg1F[1]), .o_chg(), .i_org(
        di_xanav[1]), .clk(clk), .rstz(n90), .test_si(n61), .test_so(n135), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_3 u2_xana_db ( .o_dbc(reg1F[2]), .o_chg(), .i_org(
        di_xanav[2]), .clk(clk), .rstz(n88), .test_si(n135), .test_so(n134), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_2 u3_xana_db ( .o_dbc(reg1F[3]), .o_chg(), .i_org(
        di_xanav[3]), .clk(clk), .rstz(n89), .test_si(n134), .test_so(n133), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_1 u4_xana_db ( .o_dbc(reg1F[4]), .o_chg(), .i_org(
        di_xanav[4]), .clk(clk), .rstz(n86), .test_si(n133), .test_so(n132), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_0 u5_xana_db ( .o_dbc(reg1F[5]), .o_chg(), .i_org(
        di_xanav[5]), .clk(clk), .rstz(n84), .test_si(n132), .test_so(n131), 
        .test_se(test_se) );
  dbnc_a0_1 u6_xana_db ( .o_dbc(reg1F[6]), .o_chg(), .i_org(di_xanav[0]), 
        .clk(clk_500k), .rstz(n87), .test_si(n131), .test_so(test_so1), 
        .test_se(test_se) );
  dbnc_a0_0 u0_rdet_db ( .o_dbc(reg1F[7]), .o_chg(), .i_org(di_rd_det), .clk(
        clk_500k), .rstz(n88), .test_si(n139), .test_so(n138), .test_se(
        test_se) );
  SNPS_CLOCK_GATE_HIGH_regx_a0 clk_gate_d_lt_gpi_reg ( .CLK(clk), .EN(n94), 
        .ENCLK(net8997), .TE(test_se) );
  regx_a0_DW_rightsh_1 srl_66 ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        dac_comp[9:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_sar_en[9:8], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_dac_en[9:8], 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_comp[7:0], r_sar_en[7:0], r_dac_en[7:0], dac_r_vs[63:0], 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_r_vs[79:64], reg1F, r_xana[23], r_imp_osc, r_xana[21:20], reg1E, 
        r_xana[17:0], r_do_ts[6:3], reg1B_3_, r_do_ts[2:0], r_xtm, bkpt_ena, 
        bkpt_pc, r_aopt, 1'b0, 1'b0, d_lt_aswk, sse_idle, 1'b0, n59, 
        r_i2crout[4:0], d_lt_gpi, reg14, r_dpdo_sel, r_dndo_sel, r_vpp_en, 
        r_vpp0v_en, r_otp_pwdn_en, r_otp_wpls, r_sap, r_twlb, r_bistdat, 
        reg10_7_, r_bistctl, r_sdischg, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_pwm, 
        r_adummyi, r_bck2, r_bck1, r_bck0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, r_cvofsx, r_idacsh, r_vcomp}), .DATA_TC(1'b0), .SH({
        d_regx_addr[6], n95, d_regx_addr[4:0], 1'b0, 1'b0, 1'b0}), .B({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, 
        SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, 
        SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, 
        SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, 
        SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, 
        SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, 
        SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, 
        SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, 
        SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, 
        SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, 
        SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, 
        SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, 
        SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, 
        SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, 
        SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, 
        SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, 
        SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, 
        SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, 
        SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, 
        SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, 
        SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, 
        SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, 
        SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, 
        SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, 
        SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, 
        SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, 
        SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, 
        SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, 
        SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, 
        SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, 
        SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, 
        SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, 
        SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, 
        SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, 
        SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, 
        SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, 
        SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, 
        SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, 
        SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, 
        SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, 
        SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, 
        SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, 
        SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, 
        SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, 
        SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, 
        SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, 
        SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, 
        SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, 
        SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, 
        SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, 
        SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, 
        SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, 
        SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, 
        SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, 
        SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, 
        SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, 
        SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, 
        SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, 
        SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, 
        SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, 
        SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, 
        SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, 
        SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, 
        SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, 
        SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, 
        SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, 
        SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, 
        SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, 
        SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, 
        SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, 
        SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, 
        SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, 
        SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, 
        SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, 
        SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, 
        SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, 
        SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, 
        SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, 
        SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, 
        SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, 
        SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, 
        SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, 
        SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, 
        SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, 
        SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, 
        SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, 
        SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, 
        SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, 
        SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, 
        SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, 
        SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, 
        SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, 
        SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, 
        SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, 
        SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, 
        SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, 
        SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, 
        SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, 
        SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, 
        SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, 
        SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, 
        SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, 
        SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, 
        SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, 
        SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, 
        SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, 
        SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, 
        SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, 
        SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, 
        SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, 
        SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, 
        SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, 
        SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, 
        SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, 
        SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, 
        SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, 
        SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, 
        SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, 
        SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, 
        SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, 
        SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, 
        SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, 
        SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, 
        SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, 
        SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, 
        SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, 
        SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, 
        SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, 
        SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, 
        SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, 
        SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, 
        SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, 
        SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, 
        SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, 
        SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, 
        SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, 
        SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, 
        SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, 
        SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, 
        SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, 
        SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, 
        SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, 
        SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, 
        SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, 
        SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, 
        SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, 
        SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, 
        SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, 
        SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, 
        SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, 
        SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, 
        SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, 
        SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, 
        SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, 
        SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, 
        SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, 
        SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, 
        SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, 
        SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, 
        SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, 
        SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, 
        SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, 
        SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, 
        SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, 
        SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, 
        SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, 
        SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, 
        SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, 
        SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, 
        SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, 
        SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, 
        SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, 
        SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, 
        SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, 
        SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, 
        SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, 
        SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, 
        SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, 
        SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, 
        SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, 
        SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, 
        SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, 
        SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, 
        SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, 
        SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, 
        SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, 
        SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, 
        SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, 
        SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, 
        SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, 
        SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, 
        SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, 
        SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, 
        SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, 
        SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, 
        SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, 
        SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, 
        SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, 
        SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, 
        SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, 
        SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, 
        SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, 
        SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, 
        SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, 
        SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, 
        SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, 
        SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, 
        SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, 
        SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, 
        SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, 
        SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, 
        SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, 
        SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, 
        SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, 
        SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, 
        SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, 
        SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, 
        SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, 
        SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, 
        SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, 
        SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, 
        SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, 
        SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, 
        SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, 
        SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, 
        SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, 
        SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, 
        SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, 
        SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, 
        SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, 
        SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, 
        SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, 
        SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, 
        SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, 
        SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, 
        SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, 
        SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, 
        SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, 
        SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, 
        SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, 
        SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, 
        SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, 
        SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, 
        SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, 
        SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, 
        SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, 
        SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, 
        SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, 
        SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, 
        SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, 
        SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, 
        SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, 
        SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, 
        SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, 
        SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, 
        SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, 
        SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, 
        SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, 
        SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, 
        SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, 
        SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, 
        SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, 
        SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, 
        SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, 
        SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, 
        SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, 
        SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, 
        SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, 
        SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, 
        SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, 
        SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, 
        SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, 
        SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, 
        SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, 
        SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, 
        SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, 
        SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, 
        SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, 
        SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, 
        SYNOPSYS_UNCONNECTED_1016, regx_rdat}) );
  SDFFQX1 d_regx_addr_reg_3_ ( .D(n30), .SIN(d_regx_addr[2]), .SMC(test_se), 
        .C(clk), .Q(d_regx_addr[3]) );
  SDFFQX1 d_we16_reg ( .D(N8), .SIN(d_regx_addr[6]), .SMC(test_se), .C(clk), 
        .Q(d_we16) );
  SDFFQX1 d_lt_aswk_reg_2_ ( .D(lt_aswk[2]), .SIN(d_lt_aswk[1]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[2]) );
  SDFFQX1 d_lt_aswk_reg_1_ ( .D(lt_aswk[1]), .SIN(d_lt_aswk[0]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[1]) );
  SDFFQX1 d_lt_drp_reg ( .D(lt_drp), .SIN(d_lt_aswk[5]), .SMC(test_se), .C(clk), .Q(reg14[0]) );
  SDFFQX1 d_lt_gpi_reg_0_ ( .D(lt_gpi[0]), .SIN(reg14[0]), .SMC(test_se), .C(
        net8997), .Q(d_lt_gpi[0]) );
  SDFFQX1 d_lt_aswk_reg_4_ ( .D(lt_aswk[4]), .SIN(d_lt_aswk[3]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[4]) );
  SDFFQX1 d_lt_aswk_reg_0_ ( .D(lt_aswk[0]), .SIN(reg14[3]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[0]) );
  SDFFQX1 d_regx_addr_reg_1_ ( .D(regx_addr[1]), .SIN(d_regx_addr[0]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[1]) );
  SDFFQX1 d_regx_addr_reg_0_ ( .D(regx_addr[0]), .SIN(d_lt_gpi[3]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[0]) );
  SDFFQX1 d_di_tst_reg ( .D(di_tst), .SIN(test_si1), .SMC(test_se), .C(clk), 
        .Q(reg14[3]) );
  SDFFQX1 d_lt_gpi_reg_1_ ( .D(lt_gpi[1]), .SIN(d_lt_gpi[0]), .SMC(test_se), 
        .C(net8997), .Q(d_lt_gpi[1]) );
  SDFFQX1 d_lt_aswk_reg_5_ ( .D(lt_aswk[5]), .SIN(d_lt_aswk[4]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[5]) );
  SDFFQX1 d_lt_aswk_reg_3_ ( .D(lt_aswk[3]), .SIN(d_lt_aswk[2]), .SMC(test_se), 
        .C(clk), .Q(d_lt_aswk[3]) );
  SDFFQX1 d_lt_gpi_reg_2_ ( .D(lt_gpi[2]), .SIN(d_lt_gpi[1]), .SMC(test_se), 
        .C(net8997), .Q(d_lt_gpi[2]) );
  SDFFQX1 d_lt_gpi_reg_3_ ( .D(lt_gpi[3]), .SIN(d_lt_gpi[2]), .SMC(test_se), 
        .C(net8997), .Q(d_lt_gpi[3]) );
  SDFFQX1 d_regx_addr_reg_2_ ( .D(n57), .SIN(d_regx_addr[1]), .SMC(test_se), 
        .C(clk), .Q(d_regx_addr[2]) );
  SDFFQX1 d_regx_addr_reg_4_ ( .D(n52), .SIN(d_regx_addr[3]), .SMC(test_se), 
        .C(clk), .Q(d_regx_addr[4]) );
  SDFFQX1 d_regx_addr_reg_6_ ( .D(regx_addr[6]), .SIN(d_regx_addr[5]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[6]) );
  SDFFQX1 d_regx_addr_reg_5_ ( .D(regx_addr[5]), .SIN(d_regx_addr[4]), .SMC(
        test_se), .C(clk), .Q(d_regx_addr[5]) );
  SDFFRQX1 lt_drp_reg ( .D(di_drposc), .SIN(lt_aswk[5]), .SMC(test_se), .C(
        detclk), .XR(n87), .Q(lt_drp) );
  SDFFRQX1 lt_aswk_reg_5_ ( .D(1'b1), .SIN(lt_aswk[4]), .SMC(test_se), .C(
        aswclk), .XR(n6), .Q(lt_aswk[5]) );
  SDFFRQX1 lt_aswk_reg_4_ ( .D(di_aswk[4]), .SIN(lt_aswk[3]), .SMC(test_se), 
        .C(aswclk), .XR(n6), .Q(lt_aswk[4]) );
  SDFFRQX1 lt_aswk_reg_3_ ( .D(di_aswk[3]), .SIN(lt_aswk[2]), .SMC(test_se), 
        .C(aswclk), .XR(n6), .Q(lt_aswk[3]) );
  SDFFRQX1 lt_aswk_reg_2_ ( .D(di_aswk[2]), .SIN(lt_aswk[1]), .SMC(test_se), 
        .C(aswclk), .XR(n6), .Q(lt_aswk[2]) );
  SDFFRQX1 lt_aswk_reg_1_ ( .D(di_aswk[1]), .SIN(lt_aswk[0]), .SMC(test_se), 
        .C(aswclk), .XR(n6), .Q(lt_aswk[1]) );
  SDFFRQX1 lt_aswk_reg_0_ ( .D(di_aswk[0]), .SIN(d_we16), .SMC(test_se), .C(
        aswclk), .XR(n6), .Q(lt_aswk[0]) );
  AND2X1 U4 ( .A(n67), .B(regx_addr[0]), .Y(n54) );
  INVX3 U7 ( .A(n1), .Y(n5) );
  NAND2X1 U8 ( .A(regx_addr[5]), .B(regx_w), .Y(n1) );
  INVX3 U9 ( .A(regx_addr[6]), .Y(n122) );
  AND3XL U10 ( .A(n65), .B(n145), .C(n141), .Y(regx_wrdac[0]) );
  NOR2XL U11 ( .A(regx_addr[4]), .B(n141), .Y(n62) );
  INVX4 U12 ( .A(regx_addr[2]), .Y(n28) );
  AND3X2 U13 ( .A(n146), .B(n65), .C(n141), .Y(regx_wrdac[1]) );
  NOR2X1 U14 ( .A(n129), .B(n125), .Y(n65) );
  NAND3X2 U15 ( .A(n122), .B(regx_w), .C(regx_addr[5]), .Y(n125) );
  INVX2 U16 ( .A(n62), .Y(n63) );
  NAND32X1 U17 ( .B(regx_addr[3]), .C(n125), .A(n129), .Y(n126) );
  AND2XL U18 ( .A(n146), .B(n37), .Y(regx_wrdac[3]) );
  INVX2 U19 ( .A(n115), .Y(n123) );
  NAND32X1 U20 ( .B(n107), .C(n28), .A(n53), .Y(n115) );
  AND2X1 U21 ( .A(n127), .B(n145), .Y(regx_wrdac[12]) );
  INVX1 U22 ( .A(n31), .Y(n108) );
  INVX1 U23 ( .A(n141), .Y(n30) );
  NAND2X2 U24 ( .A(n122), .B(n5), .Y(n23) );
  NOR32XL U25 ( .B(n107), .C(regx_addr[1]), .A(n57), .Y(n36) );
  AND3XL U26 ( .A(regx_addr[0]), .B(regx_addr[1]), .C(n28), .Y(n56) );
  INVXL U27 ( .A(n28), .Y(n57) );
  NAND21X2 U28 ( .B(regx_addr[0]), .A(n67), .Y(n103) );
  INVX2 U29 ( .A(regx_addr[3]), .Y(n141) );
  NOR32XL U30 ( .B(n107), .C(regx_addr[2]), .A(regx_addr[1]), .Y(n66) );
  INVX1 U31 ( .A(regx_addr[4]), .Y(n129) );
  OA21X1 U32 ( .B(atpg_en), .C(n111), .A(n85), .Y(n6) );
  INVXL U33 ( .A(regx_wdat[3]), .Y(n7) );
  INVXL U34 ( .A(n7), .Y(n8) );
  INVXL U35 ( .A(regx_wdat[5]), .Y(n9) );
  INVXL U36 ( .A(n9), .Y(n10) );
  INVXL U37 ( .A(n9), .Y(n11) );
  INVXL U38 ( .A(regx_wdat[6]), .Y(n12) );
  INVXL U39 ( .A(n12), .Y(n13) );
  INVXL U40 ( .A(n12), .Y(n14) );
  INVXL U41 ( .A(regx_wdat[7]), .Y(n15) );
  INVXL U42 ( .A(n15), .Y(n16) );
  INVXL U43 ( .A(regx_wdat[4]), .Y(n17) );
  INVXL U44 ( .A(n17), .Y(n18) );
  INVXL U45 ( .A(n17), .Y(n19) );
  INVXL U46 ( .A(regx_wdat[2]), .Y(n20) );
  INVXL U47 ( .A(n20), .Y(n21) );
  INVXL U48 ( .A(n20), .Y(n22) );
  INVX4 U49 ( .A(regx_addr[1]), .Y(n68) );
  AND2X1 U50 ( .A(n45), .B(n145), .Y(regx_wrdac[2]) );
  BUFXL U51 ( .A(n67), .Y(n25) );
  INVX2 U52 ( .A(n104), .Y(n146) );
  NAND43X1 U53 ( .B(regx_addr[6]), .C(regx_addr[5]), .D(n30), .A(n52), .Y(n144) );
  NAND21XL U54 ( .B(regx_addr[0]), .A(n25), .Y(n26) );
  AND2XL U55 ( .A(regx_addr[0]), .B(n25), .Y(n27) );
  INVX1 U56 ( .A(regx_addr[0]), .Y(n107) );
  INVX2 U57 ( .A(regx_addr[0]), .Y(n29) );
  NOR2X1 U58 ( .A(n23), .B(n63), .Y(n64) );
  AND3X2 U59 ( .A(n146), .B(n30), .C(n65), .Y(regx_wrdac[11]) );
  NOR2X2 U60 ( .A(n23), .B(n63), .Y(n45) );
  BUFXL U61 ( .A(n36), .Y(n31) );
  NOR2X2 U62 ( .A(n63), .B(n23), .Y(n37) );
  INVXL U63 ( .A(n26), .Y(n32) );
  INVX3 U64 ( .A(n103), .Y(n124) );
  BUFXL U65 ( .A(n145), .Y(n34) );
  AND3X2 U66 ( .A(n145), .B(n30), .C(n65), .Y(regx_wrdac[10]) );
  BUFXL U67 ( .A(n56), .Y(n48) );
  AND2X1 U68 ( .A(n66), .B(n64), .Y(regx_wrdac[6]) );
  BUFXL U69 ( .A(n27), .Y(n51) );
  NAND32X1 U70 ( .B(n29), .C(regx_addr[1]), .A(n28), .Y(n104) );
  INVXL U71 ( .A(n129), .Y(n52) );
  AND2X2 U72 ( .A(n56), .B(n37), .Y(regx_wrdac[5]) );
  INVXL U73 ( .A(regx_addr[1]), .Y(n53) );
  AND2X4 U74 ( .A(n123), .B(n37), .Y(regx_wrdac[7]) );
  AND2X2 U75 ( .A(n36), .B(n45), .Y(regx_wrdac[4]) );
  AND2XL U76 ( .A(n114), .B(n51), .Y(we[23]) );
  AND2XL U77 ( .A(n51), .B(n143), .Y(regx_wrcvc[3]) );
  AND2X2 U78 ( .A(n124), .B(n45), .Y(regx_wrdac[8]) );
  AND2X2 U79 ( .A(n127), .B(n146), .Y(regx_wrdac[13]) );
  BUFXL U80 ( .A(n146), .Y(n55) );
  INVX1 U81 ( .A(n148), .Y(n58) );
  INVX1 U82 ( .A(n58), .Y(n59) );
  INVX1 U83 ( .A(n58), .Y(r_i2crout[5]) );
  INVX1 U84 ( .A(n58), .Y(n61) );
  BUFX3 U85 ( .A(r_imp_osc), .Y(r_xana[22]) );
  AND2XL U86 ( .A(n34), .B(n147), .Y(regx_hitbst[0]) );
  AND2XL U87 ( .A(n128), .B(n145), .Y(regx_wrcvc[0]) );
  AND2XL U88 ( .A(n143), .B(n34), .Y(regx_wrpwm[0]) );
  AND2XL U89 ( .A(n66), .B(n128), .Y(we_4) );
  AND2XL U90 ( .A(n66), .B(n113), .Y(we[28]) );
  AND2XL U91 ( .A(n34), .B(n113), .Y(we[24]) );
  INVXL U92 ( .A(regx_wdat[0]), .Y(n99) );
  NOR2X4 U93 ( .A(n28), .B(n68), .Y(n67) );
  AND2X2 U94 ( .A(n54), .B(n37), .Y(regx_wrdac[9]) );
  INVX1 U95 ( .A(n116), .Y(n49) );
  NAND21XL U96 ( .B(n115), .A(n114), .Y(n116) );
  AND2XL U97 ( .A(n123), .B(n113), .Y(we[29]) );
  AND2X1 U98 ( .A(n48), .B(n113), .Y(we[27]) );
  AND2X1 U99 ( .A(n31), .B(n113), .Y(we[26]) );
  AND2X1 U100 ( .A(n114), .B(n48), .Y(we_19) );
  INVX1 U101 ( .A(n99), .Y(wd_twlb[0]) );
  INVX1 U102 ( .A(n102), .Y(wd_twlb[1]) );
  INVX1 U103 ( .A(n99), .Y(n98) );
  INVX1 U104 ( .A(n102), .Y(n101) );
  INVX1 U105 ( .A(n33), .Y(n130) );
  INVX1 U106 ( .A(n144), .Y(n147) );
  AND2XL U107 ( .A(n31), .B(n128), .Y(regx_wrcvc[2]) );
  AND2XL U108 ( .A(n128), .B(n55), .Y(regx_wrcvc[1]) );
  INVX1 U109 ( .A(n106), .Y(n114) );
  NAND21X1 U110 ( .B(n144), .A(regx_w), .Y(n106) );
  INVX1 U111 ( .A(n142), .Y(n143) );
  NAND32XL U112 ( .B(n141), .C(n130), .A(n129), .Y(n142) );
  INVX1 U113 ( .A(n109), .Y(we_twlb) );
  NAND21XL U114 ( .B(n108), .A(n114), .Y(n109) );
  INVX1 U115 ( .A(n24), .Y(n113) );
  INVX1 U138 ( .A(n105), .Y(n50) );
  NAND21XL U139 ( .B(n24), .A(n55), .Y(n105) );
  AND2XL U143 ( .A(n143), .B(n55), .Y(regx_wrpwm[1]) );
  AND2X1 U144 ( .A(n32), .B(n113), .Y(we[30]) );
  AND2X1 U145 ( .A(n32), .B(n128), .Y(we_6) );
  AND2XL U146 ( .A(n123), .B(n128), .Y(we_5) );
  AND2XL U147 ( .A(n128), .B(n51), .Y(we_7) );
  AND2XL U148 ( .A(n147), .B(n55), .Y(regx_hitbst[1]) );
  INVX1 U149 ( .A(regx_wdat[1]), .Y(n102) );
  INVX1 U150 ( .A(n15), .Y(n118) );
  INVX2 U151 ( .A(n112), .Y(n145) );
  INVX1 U152 ( .A(n96), .Y(n95) );
  INVX1 U153 ( .A(n121), .Y(n128) );
  NOR43XL U154 ( .B(n102), .C(n20), .D(n110), .A(n46), .Y(N8) );
  NAND3X1 U155 ( .A(n17), .B(n9), .C(n7), .Y(n46) );
  AND4XL U156 ( .A(wd_twlb[0]), .B(n47), .C(n114), .D(n32), .Y(n110) );
  AO21X1 U157 ( .B(bus_idle), .C(n120), .A(n119), .Y(i2c_mode_upd) );
  AND3X1 U158 ( .A(n49), .B(n118), .C(n12), .Y(n119) );
  NAND32X1 U159 ( .B(n38), .C(n49), .A(n117), .Y(n120) );
  NOR21XL U160 ( .B(n13), .A(n15), .Y(n47) );
  XNOR2XL U161 ( .A(reg1E[3]), .B(n35), .Y(r_xana[19]) );
  XNOR2XL U162 ( .A(reg1E[2]), .B(n35), .Y(r_xana[18]) );
  NAND2X1 U163 ( .A(r_xana[20]), .B(di_drposc), .Y(n35) );
  INVX1 U164 ( .A(d_regx_addr[5]), .Y(n96) );
  MUX2X1 U165 ( .D0(lt_reg15_5_0[2]), .D1(n21), .S(n49), .Y(i2c_mode_wdat[2])
         );
  MUX2X1 U166 ( .D0(lt_reg15_5_0[0]), .D1(n98), .S(n49), .Y(i2c_mode_wdat[0])
         );
  MUX2X1 U167 ( .D0(lt_reg15_5_0[1]), .D1(n101), .S(n49), .Y(i2c_mode_wdat[1])
         );
  MUX2BXL U168 ( .D0(lt_reg15_5_0[5]), .D1(n9), .S(n49), .Y(i2c_mode_wdat[5])
         );
  MUX2BXL U169 ( .D0(lt_reg15_5_0[4]), .D1(n17), .S(n49), .Y(i2c_mode_wdat[4])
         );
  MUX2BXL U170 ( .D0(lt_reg15_5_0[3]), .D1(n7), .S(n49), .Y(i2c_mode_wdat[3])
         );
  NAND3X1 U171 ( .A(n39), .B(n40), .C(n41), .Y(n38) );
  XNOR2XL U172 ( .A(r_i2crout[3]), .B(lt_reg15_5_0[3]), .Y(n41) );
  XNOR2XL U173 ( .A(r_i2crout[4]), .B(lt_reg15_5_0[4]), .Y(n39) );
  XNOR2XL U174 ( .A(n61), .B(lt_reg15_5_0[5]), .Y(n40) );
  AND3X1 U175 ( .A(n43), .B(n44), .C(n42), .Y(n117) );
  XNOR2XL U176 ( .A(r_i2crout[1]), .B(lt_reg15_5_0[1]), .Y(n44) );
  XNOR2XL U177 ( .A(r_i2crout[0]), .B(lt_reg15_5_0[0]), .Y(n43) );
  XNOR2XL U178 ( .A(r_i2crout[2]), .B(lt_reg15_5_0[2]), .Y(n42) );
  INVX1 U179 ( .A(d_we16), .Y(n111) );
  INVX2 U180 ( .A(n126), .Y(n127) );
  NAND3XL U181 ( .A(n33), .B(n52), .C(n30), .Y(n24) );
  NOR31XL U182 ( .C(regx_w), .A(regx_addr[6]), .B(regx_addr[5]), .Y(n33) );
  NAND32XL U183 ( .B(n30), .C(n130), .A(n129), .Y(n121) );
  NAND32X1 U184 ( .B(regx_addr[0]), .C(regx_addr[1]), .A(n28), .Y(n112) );
endmodule


module regx_a0_DW_rightsh_1 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70, n72, n74, n75,
         n77, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n151,
         n154, n155, n156, n157, n158, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n197, n198, n202, n203, n205,
         n209, n210, n211, n212, n213, n214, n215, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n243,
         n247, n251, n254, n297, n299, n302, n303, n305, n307, n310, n311,
         n312, n313, n315, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n342, n343, n345, n347, n350, n351, n353, n354, n355,
         n356, n357, n358, n359, n361, n363, n366, n367, n368, n369, n371,
         n374, n375, n376, n385, n386, n387, n388, n389, n390, n391, n392,
         n416, n425, n427, n430, n431, n433, n435, n438, n439, n440, n441,
         n443, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n465, n466, n467, n470, n471, n473, n475, n478, n479, n480, n505,
         n507, n509, n511, n513, n515, n517, n519, n521, n523, n525, n527,
         n529, n531, n533, n535, n553, n555, n557, n559, n561, n563, n565,
         n567, n569, n572, n575, n578, n581, n584, n587, n590, n593, n596,
         n599, n602, n605, n608, n611, n614, n617, n620, n623, n626, n629,
         n632, n635, n638, n689, n691, n693, n695, n697, n699, n701, n703,
         n705, n707, n709, n711, n713, n715, n717, n719, n721, n724, n727,
         n730, n733, n736, n739, n742, n745, n748, n751, n754, n757, n760,
         n763, n766, n769, n772, n775, n778, n781, n784, n787, n790, n796,
         n799, n802, n805, n808, n811, n814, n817, n820, n823, n826, n829,
         n832, n835, n838, n841, n844, n847, n850, n853, n856, n859, n862,
         n865, n868, n871, n874, n877, n880, n883, n886, n889, n892, n895,
         n898, n901, n904, n907, n910, n913, n916, n919, n922, n925, n928,
         n931, n934, n937, n940, n943, n946, n949, n952, n955, n958, n961,
         n964, n967, n970, n973, n976, n979, n982, n1033, n1035, n1037, n1039,
         n1041, n1043, n1045, n1047, n1057, n1059, n1061, n1063, n1065, n1067,
         n1069, n1071, n1073, n1076, n1079, n1082, n1085, n1088, n1091, n1094,
         n1097, n1100, n1103, n1106, n1109, n1112, n1115, n1118, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1296, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443;

  MUX2IX4 U4 ( .D0(n5), .D1(n13), .S(SH[3]), .Y(B[4]) );
  MUX2IX4 U5 ( .D0(n4), .D1(n12), .S(SH[3]), .Y(B[3]) );
  MUX2IX4 U9 ( .D0(n32), .D1(n48), .S(n3367), .Y(n16) );
  MUX2IX4 U13 ( .D0(n28), .D1(n44), .S(n3367), .Y(n12) );
  MUX2IX4 U20 ( .D0(n21), .D1(n37), .S(n3368), .Y(n5) );
  MUX2IX4 U21 ( .D0(n20), .D1(n36), .S(n3367), .Y(n4) );
  MUX2IX4 U35 ( .D0(n70), .D1(n102), .S(n3374), .Y(n38) );
  MUX2IX4 U40 ( .D0(n65), .D1(n97), .S(n3374), .Y(n33) );
  MUX2IX4 U65 ( .D0(n232), .D1(n1232), .S(n3219), .Y(n104) );
  MUX2IX4 U66 ( .D0(n231), .D1(n3202), .S(n3233), .Y(n103) );
  MUX2IX4 U72 ( .D0(n193), .D1(n225), .S(n3230), .Y(n97) );
  MUX2IX4 U241 ( .D0(n3203), .D1(n368), .S(n3241), .Y(n120) );
  NAND21X1 U548 ( .B(n3440), .A(n505), .Y(n1360) );
  NOR2X1 U550 ( .A(n3401), .B(A[247]), .Y(n505) );
  NAND21X1 U554 ( .B(SH[9]), .A(n507), .Y(n1359) );
  NOR2X1 U556 ( .A(n3401), .B(A[246]), .Y(n507) );
  NAND21X1 U560 ( .B(n3417), .A(n509), .Y(n1358) );
  NOR2X1 U562 ( .A(n3401), .B(A[245]), .Y(n509) );
  NAND21X1 U566 ( .B(n3417), .A(n511), .Y(n1357) );
  NOR2X1 U568 ( .A(n3401), .B(A[244]), .Y(n511) );
  NAND21X1 U572 ( .B(n3417), .A(n513), .Y(n1356) );
  NOR2X1 U574 ( .A(n3402), .B(A[243]), .Y(n513) );
  NAND21X1 U578 ( .B(n3417), .A(n515), .Y(n1355) );
  NOR2X1 U580 ( .A(n3402), .B(A[242]), .Y(n515) );
  NAND21X1 U584 ( .B(n3417), .A(n517), .Y(n1354) );
  NOR2X1 U586 ( .A(n3402), .B(A[241]), .Y(n517) );
  NAND21X1 U590 ( .B(n3417), .A(n519), .Y(n1353) );
  NOR2X1 U592 ( .A(n3402), .B(A[240]), .Y(n519) );
  NAND21X1 U596 ( .B(n3417), .A(n521), .Y(n1352) );
  NOR2X1 U598 ( .A(n3406), .B(A[239]), .Y(n521) );
  NAND21X1 U602 ( .B(n3417), .A(n523), .Y(n1351) );
  NOR2X1 U604 ( .A(n3406), .B(A[238]), .Y(n523) );
  NAND21X1 U608 ( .B(n3417), .A(n525), .Y(n1350) );
  NOR2X1 U610 ( .A(n3406), .B(A[237]), .Y(n525) );
  NAND21X1 U614 ( .B(n3417), .A(n527), .Y(n1349) );
  NOR2X1 U616 ( .A(n3406), .B(A[236]), .Y(n527) );
  NAND21X1 U620 ( .B(n3418), .A(n529), .Y(n1348) );
  NOR2X1 U622 ( .A(n3406), .B(A[235]), .Y(n529) );
  NAND21X1 U626 ( .B(n3418), .A(n531), .Y(n1347) );
  NOR2X1 U628 ( .A(n3407), .B(A[234]), .Y(n531) );
  NAND21X1 U632 ( .B(n3418), .A(n533), .Y(n1346) );
  NOR2X1 U634 ( .A(n3407), .B(A[233]), .Y(n533) );
  NAND21X1 U638 ( .B(n3418), .A(n535), .Y(n1345) );
  NOR2X1 U640 ( .A(n3407), .B(A[232]), .Y(n535) );
  NAND21X1 U692 ( .B(n3419), .A(n553), .Y(n1336) );
  NOR2X1 U694 ( .A(n3408), .B(A[223]), .Y(n553) );
  NAND21X1 U698 ( .B(n3419), .A(n555), .Y(n1335) );
  NOR2X1 U700 ( .A(n3408), .B(A[222]), .Y(n555) );
  NAND21X1 U704 ( .B(n3419), .A(n557), .Y(n1334) );
  NOR2X1 U706 ( .A(n3408), .B(A[221]), .Y(n557) );
  NAND21X1 U710 ( .B(n3419), .A(n559), .Y(n1333) );
  NOR2X1 U712 ( .A(n3408), .B(A[220]), .Y(n559) );
  NAND21X1 U716 ( .B(n3419), .A(n561), .Y(n1332) );
  NOR2X1 U718 ( .A(n3408), .B(A[219]), .Y(n561) );
  NAND21X1 U722 ( .B(n3419), .A(n563), .Y(n1331) );
  NOR2X1 U724 ( .A(n3408), .B(A[218]), .Y(n563) );
  NAND21X1 U728 ( .B(n3419), .A(n565), .Y(n1330) );
  NOR2X1 U730 ( .A(n3408), .B(A[217]), .Y(n565) );
  NAND21X1 U734 ( .B(n3419), .A(n567), .Y(n1329) );
  NOR2X1 U736 ( .A(n3408), .B(A[216]), .Y(n567) );
  NAND21X1 U740 ( .B(n3420), .A(n569), .Y(n1328) );
  NAND21X1 U743 ( .B(n3395), .A(A[215]), .Y(n569) );
  NAND21X1 U747 ( .B(n3420), .A(n572), .Y(n1327) );
  NAND21X1 U750 ( .B(n3395), .A(A[214]), .Y(n572) );
  NAND21X1 U754 ( .B(n3420), .A(n575), .Y(n1326) );
  NAND21X1 U757 ( .B(n3395), .A(A[213]), .Y(n575) );
  NAND21X1 U761 ( .B(n3420), .A(n578), .Y(n1325) );
  NAND21X1 U764 ( .B(n3395), .A(A[212]), .Y(n578) );
  NAND21X1 U768 ( .B(n3420), .A(n581), .Y(n1324) );
  NAND21X1 U771 ( .B(n3395), .A(A[211]), .Y(n581) );
  NAND21X1 U775 ( .B(n3420), .A(n584), .Y(n1323) );
  NAND21X1 U778 ( .B(n3396), .A(A[210]), .Y(n584) );
  NAND21X1 U782 ( .B(n3420), .A(n587), .Y(n1322) );
  NAND21X1 U789 ( .B(n3420), .A(n590), .Y(n1321) );
  NAND21X1 U796 ( .B(n3420), .A(n593), .Y(n1320) );
  NAND21X1 U799 ( .B(n3396), .A(A[207]), .Y(n593) );
  NAND21X1 U803 ( .B(n3420), .A(n596), .Y(n1319) );
  NAND21X1 U806 ( .B(n3396), .A(A[206]), .Y(n596) );
  NAND21X1 U810 ( .B(n3421), .A(n599), .Y(n1318) );
  NAND21X1 U813 ( .B(n3395), .A(A[205]), .Y(n599) );
  NAND21X1 U817 ( .B(n3421), .A(n602), .Y(n1317) );
  NAND21X1 U820 ( .B(n3396), .A(A[204]), .Y(n602) );
  NAND21X1 U824 ( .B(n3421), .A(n605), .Y(n1316) );
  NAND21X1 U827 ( .B(n3395), .A(A[203]), .Y(n605) );
  NAND21X1 U831 ( .B(n3421), .A(n608), .Y(n1315) );
  NAND21X1 U834 ( .B(n3395), .A(A[202]), .Y(n608) );
  NAND21X1 U838 ( .B(n3421), .A(n611), .Y(n1314) );
  NAND21X1 U845 ( .B(n3421), .A(n614), .Y(n1313) );
  NAND21X1 U852 ( .B(n3421), .A(n617), .Y(n1312) );
  NAND21X1 U855 ( .B(n3396), .A(A[199]), .Y(n617) );
  NAND21X1 U859 ( .B(n3421), .A(n620), .Y(n1311) );
  NAND21X1 U862 ( .B(n3396), .A(A[198]), .Y(n620) );
  NAND21X1 U866 ( .B(n3421), .A(n623), .Y(n1310) );
  NAND21X1 U869 ( .B(n3396), .A(A[197]), .Y(n623) );
  NAND21X1 U873 ( .B(n3421), .A(n626), .Y(n1309) );
  NAND21X1 U876 ( .B(n3395), .A(A[196]), .Y(n626) );
  NAND21X1 U880 ( .B(n3422), .A(n629), .Y(n1308) );
  NAND21X1 U883 ( .B(n3396), .A(A[195]), .Y(n629) );
  NAND21X1 U887 ( .B(n3422), .A(n632), .Y(n1307) );
  NAND21X1 U890 ( .B(n3395), .A(A[194]), .Y(n632) );
  NAND21X1 U894 ( .B(n3422), .A(n635), .Y(n1306) );
  NAND21X1 U901 ( .B(n3422), .A(n638), .Y(n1305) );
  NAND21X1 U956 ( .B(n3423), .A(n3414), .Y(n1296) );
  NAND21X1 U1052 ( .B(n3424), .A(n689), .Y(n1280) );
  NOR2X1 U1054 ( .A(n3410), .B(A[167]), .Y(n689) );
  NAND21X1 U1058 ( .B(n3424), .A(n691), .Y(n1279) );
  NOR2X1 U1060 ( .A(n3411), .B(A[166]), .Y(n691) );
  NAND21X1 U1064 ( .B(n3425), .A(n693), .Y(n1278) );
  NOR2X1 U1066 ( .A(n3411), .B(A[165]), .Y(n693) );
  NAND21X1 U1070 ( .B(n3425), .A(n695), .Y(n1277) );
  NOR2X1 U1072 ( .A(n3411), .B(A[164]), .Y(n695) );
  NAND21X1 U1076 ( .B(n3425), .A(n697), .Y(n1276) );
  NOR2X1 U1078 ( .A(n3411), .B(A[163]), .Y(n697) );
  NAND21X1 U1082 ( .B(n3425), .A(n699), .Y(n1275) );
  NOR2X1 U1084 ( .A(n3411), .B(A[162]), .Y(n699) );
  NAND21X1 U1088 ( .B(n3425), .A(n701), .Y(n1274) );
  NOR2X1 U1090 ( .A(n3411), .B(A[161]), .Y(n701) );
  NAND21X1 U1094 ( .B(n3425), .A(n703), .Y(n1273) );
  NOR2X1 U1096 ( .A(n3411), .B(A[160]), .Y(n703) );
  NAND21X1 U1100 ( .B(n3425), .A(n705), .Y(n1272) );
  NOR2X1 U1102 ( .A(n3411), .B(A[159]), .Y(n705) );
  NAND21X1 U1106 ( .B(n3425), .A(n707), .Y(n1271) );
  NOR2X1 U1108 ( .A(n3411), .B(A[158]), .Y(n707) );
  NAND21X1 U1112 ( .B(n3425), .A(n709), .Y(n1270) );
  NOR2X1 U1114 ( .A(n3411), .B(A[157]), .Y(n709) );
  NAND21X1 U1118 ( .B(n3425), .A(n711), .Y(n1269) );
  NOR2X1 U1120 ( .A(n3392), .B(A[156]), .Y(n711) );
  NAND21X1 U1124 ( .B(n3426), .A(n713), .Y(n1268) );
  NOR2X1 U1126 ( .A(n3392), .B(A[155]), .Y(n713) );
  NAND21X1 U1130 ( .B(n3426), .A(n715), .Y(n1267) );
  NOR2X1 U1132 ( .A(n3394), .B(A[154]), .Y(n715) );
  NAND21X1 U1136 ( .B(n3426), .A(n717), .Y(n1266) );
  NOR2X1 U1138 ( .A(n3394), .B(A[153]), .Y(n717) );
  NAND21X1 U1142 ( .B(n3426), .A(n719), .Y(n1265) );
  NOR2X1 U1144 ( .A(n3400), .B(A[152]), .Y(n719) );
  NAND21X1 U1148 ( .B(n3426), .A(n721), .Y(n1264) );
  NAND21X1 U1155 ( .B(n3426), .A(n724), .Y(n1263) );
  NAND21X1 U1162 ( .B(n3426), .A(n727), .Y(n1262) );
  NAND21X1 U1169 ( .B(n3426), .A(n730), .Y(n1261) );
  NAND21X1 U1176 ( .B(n3426), .A(n733), .Y(n1260) );
  NAND21X1 U1183 ( .B(n3426), .A(n736), .Y(n1259) );
  NAND21X1 U1190 ( .B(n3427), .A(n739), .Y(n1258) );
  NAND21X1 U1197 ( .B(n3427), .A(n742), .Y(n1257) );
  NAND21X1 U1204 ( .B(n3427), .A(n745), .Y(n1256) );
  NAND21X1 U1211 ( .B(n3427), .A(n748), .Y(n1255) );
  NAND21X1 U1218 ( .B(n3427), .A(n751), .Y(n1254) );
  NAND21X1 U1225 ( .B(n3427), .A(n754), .Y(n1253) );
  NAND21X1 U1232 ( .B(n3427), .A(n757), .Y(n1252) );
  NAND21X1 U1239 ( .B(n3427), .A(n760), .Y(n1251) );
  NAND21X1 U1246 ( .B(n3427), .A(n763), .Y(n1250) );
  NAND21X1 U1253 ( .B(n3427), .A(n766), .Y(n1249) );
  NAND21X1 U1260 ( .B(n3428), .A(n769), .Y(n1248) );
  NAND21X1 U1267 ( .B(n3428), .A(n772), .Y(n1247) );
  NAND21X1 U1274 ( .B(n3428), .A(n775), .Y(n1246) );
  NAND21X1 U1281 ( .B(n3428), .A(n778), .Y(n1245) );
  NAND21X1 U1288 ( .B(n3428), .A(n781), .Y(n1244) );
  NAND21X1 U1295 ( .B(n3428), .A(n784), .Y(n1243) );
  NAND21X1 U1302 ( .B(n3428), .A(n787), .Y(n1242) );
  NAND21X1 U1309 ( .B(n3428), .A(n790), .Y(n1241) );
  NAND21X1 U1323 ( .B(n3428), .A(n796), .Y(n1239) );
  NAND21X1 U1330 ( .B(n3429), .A(n799), .Y(n1238) );
  NAND21X1 U1337 ( .B(n3429), .A(n802), .Y(n1237) );
  NAND21X1 U1344 ( .B(n3429), .A(n805), .Y(n1236) );
  NAND21X1 U1351 ( .B(n3429), .A(n808), .Y(n1235) );
  NAND21X1 U1358 ( .B(n3429), .A(n811), .Y(n1234) );
  NAND21X1 U1365 ( .B(n3429), .A(n814), .Y(n1233) );
  NAND21X1 U1372 ( .B(n3429), .A(n817), .Y(n1232) );
  NAND21X1 U1379 ( .B(n3429), .A(n820), .Y(n1231) );
  NOR21X1 U1382 ( .B(n3400), .A(A[374]), .Y(n820) );
  NAND21X1 U1386 ( .B(n3429), .A(n823), .Y(n1230) );
  NAND21X1 U1393 ( .B(n3429), .A(n826), .Y(n1229) );
  NAND21X1 U1400 ( .B(n3430), .A(n829), .Y(n1228) );
  NAND21X1 U1407 ( .B(n3430), .A(n832), .Y(n1227) );
  NAND21X1 U1414 ( .B(n3430), .A(n835), .Y(n1226) );
  NAND21X1 U1421 ( .B(n3430), .A(n838), .Y(n1225) );
  NAND21X1 U1428 ( .B(n3430), .A(n841), .Y(n1224) );
  NAND21X1 U1435 ( .B(n3430), .A(n844), .Y(n1223) );
  NAND21X1 U1442 ( .B(n3430), .A(n847), .Y(n1222) );
  NAND21X1 U1449 ( .B(n3430), .A(n850), .Y(n1221) );
  NAND21X1 U1456 ( .B(n3430), .A(n853), .Y(n1220) );
  NAND21X1 U1463 ( .B(n3430), .A(n856), .Y(n1219) );
  NAND21X1 U1470 ( .B(n3431), .A(n859), .Y(n1218) );
  NAND21X1 U1477 ( .B(n3431), .A(n862), .Y(n1217) );
  NAND21X1 U1484 ( .B(n3431), .A(n865), .Y(n1216) );
  NAND21X1 U1491 ( .B(n3431), .A(n868), .Y(n1215) );
  NAND21X1 U1498 ( .B(n3431), .A(n871), .Y(n1214) );
  NAND21X1 U1505 ( .B(n3431), .A(n874), .Y(n1213) );
  NOR21X1 U1508 ( .B(n3400), .A(A[356]), .Y(n874) );
  NAND21X1 U1512 ( .B(n3431), .A(n877), .Y(n1212) );
  NOR21X1 U1515 ( .B(n3397), .A(A[355]), .Y(n877) );
  NAND21X1 U1519 ( .B(n3431), .A(n880), .Y(n1211) );
  NAND21X1 U1526 ( .B(n3431), .A(n883), .Y(n1210) );
  NAND21X1 U1533 ( .B(n3431), .A(n886), .Y(n1209) );
  NAND21X1 U1540 ( .B(n3432), .A(n889), .Y(n1208) );
  NOR21X1 U1543 ( .B(n3399), .A(A[351]), .Y(n889) );
  NAND21X1 U1547 ( .B(n3432), .A(n892), .Y(n1207) );
  NAND21X1 U1554 ( .B(n3432), .A(n895), .Y(n1206) );
  NAND21X1 U1561 ( .B(n3432), .A(n898), .Y(n1205) );
  NAND21X1 U1568 ( .B(n3432), .A(n901), .Y(n1204) );
  NOR21X1 U1571 ( .B(n3399), .A(A[347]), .Y(n901) );
  NAND21X1 U1575 ( .B(n3432), .A(n904), .Y(n1203) );
  NAND21X1 U1582 ( .B(n3432), .A(n907), .Y(n1202) );
  NAND21X1 U1589 ( .B(n3432), .A(n910), .Y(n1201) );
  NAND21X1 U1596 ( .B(n3432), .A(n913), .Y(n1200) );
  NAND21X1 U1603 ( .B(n3432), .A(n916), .Y(n1199) );
  NAND21X1 U1610 ( .B(n3433), .A(n919), .Y(n1198) );
  NAND21X1 U1617 ( .B(n3433), .A(n922), .Y(n1197) );
  NAND21X1 U1624 ( .B(n3433), .A(n925), .Y(n1196) );
  NAND21X1 U1631 ( .B(n3433), .A(n928), .Y(n1195) );
  NAND21X1 U1638 ( .B(n3433), .A(n931), .Y(n1194) );
  NAND21X1 U1645 ( .B(n3433), .A(n934), .Y(n1193) );
  NAND21X1 U1652 ( .B(n3433), .A(n937), .Y(n1192) );
  NAND21X1 U1659 ( .B(n3433), .A(n940), .Y(n1191) );
  NAND21X1 U1666 ( .B(n3433), .A(n943), .Y(n1190) );
  NAND21X1 U1673 ( .B(n3433), .A(n946), .Y(n1189) );
  NAND21X1 U1680 ( .B(n3434), .A(n949), .Y(n1188) );
  NAND21X1 U1687 ( .B(n3434), .A(n952), .Y(n1187) );
  NAND21X1 U1694 ( .B(n3434), .A(n955), .Y(n1186) );
  NAND21X1 U1701 ( .B(n3434), .A(n958), .Y(n1185) );
  NAND21X1 U1708 ( .B(n3434), .A(n961), .Y(n1184) );
  NAND21X1 U1715 ( .B(n3434), .A(n964), .Y(n1183) );
  NAND21X1 U1722 ( .B(n3434), .A(n967), .Y(n1182) );
  NAND21X1 U1729 ( .B(n3434), .A(n970), .Y(n1181) );
  NAND21X1 U1736 ( .B(n3434), .A(n973), .Y(n1180) );
  NAND21X1 U1743 ( .B(n3434), .A(n976), .Y(n1179) );
  NAND21X1 U1750 ( .B(n3435), .A(n979), .Y(n1178) );
  NAND21X1 U1757 ( .B(n3435), .A(n982), .Y(n1177) );
  NAND21X1 U1908 ( .B(n3437), .A(n1033), .Y(n1152) );
  NOR2X1 U1910 ( .A(n3403), .B(A[39]), .Y(n1033) );
  NAND21X1 U1914 ( .B(n3437), .A(n1035), .Y(n1151) );
  NOR2X1 U1916 ( .A(n3403), .B(A[38]), .Y(n1035) );
  NAND21X1 U1920 ( .B(n3437), .A(n1037), .Y(n1150) );
  NOR2X1 U1922 ( .A(n3403), .B(A[37]), .Y(n1037) );
  NAND21X1 U1926 ( .B(n3437), .A(n1039), .Y(n1149) );
  NOR2X1 U1928 ( .A(n3403), .B(A[36]), .Y(n1039) );
  NAND21X1 U1932 ( .B(n3438), .A(n1041), .Y(n1148) );
  NOR2X1 U1934 ( .A(n3403), .B(A[35]), .Y(n1041) );
  NAND21X1 U1938 ( .B(n3438), .A(n1043), .Y(n1147) );
  NOR2X1 U1940 ( .A(n3403), .B(A[34]), .Y(n1043) );
  NAND21X1 U1944 ( .B(n3438), .A(n1045), .Y(n1146) );
  NOR2X1 U1946 ( .A(n3403), .B(A[33]), .Y(n1045) );
  NAND21X1 U1950 ( .B(n3438), .A(n1047), .Y(n1145) );
  NOR2X1 U1952 ( .A(n3403), .B(A[32]), .Y(n1047) );
  NAND21X1 U1988 ( .B(n3438), .A(n1057), .Y(n1144) );
  NOR2X1 U1990 ( .A(n3403), .B(A[23]), .Y(n1057) );
  NAND21X1 U1994 ( .B(n3438), .A(n1059), .Y(n1143) );
  NOR2X1 U1996 ( .A(n3403), .B(A[22]), .Y(n1059) );
  NAND21X1 U2000 ( .B(n3438), .A(n1061), .Y(n1142) );
  NOR2X1 U2002 ( .A(n3402), .B(A[21]), .Y(n1061) );
  NAND21X1 U2006 ( .B(n3438), .A(n1063), .Y(n1141) );
  NOR2X1 U2008 ( .A(n3402), .B(A[20]), .Y(n1063) );
  NAND21X1 U2012 ( .B(n3438), .A(n1065), .Y(n1140) );
  NOR2X1 U2014 ( .A(n3402), .B(A[19]), .Y(n1065) );
  NAND21X1 U2018 ( .B(n3438), .A(n1067), .Y(n1139) );
  NOR2X1 U2020 ( .A(n3402), .B(A[18]), .Y(n1067) );
  NAND21X1 U2024 ( .B(n3439), .A(n1069), .Y(n1138) );
  NOR2X1 U2026 ( .A(n3402), .B(A[17]), .Y(n1069) );
  NAND21X1 U2030 ( .B(n3439), .A(n1071), .Y(n1137) );
  NOR2X1 U2032 ( .A(n3402), .B(A[16]), .Y(n1071) );
  NAND21X1 U2036 ( .B(n3439), .A(n1073), .Y(n1136) );
  NAND21X1 U2043 ( .B(n3439), .A(n1076), .Y(n1135) );
  NAND21X1 U2050 ( .B(n3439), .A(n1079), .Y(n1134) );
  NAND21X1 U2057 ( .B(n3439), .A(n1082), .Y(n1133) );
  NAND21X1 U2064 ( .B(n3439), .A(n1085), .Y(n1132) );
  NAND21X1 U2071 ( .B(n3439), .A(n1088), .Y(n1131) );
  NAND21X1 U2078 ( .B(n3439), .A(n1091), .Y(n1130) );
  NAND21X1 U2085 ( .B(n3439), .A(n1094), .Y(n1129) );
  NAND21X1 U2099 ( .B(n3440), .A(n1100), .Y(n1127) );
  NAND21X1 U2106 ( .B(n3440), .A(n1103), .Y(n1126) );
  NAND21X1 U2113 ( .B(n3440), .A(n1106), .Y(n1125) );
  NAND21X1 U2120 ( .B(n3440), .A(n1109), .Y(n1124) );
  NAND21X1 U2127 ( .B(n3440), .A(n1112), .Y(n1123) );
  NAND21X1 U2134 ( .B(n3440), .A(n1115), .Y(n1122) );
  NAND21X1 U2141 ( .B(n3440), .A(n1118), .Y(n1121) );
  MUX2IX4 U2149 ( .D0(n96), .D1(n64), .S(n3375), .Y(n32) );
  MUX2IX2 U2150 ( .D0(n3201), .D1(n228), .S(n3374), .Y(n100) );
  MUX2BX2 U2151 ( .D0(n3186), .D1(n156), .S(n3372), .Y(n60) );
  MUX2IX1 U2152 ( .D0(n1132), .D1(n1252), .S(n3385), .Y(n3186) );
  MUX2IX1 U2153 ( .D0(n3196), .D1(n100), .S(n3226), .Y(n36) );
  MUX2IX4 U2154 ( .D0(n313), .D1(n441), .S(n3381), .Y(n193) );
  INVX2 U2155 ( .A(n1193), .Y(n313) );
  MUX2X2 U2156 ( .D0(n1124), .D1(n1244), .S(n3380), .Y(n116) );
  MUX2IX2 U2157 ( .D0(n116), .D1(n148), .S(n3230), .Y(n52) );
  MUX2IX2 U2158 ( .D0(n1136), .D1(n128), .S(n3237), .Y(n64) );
  MUX2IX2 U2159 ( .D0(n112), .D1(n3229), .S(n3242), .Y(n48) );
  MUX2IX4 U2160 ( .D0(n3235), .D1(n88), .S(n3240), .Y(n24) );
  MUX2IX2 U2161 ( .D0(n29), .D1(n45), .S(n3368), .Y(n13) );
  MUX2IX2 U2162 ( .D0(A[263]), .D1(A[7]), .S(n3414), .Y(n1097) );
  MUX2IX4 U2163 ( .D0(n69), .D1(n101), .S(n3374), .Y(n37) );
  MUX2IX4 U2164 ( .D0(n197), .D1(n229), .S(SH[5]), .Y(n101) );
  NOR21XL U2165 ( .B(n3400), .A(A[336]), .Y(n934) );
  INVX1 U2166 ( .A(n3210), .Y(n3187) );
  NOR21XL U2167 ( .B(n3398), .A(A[338]), .Y(n928) );
  NOR21XL U2168 ( .B(n3399), .A(A[337]), .Y(n931) );
  INVX1 U2169 ( .A(n3387), .Y(n3210) );
  MUX2IX2 U2170 ( .D0(n1), .D1(n9), .S(SH[3]), .Y(B[0]) );
  MUX2IX1 U2171 ( .D0(n25), .D1(n41), .S(n3368), .Y(n9) );
  MUX2IX1 U2172 ( .D0(n17), .D1(n33), .S(n3368), .Y(n1) );
  MUX2IX1 U2173 ( .D0(n3191), .D1(n105), .S(n3232), .Y(n41) );
  MUX2IX2 U2174 ( .D0(n198), .D1(n230), .S(SH[5]), .Y(n102) );
  MUX2IX1 U2175 ( .D0(n31), .D1(n47), .S(n3368), .Y(n15) );
  MUX2IX1 U2176 ( .D0(n3195), .D1(n111), .S(n3236), .Y(n47) );
  NOR21XL U2177 ( .B(n3400), .A(A[368]), .Y(n838) );
  NOR21XL U2178 ( .B(n3398), .A(A[360]), .Y(n862) );
  NOR21XL U2179 ( .B(n3398), .A(A[366]), .Y(n844) );
  NOR21XL U2180 ( .B(n3397), .A(A[346]), .Y(n904) );
  NOR21XL U2181 ( .B(n3397), .A(A[345]), .Y(n907) );
  NOR21XL U2182 ( .B(n3396), .A(A[344]), .Y(n910) );
  NOR21XL U2183 ( .B(n3397), .A(A[352]), .Y(n886) );
  NOR21XL U2184 ( .B(n3397), .A(A[348]), .Y(n898) );
  NOR21XL U2185 ( .B(n3399), .A(A[359]), .Y(n865) );
  NOR21XL U2186 ( .B(n3398), .A(A[367]), .Y(n841) );
  NOR21XL U2187 ( .B(n3397), .A(A[341]), .Y(n919) );
  NOR21XL U2188 ( .B(n3397), .A(A[357]), .Y(n871) );
  NOR21XL U2189 ( .B(n3399), .A(A[350]), .Y(n892) );
  INVX1 U2190 ( .A(n1199), .Y(n319) );
  NOR21XL U2191 ( .B(n3399), .A(A[342]), .Y(n916) );
  MUX2IX1 U2192 ( .D0(n247), .D1(n367), .S(n3210), .Y(n119) );
  NOR21XL U2193 ( .B(n3399), .A(A[362]), .Y(n856) );
  NOR21XL U2194 ( .B(n3397), .A(A[354]), .Y(n880) );
  INVX1 U2195 ( .A(n3190), .Y(n212) );
  NAND2X1 U2196 ( .A(n3279), .B(n3210), .Y(n3189) );
  NOR21XL U2197 ( .B(n3399), .A(A[353]), .Y(n883) );
  MUX2X1 U2198 ( .D0(n1122), .D1(n1242), .S(n3379), .Y(n114) );
  MUX2X1 U2199 ( .D0(n1178), .D1(n1306), .S(n3379), .Y(n178) );
  INVX1 U2200 ( .A(n1200), .Y(n320) );
  NOR21XL U2201 ( .B(n3396), .A(A[343]), .Y(n913) );
  MUX2IX1 U2202 ( .D0(n480), .D1(n72), .S(n3375), .Y(n232) );
  NOR21XL U2203 ( .B(n3397), .A(A[349]), .Y(n895) );
  NOR21XL U2204 ( .B(n3400), .A(A[365]), .Y(n847) );
  MUX2IX1 U2205 ( .D0(n95), .D1(n63), .S(n3233), .Y(n31) );
  MUX2IX1 U2206 ( .D0(n1135), .D1(n127), .S(n3225), .Y(n63) );
  MUX2IX1 U2207 ( .D0(n191), .D1(n223), .S(n3369), .Y(n95) );
  MUX2IX1 U2208 ( .D0(n3199), .D1(n375), .S(n3238), .Y(n127) );
  MUX2IX1 U2209 ( .D0(n195), .D1(n227), .S(SH[5]), .Y(n99) );
  MUX2IX1 U2210 ( .D0(n75), .D1(n107), .S(n3212), .Y(n43) );
  MUX2X1 U2211 ( .D0(n1188), .D1(n1316), .S(n3380), .Y(n188) );
  MUX2IX1 U2212 ( .D0(n3192), .D1(n108), .S(n3234), .Y(n44) );
  MUX2IX1 U2213 ( .D0(n194), .D1(n226), .S(SH[5]), .Y(n98) );
  MUX2X1 U2214 ( .D0(n1226), .D1(n1354), .S(n3210), .Y(n226) );
  MUX2X1 U2215 ( .D0(n1194), .D1(n1322), .S(n3381), .Y(n194) );
  MUX2IX1 U2216 ( .D0(n74), .D1(n106), .S(n3213), .Y(n42) );
  MUX2X1 U2217 ( .D0(n1186), .D1(n1314), .S(n3380), .Y(n186) );
  MUX2IX1 U2218 ( .D0(n181), .D1(n213), .S(n3372), .Y(n85) );
  MUX2X1 U2219 ( .D0(n1181), .D1(n1309), .S(n3380), .Y(n181) );
  MUX2X1 U2220 ( .D0(n1125), .D1(n1245), .S(n3210), .Y(n117) );
  MUX2X1 U2221 ( .D0(n1221), .D1(n1349), .S(n3383), .Y(n221) );
  MUX2IX1 U2222 ( .D0(n77), .D1(n109), .S(n3212), .Y(n45) );
  MUX2IX1 U2223 ( .D0(n1208), .D1(n1336), .S(n3382), .Y(n3229) );
  MUX2IX1 U2224 ( .D0(n240), .D1(n3197), .S(n3214), .Y(n112) );
  MUX2IX1 U2225 ( .D0(n1184), .D1(n1312), .S(n3210), .Y(n3235) );
  MUX2IX1 U2226 ( .D0(n3200), .D1(n376), .S(n3238), .Y(n128) );
  INVX1 U2227 ( .A(n3367), .Y(n3224) );
  MUX2IX1 U2228 ( .D0(n3), .D1(n11), .S(SH[3]), .Y(B[2]) );
  MUX2IX1 U2229 ( .D0(n19), .D1(n35), .S(n3368), .Y(n3) );
  MUX2IX1 U2230 ( .D0(n27), .D1(n43), .S(n3368), .Y(n11) );
  MUX2IX1 U2231 ( .D0(n67), .D1(n99), .S(n3374), .Y(n35) );
  MUX2IX2 U2232 ( .D0(n2), .D1(n10), .S(SH[3]), .Y(B[1]) );
  MUX2IX1 U2233 ( .D0(n18), .D1(n34), .S(n3367), .Y(n2) );
  MUX2IX2 U2234 ( .D0(n26), .D1(n42), .S(n3367), .Y(n10) );
  MUX2IX1 U2235 ( .D0(n66), .D1(n98), .S(n3374), .Y(n34) );
  MUX2IX2 U2236 ( .D0(n6), .D1(n14), .S(SH[3]), .Y(B[5]) );
  MUX2IX1 U2237 ( .D0(n30), .D1(n46), .S(n3367), .Y(n14) );
  MUX2IX1 U2238 ( .D0(n3193), .D1(n110), .S(n3220), .Y(n46) );
  MUX2IX1 U2239 ( .D0(n15), .D1(n7), .S(n3231), .Y(B[6]) );
  MUX2IX2 U2240 ( .D0(n39), .D1(n23), .S(n3224), .Y(n7) );
  MUX2IX4 U2241 ( .D0(n103), .D1(n3194), .S(n3222), .Y(n39) );
  INVX2 U2242 ( .A(n1231), .Y(n351) );
  NAND2X1 U2243 ( .A(n332), .B(n3187), .Y(n3188) );
  NAND2X1 U2244 ( .A(n3188), .B(n3189), .Y(n3190) );
  INVX1 U2245 ( .A(n1212), .Y(n332) );
  INVX2 U2246 ( .A(n1192), .Y(n312) );
  MUX2IX4 U2247 ( .D0(n119), .D1(n151), .S(n3372), .Y(n55) );
  MUX2IX4 U2248 ( .D0(n431), .D1(n303), .S(n3227), .Y(n183) );
  INVX2 U2249 ( .A(n1183), .Y(n303) );
  NAND2X2 U2250 ( .A(n183), .B(n3238), .Y(n3215) );
  MUX2IX4 U2251 ( .D0(n55), .D1(n87), .S(n3212), .Y(n23) );
  INVX1 U2252 ( .A(n3372), .Y(n3241) );
  INVX1 U2253 ( .A(n3371), .Y(n3238) );
  INVX1 U2254 ( .A(n3393), .Y(n3221) );
  INVX1 U2255 ( .A(n3374), .Y(n3233) );
  MUX2X1 U2256 ( .D0(n321), .D1(n449), .S(n3382), .Y(n3191) );
  MUX2X1 U2257 ( .D0(n324), .D1(n452), .S(n3382), .Y(n3192) );
  MUX2X1 U2258 ( .D0(n326), .D1(n454), .S(n3382), .Y(n3193) );
  MUX2X1 U2259 ( .D0(n447), .D1(n319), .S(n3227), .Y(n3194) );
  MUX2X1 U2260 ( .D0(n327), .D1(n455), .S(n3382), .Y(n3195) );
  MUX2IX1 U2261 ( .D0(n1196), .D1(n1324), .S(n3381), .Y(n3196) );
  OR2X1 U2262 ( .A(n3428), .B(n3246), .Y(n3197) );
  MUX2X2 U2263 ( .D0(n320), .D1(n448), .S(n3382), .Y(n3198) );
  MUX2X1 U2264 ( .D0(n3295), .D1(n416), .S(n3377), .Y(n3199) );
  MUX2X1 U2265 ( .D0(n3299), .D1(n3244), .S(n3377), .Y(n3200) );
  MUX2X1 U2266 ( .D0(n132), .D1(n164), .S(n3371), .Y(n3201) );
  MUX2X1 U2267 ( .D0(n135), .D1(n167), .S(n3371), .Y(n3202) );
  MUX2IX1 U2268 ( .D0(n1152), .D1(n1280), .S(n3377), .Y(n3203) );
  MUX2X1 U2269 ( .D0(n3275), .D1(n3257), .S(n3377), .Y(n3204) );
  MUX2X1 U2270 ( .D0(n143), .D1(n175), .S(n3370), .Y(n3205) );
  MUX2X1 U2271 ( .D0(n137), .D1(n169), .S(n3370), .Y(n3206) );
  MUX2X1 U2272 ( .D0(n142), .D1(n174), .S(n3370), .Y(n3207) );
  MUX2X1 U2273 ( .D0(n140), .D1(n172), .S(n3370), .Y(n3208) );
  MUX2IX1 U2274 ( .D0(n1150), .D1(n1278), .S(n3376), .Y(n3209) );
  INVX1 U2275 ( .A(n3381), .Y(n3227) );
  INVX1 U2276 ( .A(SH[3]), .Y(n3231) );
  INVXL U2277 ( .A(n3387), .Y(n3211) );
  INVXL U2278 ( .A(n3375), .Y(n3212) );
  INVXL U2279 ( .A(n3375), .Y(n3213) );
  NOR2X1 U2280 ( .A(n3375), .B(n3210), .Y(n3214) );
  NOR21XL U2281 ( .B(n3399), .A(A[375]), .Y(n817) );
  MUX2IX1 U2282 ( .D0(A[335]), .D1(A[79]), .S(n3415), .Y(n937) );
  NAND2X1 U2283 ( .A(n215), .B(n3230), .Y(n3216) );
  NAND2X2 U2284 ( .A(n3215), .B(n3216), .Y(n3217) );
  INVX2 U2285 ( .A(n3217), .Y(n87) );
  INVX1 U2286 ( .A(n3238), .Y(n3230) );
  NOR21XL U2287 ( .B(n3400), .A(A[358]), .Y(n868) );
  MUX2IX4 U2288 ( .D0(n351), .D1(n479), .S(n3384), .Y(n231) );
  MUX2IX4 U2289 ( .D0(n3339), .D1(n336), .S(n3387), .Y(n3243) );
  MUX2IX4 U2290 ( .D0(n104), .D1(n3198), .S(n3218), .Y(n40) );
  NOR2X4 U2291 ( .A(n3233), .B(n3369), .Y(n3218) );
  MUX2IX4 U2292 ( .D0(n92), .D1(n60), .S(n3233), .Y(n28) );
  MUX2IX1 U2293 ( .D0(n94), .D1(n62), .S(n3233), .Y(n30) );
  NOR2X1 U2294 ( .A(n3375), .B(n3384), .Y(n3219) );
  NAND2X1 U2295 ( .A(n3213), .B(n3241), .Y(n3220) );
  MUX2IX1 U2296 ( .D0(A[267]), .D1(A[11]), .S(n3221), .Y(n1085) );
  MUX2IX4 U2297 ( .D0(n440), .D1(n312), .S(n3387), .Y(n192) );
  NOR2X1 U2298 ( .A(n3233), .B(n3369), .Y(n3222) );
  MUX2IX4 U2299 ( .D0(n1128), .D1(n120), .S(n3237), .Y(n56) );
  MUX2IX1 U2300 ( .D0(n93), .D1(n61), .S(n3233), .Y(n29) );
  NAND2X1 U2301 ( .A(n3241), .B(n3227), .Y(n3223) );
  MUX2IX4 U2302 ( .D0(n40), .D1(n24), .S(n3224), .Y(n8) );
  MUX2IX1 U2303 ( .D0(n1129), .D1(n121), .S(n3223), .Y(n57) );
  NAND2X1 U2304 ( .A(n3238), .B(n3227), .Y(n3225) );
  NAND2X1 U2305 ( .A(n3374), .B(n3241), .Y(n3226) );
  MUX2IX1 U2306 ( .D0(A[264]), .D1(A[8]), .S(n3221), .Y(n1094) );
  NAND2X1 U2307 ( .A(n3241), .B(n3386), .Y(n3228) );
  MUX2IX1 U2308 ( .D0(A[270]), .D1(A[14]), .S(n3221), .Y(n1076) );
  MUX2IX1 U2309 ( .D0(n1126), .D1(n118), .S(n3228), .Y(n54) );
  NOR21XL U2310 ( .B(n3398), .A(A[370]), .Y(n832) );
  NOR21XL U2311 ( .B(n3398), .A(A[369]), .Y(n835) );
  NOR21XL U2312 ( .B(n3399), .A(A[373]), .Y(n823) );
  MUX2IX1 U2313 ( .D0(n209), .D1(n177), .S(n3238), .Y(n81) );
  MUX2IX1 U2314 ( .D0(n425), .D1(n297), .S(n3227), .Y(n177) );
  MUX2IX4 U2315 ( .D0(n52), .D1(n84), .S(n3212), .Y(n20) );
  MUX2IX2 U2316 ( .D0(n180), .D1(n212), .S(n3369), .Y(n84) );
  MUX2IX1 U2317 ( .D0(A[320]), .D1(A[64]), .S(n3221), .Y(n982) );
  NAND2X1 U2318 ( .A(n3213), .B(n3238), .Y(n3232) );
  MUX2IX1 U2319 ( .D0(A[261]), .D1(A[5]), .S(n3221), .Y(n1103) );
  NAND2X1 U2320 ( .A(n3212), .B(n3241), .Y(n3234) );
  MUX2IX1 U2321 ( .D0(A[326]), .D1(A[70]), .S(n3221), .Y(n964) );
  MUX2IX4 U2322 ( .D0(n192), .D1(n224), .S(n3369), .Y(n96) );
  MUX2X2 U2323 ( .D0(n1224), .D1(n1352), .S(n3383), .Y(n224) );
  MUX2IX1 U2324 ( .D0(n86), .D1(n54), .S(n3375), .Y(n22) );
  MUX2IX2 U2325 ( .D0(n22), .D1(n38), .S(n3367), .Y(n6) );
  NAND2X1 U2326 ( .A(n3213), .B(n3241), .Y(n3236) );
  INVX2 U2327 ( .A(n1216), .Y(n336) );
  NAND2X1 U2328 ( .A(n3238), .B(n3386), .Y(n3237) );
  INVX4 U2329 ( .A(n56), .Y(n3239) );
  NAND21X2 U2330 ( .B(n3440), .A(n1097), .Y(n1128) );
  MUX2IX1 U2331 ( .D0(A[271]), .D1(A[15]), .S(n3416), .Y(n1073) );
  NAND2X1 U2332 ( .A(n3213), .B(n3238), .Y(n3240) );
  MUX2IX4 U2333 ( .D0(n16), .D1(n8), .S(n3231), .Y(B[7]) );
  NOR2X1 U2334 ( .A(n3375), .B(n3369), .Y(n3242) );
  MUX2IX4 U2335 ( .D0(n3239), .D1(n3243), .S(n3212), .Y(n88) );
  MUX2IX1 U2336 ( .D0(A[327]), .D1(A[71]), .S(n3221), .Y(n961) );
  INVXL U2337 ( .A(n1218), .Y(n338) );
  INVX1 U2338 ( .A(n1213), .Y(n333) );
  MUX2IX2 U2339 ( .D0(n53), .D1(n85), .S(SH[6]), .Y(n21) );
  INVXL U2340 ( .A(n1237), .Y(n357) );
  MUX2IX1 U2341 ( .D0(n58), .D1(n90), .S(n3213), .Y(n26) );
  INVX1 U2342 ( .A(n1204), .Y(n324) );
  INVX1 U2343 ( .A(n1205), .Y(n325) );
  INVX1 U2344 ( .A(n1210), .Y(n330) );
  MUX2X1 U2345 ( .D0(A[127]), .D1(A[383]), .S(n3388), .Y(n3246) );
  INVX1 U2346 ( .A(n1236), .Y(n356) );
  MUX2X2 U2347 ( .D0(n1197), .D1(n1325), .S(n3381), .Y(n197) );
  MUX2X2 U2348 ( .D0(n1228), .D1(n1356), .S(n3384), .Y(n228) );
  MUX2X2 U2349 ( .D0(n1189), .D1(n1317), .S(n3380), .Y(n189) );
  MUX2X2 U2350 ( .D0(n1130), .D1(n1250), .S(n3383), .Y(n122) );
  MUX2X2 U2351 ( .D0(n1220), .D1(n1348), .S(n3383), .Y(n220) );
  MUX2X2 U2352 ( .D0(n1133), .D1(n1253), .S(SH[7]), .Y(n125) );
  MUX2X2 U2353 ( .D0(n1180), .D1(n1308), .S(n3379), .Y(n180) );
  NOR21XL U2354 ( .B(n3397), .A(A[340]), .Y(n922) );
  NOR21XL U2355 ( .B(n3398), .A(A[339]), .Y(n925) );
  NOR21XL U2356 ( .B(n3398), .A(A[363]), .Y(n853) );
  NOR21XL U2357 ( .B(n3398), .A(A[361]), .Y(n859) );
  NOR21XL U2358 ( .B(n3400), .A(A[372]), .Y(n826) );
  NOR21XL U2359 ( .B(n3400), .A(A[371]), .Y(n829) );
  NOR21XL U2360 ( .B(n3398), .A(A[364]), .Y(n850) );
  MUX2X2 U2361 ( .D0(n1229), .D1(n1357), .S(n3383), .Y(n229) );
  INVX1 U2362 ( .A(n3413), .Y(n3392) );
  INVX1 U2363 ( .A(n3412), .Y(n3389) );
  INVX1 U2364 ( .A(n3412), .Y(n3390) );
  INVX1 U2365 ( .A(n3413), .Y(n3393) );
  INVX1 U2366 ( .A(n3414), .Y(n3394) );
  INVX1 U2367 ( .A(n3412), .Y(n3388) );
  INVX1 U2368 ( .A(n3414), .Y(n3395) );
  INVX1 U2369 ( .A(n3414), .Y(n3396) );
  INVX1 U2370 ( .A(n3415), .Y(n3398) );
  INVX1 U2371 ( .A(n3415), .Y(n3399) );
  INVX1 U2372 ( .A(n3413), .Y(n3391) );
  INVX1 U2373 ( .A(n3415), .Y(n3397) );
  INVX1 U2374 ( .A(n3416), .Y(n3400) );
  INVX1 U2375 ( .A(n3414), .Y(n3407) );
  INVX1 U2376 ( .A(n3414), .Y(n3404) );
  INVX1 U2377 ( .A(n3416), .Y(n3402) );
  INVX1 U2378 ( .A(n3413), .Y(n3410) );
  INVX1 U2379 ( .A(n3415), .Y(n3409) );
  INVX1 U2380 ( .A(n3416), .Y(n3401) );
  INVX1 U2381 ( .A(n3413), .Y(n3403) );
  INVX1 U2382 ( .A(n3413), .Y(n3405) );
  INVX1 U2383 ( .A(n3416), .Y(n3408) );
  INVX1 U2384 ( .A(n3415), .Y(n3406) );
  INVX1 U2385 ( .A(n3413), .Y(n3411) );
  INVX1 U2386 ( .A(SH[8]), .Y(n3412) );
  INVX1 U2387 ( .A(SH[8]), .Y(n3413) );
  INVX1 U2388 ( .A(SH[8]), .Y(n3415) );
  INVX1 U2389 ( .A(SH[8]), .Y(n3414) );
  NOR2X1 U2390 ( .A(n3424), .B(n3245), .Y(n3244) );
  OR2X1 U2391 ( .A(A[175]), .B(n3393), .Y(n3245) );
  INVX1 U2392 ( .A(n1296), .Y(n416) );
  INVX1 U2393 ( .A(SH[8]), .Y(n3416) );
  MUX2IX1 U2394 ( .D0(n3337), .D1(n80), .S(n3375), .Y(n240) );
  INVX1 U2395 ( .A(n1248), .Y(n368) );
  INVX1 U2396 ( .A(n1320), .Y(n440) );
  INVX1 U2397 ( .A(n1328), .Y(n448) );
  MUX2IX1 U2398 ( .D0(n122), .D1(n154), .S(n3372), .Y(n58) );
  MUX2IX1 U2399 ( .D0(n186), .D1(n218), .S(n3230), .Y(n90) );
  MUX2IX1 U2400 ( .D0(n3271), .D1(n3331), .S(n3377), .Y(n154) );
  MUX2IX1 U2401 ( .D0(n335), .D1(n3293), .S(n3211), .Y(n215) );
  MUX2IX1 U2402 ( .D0(n57), .D1(n89), .S(n3213), .Y(n25) );
  MUX2IX1 U2403 ( .D0(n185), .D1(n217), .S(n3230), .Y(n89) );
  MUX2IX1 U2404 ( .D0(n117), .D1(n149), .S(n3372), .Y(n53) );
  MUX2IX1 U2405 ( .D0(n333), .D1(n3283), .S(n3211), .Y(n213) );
  MUX2IX1 U2406 ( .D0(n125), .D1(n157), .S(n3372), .Y(n61) );
  MUX2IX1 U2407 ( .D0(n189), .D1(n221), .S(n3372), .Y(n93) );
  MUX2IX1 U2408 ( .D0(n3285), .D1(n3255), .S(n3377), .Y(n157) );
  MUX2IX1 U2409 ( .D0(n59), .D1(n91), .S(SH[6]), .Y(n27) );
  MUX2IX1 U2410 ( .D0(n123), .D1(n155), .S(n3372), .Y(n59) );
  MUX2IX1 U2411 ( .D0(n187), .D1(n219), .S(SH[5]), .Y(n91) );
  MUX2IX1 U2412 ( .D0(n3357), .D1(n3351), .S(n3377), .Y(n155) );
  MUX2IX1 U2413 ( .D0(n182), .D1(n214), .S(n3369), .Y(n86) );
  MUX2IX1 U2414 ( .D0(n334), .D1(n3289), .S(n3210), .Y(n214) );
  MUX2IX1 U2415 ( .D0(n126), .D1(n158), .S(n3372), .Y(n62) );
  MUX2IX1 U2416 ( .D0(n190), .D1(n222), .S(SH[5]), .Y(n94) );
  MUX2IX1 U2417 ( .D0(n3291), .D1(n3329), .S(n3377), .Y(n158) );
  MUX2IX1 U2418 ( .D0(n188), .D1(n220), .S(n3230), .Y(n92) );
  MUX2IX1 U2419 ( .D0(n3281), .D1(n3333), .S(n3377), .Y(n156) );
  INVX1 U2420 ( .A(n1327), .Y(n447) );
  MUX2IX1 U2421 ( .D0(n318), .D1(n446), .S(n3381), .Y(n198) );
  INVX1 U2422 ( .A(n1326), .Y(n446) );
  INVX1 U2423 ( .A(n1198), .Y(n318) );
  MUX2IX1 U2424 ( .D0(n136), .D1(n168), .S(n3371), .Y(n72) );
  MUX2IX1 U2425 ( .D0(n3325), .D1(n416), .S(n3378), .Y(n168) );
  INVX1 U2426 ( .A(n1360), .Y(n480) );
  MUX2IX1 U2427 ( .D0(n202), .D1(n234), .S(n3369), .Y(n106) );
  MUX2IX1 U2428 ( .D0(n322), .D1(n450), .S(n3382), .Y(n202) );
  MUX2IX1 U2429 ( .D0(n354), .D1(n3247), .S(n3384), .Y(n234) );
  INVX1 U2430 ( .A(n1330), .Y(n450) );
  MUX2IX1 U2431 ( .D0(n3205), .D1(n239), .S(n3212), .Y(n111) );
  MUX2IX1 U2432 ( .D0(n359), .D1(n3253), .S(n3211), .Y(n239) );
  INVX1 U2433 ( .A(n1335), .Y(n455) );
  MUX2IX1 U2434 ( .D0(n3206), .D1(n233), .S(n3212), .Y(n105) );
  MUX2IX1 U2435 ( .D0(n353), .D1(n3259), .S(n3384), .Y(n233) );
  INVX1 U2436 ( .A(n1329), .Y(n449) );
  MUX2IX1 U2437 ( .D0(n3321), .D1(n416), .S(n3378), .Y(n167) );
  MUX2IX1 U2438 ( .D0(n205), .D1(n237), .S(n3369), .Y(n109) );
  MUX2IX1 U2439 ( .D0(n325), .D1(n453), .S(n3382), .Y(n205) );
  MUX2IX1 U2440 ( .D0(n357), .D1(n3263), .S(n3384), .Y(n237) );
  INVX1 U2441 ( .A(n1333), .Y(n453) );
  MUX2IX1 U2442 ( .D0(n133), .D1(n165), .S(n3371), .Y(n69) );
  MUX2IX1 U2443 ( .D0(n3315), .D1(n3347), .S(n3378), .Y(n165) );
  MUX2IX1 U2444 ( .D0(n3207), .D1(n238), .S(n3212), .Y(n110) );
  MUX2IX1 U2445 ( .D0(n358), .D1(n3265), .S(n3384), .Y(n238) );
  INVX1 U2446 ( .A(n1334), .Y(n454) );
  MUX2IX1 U2447 ( .D0(n3208), .D1(n236), .S(n3213), .Y(n108) );
  MUX2IX1 U2448 ( .D0(n356), .D1(n3261), .S(n3384), .Y(n236) );
  INVX1 U2449 ( .A(n1332), .Y(n452) );
  MUX2IX1 U2450 ( .D0(n134), .D1(n166), .S(n3371), .Y(n70) );
  MUX2IX1 U2451 ( .D0(n3317), .D1(n3349), .S(n3378), .Y(n166) );
  MUX2IX1 U2452 ( .D0(n3311), .D1(n3345), .S(n3378), .Y(n164) );
  INVX1 U2453 ( .A(n1359), .Y(n479) );
  MUX2IX1 U2454 ( .D0(n350), .D1(n478), .S(n3384), .Y(n230) );
  INVX1 U2455 ( .A(n1358), .Y(n478) );
  INVX1 U2456 ( .A(n1230), .Y(n350) );
  MUX2IX1 U2457 ( .D0(n343), .D1(n471), .S(n3383), .Y(n223) );
  INVX1 U2458 ( .A(n1351), .Y(n471) );
  INVX1 U2459 ( .A(n1223), .Y(n343) );
  MUX2IX1 U2460 ( .D0(n342), .D1(n470), .S(n3383), .Y(n222) );
  INVX1 U2461 ( .A(n1350), .Y(n470) );
  INVX1 U2462 ( .A(n1222), .Y(n342) );
  MUX2IX1 U2463 ( .D0(n50), .D1(n82), .S(n3374), .Y(n18) );
  MUX2IX1 U2464 ( .D0(n178), .D1(n210), .S(n3370), .Y(n82) );
  MUX2IX1 U2465 ( .D0(n114), .D1(n146), .S(n3230), .Y(n50) );
  MUX2IX1 U2466 ( .D0(n330), .D1(n3269), .S(n3211), .Y(n210) );
  MUX2IX1 U2467 ( .D0(n49), .D1(n81), .S(n3212), .Y(n17) );
  MUX2IX1 U2468 ( .D0(n113), .D1(n145), .S(n3230), .Y(n49) );
  MUX2IX1 U2469 ( .D0(n329), .D1(n3249), .S(n3382), .Y(n209) );
  MUX2IX1 U2470 ( .D0(n51), .D1(n83), .S(n3213), .Y(n19) );
  MUX2IX1 U2471 ( .D0(n179), .D1(n211), .S(n3230), .Y(n83) );
  MUX2IX1 U2472 ( .D0(n115), .D1(n147), .S(n3230), .Y(n51) );
  MUX2IX1 U2473 ( .D0(n331), .D1(n3355), .S(n3210), .Y(n211) );
  INVX1 U2474 ( .A(n1256), .Y(n376) );
  MUX2IX1 U2475 ( .D0(n241), .D1(n361), .S(n3380), .Y(n113) );
  INVX1 U2476 ( .A(n1241), .Y(n361) );
  INVX1 U2477 ( .A(n1121), .Y(n241) );
  INVX1 U2478 ( .A(n1247), .Y(n367) );
  INVX1 U2479 ( .A(n1127), .Y(n247) );
  MUX2IX1 U2480 ( .D0(n305), .D1(n433), .S(n3380), .Y(n185) );
  INVX1 U2481 ( .A(n1313), .Y(n433) );
  INVX1 U2482 ( .A(n1185), .Y(n305) );
  MUX2IX1 U2483 ( .D0(n311), .D1(n439), .S(n3381), .Y(n191) );
  INVX1 U2484 ( .A(n1319), .Y(n439) );
  INVX1 U2485 ( .A(n1191), .Y(n311) );
  INVX1 U2486 ( .A(n1311), .Y(n431) );
  INVX1 U2487 ( .A(n1305), .Y(n425) );
  INVX1 U2488 ( .A(n1177), .Y(n297) );
  INVX1 U2489 ( .A(n1255), .Y(n375) );
  MUX2IX1 U2490 ( .D0(n3204), .D1(n369), .S(n3241), .Y(n121) );
  INVX1 U2491 ( .A(n1249), .Y(n369) );
  MUX2IX1 U2492 ( .D0(n243), .D1(n363), .S(n3381), .Y(n115) );
  INVX1 U2493 ( .A(n1243), .Y(n363) );
  INVX1 U2494 ( .A(n1123), .Y(n243) );
  MUX2IX1 U2495 ( .D0(n307), .D1(n435), .S(n3380), .Y(n187) );
  INVX1 U2496 ( .A(n1315), .Y(n435) );
  INVX1 U2497 ( .A(n1187), .Y(n307) );
  MUX2IX1 U2498 ( .D0(n3209), .D1(n366), .S(n3241), .Y(n118) );
  INVX1 U2499 ( .A(n1246), .Y(n366) );
  MUX2IX1 U2500 ( .D0(n310), .D1(n438), .S(n3381), .Y(n190) );
  INVX1 U2501 ( .A(n1318), .Y(n438) );
  INVX1 U2502 ( .A(n1190), .Y(n310) );
  MUX2IX1 U2503 ( .D0(n302), .D1(n430), .S(n3380), .Y(n182) );
  INVX1 U2504 ( .A(n1310), .Y(n430) );
  INVX1 U2505 ( .A(n1182), .Y(n302) );
  MUX2IX1 U2506 ( .D0(n254), .D1(n374), .S(SH[7]), .Y(n126) );
  INVX1 U2507 ( .A(n1254), .Y(n374) );
  INVX1 U2508 ( .A(n1134), .Y(n254) );
  INVX1 U2509 ( .A(n1207), .Y(n327) );
  INVX1 U2510 ( .A(n1206), .Y(n326) );
  INVX1 U2511 ( .A(n1215), .Y(n335) );
  INVX1 U2512 ( .A(n1214), .Y(n334) );
  INVX1 U2513 ( .A(n1321), .Y(n441) );
  MUX2IX1 U2514 ( .D0(n315), .D1(n443), .S(n3381), .Y(n195) );
  INVX1 U2515 ( .A(n1323), .Y(n443) );
  INVX1 U2516 ( .A(n1195), .Y(n315) );
  MUX2IX1 U2517 ( .D0(n130), .D1(n162), .S(n3371), .Y(n66) );
  MUX2IX1 U2518 ( .D0(n3303), .D1(n3341), .S(n3378), .Y(n162) );
  MUX2IX1 U2519 ( .D0(n129), .D1(n161), .S(n3371), .Y(n65) );
  MUX2IX1 U2520 ( .D0(n3305), .D1(n3343), .S(n3378), .Y(n161) );
  MUX2IX1 U2521 ( .D0(n203), .D1(n235), .S(n3369), .Y(n107) );
  MUX2IX1 U2522 ( .D0(n323), .D1(n451), .S(n3382), .Y(n203) );
  MUX2IX1 U2523 ( .D0(n355), .D1(n3353), .S(n3384), .Y(n235) );
  INVX1 U2524 ( .A(n1331), .Y(n451) );
  MUX2IX1 U2525 ( .D0(n131), .D1(n163), .S(n3371), .Y(n67) );
  MUX2IX1 U2526 ( .D0(n3361), .D1(n3365), .S(n3378), .Y(n163) );
  MUX2IX1 U2527 ( .D0(n345), .D1(n473), .S(n3383), .Y(n225) );
  INVX1 U2528 ( .A(n1353), .Y(n473) );
  INVX1 U2529 ( .A(n1225), .Y(n345) );
  MUX2IX1 U2530 ( .D0(n338), .D1(n466), .S(n3383), .Y(n218) );
  INVX1 U2531 ( .A(n1346), .Y(n466) );
  MUX2IX1 U2532 ( .D0(n347), .D1(n475), .S(n3383), .Y(n227) );
  INVX1 U2533 ( .A(n1355), .Y(n475) );
  INVX1 U2534 ( .A(n1227), .Y(n347) );
  MUX2IX1 U2535 ( .D0(n337), .D1(n465), .S(n3210), .Y(n217) );
  INVX1 U2536 ( .A(n1345), .Y(n465) );
  INVX1 U2537 ( .A(n1217), .Y(n337) );
  MUX2IX1 U2538 ( .D0(n339), .D1(n467), .S(n3211), .Y(n219) );
  INVX1 U2539 ( .A(n1347), .Y(n467) );
  INVX1 U2540 ( .A(n1219), .Y(n339) );
  MUX2IX1 U2541 ( .D0(n299), .D1(n427), .S(n3379), .Y(n179) );
  INVX1 U2542 ( .A(n1307), .Y(n427) );
  INVX1 U2543 ( .A(n1179), .Y(n299) );
  MUX2IX1 U2544 ( .D0(n251), .D1(n371), .S(SH[7]), .Y(n123) );
  INVX1 U2545 ( .A(n1251), .Y(n371) );
  INVX1 U2546 ( .A(n1131), .Y(n251) );
  INVX1 U2547 ( .A(n1202), .Y(n322) );
  INVX1 U2548 ( .A(n1201), .Y(n321) );
  INVX1 U2549 ( .A(n1203), .Y(n323) );
  INVX1 U2550 ( .A(n1209), .Y(n329) );
  INVX1 U2551 ( .A(n1211), .Y(n331) );
  MUX2X1 U2552 ( .D0(n1144), .D1(n1264), .S(n3376), .Y(n136) );
  MUX2X1 U2553 ( .D0(n1138), .D1(n1258), .S(SH[7]), .Y(n130) );
  MUX2IX1 U2554 ( .D0(n138), .D1(n170), .S(n3370), .Y(n74) );
  NAND2X1 U2555 ( .A(n386), .B(n3385), .Y(n138) );
  MUX2IX1 U2556 ( .D0(n3307), .D1(n3273), .S(n3378), .Y(n170) );
  INVX1 U2557 ( .A(n1266), .Y(n386) );
  NAND2X1 U2558 ( .A(n385), .B(n3385), .Y(n137) );
  MUX2IX1 U2559 ( .D0(n3309), .D1(n3277), .S(n3378), .Y(n169) );
  INVX1 U2560 ( .A(n1265), .Y(n385) );
  MUX2X1 U2561 ( .D0(n1143), .D1(n1263), .S(n3376), .Y(n135) );
  NAND2X1 U2562 ( .A(n388), .B(n3385), .Y(n140) );
  MUX2IX1 U2563 ( .D0(n3313), .D1(n3267), .S(n3379), .Y(n172) );
  INVX1 U2564 ( .A(n1268), .Y(n388) );
  MUX2IX1 U2565 ( .D0(n141), .D1(n173), .S(n3370), .Y(n77) );
  NAND2X1 U2566 ( .A(n389), .B(n3385), .Y(n141) );
  MUX2IX1 U2567 ( .D0(n3251), .D1(n3287), .S(n3379), .Y(n173) );
  INVX1 U2568 ( .A(n1269), .Y(n389) );
  NAND2X1 U2569 ( .A(n390), .B(n3385), .Y(n142) );
  MUX2IX1 U2570 ( .D0(n3319), .D1(n3335), .S(n3379), .Y(n174) );
  INVX1 U2571 ( .A(n1270), .Y(n390) );
  NAND2X1 U2572 ( .A(n391), .B(n3385), .Y(n143) );
  MUX2IX1 U2573 ( .D0(n3323), .D1(n3297), .S(n3379), .Y(n175) );
  INVX1 U2574 ( .A(n1271), .Y(n391) );
  MUX2IX1 U2575 ( .D0(n144), .D1(n176), .S(n3370), .Y(n80) );
  NAND2X1 U2576 ( .A(n392), .B(n3385), .Y(n144) );
  MUX2IX1 U2577 ( .D0(n3327), .D1(n3301), .S(n3379), .Y(n176) );
  INVX1 U2578 ( .A(n1272), .Y(n392) );
  MUX2X1 U2579 ( .D0(n1148), .D1(n1276), .S(n3376), .Y(n148) );
  MUX2X1 U2580 ( .D0(n1137), .D1(n1257), .S(SH[7]), .Y(n129) );
  MUX2X1 U2581 ( .D0(n1139), .D1(n1259), .S(SH[7]), .Y(n131) );
  MUX2X1 U2582 ( .D0(n1140), .D1(n1260), .S(n3385), .Y(n132) );
  MUX2X1 U2583 ( .D0(n1141), .D1(n1261), .S(n3376), .Y(n133) );
  MUX2X1 U2584 ( .D0(n1142), .D1(n1262), .S(n3376), .Y(n134) );
  MUX2X1 U2585 ( .D0(n1149), .D1(n1277), .S(n3376), .Y(n149) );
  MUX2X1 U2586 ( .D0(n1146), .D1(n1274), .S(n3376), .Y(n146) );
  MUX2X1 U2587 ( .D0(n1145), .D1(n1273), .S(n3376), .Y(n145) );
  MUX2X1 U2588 ( .D0(n1151), .D1(n1279), .S(n3377), .Y(n151) );
  INVX1 U2589 ( .A(n3442), .Y(n3435) );
  INVX1 U2590 ( .A(n3443), .Y(n3419) );
  INVX1 U2591 ( .A(n3441), .Y(n3439) );
  INVX1 U2592 ( .A(n3443), .Y(n3431) );
  INVX1 U2593 ( .A(n3441), .Y(n3423) );
  INVX1 U2594 ( .A(n3443), .Y(n3434) );
  INVX1 U2595 ( .A(n3443), .Y(n3430) );
  INVX1 U2596 ( .A(n3441), .Y(n3426) );
  INVX1 U2597 ( .A(n3442), .Y(n3422) );
  INVX1 U2598 ( .A(n3443), .Y(n3418) );
  INVX1 U2599 ( .A(n3442), .Y(n3437) );
  INVX1 U2600 ( .A(n3441), .Y(n3421) );
  INVX1 U2601 ( .A(n3443), .Y(n3429) );
  INVX1 U2602 ( .A(n3441), .Y(n3438) );
  INVX1 U2603 ( .A(n3443), .Y(n3433) );
  INVX1 U2604 ( .A(n3442), .Y(n3420) );
  INVX1 U2605 ( .A(n3443), .Y(n3417) );
  INVX1 U2606 ( .A(n3442), .Y(n3427) );
  INVX1 U2607 ( .A(n3441), .Y(n3424) );
  INVX1 U2608 ( .A(n3442), .Y(n3436) );
  INVX1 U2609 ( .A(n3442), .Y(n3428) );
  INVX1 U2610 ( .A(n3443), .Y(n3432) );
  INVX1 U2611 ( .A(n3442), .Y(n3425) );
  INVX1 U2612 ( .A(n3441), .Y(n3440) );
  MUX2IX1 U2613 ( .D0(n139), .D1(n171), .S(n3370), .Y(n75) );
  NAND2X1 U2614 ( .A(n387), .B(n3385), .Y(n139) );
  MUX2IX1 U2615 ( .D0(n3363), .D1(n3359), .S(n3379), .Y(n171) );
  INVX1 U2616 ( .A(n1267), .Y(n387) );
  MUX2X1 U2617 ( .D0(n1147), .D1(n1275), .S(n3376), .Y(n147) );
  INVX1 U2618 ( .A(n3373), .Y(n3370) );
  INVX1 U2619 ( .A(n3387), .Y(n3382) );
  INVX1 U2620 ( .A(n3386), .Y(n3380) );
  INVX1 U2621 ( .A(n3387), .Y(n3384) );
  INVX1 U2622 ( .A(n3386), .Y(n3376) );
  INVX1 U2623 ( .A(n3386), .Y(n3378) );
  INVX1 U2624 ( .A(n3387), .Y(n3381) );
  INVX1 U2625 ( .A(n3387), .Y(n3383) );
  INVX1 U2626 ( .A(n3386), .Y(n3377) );
  INVX1 U2627 ( .A(n3386), .Y(n3379) );
  INVX1 U2628 ( .A(n3373), .Y(n3372) );
  INVX1 U2629 ( .A(n3373), .Y(n3371) );
  INVX1 U2630 ( .A(n3375), .Y(n3374) );
  INVX1 U2631 ( .A(n3387), .Y(n3385) );
  MUX2IX1 U2632 ( .D0(A[73]), .D1(A[329]), .S(n3393), .Y(n955) );
  MUX2IX1 U2633 ( .D0(A[72]), .D1(A[328]), .S(n3393), .Y(n958) );
  MUX2IX1 U2634 ( .D0(A[78]), .D1(A[334]), .S(n3392), .Y(n940) );
  MUX2IX1 U2635 ( .D0(A[76]), .D1(A[332]), .S(n3393), .Y(n946) );
  MUX2IX1 U2636 ( .D0(A[74]), .D1(A[330]), .S(n3392), .Y(n952) );
  MUX2IX1 U2637 ( .D0(A[77]), .D1(A[333]), .S(n3392), .Y(n943) );
  MUX2IX1 U2638 ( .D0(A[75]), .D1(A[331]), .S(n3393), .Y(n949) );
  INVX1 U2639 ( .A(n1234), .Y(n354) );
  MUX2IX1 U2640 ( .D0(A[121]), .D1(A[377]), .S(n3391), .Y(n811) );
  INVX1 U2641 ( .A(n1239), .Y(n359) );
  MUX2IX1 U2642 ( .D0(A[126]), .D1(A[382]), .S(n3391), .Y(n796) );
  INVX1 U2643 ( .A(n1233), .Y(n353) );
  MUX2IX1 U2644 ( .D0(A[120]), .D1(A[376]), .S(n3391), .Y(n814) );
  MUX2IX1 U2645 ( .D0(A[1]), .D1(A[257]), .S(n3388), .Y(n1115) );
  MUX2IX1 U2646 ( .D0(A[124]), .D1(A[380]), .S(n3390), .Y(n802) );
  INVX1 U2647 ( .A(n1238), .Y(n358) );
  MUX2IX1 U2648 ( .D0(A[125]), .D1(A[381]), .S(n3390), .Y(n799) );
  MUX2IX1 U2649 ( .D0(A[123]), .D1(A[379]), .S(n3390), .Y(n805) );
  MUX2IX1 U2650 ( .D0(A[0]), .D1(A[256]), .S(n3391), .Y(n1118) );
  MUX2IX1 U2651 ( .D0(A[6]), .D1(A[262]), .S(n3394), .Y(n1100) );
  MUX2IX1 U2652 ( .D0(A[4]), .D1(A[260]), .S(n3394), .Y(n1106) );
  MUX2IX1 U2653 ( .D0(A[2]), .D1(A[258]), .S(n3392), .Y(n1112) );
  MUX2IX1 U2654 ( .D0(A[3]), .D1(A[259]), .S(n3394), .Y(n1109) );
  MUX2IX1 U2655 ( .D0(A[65]), .D1(A[321]), .S(n3392), .Y(n979) );
  MUX2IX1 U2656 ( .D0(A[9]), .D1(A[265]), .S(n3392), .Y(n1091) );
  MUX2IX1 U2657 ( .D0(A[68]), .D1(A[324]), .S(n3392), .Y(n970) );
  MUX2IX1 U2658 ( .D0(A[12]), .D1(A[268]), .S(n3394), .Y(n1082) );
  MUX2IX1 U2659 ( .D0(A[69]), .D1(A[325]), .S(n3394), .Y(n967) );
  MUX2IX1 U2660 ( .D0(A[13]), .D1(A[269]), .S(n3394), .Y(n1079) );
  MUX2IX1 U2661 ( .D0(A[67]), .D1(A[323]), .S(n3392), .Y(n973) );
  INVX1 U2662 ( .A(n1235), .Y(n355) );
  MUX2IX1 U2663 ( .D0(A[122]), .D1(A[378]), .S(n3390), .Y(n808) );
  MUX2IX1 U2664 ( .D0(A[66]), .D1(A[322]), .S(n3394), .Y(n976) );
  MUX2IX1 U2665 ( .D0(A[10]), .D1(A[266]), .S(n3394), .Y(n1088) );
  MUX2IX1 U2666 ( .D0(A[151]), .D1(A[407]), .S(n3390), .Y(n721) );
  MUX2IX1 U2667 ( .D0(A[128]), .D1(A[384]), .S(n3388), .Y(n790) );
  MUX2IX1 U2668 ( .D0(A[135]), .D1(A[391]), .S(n3388), .Y(n769) );
  MUX2IX1 U2669 ( .D0(A[143]), .D1(A[399]), .S(n3389), .Y(n745) );
  MUX2IX1 U2670 ( .D0(A[145]), .D1(A[401]), .S(n3389), .Y(n739) );
  NOR2X1 U2671 ( .A(SH[9]), .B(n3248), .Y(n3247) );
  OR2X1 U2672 ( .A(n3401), .B(A[249]), .Y(n3248) );
  MUX2IX1 U2673 ( .D0(A[144]), .D1(A[400]), .S(n3389), .Y(n742) );
  NOR2X1 U2674 ( .A(n3419), .B(n3250), .Y(n3249) );
  OR2X1 U2675 ( .A(n3408), .B(A[224]), .Y(n3250) );
  MUX2IX1 U2676 ( .D0(A[146]), .D1(A[402]), .S(n3390), .Y(n736) );
  MUX2IX1 U2677 ( .D0(A[147]), .D1(A[403]), .S(n3390), .Y(n733) );
  MUX2IX1 U2678 ( .D0(A[148]), .D1(A[404]), .S(n3390), .Y(n730) );
  MUX2IX1 U2679 ( .D0(A[149]), .D1(A[405]), .S(n3390), .Y(n727) );
  MUX2IX1 U2680 ( .D0(A[150]), .D1(A[406]), .S(n3390), .Y(n724) );
  NOR2X1 U2681 ( .A(n3435), .B(n3252), .Y(n3251) );
  OR2X1 U2682 ( .A(n3406), .B(A[60]), .Y(n3252) );
  NOR2X1 U2683 ( .A(n3424), .B(n3254), .Y(n3253) );
  OR2X1 U2684 ( .A(n3400), .B(A[254]), .Y(n3254) );
  MUX2IX1 U2685 ( .D0(A[129]), .D1(A[385]), .S(n3388), .Y(n787) );
  MUX2IX1 U2686 ( .D0(A[193]), .D1(A[449]), .S(n3391), .Y(n635) );
  MUX2IX1 U2687 ( .D0(A[209]), .D1(A[465]), .S(n3391), .Y(n587) );
  MUX2IX1 U2688 ( .D0(A[201]), .D1(A[457]), .S(n3391), .Y(n611) );
  MUX2IX1 U2689 ( .D0(A[137]), .D1(A[393]), .S(n3389), .Y(n763) );
  MUX2IX1 U2690 ( .D0(A[192]), .D1(A[448]), .S(n3391), .Y(n638) );
  MUX2IX1 U2691 ( .D0(A[208]), .D1(A[464]), .S(n3391), .Y(n590) );
  MUX2IX1 U2692 ( .D0(A[200]), .D1(A[456]), .S(n3391), .Y(n614) );
  MUX2IX1 U2693 ( .D0(A[136]), .D1(A[392]), .S(n3389), .Y(n766) );
  MUX2IX1 U2694 ( .D0(A[130]), .D1(A[386]), .S(n3388), .Y(n784) );
  MUX2IX1 U2695 ( .D0(A[138]), .D1(A[394]), .S(n3389), .Y(n760) );
  MUX2IX1 U2696 ( .D0(A[131]), .D1(A[387]), .S(n3388), .Y(n781) );
  MUX2IX1 U2697 ( .D0(A[139]), .D1(A[395]), .S(n3389), .Y(n757) );
  MUX2IX1 U2698 ( .D0(A[132]), .D1(A[388]), .S(n3388), .Y(n778) );
  MUX2IX1 U2699 ( .D0(A[140]), .D1(A[396]), .S(n3389), .Y(n754) );
  MUX2IX1 U2700 ( .D0(A[133]), .D1(A[389]), .S(n3388), .Y(n775) );
  MUX2IX1 U2701 ( .D0(A[141]), .D1(A[397]), .S(n3389), .Y(n751) );
  MUX2IX1 U2702 ( .D0(A[134]), .D1(A[390]), .S(n3388), .Y(n772) );
  MUX2IX1 U2703 ( .D0(A[142]), .D1(A[398]), .S(n3389), .Y(n748) );
  NOR2X1 U2704 ( .A(n3424), .B(n3256), .Y(n3255) );
  OR2X1 U2705 ( .A(n3410), .B(A[172]), .Y(n3256) );
  NOR2X1 U2706 ( .A(n3424), .B(n3258), .Y(n3257) );
  OR2X1 U2707 ( .A(n3410), .B(A[168]), .Y(n3258) );
  NOR2X1 U2708 ( .A(SH[9]), .B(n3260), .Y(n3259) );
  OR2X1 U2709 ( .A(n3401), .B(A[248]), .Y(n3260) );
  NOR2X1 U2710 ( .A(n3423), .B(n3262), .Y(n3261) );
  OR2X1 U2711 ( .A(n3401), .B(A[251]), .Y(n3262) );
  NOR2X1 U2712 ( .A(SH[9]), .B(n3264), .Y(n3263) );
  OR2X1 U2713 ( .A(n3401), .B(A[252]), .Y(n3264) );
  NOR2X1 U2714 ( .A(SH[9]), .B(n3266), .Y(n3265) );
  OR2X1 U2715 ( .A(n3401), .B(A[253]), .Y(n3266) );
  NOR2X1 U2716 ( .A(n3422), .B(n3268), .Y(n3267) );
  OR2X1 U2717 ( .A(n3409), .B(A[187]), .Y(n3268) );
  NOR2X1 U2718 ( .A(n3419), .B(n3270), .Y(n3269) );
  OR2X1 U2719 ( .A(n3407), .B(A[225]), .Y(n3270) );
  NOR2X1 U2720 ( .A(n3437), .B(n3272), .Y(n3271) );
  OR2X1 U2721 ( .A(n3404), .B(A[41]), .Y(n3272) );
  NOR2X1 U2722 ( .A(n3423), .B(n3274), .Y(n3273) );
  OR2X1 U2723 ( .A(n3409), .B(A[185]), .Y(n3274) );
  NOR2X1 U2724 ( .A(n3437), .B(n3276), .Y(n3275) );
  OR2X1 U2725 ( .A(n3404), .B(A[40]), .Y(n3276) );
  NOR2X1 U2726 ( .A(n3423), .B(n3278), .Y(n3277) );
  OR2X1 U2727 ( .A(n3409), .B(A[184]), .Y(n3278) );
  NOR2X1 U2728 ( .A(n3418), .B(n3280), .Y(n3279) );
  OR2X1 U2729 ( .A(n3407), .B(A[227]), .Y(n3280) );
  NOR2X1 U2730 ( .A(n3437), .B(n3282), .Y(n3281) );
  OR2X1 U2731 ( .A(n3404), .B(A[43]), .Y(n3282) );
  NOR2X1 U2732 ( .A(n3418), .B(n3284), .Y(n3283) );
  OR2X1 U2733 ( .A(n3407), .B(A[228]), .Y(n3284) );
  NOR2X1 U2734 ( .A(n3437), .B(n3286), .Y(n3285) );
  OR2X1 U2735 ( .A(n3404), .B(A[44]), .Y(n3286) );
  NOR2X1 U2736 ( .A(n3422), .B(n3288), .Y(n3287) );
  OR2X1 U2737 ( .A(n3409), .B(A[188]), .Y(n3288) );
  NOR2X1 U2738 ( .A(n3418), .B(n3290), .Y(n3289) );
  OR2X1 U2739 ( .A(n3407), .B(A[229]), .Y(n3290) );
  NOR2X1 U2740 ( .A(n3437), .B(n3292), .Y(n3291) );
  OR2X1 U2741 ( .A(n3404), .B(A[45]), .Y(n3292) );
  NOR2X1 U2742 ( .A(n3418), .B(n3294), .Y(n3293) );
  OR2X1 U2743 ( .A(n3407), .B(A[230]), .Y(n3294) );
  NOR2X1 U2744 ( .A(n3436), .B(n3296), .Y(n3295) );
  OR2X1 U2745 ( .A(n3404), .B(A[46]), .Y(n3296) );
  NOR2X1 U2746 ( .A(n3422), .B(n3298), .Y(n3297) );
  OR2X1 U2747 ( .A(n3409), .B(A[190]), .Y(n3298) );
  NOR2X1 U2748 ( .A(n3436), .B(n3300), .Y(n3299) );
  OR2X1 U2749 ( .A(n3404), .B(A[47]), .Y(n3300) );
  NOR2X1 U2750 ( .A(n3422), .B(n3302), .Y(n3301) );
  OR2X1 U2751 ( .A(n3408), .B(A[191]), .Y(n3302) );
  NOR2X1 U2752 ( .A(n3436), .B(n3304), .Y(n3303) );
  OR2X1 U2753 ( .A(n3404), .B(A[49]), .Y(n3304) );
  NOR2X1 U2754 ( .A(n3436), .B(n3306), .Y(n3305) );
  OR2X1 U2755 ( .A(n3404), .B(A[48]), .Y(n3306) );
  NOR2X1 U2756 ( .A(n3435), .B(n3308), .Y(n3307) );
  OR2X1 U2757 ( .A(n3405), .B(A[57]), .Y(n3308) );
  NOR2X1 U2758 ( .A(n3435), .B(n3310), .Y(n3309) );
  OR2X1 U2759 ( .A(n3405), .B(A[56]), .Y(n3310) );
  NOR2X1 U2760 ( .A(n3436), .B(n3312), .Y(n3311) );
  OR2X1 U2761 ( .A(n3405), .B(A[51]), .Y(n3312) );
  NOR2X1 U2762 ( .A(n3435), .B(n3314), .Y(n3313) );
  OR2X1 U2763 ( .A(n3405), .B(A[59]), .Y(n3314) );
  NOR2X1 U2764 ( .A(n3436), .B(n3316), .Y(n3315) );
  OR2X1 U2765 ( .A(n3405), .B(A[52]), .Y(n3316) );
  NOR2X1 U2766 ( .A(n3436), .B(n3318), .Y(n3317) );
  OR2X1 U2767 ( .A(n3405), .B(A[53]), .Y(n3318) );
  NOR2X1 U2768 ( .A(n3435), .B(n3320), .Y(n3319) );
  OR2X1 U2769 ( .A(n3406), .B(A[61]), .Y(n3320) );
  NOR2X1 U2770 ( .A(n3436), .B(n3322), .Y(n3321) );
  OR2X1 U2771 ( .A(n3405), .B(A[54]), .Y(n3322) );
  NOR2X1 U2772 ( .A(n3435), .B(n3324), .Y(n3323) );
  OR2X1 U2773 ( .A(n3406), .B(A[62]), .Y(n3324) );
  NOR2X1 U2774 ( .A(n3436), .B(n3326), .Y(n3325) );
  OR2X1 U2775 ( .A(n3405), .B(A[55]), .Y(n3326) );
  NOR2X1 U2776 ( .A(n3435), .B(n3328), .Y(n3327) );
  OR2X1 U2777 ( .A(n3406), .B(A[63]), .Y(n3328) );
  NOR2X1 U2778 ( .A(n3424), .B(n3330), .Y(n3329) );
  OR2X1 U2779 ( .A(n3410), .B(A[173]), .Y(n3330) );
  NOR2X1 U2780 ( .A(n3424), .B(n3332), .Y(n3331) );
  OR2X1 U2781 ( .A(n3410), .B(A[169]), .Y(n3332) );
  NOR2X1 U2782 ( .A(n3424), .B(n3334), .Y(n3333) );
  OR2X1 U2783 ( .A(n3410), .B(A[171]), .Y(n3334) );
  NOR2X1 U2784 ( .A(n3422), .B(n3336), .Y(n3335) );
  OR2X1 U2785 ( .A(n3409), .B(A[189]), .Y(n3336) );
  NOR2X1 U2786 ( .A(n3440), .B(n3338), .Y(n3337) );
  OR2X1 U2787 ( .A(n3406), .B(A[255]), .Y(n3338) );
  NOR2X1 U2788 ( .A(n3418), .B(n3340), .Y(n3339) );
  OR2X1 U2789 ( .A(n3407), .B(A[231]), .Y(n3340) );
  NOR2X1 U2790 ( .A(n3423), .B(n3342), .Y(n3341) );
  OR2X1 U2791 ( .A(n3410), .B(A[177]), .Y(n3342) );
  NOR2X1 U2792 ( .A(n3423), .B(n3344), .Y(n3343) );
  OR2X1 U2793 ( .A(n3410), .B(A[176]), .Y(n3344) );
  NOR2X1 U2794 ( .A(n3423), .B(n3346), .Y(n3345) );
  OR2X1 U2795 ( .A(n3409), .B(A[179]), .Y(n3346) );
  NOR2X1 U2796 ( .A(n3423), .B(n3348), .Y(n3347) );
  OR2X1 U2797 ( .A(n3409), .B(A[180]), .Y(n3348) );
  NOR2X1 U2798 ( .A(n3423), .B(n3350), .Y(n3349) );
  OR2X1 U2799 ( .A(n3409), .B(A[181]), .Y(n3350) );
  INVX1 U2800 ( .A(SH[9]), .Y(n3442) );
  INVX1 U2801 ( .A(SH[9]), .Y(n3441) );
  INVX1 U2802 ( .A(SH[9]), .Y(n3443) );
  NOR2X1 U2803 ( .A(n3424), .B(n3352), .Y(n3351) );
  OR2X1 U2804 ( .A(n3410), .B(A[170]), .Y(n3352) );
  NOR2X1 U2805 ( .A(SH[9]), .B(n3354), .Y(n3353) );
  OR2X1 U2806 ( .A(n3401), .B(A[250]), .Y(n3354) );
  NOR2X1 U2807 ( .A(n3418), .B(n3356), .Y(n3355) );
  OR2X1 U2808 ( .A(n3407), .B(A[226]), .Y(n3356) );
  NOR2X1 U2809 ( .A(n3437), .B(n3358), .Y(n3357) );
  OR2X1 U2810 ( .A(n3404), .B(A[42]), .Y(n3358) );
  NOR2X1 U2811 ( .A(n3422), .B(n3360), .Y(n3359) );
  OR2X1 U2812 ( .A(n3409), .B(A[186]), .Y(n3360) );
  INVX1 U2813 ( .A(SH[7]), .Y(n3387) );
  INVX1 U2814 ( .A(n3238), .Y(n3369) );
  NOR2X1 U2815 ( .A(n3436), .B(n3362), .Y(n3361) );
  OR2X1 U2816 ( .A(n3405), .B(A[50]), .Y(n3362) );
  NOR2X1 U2817 ( .A(n3435), .B(n3364), .Y(n3363) );
  OR2X1 U2818 ( .A(n3405), .B(A[58]), .Y(n3364) );
  NOR2X1 U2819 ( .A(n3423), .B(n3366), .Y(n3365) );
  OR2X1 U2820 ( .A(n3410), .B(A[178]), .Y(n3366) );
  INVX1 U2821 ( .A(SH[6]), .Y(n3375) );
  INVX1 U2822 ( .A(SH[7]), .Y(n3386) );
  INVX1 U2823 ( .A(SH[5]), .Y(n3373) );
  BUFX3 U2824 ( .A(SH[4]), .Y(n3368) );
  BUFX3 U2825 ( .A(SH[4]), .Y(n3367) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regx_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N16, N17, N18, N19, N20,
         net9015, n12, n5, n7, n1, n2, n3, n4, n6, n8, n9, n10, n11, n13, n14,
         n15, n16, n17;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9015), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N20), .SIN(db_cnt_2_), .SMC(test_se), .C(net9015), .XR(rstz), .Q(test_so) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N18), .SIN(db_cnt_0_), .SMC(test_se), .C(net9015), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N17), .SIN(o_dbc), .SMC(test_se), .C(net9015), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N19), .SIN(db_cnt_1_), .SMC(test_se), .C(net9015), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n12), .SIN(d_org_0_), .SMC(test_se), .C(net9015), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n17), .Y(n16) );
  NAND32X1 U4 ( .B(n13), .C(n11), .A(n15), .Y(n3) );
  NAND21X1 U5 ( .B(n10), .A(n3), .Y(n17) );
  NAND21X1 U6 ( .B(n17), .A(n15), .Y(n5) );
  XNOR2XL U7 ( .A(d_org_0_), .B(o_dbc), .Y(n10) );
  INVX1 U8 ( .A(n1), .Y(n15) );
  NAND21X1 U9 ( .B(n9), .A(db_cnt_0_), .Y(n1) );
  OAI22X1 U10 ( .A(db_cnt_2_), .B(n5), .C(n7), .D(n11), .Y(N19) );
  AOI21BBXL U11 ( .B(n17), .C(db_cnt_1_), .A(N17), .Y(n7) );
  INVX1 U12 ( .A(n8), .Y(N17) );
  NAND21X1 U13 ( .B(db_cnt_0_), .A(n16), .Y(n8) );
  INVX1 U14 ( .A(db_cnt_2_), .Y(n11) );
  ENOX1 U15 ( .A(n11), .B(n5), .C(test_so), .D(n16), .Y(N20) );
  INVX1 U16 ( .A(db_cnt_1_), .Y(n9) );
  INVX1 U17 ( .A(test_so), .Y(n13) );
  MUX2X1 U18 ( .D0(o_dbc), .D1(d_org_0_), .S(o_chg), .Y(n12) );
  INVX1 U19 ( .A(n6), .Y(o_chg) );
  NAND21X1 U20 ( .B(n10), .A(n4), .Y(n6) );
  INVX1 U21 ( .A(n3), .Y(n4) );
  NAND5XL U22 ( .A(n14), .B(n13), .C(n11), .D(n10), .E(n9), .Y(N16) );
  INVX1 U23 ( .A(db_cnt_0_), .Y(n14) );
  AND2X1 U24 ( .A(n2), .B(n16), .Y(N18) );
  XOR2X1 U25 ( .A(db_cnt_0_), .B(db_cnt_1_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N16, N17, N18, N19, N20,
         net9033, n12, n3, n4, n5, n6, n7, n8, n9, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9033), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N20), .SIN(db_cnt_2_), .SMC(test_se), .C(net9033), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N18), .SIN(db_cnt_0_), .SMC(test_se), .C(net9033), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N17), .SIN(o_dbc), .SMC(test_se), .C(net9033), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N19), .SIN(db_cnt_1_), .SMC(test_se), .C(net9033), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n12), .SIN(d_org_0_), .SMC(test_se), .C(net9033), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n6), .Y(n1) );
  NOR21XL U4 ( .B(n3), .A(n4), .Y(n6) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  OAI22X1 U6 ( .A(db_cnt_2_), .B(n5), .C(n7), .D(n2), .Y(N19) );
  AOI21BBXL U7 ( .B(n1), .C(db_cnt_1_), .A(N17), .Y(n7) );
  AO22AXL U8 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR2X1 U9 ( .A(n3), .B(n4), .Y(o_chg) );
  NOR2X1 U10 ( .A(n1), .B(db_cnt_0_), .Y(N17) );
  NAND4X1 U11 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_1_), .D(db_cnt_0_), .Y(
        n3) );
  NAND3X1 U12 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(n6), .Y(n5) );
  ENOX1 U13 ( .A(n2), .B(n5), .C(test_so), .D(n6), .Y(N20) );
  NOR2X1 U14 ( .A(n8), .B(n1), .Y(N18) );
  XNOR2XL U15 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n8) );
  NAND31X1 U16 ( .C(db_cnt_0_), .A(n4), .B(n9), .Y(N16) );
  NOR3XL U17 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n9) );
  INVX1 U18 ( .A(db_cnt_2_), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_4 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_5 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_6 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_7 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module glreg_a0_7 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9051;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_7 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9051), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9051), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9051), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9051), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9051), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9051), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9051), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9051), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9051), 
        .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_8 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9069;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_8 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9069), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9069), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9069), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9069), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9069), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9069), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9069), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9069), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9069), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_9 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9087;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_9 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9087), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9087), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9087), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9087), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9087), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9087), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9087), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9087), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9087), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH7_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9105;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9105), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9105), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9105), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9105), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9105), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9105), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9105), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9105), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_8 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n7, n8, n9, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n7) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n8) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module glreg_a0_10 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9123;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_10 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9123), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9123), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9123), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9123), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9123), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9123), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9123), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9123), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9123), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_11 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9141;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_11 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9141), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9141), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9141), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9141), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9141), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9141), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9141), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9141), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9141), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_12 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9159;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_12 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9159), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9159), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9159), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9159), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9159), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9159), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9159), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9159), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9159), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_13 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9177;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_13 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9177), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9177), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9177), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9177), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9177), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9177), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9177), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9177), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9177), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_14 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9195;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_14 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9195), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9195), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9195), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9195), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9195), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9195), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9195), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9195), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9195), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9213;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9213), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9213), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9213), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9213), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9213), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9213), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9213), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9231;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9231), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9231), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9231), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9231), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9231), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9231), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9231), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_15 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9249;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_15 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9249), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9249), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9249), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9249), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9249), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9249), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9249), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9249), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9249), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_6_00000002 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9267;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9267), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9267), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9267), 
        .XS(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9267), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9267), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9267), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9267), 
        .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  MUX2X1 U2 ( .D0(rdat[0]), .D1(wdat[0]), .S(we), .Y(n2) );
endmodule


module glreg_a0_16 ( clk, arstz, we, wdat, rdat, test_si2, test_si1, test_se
 );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si2, test_si1, test_se;
  wire   net9285;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_16 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9285), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(test_si2), .SMC(test_se), .C(net9285), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9285), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9285), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si1), .SMC(test_se), .C(net9285), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9285), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[3]), .SMC(test_se), .C(net9285), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9285), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9285), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_17 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9303;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_17 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9303), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9303), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9303), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9303), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9303), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9303), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9303), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9303), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9303), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_18 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9321;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_18 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9321), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9321), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9321), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9321), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9321), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9321), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9321), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9321), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9321), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_19 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9339;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_19 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9339), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9339), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9339), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9339), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9339), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9339), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9339), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9339), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9339), 
        .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module cvctl_a0 ( r_cvcwr, wdat, r_sdischg, r_vcomp, r_idacsh, r_cvofsx, 
        r_cvofs, sdischg_duty, r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, 
        r_fw_pwrv, r_dac0, r_dac3, clk_100k, clk, srstz, test_si, test_se );
  input [5:0] r_cvcwr;
  input [7:0] wdat;
  output [7:0] r_sdischg;
  output [7:0] r_vcomp;
  output [7:0] r_idacsh;
  output [7:0] r_cvofsx;
  output [15:0] r_cvofs;
  input [11:0] r_fw_pwrv;
  output [10:0] r_dac0;
  output [5:0] r_dac3;
  input r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, clk_100k, clk, srstz,
         test_si, test_se;
  output sdischg_duty;
  wire   clk_5k, N29, N34, N35, N36, N38, N39, N40, N41, N42, N47, N84, N94,
         N95, N96, N97, N98, N99, N106, N107, N108, N109, N115, N121, N122,
         N123, N126, N127, N128, N129, N130, net9357, n81, N68, N67, N66, N65,
         N64, N63, N62, N61, N60, n2, n4, n5, n6, n7, n8, n9, N83, N82, N81,
         N80, N79, N78, N77, N76, N75, N74, N73, N72, N59, N58, N57, N56, N55,
         N54, N53, N52, N51, N50, N49, N48, n34, n35, n36, n37, n38, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, add_62_carry_1_, add_62_carry_2_, add_62_carry_3_,
         add_62_carry_4_, add_62_carry_5_, n3, n12, n17, n18, n19, n20, n21,
         n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33;
  wire   [4:0] div20_cnt;
  wire   [10:1] cv_code;
  wire   [4:0] sdischg_cnt;
  wire   [4:2] add_81_carry;
  wire   [4:2] add_41_carry;
  wire   [2:1] add_3_root_sub_0_root_add_46_3_carry;

  HAD1X1 add_81_U1_1_1 ( .A(sdischg_cnt[1]), .B(sdischg_cnt[0]), .CO(
        add_81_carry[2]), .SO(N121) );
  HAD1X1 add_81_U1_1_2 ( .A(sdischg_cnt[2]), .B(add_81_carry[2]), .CO(
        add_81_carry[3]), .SO(N122) );
  HAD1X1 add_81_U1_1_3 ( .A(sdischg_cnt[3]), .B(add_81_carry[3]), .CO(
        add_81_carry[4]), .SO(N123) );
  HAD1X1 add_41_U1_1_1 ( .A(div20_cnt[1]), .B(div20_cnt[0]), .CO(
        add_41_carry[2]), .SO(N34) );
  HAD1X1 add_41_U1_1_2 ( .A(div20_cnt[2]), .B(add_41_carry[2]), .CO(
        add_41_carry[3]), .SO(N35) );
  HAD1X1 add_41_U1_1_3 ( .A(div20_cnt[3]), .B(add_41_carry[3]), .CO(
        add_41_carry[4]), .SO(N36) );
  FAD1X1 add_3_root_sub_0_root_add_46_3_U1_1 ( .A(N47), .B(r_vcomp[1]), .CI(
        add_3_root_sub_0_root_add_46_3_carry[1]), .CO(
        add_3_root_sub_0_root_add_46_3_carry[2]), .SO(N61) );
  INVX1 U4 ( .A(n9), .Y(n8) );
  INVX1 U5 ( .A(n9), .Y(n4) );
  INVX1 U6 ( .A(n9), .Y(n5) );
  INVX1 U7 ( .A(n9), .Y(n6) );
  INVX1 U8 ( .A(n9), .Y(n7) );
  INVX1 U9 ( .A(n9), .Y(n2) );
  INVX1 U10 ( .A(srstz), .Y(n9) );
  glreg_a0_25 u0_v_comp ( .clk(clk), .arstz(n8), .we(r_cvcwr[3]), .wdat(wdat), 
        .rdat(r_vcomp), .test_si(r_sdischg[7]), .test_se(test_se) );
  glreg_a0_24 u0_idac_shift ( .clk(clk), .arstz(n7), .we(r_cvcwr[4]), .wdat(
        wdat), .rdat(r_idacsh), .test_si(r_cvofs[15]), .test_se(test_se) );
  glreg_a0_23 u0_cv_ofsx ( .clk(clk), .arstz(n6), .we(r_cvcwr[5]), .wdat(wdat), 
        .rdat(r_cvofsx), .test_si(sdischg_duty), .test_se(test_se) );
  glreg_a0_22 u0_cvofs01 ( .clk(clk), .arstz(n5), .we(r_cvcwr[0]), .wdat(wdat), 
        .rdat(r_cvofs[7:0]), .test_si(r_cvofsx[7]), .test_se(test_se) );
  glreg_a0_21 u0_cvofs23 ( .clk(clk), .arstz(n4), .we(r_cvcwr[1]), .wdat(wdat), 
        .rdat(r_cvofs[15:8]), .test_si(r_cvofs[7]), .test_se(test_se) );
  glreg_a0_20 u0_sdischg ( .clk(clk), .arstz(n2), .we(r_cvcwr[2]), .wdat(wdat), 
        .rdat(r_sdischg), .test_si(r_idacsh[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_cvctl_a0 clk_gate_sdischg_cnt_reg ( .CLK(clk_100k), 
        .EN(N115), .ENCLK(net9357), .TE(test_se) );
  cvctl_a0_DW01_sub_1 sub_2_root_sub_0_root_add_46_3 ( .A(r_fw_pwrv), .B({1'b0, 
        1'b0, 1'b0, 1'b0, r_idacsh}), .CI(1'b0), .DIFF({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .CO() );
  cvctl_a0_DW01_add_2 add_1_root_sub_0_root_add_46_3 ( .A({r_cvofsx[7], 
        r_cvofsx[7], r_cvofsx[7], r_cvofsx[7], r_cvofsx}), .B({1'b0, 1'b0, 
        1'b0, N68, N67, N66, N65, N64, N63, N62, N61, N60}), .CI(1'b0), .SUM({
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}), .CO() );
  cvctl_a0_DW01_add_1 add_0_root_sub_0_root_add_46_3 ( .A({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .B({N83, N82, N81, N80, N79, 
        N78, N77, N76, N75, N74, N73, N72}), .CI(1'b0), .SUM({N84, cv_code, 
        r_dac0[0]}), .CO() );
  FAD1X1 add_62_U1_1 ( .A(N95), .B(N107), .CI(add_62_carry_1_), .CO(
        add_62_carry_2_), .SO(r_dac3[1]) );
  FAD1X1 add_62_U1_2 ( .A(N96), .B(N108), .CI(add_62_carry_2_), .CO(
        add_62_carry_3_), .SO(r_dac3[2]) );
  FAD1X1 add_62_U1_3 ( .A(N97), .B(N109), .CI(add_62_carry_3_), .CO(
        add_62_carry_4_), .SO(r_dac3[3]) );
  SDFFRQX1 sdischg_cnt_reg_0_ ( .D(N126), .SIN(div20_cnt[4]), .SMC(test_se), 
        .C(net9357), .XR(srstz), .Q(sdischg_cnt[0]) );
  SDFFRQX1 sdischg_cnt_reg_4_ ( .D(N130), .SIN(sdischg_cnt[3]), .SMC(test_se), 
        .C(net9357), .XR(n6), .Q(sdischg_cnt[4]) );
  SDFFRQX1 sdischg_cnt_reg_1_ ( .D(N127), .SIN(sdischg_cnt[0]), .SMC(test_se), 
        .C(net9357), .XR(srstz), .Q(sdischg_cnt[1]) );
  SDFFRQX1 sdischg_cnt_reg_2_ ( .D(N128), .SIN(sdischg_cnt[1]), .SMC(test_se), 
        .C(net9357), .XR(n4), .Q(sdischg_cnt[2]) );
  SDFFRQX1 div20_cnt_reg_2_ ( .D(N40), .SIN(div20_cnt[1]), .SMC(test_se), .C(
        clk_100k), .XR(n2), .Q(div20_cnt[2]) );
  SDFFRQX1 div20_cnt_reg_1_ ( .D(N39), .SIN(div20_cnt[0]), .SMC(test_se), .C(
        clk_100k), .XR(n5), .Q(div20_cnt[1]) );
  SDFFRQX1 div20_cnt_reg_3_ ( .D(N41), .SIN(div20_cnt[2]), .SMC(test_se), .C(
        clk_100k), .XR(n4), .Q(div20_cnt[3]) );
  SDFFRQX1 div20_cnt_reg_0_ ( .D(N38), .SIN(clk_5k), .SMC(test_se), .C(
        clk_100k), .XR(n8), .Q(div20_cnt[0]) );
  SDFFRQX1 div20_cnt_reg_4_ ( .D(N42), .SIN(div20_cnt[3]), .SMC(test_se), .C(
        clk_100k), .XR(n8), .Q(div20_cnt[4]) );
  SDFFRQX1 sdischg_cnt_reg_3_ ( .D(N129), .SIN(sdischg_cnt[2]), .SMC(test_se), 
        .C(net9357), .XR(n6), .Q(sdischg_cnt[3]) );
  SDFFRQX1 sdischg_reg ( .D(n81), .SIN(sdischg_cnt[4]), .SMC(test_se), .C(
        net9357), .XR(n7), .Q(sdischg_duty) );
  SDFFRQX1 clk_5k_reg ( .D(N29), .SIN(test_si), .SMC(test_se), .C(clk_100k), 
        .XR(n5), .Q(clk_5k) );
  INVX1 U11 ( .A(N84), .Y(n3) );
  INVX1 U14 ( .A(N98), .Y(n12) );
  NOR2X1 U19 ( .A(n26), .B(n52), .Y(n50) );
  NOR2X1 U20 ( .A(n72), .B(r_dac0[10]), .Y(n75) );
  NOR2X1 U21 ( .A(n76), .B(r_dac0[9]), .Y(n73) );
  INVX1 U22 ( .A(n76), .Y(r_dac0[10]) );
  NOR2X1 U23 ( .A(n23), .B(cv_code[1]), .Y(N94) );
  NOR2X1 U24 ( .A(n51), .B(n23), .Y(N98) );
  XNOR2XL U25 ( .A(cv_code[5]), .B(n50), .Y(n51) );
  NAND2X1 U26 ( .A(n28), .B(n23), .Y(r_dac0[1]) );
  NAND2X1 U27 ( .A(n27), .B(n23), .Y(r_dac0[2]) );
  NAND2X1 U28 ( .A(n26), .B(n3), .Y(r_dac0[4]) );
  NAND2X1 U29 ( .A(n25), .B(n3), .Y(r_dac0[6]) );
  INVX1 U30 ( .A(cv_code[6]), .Y(n25) );
  INVX1 U31 ( .A(cv_code[2]), .Y(n27) );
  INVX1 U32 ( .A(cv_code[4]), .Y(n26) );
  XNOR2XL U33 ( .A(cv_code[2]), .B(cv_code[1]), .Y(n55) );
  NAND3X1 U34 ( .A(cv_code[2]), .B(cv_code[1]), .C(cv_code[3]), .Y(n52) );
  NAND2X1 U35 ( .A(cv_code[5]), .B(n50), .Y(n49) );
  INVX1 U36 ( .A(cv_code[1]), .Y(n28) );
  INVX1 U37 ( .A(N84), .Y(n23) );
  NOR2X1 U38 ( .A(N84), .B(cv_code[10]), .Y(n76) );
  NAND21X1 U39 ( .B(cv_code[9]), .A(n23), .Y(r_dac0[9]) );
  XOR2X1 U40 ( .A(add_62_carry_4_), .B(N98), .Y(r_dac3[4]) );
  XOR2X1 U41 ( .A(N99), .B(add_62_carry_5_), .Y(r_dac3[5]) );
  NOR2X1 U42 ( .A(n48), .B(n23), .Y(N99) );
  NOR21XL U43 ( .B(add_62_carry_4_), .A(n12), .Y(add_62_carry_5_) );
  XNOR2XL U44 ( .A(n49), .B(n25), .Y(n48) );
  OAI21BBX1 U45 ( .A(cv_code[10]), .B(cv_code[9]), .C(n23), .Y(n74) );
  INVX1 U46 ( .A(N106), .Y(n17) );
  NOR2X1 U47 ( .A(r_dac0[10]), .B(cv_code[9]), .Y(n72) );
  NOR3XL U48 ( .A(n30), .B(n58), .C(n29), .Y(n56) );
  XOR2X1 U49 ( .A(N94), .B(N106), .Y(r_dac3[0]) );
  OR2X1 U50 ( .A(cv_code[3]), .B(N84), .Y(r_dac0[3]) );
  OR2X1 U51 ( .A(cv_code[5]), .B(N84), .Y(r_dac0[5]) );
  OR2X1 U52 ( .A(cv_code[8]), .B(N84), .Y(r_dac0[8]) );
  OR2X1 U53 ( .A(cv_code[7]), .B(N84), .Y(r_dac0[7]) );
  NOR21XL U54 ( .B(N35), .A(n62), .Y(N40) );
  NOR21XL U55 ( .B(N36), .A(n62), .Y(N41) );
  NOR21XL U56 ( .B(N34), .A(n62), .Y(N39) );
  INVX1 U57 ( .A(n37), .Y(n19) );
  NOR21XL U58 ( .B(N123), .A(n37), .Y(N129) );
  NOR21XL U59 ( .B(N122), .A(n37), .Y(N128) );
  NOR21XL U60 ( .B(N121), .A(n37), .Y(N127) );
  NOR2X1 U61 ( .A(n53), .B(n23), .Y(N97) );
  AO2222XL U62 ( .A(r_cvofs[7]), .B(n72), .C(r_cvofs[15]), .D(n73), .E(
        r_cvofs[14]), .F(n74), .G(r_cvofs[6]), .H(n75), .Y(N109) );
  XNOR2XL U63 ( .A(n52), .B(n26), .Y(n53) );
  XOR2X1 U64 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .Y(N62) );
  XNOR2XL U65 ( .A(r_vcomp[3]), .B(n60), .Y(N63) );
  NAND2X1 U66 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .Y(n60) );
  XNOR2XL U67 ( .A(r_vcomp[4]), .B(n58), .Y(N64) );
  XNOR2XL U68 ( .A(n59), .B(n29), .Y(N65) );
  NOR2X1 U69 ( .A(n58), .B(n30), .Y(n59) );
  XOR2X1 U70 ( .A(n56), .B(r_vcomp[6]), .Y(N66) );
  XNOR2XL U71 ( .A(r_vcomp[7]), .B(n57), .Y(N67) );
  NAND2X1 U72 ( .A(r_vcomp[6]), .B(n56), .Y(n57) );
  GEN2XL U73 ( .D(N84), .E(n27), .C(N94), .B(cv_code[3]), .A(n54), .Y(N96) );
  AO2222XL U74 ( .A(r_cvofs[2]), .B(n72), .C(r_cvofs[10]), .D(n73), .E(
        r_cvofs[13]), .F(n74), .G(r_cvofs[5]), .H(n75), .Y(N108) );
  NOR4XL U75 ( .A(cv_code[3]), .B(n28), .C(n27), .D(n23), .Y(n54) );
  NOR32XL U76 ( .B(r_hlsb_en), .C(clk_5k), .A(r_hlsb_sel), .Y(N47) );
  NOR21XL U77 ( .B(r_vcomp[0]), .A(n47), .Y(
        add_3_root_sub_0_root_add_46_3_carry[1]) );
  AND3X1 U78 ( .A(r_vcomp[7]), .B(n56), .C(r_vcomp[6]), .Y(N68) );
  AO2222XL U79 ( .A(r_cvofs[0]), .B(n72), .C(r_cvofs[8]), .D(n73), .E(
        r_cvofs[11]), .F(n74), .G(r_cvofs[3]), .H(n75), .Y(N106) );
  NOR2X1 U80 ( .A(n55), .B(n23), .Y(N95) );
  AO2222XL U81 ( .A(r_cvofs[1]), .B(n72), .C(r_cvofs[9]), .D(n73), .E(
        r_cvofs[12]), .F(n74), .G(r_cvofs[4]), .H(n75), .Y(N107) );
  NOR21XL U82 ( .B(N94), .A(n17), .Y(add_62_carry_1_) );
  XNOR2XL U83 ( .A(r_vcomp[0]), .B(n47), .Y(N60) );
  NAND3X1 U84 ( .A(r_hlsb_en), .B(clk_5k), .C(r_hlsb_sel), .Y(n47) );
  NAND3X1 U85 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .C(r_vcomp[3]), .Y(n58) );
  INVX1 U86 ( .A(r_vcomp[4]), .Y(n30) );
  INVX1 U87 ( .A(r_vcomp[5]), .Y(n29) );
  NOR21XL U88 ( .B(sdischg_cnt[3]), .A(r_sdischg[3]), .Y(n46) );
  OAI32X1 U89 ( .A(n22), .B(sdischg_cnt[2]), .C(n46), .D(sdischg_cnt[3]), .E(
        n21), .Y(n44) );
  INVX1 U90 ( .A(r_sdischg[3]), .Y(n21) );
  AO222X1 U91 ( .A(n34), .B(n19), .C(n35), .D(n36), .E(sdischg_duty), .F(n37), 
        .Y(n81) );
  AOI22BXL U92 ( .B(N126), .A(n38), .D(r_sdischg[1]), .C(sdischg_cnt[1]), .Y(
        n35) );
  OAI22AX1 U93 ( .D(n36), .C(n43), .A(sdischg_cnt[4]), .B(n20), .Y(n34) );
  EORX1 U94 ( .A(n20), .B(sdischg_cnt[4]), .C(n45), .D(n44), .Y(n36) );
  AOI21X1 U95 ( .B(sdischg_cnt[2]), .C(n22), .A(n46), .Y(n45) );
  AOI21BX1 U96 ( .C(sdischg_cnt[1]), .B(r_sdischg[1]), .A(n44), .Y(n43) );
  OAI221X1 U97 ( .A(n63), .B(n18), .C(n64), .D(n33), .E(r_hlsb_en), .Y(n62) );
  INVX1 U98 ( .A(r_hlsb_freq), .Y(n18) );
  AOI211X1 U99 ( .C(div20_cnt[1]), .D(div20_cnt[0]), .A(div20_cnt[3]), .B(
        div20_cnt[2]), .Y(n64) );
  AOI21X1 U100 ( .B(div20_cnt[0]), .C(div20_cnt[3]), .A(n65), .Y(n63) );
  NOR2X1 U101 ( .A(r_sdischg[6]), .B(r_sdischg[5]), .Y(n37) );
  NAND2X1 U102 ( .A(n33), .B(n68), .Y(n65) );
  OAI21X1 U103 ( .B(div20_cnt[1]), .C(div20_cnt[2]), .A(div20_cnt[3]), .Y(n68)
         );
  INVX1 U104 ( .A(div20_cnt[4]), .Y(n33) );
  INVX1 U105 ( .A(r_sdischg[4]), .Y(n20) );
  NOR2X1 U106 ( .A(n37), .B(sdischg_cnt[0]), .Y(N126) );
  INVX1 U107 ( .A(r_sdischg[2]), .Y(n22) );
  NAND2X1 U108 ( .A(r_sdischg[0]), .B(n19), .Y(n38) );
  NOR2X1 U109 ( .A(n61), .B(n62), .Y(N42) );
  XNOR2XL U110 ( .A(div20_cnt[4]), .B(add_41_carry[4]), .Y(n61) );
  NOR2X1 U111 ( .A(div20_cnt[0]), .B(n62), .Y(N38) );
  NOR2X1 U112 ( .A(n37), .B(n70), .Y(N130) );
  XNOR2XL U113 ( .A(sdischg_cnt[4]), .B(add_81_carry[4]), .Y(n70) );
  OAI21BX1 U114 ( .C(n69), .B(div20_cnt[3]), .A(r_hlsb_freq), .Y(n66) );
  OAI31XL U115 ( .A(div20_cnt[1]), .B(r_hlsb_duty), .C(div20_cnt[0]), .D(
        div20_cnt[2]), .Y(n69) );
  AOI31X1 U116 ( .A(n66), .B(n67), .C(n32), .D(n31), .Y(N29) );
  INVX1 U117 ( .A(r_hlsb_en), .Y(n31) );
  NAND3X1 U118 ( .A(div20_cnt[0]), .B(div20_cnt[3]), .C(r_hlsb_duty), .Y(n67)
         );
  INVX1 U119 ( .A(n65), .Y(n32) );
  NAND42X1 U120 ( .C(sdischg_cnt[0]), .D(sdischg_cnt[1]), .A(n37), .B(n71), 
        .Y(N115) );
  NOR3XL U121 ( .A(sdischg_cnt[2]), .B(sdischg_cnt[4]), .C(sdischg_cnt[3]), 
        .Y(n71) );
endmodule


module cvctl_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module cvctl_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  XOR2X1 U2 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U4 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  XOR2X1 U5 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U6 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  AND2X1 U7 ( .A(carry[10]), .B(A[10]), .Y(carry[11]) );
endmodule


module cvctl_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n11, n12, n13, n14, n15, n16, n17, n18, n19;
  wire   [10:1] carry;

  FAD1X1 U2_7 ( .A(A[7]), .B(n18), .CI(carry[7]), .CO(carry[8]), .SO(DIFF[7])
         );
  FAD1X1 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR2X1 U1 ( .A(n1), .B(A[11]), .Y(DIFF[11]) );
  NOR2X1 U2 ( .A(A[10]), .B(carry[10]), .Y(n1) );
  XNOR2XL U3 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2XL U4 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2XL U5 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  INVX1 U6 ( .A(B[2]), .Y(n15) );
  INVX1 U7 ( .A(B[3]), .Y(n14) );
  INVX1 U8 ( .A(B[4]), .Y(n13) );
  INVX1 U9 ( .A(B[5]), .Y(n12) );
  INVX1 U10 ( .A(B[6]), .Y(n11) );
  INVX1 U11 ( .A(B[1]), .Y(n16) );
  NAND21X1 U12 ( .B(n17), .A(n19), .Y(carry[1]) );
  INVX1 U13 ( .A(A[0]), .Y(n19) );
  INVX1 U14 ( .A(B[7]), .Y(n18) );
  XNOR2XL U15 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  OR2X1 U16 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  INVX1 U17 ( .A(B[0]), .Y(n17) );
  OR2X1 U18 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_cvctl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_20 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9375;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_20 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9375), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9375), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9375), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9375), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9375), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9375), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9375), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9375), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9375), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_21 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9393;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_21 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9393), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9393), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9393), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9393), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9393), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9393), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9393), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9393), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9393), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_22 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9411;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_22 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9411), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9411), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9411), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9411), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9411), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9411), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9411), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9411), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9411), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_23 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9429;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_23 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9429), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9429), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9429), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9429), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9429), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9429), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9429), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9429), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9429), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_24 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9447;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_24 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9447), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9447), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9447), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9447), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9447), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9447), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9447), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9447), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9447), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_25 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9465;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_25 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9465), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9465), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9465), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9465), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9465), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9465), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9465), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9465), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9465), 
        .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcp_a0 ( dp_comp, dm_comp, id_comp, intr, tx_en, tx_dat, r_dat, r_sta, 
        r_ctl, r_msk, r_crc, r_acc, r_dpdmsta, r_wdat, r_wr, r_re, clk, srstz, 
        r_tui, test_si, test_so, test_se );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  output [7:0] r_crc;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input [7:0] r_wdat;
  input [6:0] r_wr;
  output [7:0] r_tui;
  input dp_comp, dm_comp, id_comp, r_re, clk, srstz, test_si, test_se;
  output intr, tx_en, tx_dat, test_so;
  wire   r_dm, r_dmchg, r_acc_int, r_wr_last, r_wr_other, n2, n3, n1, n4;

  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(srstz), .Y(n3) );
  dpdmacc_a0 u0_dpdmacc ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(
        id_comp), .r_re_0(r_re), .r_wr_1(r_wr[6]), .r_wdat(r_wdat), .r_acc(
        r_acc), .r_dpdmsta(r_dpdmsta), .r_dm(r_dm), .r_dmchg(r_dmchg), .r_int(
        r_acc_int), .clk(clk), .rstz(srstz), .test_si(test_si), .test_se(
        test_se) );
  fcpegn_a0 u0_fcpegn ( .intr(intr), .tx_en(tx_en), .tx_dat(tx_dat), .r_dat(
        r_dat), .r_sta(r_sta), .r_ctl(r_ctl), .r_msk(r_msk), .r_wr(r_wr[4:0]), 
        .r_wdat(r_wdat), .ff_idn(n4), .ff_chg(n1), .r_acc_int(r_acc_int), 
        .clk(clk), .srstz(n2), .r_tui(r_tui), .test_si(r_crc[7]), .test_so(
        test_so), .test_se(test_se) );
  fcpcrc_a0 u0_fcpcrc ( .tx_crc(r_crc), .crc_din(r_wdat), .crc_en(r_ctl[2]), 
        .crc_shfi(r_wr_other), .crc_shfl(r_wr_last), .clk(clk), .srstz(n2), 
        .test_si(r_dpdmsta[5]), .test_se(test_se) );
  BUFX3 U1 ( .A(r_dmchg), .Y(n1) );
  BUFX3 U4 ( .A(r_dm), .Y(n4) );
  AND2X1 U5 ( .A(r_wr[5]), .B(r_ctl[3]), .Y(r_wr_last) );
  NOR21XL U6 ( .B(r_wr[5]), .A(r_ctl[3]), .Y(r_wr_other) );
endmodule


module fcpcrc_a0 ( tx_crc, crc_din, crc_en, crc_shfi, crc_shfl, clk, srstz, 
        test_si, test_se );
  output [7:0] tx_crc;
  input [7:0] crc_din;
  input crc_en, crc_shfi, crc_shfl, clk, srstz, test_si, test_se;
  wire   N81, N82, N83, N84, N85, N86, N87, N88, N89, net9483, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n1, n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 clk_gate_crc8_r_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net9483), .TE(test_se) );
  SDFFRQX1 crc8_r_reg_6_ ( .D(N88), .SIN(tx_crc[5]), .SMC(test_se), .C(net9483), .XR(srstz), .Q(tx_crc[6]) );
  SDFFRQX1 crc8_r_reg_7_ ( .D(N89), .SIN(tx_crc[6]), .SMC(test_se), .C(net9483), .XR(srstz), .Q(tx_crc[7]) );
  SDFFRQX1 crc8_r_reg_4_ ( .D(N86), .SIN(tx_crc[3]), .SMC(test_se), .C(net9483), .XR(srstz), .Q(tx_crc[4]) );
  SDFFRQX1 crc8_r_reg_5_ ( .D(N87), .SIN(tx_crc[4]), .SMC(test_se), .C(net9483), .XR(srstz), .Q(tx_crc[5]) );
  SDFFRQX1 crc8_r_reg_3_ ( .D(N85), .SIN(tx_crc[2]), .SMC(test_se), .C(net9483), .XR(srstz), .Q(tx_crc[3]) );
  SDFFRQX1 crc8_r_reg_2_ ( .D(N84), .SIN(tx_crc[1]), .SMC(test_se), .C(net9483), .XR(srstz), .Q(tx_crc[2]) );
  SDFFRQX1 crc8_r_reg_1_ ( .D(N83), .SIN(tx_crc[0]), .SMC(test_se), .C(net9483), .XR(srstz), .Q(tx_crc[1]) );
  SDFFRQX1 crc8_r_reg_0_ ( .D(N82), .SIN(test_si), .SMC(test_se), .C(net9483), 
        .XR(srstz), .Q(tx_crc[0]) );
  XNOR2XL U3 ( .A(n16), .B(n25), .Y(n10) );
  XNOR2XL U4 ( .A(n30), .B(n26), .Y(n16) );
  XNOR2XL U5 ( .A(n3), .B(n29), .Y(n11) );
  XNOR2XL U6 ( .A(n30), .B(n28), .Y(n29) );
  XOR2X1 U7 ( .A(n21), .B(n11), .Y(n14) );
  XNOR2XL U8 ( .A(n22), .B(n2), .Y(n25) );
  XNOR2XL U9 ( .A(n2), .B(n12), .Y(n30) );
  XNOR2XL U10 ( .A(n37), .B(n36), .Y(n20) );
  XNOR2XL U11 ( .A(n10), .B(n17), .Y(n37) );
  OAI22X1 U12 ( .A(n26), .B(n9), .C(n27), .D(n5), .Y(N85) );
  XOR2X1 U13 ( .A(n20), .B(n16), .Y(n27) );
  OAI22X1 U14 ( .A(n17), .B(n9), .C(n18), .D(n5), .Y(N87) );
  XNOR2XL U15 ( .A(n19), .B(n20), .Y(n18) );
  XNOR2XL U16 ( .A(n14), .B(n3), .Y(n19) );
  OAI22X1 U17 ( .A(n22), .B(n9), .C(n23), .D(n5), .Y(N86) );
  XOR2X1 U18 ( .A(n20), .B(n24), .Y(n23) );
  XNOR2XL U19 ( .A(n21), .B(n25), .Y(n24) );
  XNOR2XL U20 ( .A(n33), .B(n34), .Y(n21) );
  XNOR2XL U21 ( .A(n3), .B(n12), .Y(n33) );
  XNOR2XL U22 ( .A(n25), .B(n32), .Y(n34) );
  XOR2X1 U23 ( .A(n40), .B(n41), .Y(n22) );
  XNOR2XL U24 ( .A(crc_din[4]), .B(n42), .Y(n41) );
  OAI32X1 U25 ( .A(n5), .B(n6), .C(n2), .D(n7), .E(n8), .Y(N89) );
  OA21X1 U26 ( .B(n1), .C(n5), .A(n9), .Y(n7) );
  INVX1 U27 ( .A(n6), .Y(n1) );
  XNOR2XL U28 ( .A(n10), .B(n11), .Y(n6) );
  INVX1 U29 ( .A(n8), .Y(n2) );
  OAI22X1 U30 ( .A(n36), .B(n9), .C(n20), .D(n5), .Y(N82) );
  OAI22X1 U31 ( .A(n32), .B(n9), .C(n21), .D(n5), .Y(N83) );
  OAI22X1 U32 ( .A(n28), .B(n9), .C(n11), .D(n5), .Y(N84) );
  OAI22X1 U33 ( .A(n12), .B(n9), .C(n13), .D(n5), .Y(N88) );
  XNOR2XL U34 ( .A(n14), .B(n15), .Y(n13) );
  XNOR2XL U35 ( .A(n16), .B(n12), .Y(n15) );
  XNOR2XL U36 ( .A(n43), .B(n44), .Y(n26) );
  XNOR2XL U37 ( .A(crc_din[3]), .B(n45), .Y(n44) );
  INVX1 U38 ( .A(n17), .Y(n3) );
  XNOR2XL U39 ( .A(crc_din[2]), .B(n31), .Y(n28) );
  XNOR2XL U40 ( .A(crc_din[1]), .B(n35), .Y(n32) );
  XNOR2XL U41 ( .A(crc_din[0]), .B(n43), .Y(n36) );
  XOR2X1 U42 ( .A(n45), .B(n42), .Y(n53) );
  XNOR2XL U43 ( .A(n43), .B(n35), .Y(n40) );
  XNOR2XL U44 ( .A(n46), .B(n47), .Y(n12) );
  XNOR2XL U45 ( .A(n35), .B(n45), .Y(n47) );
  XNOR2XL U46 ( .A(n31), .B(n50), .Y(n46) );
  XNOR2XL U47 ( .A(tx_crc[6]), .B(crc_din[6]), .Y(n50) );
  NAND21X1 U48 ( .B(crc_shfl), .A(crc_en), .Y(n9) );
  XNOR2XL U49 ( .A(n51), .B(n52), .Y(n8) );
  XNOR2XL U50 ( .A(n53), .B(n31), .Y(n51) );
  XNOR2XL U51 ( .A(tx_crc[7]), .B(crc_din[7]), .Y(n52) );
  NAND2X1 U52 ( .A(crc_shfl), .B(crc_en), .Y(n5) );
  OR2X1 U53 ( .A(crc_shfi), .B(n9), .Y(N81) );
  XNOR2XL U54 ( .A(n38), .B(n39), .Y(n17) );
  XOR2X1 U55 ( .A(n40), .B(n31), .Y(n38) );
  XNOR2XL U56 ( .A(tx_crc[5]), .B(crc_din[5]), .Y(n39) );
  XOR2X1 U57 ( .A(n53), .B(n56), .Y(n43) );
  XNOR2XL U58 ( .A(tx_crc[0]), .B(n4), .Y(n56) );
  XNOR2XL U59 ( .A(tx_crc[3]), .B(n55), .Y(n45) );
  XOR2X1 U60 ( .A(tx_crc[7]), .B(tx_crc[6]), .Y(n55) );
  XNOR2XL U61 ( .A(n54), .B(n55), .Y(n31) );
  XNOR2XL U62 ( .A(tx_crc[5]), .B(tx_crc[2]), .Y(n54) );
  XOR2X1 U63 ( .A(n48), .B(n49), .Y(n35) );
  XNOR2XL U64 ( .A(n4), .B(tx_crc[6]), .Y(n48) );
  XNOR2XL U65 ( .A(tx_crc[1]), .B(n42), .Y(n49) );
  XNOR2XL U66 ( .A(tx_crc[7]), .B(tx_crc[4]), .Y(n42) );
  INVX1 U67 ( .A(tx_crc[5]), .Y(n4) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcpegn_a0 ( intr, tx_en, tx_dat, r_dat, r_sta, r_ctl, r_msk, r_wr, 
        r_wdat, ff_idn, ff_chg, r_acc_int, clk, srstz, r_tui, test_si, test_so, 
        test_se );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  input [4:0] r_wr;
  input [7:0] r_wdat;
  output [7:0] r_tui;
  input ff_idn, ff_chg, r_acc_int, clk, srstz, test_si, test_se;
  output intr, tx_en, tx_dat, test_so;
  wire   N22, upd_dbuf_en, us_cnt_2_, us_cnt_1_, us_cnt_0_, N85, N87, N88,
         N141, N142, N144, N145, N172, N173, adp_tx_ui_7_, adp_tx_ui_6_, N205,
         N221, N222, N223, N224, N225, N226, N227, N228, N260, N261, N348,
         N349, N356, N362, N363, N444, rx_trans_8_chg, N1005, N1006, N1007,
         N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1043,
         net9505, net9509, net9512, net9513, net9514, net9515, net9516,
         net9517, net9520, net9523, net9528, net9533, net9538, n26, n27, n28,
         n29, n30, n31, n32, n516, n525, N1259, N1258, N1257, N1256, N1255,
         N1254, N1253, N1252, N161, N160, N159, N108, N107, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n506, n509, n2, n80, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n508,
         n510, n511, n512, n513, n514, n515, n517, n518, n519, n520, n521,
         n522, n523, n524, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n18, n19, n20, n21, n22, n23, n24, n25,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3;
  wire   [6:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;
  wire   [7:0] upd_dbuf;
  wire   [10:0] rxtx_buf;
  wire   [4:1] rx_ui_3_8;
  wire   [4:1] rx_ui_5_8;
  wire   [5:0] catch_sync;
  wire   [7:0] ui_intv_cnt;
  wire   [6:2] symb_cnt;
  wire   [6:0] adp_tx_1_4;
  wire   [7:0] tui_wdat;
  wire   [11:0] trans_buf;
  wire   [1:0] new_rx_sync_cnt;
  wire   [3:0] fcp_state;
  wire   [5:1] add_264_carry;
  wire   [5:1] add_263_carry;
  wire   [8:6] add_274_2_carry;
  wire   [8:6] add_274_carry;

  FAD1X1 add_264_U1_1 ( .A(n69), .B(n66), .CI(add_264_carry[1]), .CO(
        add_264_carry[2]), .SO(rx_ui_5_8[1]) );
  FAD1X1 add_264_U1_2 ( .A(n67), .B(n65), .CI(add_264_carry[2]), .CO(
        add_264_carry[3]), .SO(rx_ui_5_8[2]) );
  FAD1X1 add_264_U1_3 ( .A(n66), .B(n61), .CI(add_264_carry[3]), .CO(
        add_264_carry[4]), .SO(rx_ui_5_8[3]) );
  FAD1X1 add_264_U1_4 ( .A(n65), .B(n63), .CI(add_264_carry[4]), .CO(
        add_264_carry[5]), .SO(rx_ui_5_8[4]) );
  FAD1X1 add_263_U1_1 ( .A(n67), .B(n66), .CI(add_263_carry[1]), .CO(
        add_263_carry[2]), .SO(rx_ui_3_8[1]) );
  FAD1X1 add_263_U1_2 ( .A(n66), .B(n65), .CI(add_263_carry[2]), .CO(
        add_263_carry[3]), .SO(rx_ui_3_8[2]) );
  FAD1X1 add_263_U1_3 ( .A(n65), .B(n61), .CI(add_263_carry[3]), .CO(
        add_263_carry[4]), .SO(rx_ui_3_8[3]) );
  FAD1X1 add_263_U1_4 ( .A(n61), .B(n63), .CI(add_263_carry[4]), .CO(
        add_263_carry[5]), .SO(rx_ui_3_8[4]) );
  FAD1X1 add_274_2_U1_6 ( .A(N160), .B(ui_intv_cnt[6]), .CI(add_274_2_carry[6]), .CO(add_274_2_carry[7]), .SO(N172) );
  FAD1X1 add_274_2_U1_7 ( .A(N161), .B(ui_intv_cnt[7]), .CI(add_274_2_carry[7]), .CO(add_274_2_carry[8]), .SO(N173) );
  FAD1X1 add_274_U1_6 ( .A(N107), .B(ui_intv_cnt[6]), .CI(add_274_carry[6]), 
        .CO(add_274_carry[7]), .SO(N144) );
  FAD1X1 add_274_U1_7 ( .A(N108), .B(ui_intv_cnt[7]), .CI(add_274_carry[7]), 
        .CO(add_274_carry[8]), .SO(N145) );
  INVX1 U26 ( .A(n56), .Y(n51) );
  INVX1 U27 ( .A(n56), .Y(n52) );
  INVX1 U28 ( .A(n56), .Y(n53) );
  INVX1 U29 ( .A(n56), .Y(n54) );
  INVX1 U30 ( .A(n56), .Y(n55) );
  INVX1 U31 ( .A(n56), .Y(n50) );
  INVX1 U32 ( .A(n56), .Y(n48) );
  INVX1 U33 ( .A(n56), .Y(n49) );
  INVX1 U34 ( .A(n56), .Y(n47) );
  INVX1 U35 ( .A(srstz), .Y(n56) );
  glreg_8_00000000 u0_fcpctl ( .clk(clk), .arstz(n51), .we(r_wr[0]), .wdat({
        n34, r_wdat[6:3], n21, r_wdat[1:0]}), .rdat({n509, 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, r_ctl[4:0]}), 
        .test_si(r_ctl[7]), .test_se(test_se) );
  glsta_a0_0 u0_fcpsta ( .clk(clk), .arstz(n50), .rst0(1'b0), .set2({r_acc_int, 
        setsta[6:5], n539, setsta[3], n525, n2, setsta[0]}), .clr1(clrsta), 
        .rdat(r_sta), .irq(r_irq), .test_si(r_msk[7]), .test_se(test_se) );
  glreg_a0_4 u0_fcpmsk ( .clk(clk), .arstz(n49), .we(r_wr[2]), .wdat({n34, 
        r_wdat[6:3], n21, r_wdat[1:0]}), .rdat(r_msk), .test_si(r_dat[7]), 
        .test_se(test_se) );
  glreg_a0_3 u0_fcpdat ( .clk(clk), .arstz(n48), .we(upd_dbuf_en), .wdat(
        upd_dbuf), .rdat(r_dat), .test_si(n509), .test_se(test_se) );
  glreg_a0_2 u0_fcptui ( .clk(clk), .arstz(n47), .we(n80), .wdat(tui_wdat), 
        .rdat(r_tui), .test_si(r_sta[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 clk_gate_catch_sync_reg ( .CLK(clk), .EN(
        n540), .ENCLK(net9505), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 clk_gate_ui_intv_cnt_reg ( .CLK(clk), .EN(
        N205), .ENCLK(net9523), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 clk_gate_rxtx_buf_reg ( .CLK(clk), .EN(N22), 
        .ENCLK(net9528), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 clk_gate_fcp_state_reg ( .CLK(clk), .EN(
        N1005), .ENCLK(net9533), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 clk_gate_symb_cnt_reg ( .CLK(clk), .EN(
        N1043), .ENCLK(net9538), .TE(test_se) );
  fcpegn_a0_DW01_inc_0 r611 ( .A({symb_cnt[6:4], n12, symb_cnt[2], n11, n15}), 
        .SUM({n26, n27, n28, n29, n30, n31, n32}) );
  fcpegn_a0_DW01_inc_1 add_283_round ( .A({1'b0, adp_tx_ui_7_, adp_tx_ui_6_, 
        n71, r_tui[4:1]}), .SUM({adp_tx_1_4, SYNOPSYS_UNCONNECTED_3}) );
  fcpegn_a0_DW01_inc_2 add_316_aco ( .A({N1259, N1258, N1257, N1256, N1255, 
        N1254, N1253, N1252}), .SUM({N228, N227, N226, N225, N224, N223, N222, 
        N221}) );
  SDFFRQX1 rxtx_buf_reg_8_ ( .D(trans_buf[8]), .SIN(rxtx_buf[7]), .SMC(test_se), .C(net9528), .XR(n52), .Q(rxtx_buf[8]) );
  SDFFRQX1 rxtx_buf_reg_10_ ( .D(trans_buf[10]), .SIN(rxtx_buf[9]), .SMC(
        test_se), .C(net9528), .XR(n52), .Q(rxtx_buf[10]) );
  SDFFRQX1 rxtx_buf_reg_9_ ( .D(trans_buf[9]), .SIN(rxtx_buf[8]), .SMC(test_se), .C(net9528), .XR(n52), .Q(rxtx_buf[9]) );
  SDFFRQX1 rxtx_buf_reg_0_ ( .D(trans_buf[0]), .SIN(rx_trans_8_chg), .SMC(
        test_se), .C(net9528), .XR(n53), .Q(rxtx_buf[0]) );
  SDFFRQX1 rxtx_buf_reg_4_ ( .D(trans_buf[4]), .SIN(rxtx_buf[3]), .SMC(test_se), .C(net9528), .XR(n52), .Q(rxtx_buf[4]) );
  SDFFRQX1 rxtx_buf_reg_6_ ( .D(trans_buf[6]), .SIN(rxtx_buf[5]), .SMC(test_se), .C(net9528), .XR(n52), .Q(rxtx_buf[6]) );
  SDFFRQX1 rxtx_buf_reg_7_ ( .D(trans_buf[7]), .SIN(rxtx_buf[6]), .SMC(test_se), .C(net9528), .XR(n52), .Q(rxtx_buf[7]) );
  SDFFRQX1 rxtx_buf_reg_3_ ( .D(trans_buf[3]), .SIN(rxtx_buf[2]), .SMC(test_se), .C(net9528), .XR(n53), .Q(rxtx_buf[3]) );
  SDFFRQX1 rxtx_buf_reg_5_ ( .D(trans_buf[5]), .SIN(rxtx_buf[4]), .SMC(test_se), .C(net9528), .XR(n52), .Q(rxtx_buf[5]) );
  SDFFRQX1 rx_byte_pchk_reg ( .D(N356), .SIN(new_rx_sync_cnt[1]), .SMC(test_se), .C(clk), .XR(n55), .Q(setsta[5]) );
  SDFFRQX1 rxtx_buf_reg_2_ ( .D(trans_buf[2]), .SIN(rxtx_buf[1]), .SMC(test_se), .C(net9528), .XR(n52), .Q(rxtx_buf[2]) );
  SDFFRQX1 rxtx_buf_reg_1_ ( .D(trans_buf[1]), .SIN(rxtx_buf[0]), .SMC(test_se), .C(net9528), .XR(n54), .Q(rxtx_buf[1]) );
  SDFFRQX1 new_rx_sync_cnt_reg_1_ ( .D(N349), .SIN(new_rx_sync_cnt[0]), .SMC(
        test_se), .C(clk), .XR(n49), .Q(new_rx_sync_cnt[1]) );
  SDFFRQX1 new_rx_sync_cnt_reg_0_ ( .D(N348), .SIN(fcp_state[3]), .SMC(test_se), .C(clk), .XR(n47), .Q(new_rx_sync_cnt[0]) );
  SDFFQX1 rx_trans_8_chg_reg ( .D(n516), .SIN(setsta[5]), .SMC(test_se), .C(
        clk), .Q(rx_trans_8_chg) );
  SDFFRQX1 us_cnt_reg_2_ ( .D(N87), .SIN(us_cnt_1_), .SMC(test_se), .C(clk), 
        .XR(n50), .Q(us_cnt_2_) );
  SDFFRQX1 us_cnt_reg_3_ ( .D(N88), .SIN(us_cnt_2_), .SMC(test_se), .C(clk), 
        .XR(srstz), .Q(test_so) );
  SDFFRQX1 us_cnt_reg_1_ ( .D(n506), .SIN(us_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(n48), .Q(us_cnt_1_) );
  SDFFRQX1 us_cnt_reg_0_ ( .D(N85), .SIN(ui_intv_cnt[7]), .SMC(test_se), .C(
        clk), .XR(n52), .Q(us_cnt_0_) );
  SDFFRQX1 ui_intv_cnt_reg_7_ ( .D(net9509), .SIN(ui_intv_cnt[6]), .SMC(
        test_se), .C(net9523), .XR(n54), .Q(ui_intv_cnt[7]) );
  SDFFRQX1 ui_intv_cnt_reg_6_ ( .D(net9512), .SIN(n13), .SMC(test_se), .C(
        net9523), .XR(n54), .Q(ui_intv_cnt[6]) );
  SDFFSQX1 catch_sync_reg_5_ ( .D(n13), .SIN(catch_sync[4]), .SMC(test_se), 
        .C(net9505), .XS(n51), .Q(catch_sync[5]) );
  SDFFRQX1 symb_cnt_reg_6_ ( .D(N1016), .SIN(symb_cnt[5]), .SMC(test_se), .C(
        net9538), .XR(n54), .Q(symb_cnt[6]) );
  SDFFRQX1 symb_cnt_reg_4_ ( .D(N1014), .SIN(n12), .SMC(test_se), .C(net9538), 
        .XR(n55), .Q(symb_cnt[4]) );
  SDFFRQX1 ui_intv_cnt_reg_1_ ( .D(net9517), .SIN(ui_intv_cnt[0]), .SMC(
        test_se), .C(net9523), .XR(n53), .Q(ui_intv_cnt[1]) );
  SDFFRQX1 ui_intv_cnt_reg_0_ ( .D(net9520), .SIN(r_tui[7]), .SMC(test_se), 
        .C(net9523), .XR(n53), .Q(ui_intv_cnt[0]) );
  SDFFRQX1 symb_cnt_reg_5_ ( .D(N1015), .SIN(symb_cnt[4]), .SMC(test_se), .C(
        net9538), .XR(n55), .Q(symb_cnt[5]) );
  SDFFRQX1 ui_intv_cnt_reg_2_ ( .D(net9516), .SIN(ui_intv_cnt[1]), .SMC(
        test_se), .C(net9523), .XR(n53), .Q(ui_intv_cnt[2]) );
  SDFFRQX1 ui_intv_cnt_reg_4_ ( .D(net9514), .SIN(n10), .SMC(test_se), .C(
        net9523), .XR(n54), .Q(N142) );
  SDFFRQX1 ui_intv_cnt_reg_5_ ( .D(net9513), .SIN(N142), .SMC(test_se), .C(
        net9523), .XR(n54), .Q(ui_intv_cnt[5]) );
  SDFFRQX1 ui_intv_cnt_reg_3_ ( .D(net9515), .SIN(ui_intv_cnt[2]), .SMC(
        test_se), .C(net9523), .XR(n53), .Q(N141) );
  SDFFRQX1 catch_sync_reg_4_ ( .D(N142), .SIN(catch_sync[3]), .SMC(test_se), 
        .C(net9505), .XR(n53), .Q(catch_sync[4]) );
  SDFFRQX1 sync_length_reg_1_ ( .D(N261), .SIN(N362), .SMC(test_se), .C(
        net9523), .XR(n54), .Q(N363) );
  SDFFRQX1 sync_length_reg_0_ ( .D(N260), .SIN(symb_cnt[6]), .SMC(test_se), 
        .C(net9523), .XR(n54), .Q(N362) );
  SDFFRQX1 symb_cnt_reg_3_ ( .D(N1013), .SIN(symb_cnt[2]), .SMC(test_se), .C(
        net9538), .XR(n55), .Q(symb_cnt[3]) );
  SDFFSQX1 catch_sync_reg_3_ ( .D(n10), .SIN(catch_sync[2]), .SMC(test_se), 
        .C(net9505), .XS(n51), .Q(catch_sync[3]) );
  SDFFRQX1 catch_sync_reg_0_ ( .D(ui_intv_cnt[0]), .SIN(test_si), .SMC(test_se), .C(net9505), .XR(n53), .Q(catch_sync[0]) );
  SDFFRQX1 catch_sync_reg_2_ ( .D(ui_intv_cnt[2]), .SIN(catch_sync[1]), .SMC(
        test_se), .C(net9505), .XR(n53), .Q(catch_sync[2]) );
  SDFFRQX1 symb_cnt_reg_2_ ( .D(N1012), .SIN(n11), .SMC(test_se), .C(net9538), 
        .XR(n55), .Q(symb_cnt[2]) );
  SDFFRQX1 symb_cnt_reg_1_ ( .D(N1011), .SIN(n15), .SMC(test_se), .C(net9538), 
        .XR(n55), .Q(N160) );
  SDFFRQX1 symb_cnt_reg_0_ ( .D(N1010), .SIN(tx_dat), .SMC(test_se), .C(
        net9538), .XR(n55), .Q(N159) );
  SDFFRQX1 catch_sync_reg_1_ ( .D(ui_intv_cnt[1]), .SIN(catch_sync[0]), .SMC(
        test_se), .C(net9505), .XR(n53), .Q(catch_sync[1]) );
  SDFFSQX1 tx_dbuf_keep_empty_reg ( .D(N444), .SIN(N363), .SMC(test_se), .C(
        clk), .XS(n52), .Q(r_ctl[7]) );
  SDFFRQX1 rxtx_buf_reg_11_ ( .D(trans_buf[11]), .SIN(rxtx_buf[10]), .SMC(
        test_se), .C(net9528), .XR(n54), .Q(tx_dat) );
  SDFFRQX1 fcp_state_reg_2_ ( .D(N1008), .SIN(fcp_state[1]), .SMC(test_se), 
        .C(net9533), .XR(n55), .Q(fcp_state[2]) );
  SDFFRQX1 fcp_state_reg_0_ ( .D(N1006), .SIN(catch_sync[5]), .SMC(test_se), 
        .C(net9533), .XR(n55), .Q(fcp_state[0]) );
  SDFFRQX1 fcp_state_reg_3_ ( .D(N1009), .SIN(fcp_state[2]), .SMC(test_se), 
        .C(net9533), .XR(n54), .Q(fcp_state[3]) );
  SDFFRQX1 fcp_state_reg_1_ ( .D(N1007), .SIN(fcp_state[0]), .SMC(test_se), 
        .C(net9533), .XR(n55), .Q(fcp_state[1]) );
  INVX1 U4 ( .A(n41), .Y(n3) );
  INVX1 U5 ( .A(n106), .Y(n4) );
  BUFX3 U6 ( .A(n108), .Y(n5) );
  INVX1 U7 ( .A(n15), .Y(n6) );
  INVX1 U8 ( .A(n127), .Y(n7) );
  INVX1 U9 ( .A(n258), .Y(n8) );
  INVX1 U10 ( .A(n151), .Y(n9) );
  BUFX3 U11 ( .A(N141), .Y(n10) );
  INVX1 U12 ( .A(n542), .Y(n11) );
  BUFX3 U13 ( .A(symb_cnt[3]), .Y(n12) );
  INVX1 U14 ( .A(n122), .Y(n13) );
  INVX1 U15 ( .A(r_wr[3]), .Y(n14) );
  BUFX3 U16 ( .A(N159), .Y(n15) );
  XNOR2XL U17 ( .A(n184), .B(n185), .Y(n159) );
  OAI222XL U18 ( .A(n275), .B(n117), .C(n314), .D(n315), .E(n75), .F(n295), 
        .Y(n312) );
  AOI22AXL U19 ( .A(n471), .B(n115), .D(n472), .C(N363), .Y(n417) );
  INVX1 U20 ( .A(r_wr[4]), .Y(n81) );
  INVX1 U21 ( .A(n35), .Y(n34) );
  INVX1 U22 ( .A(n22), .Y(n21) );
  INVX1 U23 ( .A(n269), .Y(n79) );
  INVX1 U24 ( .A(n258), .Y(n43) );
  INVX1 U25 ( .A(r_wr[3]), .Y(n78) );
  NOR2X1 U36 ( .A(n25), .B(n77), .Y(clrsta[5]) );
  NOR2X1 U37 ( .A(n20), .B(n77), .Y(clrsta[1]) );
  NOR2X1 U38 ( .A(n24), .B(n77), .Y(clrsta[4]) );
  NOR2X1 U39 ( .A(n19), .B(n77), .Y(clrsta[0]) );
  NOR2X1 U40 ( .A(n33), .B(n77), .Y(clrsta[6]) );
  NOR2X1 U41 ( .A(n22), .B(n77), .Y(clrsta[2]) );
  NOR2X1 U42 ( .A(n35), .B(n77), .Y(clrsta[7]) );
  NOR2X1 U43 ( .A(n23), .B(n77), .Y(clrsta[3]) );
  INVX1 U44 ( .A(r_wdat[4]), .Y(n24) );
  INVX1 U45 ( .A(r_wdat[7]), .Y(n35) );
  INVX1 U46 ( .A(r_wdat[6]), .Y(n33) );
  INVX1 U47 ( .A(r_wdat[3]), .Y(n23) );
  INVX1 U48 ( .A(r_wdat[5]), .Y(n25) );
  INVX1 U49 ( .A(r_wdat[2]), .Y(n22) );
  INVX1 U50 ( .A(r_wdat[1]), .Y(n20) );
  INVX1 U51 ( .A(r_wdat[0]), .Y(n19) );
  INVX1 U52 ( .A(n444), .Y(n113) );
  NAND2X1 U53 ( .A(n553), .B(r_wr[3]), .Y(n269) );
  NAND2X1 U54 ( .A(n269), .B(n347), .Y(n258) );
  INVX1 U55 ( .A(n257), .Y(n42) );
  INVX1 U56 ( .A(r_wr[1]), .Y(n77) );
  OAI221X1 U57 ( .A(n102), .B(n155), .C(n23), .D(n81), .E(n158), .Y(
        tui_wdat[3]) );
  INVX1 U58 ( .A(n159), .Y(n102) );
  OAI221X1 U59 ( .A(n155), .B(n101), .C(n24), .D(n81), .E(n158), .Y(
        tui_wdat[4]) );
  OAI221X1 U60 ( .A(n100), .B(n155), .C(n25), .D(n81), .E(n158), .Y(
        tui_wdat[5]) );
  INVX1 U61 ( .A(rx_ui_3_8[3]), .Y(n59) );
  INVX1 U62 ( .A(n168), .Y(n99) );
  INVX1 U63 ( .A(n173), .Y(n100) );
  INVX1 U64 ( .A(n172), .Y(n101) );
  INVX1 U65 ( .A(n347), .Y(n40) );
  NOR2X1 U66 ( .A(n114), .B(n406), .Y(n444) );
  NAND2X1 U67 ( .A(n159), .B(n160), .Y(n179) );
  INVX1 U68 ( .A(n352), .Y(n546) );
  INVX1 U69 ( .A(n425), .Y(n550) );
  XNOR2XL U70 ( .A(n37), .B(n36), .Y(n268) );
  NAND2X1 U71 ( .A(n254), .B(n258), .Y(n257) );
  OAI21BBX1 U72 ( .A(N221), .B(n88), .C(n280), .Y(net9520) );
  NAND32X1 U73 ( .B(n162), .C(r_wr[4]), .A(n154), .Y(n155) );
  NOR21XL U74 ( .B(N224), .A(n281), .Y(net9515) );
  NOR21XL U75 ( .B(N226), .A(n281), .Y(net9513) );
  NOR21XL U76 ( .B(N223), .A(n281), .Y(net9516) );
  NOR21XL U77 ( .B(N222), .A(n281), .Y(net9517) );
  NAND2X1 U78 ( .A(n280), .B(n88), .Y(n281) );
  OAI222XL U79 ( .A(r_wr[4]), .B(n154), .C(n155), .D(n156), .E(n33), .F(n81), 
        .Y(tui_wdat[6]) );
  XNOR2XL U80 ( .A(n157), .B(n100), .Y(n156) );
  OAI2B11X1 U81 ( .D(n160), .C(n155), .A(n158), .B(n161), .Y(tui_wdat[2]) );
  AOI22AXL U82 ( .A(r_wr[4]), .B(n21), .D(n154), .C(n81), .Y(n161) );
  NAND2X1 U83 ( .A(n162), .B(n81), .Y(n158) );
  XNOR2XL U84 ( .A(n63), .B(add_263_carry[5]), .Y(n461) );
  XNOR2XL U85 ( .A(n177), .B(n176), .Y(n157) );
  AOI21X1 U86 ( .B(n176), .C(n177), .A(n175), .Y(n168) );
  OAI21BBX1 U87 ( .A(n216), .B(n233), .C(n239), .Y(n231) );
  OAI21X1 U88 ( .B(n216), .C(n233), .A(n235), .Y(n239) );
  INVX1 U89 ( .A(n404), .Y(n541) );
  NOR32XL U90 ( .B(n186), .C(n181), .A(n180), .Y(n177) );
  XNOR2XL U91 ( .A(n186), .B(n187), .Y(n173) );
  NOR21XL U92 ( .B(n181), .A(n180), .Y(n187) );
  XNOR2XL U93 ( .A(n180), .B(n181), .Y(n172) );
  XNOR2XL U94 ( .A(n233), .B(n234), .Y(n196) );
  XOR2X1 U95 ( .A(n235), .B(n216), .Y(n234) );
  NAND2X1 U96 ( .A(n45), .B(n276), .Y(n347) );
  INVX1 U97 ( .A(n515), .Y(n93) );
  NOR21XL U98 ( .B(n183), .A(n182), .Y(n185) );
  NAND32X1 U99 ( .B(n184), .C(n182), .A(n183), .Y(n180) );
  XNOR2XL U100 ( .A(n343), .B(n63), .Y(n336) );
  NAND2X1 U101 ( .A(n65), .B(n61), .Y(n343) );
  NOR2X1 U102 ( .A(n404), .B(n380), .Y(n406) );
  NOR2X1 U103 ( .A(n545), .B(n246), .Y(n392) );
  INVX1 U104 ( .A(n325), .Y(n62) );
  INVX1 U105 ( .A(n278), .Y(n2) );
  INVX1 U106 ( .A(n379), .Y(n95) );
  INVX1 U107 ( .A(n349), .Y(n114) );
  INVX1 U108 ( .A(n494), .Y(n45) );
  XNOR2XL U109 ( .A(n182), .B(n183), .Y(n160) );
  NAND21X1 U110 ( .B(n421), .A(n545), .Y(n310) );
  OAI21X1 U111 ( .B(n65), .C(n61), .A(n63), .Y(n321) );
  NOR2X1 U112 ( .A(n547), .B(n549), .Y(n352) );
  NAND2X1 U113 ( .A(n549), .B(n93), .Y(n418) );
  NAND2X1 U114 ( .A(n61), .B(add_264_carry[5]), .Y(n139) );
  INVX1 U115 ( .A(n300), .Y(n547) );
  INVX1 U116 ( .A(n298), .Y(n115) );
  INVX1 U117 ( .A(n295), .Y(n553) );
  INVX1 U118 ( .A(n491), .Y(n110) );
  NOR2X1 U119 ( .A(n496), .B(n497), .Y(n485) );
  INVX1 U120 ( .A(n519), .Y(n126) );
  INVX1 U121 ( .A(n241), .Y(n125) );
  INVX1 U122 ( .A(tx_en), .Y(n548) );
  NAND2X1 U123 ( .A(n492), .B(n493), .Y(n300) );
  NAND2X1 U124 ( .A(n360), .B(n535), .Y(n425) );
  XNOR2XL U125 ( .A(n265), .B(n266), .Y(n262) );
  XNOR2XL U126 ( .A(n270), .B(n271), .Y(n265) );
  XNOR2XL U127 ( .A(n267), .B(n268), .Y(n266) );
  XNOR2XL U128 ( .A(n252), .B(n250), .Y(n271) );
  XNOR2XL U129 ( .A(n253), .B(n255), .Y(n267) );
  XNOR2XL U130 ( .A(n249), .B(n264), .Y(n270) );
  OAI21X1 U131 ( .B(n86), .C(n258), .A(n260), .Y(trans_buf[1]) );
  AOI32X1 U132 ( .A(n42), .B(n261), .C(n262), .D(n251), .E(n37), .Y(n260) );
  INVX1 U133 ( .A(n259), .Y(n37) );
  INVX1 U134 ( .A(n256), .Y(n36) );
  AOI221XL U135 ( .A(n544), .B(n497), .C(n45), .D(n496), .E(n495), .Y(n501) );
  NOR2X1 U136 ( .A(n74), .B(n3), .Y(n254) );
  OAI222XL U137 ( .A(n255), .B(n41), .C(n256), .D(n257), .E(n83), .F(n258), 
        .Y(trans_buf[3]) );
  OAI222XL U138 ( .A(n256), .B(n41), .C(n259), .D(n257), .E(n82), .F(n258), 
        .Y(trans_buf[2]) );
  OAI211X1 U139 ( .C(tx_en), .D(n75), .A(n269), .B(n350), .Y(n283) );
  AOI22X1 U140 ( .A(n264), .B(n251), .C(n39), .D(n254), .Y(n248) );
  NOR2X1 U141 ( .A(n283), .B(n284), .Y(n280) );
  INVX1 U142 ( .A(n251), .Y(n41) );
  INVX1 U143 ( .A(n264), .Y(n39) );
  INVX1 U144 ( .A(n255), .Y(n38) );
  INVX1 U145 ( .A(n495), .Y(n46) );
  NOR21XL U146 ( .B(N228), .A(n281), .Y(net9509) );
  NOR2X1 U147 ( .A(n382), .B(n118), .Y(N1259) );
  OAI22X1 U148 ( .A(r_wr[3]), .B(n82), .C(n78), .D(n20), .Y(upd_dbuf[1]) );
  OAI22X1 U149 ( .A(r_wr[3]), .B(n86), .C(n78), .D(n19), .Y(upd_dbuf[0]) );
  OAI22X1 U150 ( .A(r_wr[3]), .B(n83), .C(n78), .D(n22), .Y(upd_dbuf[2]) );
  OAI22X1 U151 ( .A(n106), .B(n258), .C(n348), .D(n74), .Y(N260) );
  AOI22X1 U152 ( .A(n40), .B(n344), .C(n79), .D(n346), .Y(n348) );
  OAI211X1 U153 ( .C(n349), .D(n310), .A(n8), .B(n350), .Y(N22) );
  NOR2X1 U154 ( .A(n282), .B(n283), .Y(net9514) );
  AOI21X1 U155 ( .B(N225), .C(n88), .A(n284), .Y(n282) );
  NOR2X1 U156 ( .A(n285), .B(n283), .Y(net9512) );
  AOI21X1 U157 ( .B(N227), .C(n88), .A(n284), .Y(n285) );
  NAND2X1 U158 ( .A(n280), .B(n150), .Y(N205) );
  NAND3X1 U159 ( .A(n46), .B(n481), .C(n482), .Y(N1009) );
  AOI221XL U160 ( .A(n116), .B(n544), .C(n554), .D(n483), .E(n484), .Y(n482)
         );
  INVX1 U161 ( .A(n485), .Y(n116) );
  INVX1 U162 ( .A(n244), .Y(n80) );
  AOI31X1 U163 ( .A(ff_chg), .B(n245), .C(n246), .D(r_wr[4]), .Y(n244) );
  XNOR2XL U164 ( .A(n34), .B(n76), .Y(n346) );
  OAI22X1 U165 ( .A(n35), .B(n81), .C(r_wr[4]), .D(n70), .Y(tui_wdat[7]) );
  OAI21X1 U166 ( .B(n130), .C(n131), .A(n14), .Y(upd_dbuf_en) );
  NAND4X1 U167 ( .A(n145), .B(n146), .C(n147), .D(n148), .Y(n130) );
  NAND4X1 U168 ( .A(n132), .B(n133), .C(n134), .D(n135), .Y(n131) );
  NOR3XL U169 ( .A(n149), .B(n150), .C(n151), .Y(n148) );
  AOI21X1 U170 ( .B(n544), .C(n278), .A(r_wr[3]), .Y(N444) );
  AOI31X1 U171 ( .A(n547), .B(n129), .C(n277), .D(n409), .Y(n407) );
  INVX1 U172 ( .A(n331), .Y(n66) );
  INVX1 U173 ( .A(n142), .Y(n67) );
  OAI221X1 U174 ( .A(n422), .B(n76), .C(n57), .D(n423), .E(n424), .Y(n409) );
  AOI221XL U175 ( .A(n417), .B(n425), .C(n547), .D(n125), .E(n551), .Y(n423)
         );
  AOI211X1 U176 ( .C(n473), .D(n555), .A(n474), .B(n475), .Y(n422) );
  AOI33X1 U177 ( .A(n410), .B(n421), .C(n545), .D(n301), .E(n425), .F(n97), 
        .Y(n424) );
  NOR2X1 U178 ( .A(n342), .B(n142), .Y(add_263_carry[1]) );
  ENOX1 U179 ( .A(n407), .B(n123), .C(n27), .D(n408), .Y(N1015) );
  ENOX1 U180 ( .A(n407), .B(n121), .C(n28), .D(n408), .Y(N1014) );
  ENOX1 U181 ( .A(n407), .B(n542), .C(n31), .D(n408), .Y(N1011) );
  ENOX1 U182 ( .A(n407), .B(n127), .C(n30), .D(n408), .Y(N1012) );
  NOR32XL U183 ( .B(n204), .C(n205), .A(n208), .Y(n213) );
  NAND31X1 U184 ( .C(n171), .A(n170), .B(n174), .Y(n162) );
  AOI33X1 U185 ( .A(n175), .B(n176), .C(n177), .D(n98), .E(n99), .F(n178), .Y(
        n174) );
  AOI22X1 U186 ( .A(n173), .B(n179), .C(n101), .D(n173), .Y(n178) );
  INVX1 U187 ( .A(n157), .Y(n98) );
  AOI21BBXL U188 ( .B(n108), .C(rx_ui_3_8[4]), .A(n463), .Y(n459) );
  INVX1 U189 ( .A(n339), .Y(n65) );
  XNOR2XL U190 ( .A(n218), .B(n238), .Y(n204) );
  XNOR2XL U191 ( .A(n231), .B(n232), .Y(n238) );
  OAI22X1 U192 ( .A(n206), .B(n18), .C(n103), .D(n207), .Y(n175) );
  AOI21X1 U193 ( .B(n203), .C(n202), .A(n210), .Y(n206) );
  XNOR2XL U194 ( .A(n208), .B(n209), .Y(n207) );
  NAND2X1 U195 ( .A(n205), .B(n204), .Y(n209) );
  INVX1 U196 ( .A(n153), .Y(n61) );
  OAI211X1 U197 ( .C(n157), .D(n167), .A(n168), .B(n169), .Y(n154) );
  OAI31XL U198 ( .A(n172), .B(n159), .C(n160), .D(n100), .Y(n167) );
  NOR21XL U199 ( .B(n170), .A(n171), .Y(n169) );
  NAND2X1 U200 ( .A(n6), .B(n542), .Y(n404) );
  OAI21X1 U201 ( .B(n232), .C(n237), .A(n240), .Y(n233) );
  OAI21BBX1 U202 ( .A(n237), .B(n232), .C(N107), .Y(n240) );
  OAI22X1 U203 ( .A(n103), .B(n200), .C(n18), .D(n201), .Y(n176) );
  XNOR2XL U204 ( .A(n202), .B(n203), .Y(n201) );
  XNOR2XL U205 ( .A(n204), .B(n205), .Y(n200) );
  NAND2X1 U206 ( .A(n541), .B(n127), .Y(n241) );
  NAND2X1 U207 ( .A(n241), .B(n403), .Y(n235) );
  NAND2X1 U208 ( .A(n235), .B(n543), .Y(n237) );
  NOR32XL U209 ( .B(add_274_carry[8]), .C(n193), .A(n196), .Y(n205) );
  NOR21XL U210 ( .B(n231), .A(n232), .Y(n215) );
  XNOR2XL U211 ( .A(N107), .B(n236), .Y(n193) );
  XNOR2XL U212 ( .A(n232), .B(n237), .Y(n236) );
  OAI21X1 U213 ( .B(n242), .C(n121), .A(n230), .Y(n216) );
  OAI22X1 U214 ( .A(n103), .B(n190), .C(n18), .D(n191), .Y(n181) );
  XNOR2XL U215 ( .A(add_274_2_carry[8]), .B(n192), .Y(n191) );
  XNOR2XL U216 ( .A(add_274_carry[8]), .B(n193), .Y(n190) );
  INVX1 U217 ( .A(n144), .Y(n63) );
  OAI22X1 U218 ( .A(n18), .B(n194), .C(n103), .D(n195), .Y(n186) );
  XNOR2XL U219 ( .A(n198), .B(n199), .Y(n194) );
  XNOR2XL U220 ( .A(n196), .B(n197), .Y(n195) );
  NAND2X1 U221 ( .A(add_274_2_carry[8]), .B(n192), .Y(n199) );
  NAND2X1 U222 ( .A(rx_ui_3_8[2]), .B(n119), .Y(n470) );
  NAND2X1 U223 ( .A(n371), .B(n106), .Y(n379) );
  OAI21X1 U224 ( .B(n533), .C(n129), .A(n288), .Y(n515) );
  NOR2X1 U225 ( .A(n534), .B(n95), .Y(n533) );
  AOI22AXL U226 ( .A(n371), .B(n378), .D(n358), .C(n542), .Y(n534) );
  OAI22X1 U227 ( .A(rx_ui_3_8[2]), .B(n119), .C(rx_ui_3_8[1]), .D(n105), .Y(
        n467) );
  NAND2X1 U228 ( .A(n404), .B(n378), .Y(N107) );
  OAI31XL U229 ( .A(n351), .B(n96), .C(n352), .D(n353), .Y(n276) );
  AOI32X1 U230 ( .A(n93), .B(n354), .C(n551), .D(n355), .E(n356), .Y(n353) );
  NOR31X1 U231 ( .C(n357), .A(n358), .B(n359), .Y(n356) );
  NOR3XL U232 ( .A(n360), .B(n112), .C(n361), .Y(n355) );
  AOI22X1 U233 ( .A(rx_ui_3_8[1]), .B(n105), .C(n469), .D(n104), .Y(n468) );
  XNOR2XL U234 ( .A(n69), .B(n142), .Y(n469) );
  NAND2X1 U235 ( .A(n242), .B(n121), .Y(n230) );
  NOR2X1 U236 ( .A(n106), .B(n543), .Y(n358) );
  NAND2X1 U237 ( .A(add_274_carry[8]), .B(n193), .Y(n197) );
  NAND2X1 U238 ( .A(n453), .B(n153), .Y(n452) );
  INVX1 U239 ( .A(n454), .Y(n68) );
  INVX1 U240 ( .A(n463), .Y(n58) );
  XNOR2XL U241 ( .A(n339), .B(n153), .Y(n325) );
  XNOR2XL U242 ( .A(n225), .B(n129), .Y(n202) );
  XNOR2XL U243 ( .A(n18), .B(n189), .Y(n164) );
  AOI21X1 U244 ( .B(n543), .C(n122), .A(add_274_2_carry[6]), .Y(n189) );
  XNOR2XL U245 ( .A(adp_tx_1_4[5]), .B(n122), .Y(n432) );
  NOR2X1 U246 ( .A(n382), .B(n119), .Y(N1254) );
  NOR2X1 U247 ( .A(n382), .B(n124), .Y(N1255) );
  NOR2X1 U248 ( .A(n382), .B(n5), .Y(N1256) );
  NOR2X1 U249 ( .A(n382), .B(n122), .Y(N1257) );
  NOR2X1 U250 ( .A(n382), .B(n105), .Y(N1253) );
  XNOR2XL U251 ( .A(adp_tx_1_4[6]), .B(n107), .Y(n433) );
  XNOR2XL U252 ( .A(adp_tx_1_4[4]), .B(n108), .Y(n431) );
  NOR2X1 U253 ( .A(n382), .B(n107), .Y(N1258) );
  AND2X1 U254 ( .A(n489), .B(n493), .Y(n246) );
  NAND2X1 U255 ( .A(n374), .B(n129), .Y(n349) );
  AOI22X1 U256 ( .A(N172), .B(n103), .C(N144), .D(n18), .Y(n182) );
  XNOR2XL U257 ( .A(adp_tx_ui_7_), .B(n118), .Y(n530) );
  XNOR2XL U258 ( .A(n107), .B(adp_tx_ui_6_), .Y(n528) );
  INVX1 U259 ( .A(n151), .Y(n545) );
  NOR2X1 U260 ( .A(n382), .B(n104), .Y(N1252) );
  NOR3XL U261 ( .A(n124), .B(n108), .C(n164), .Y(n183) );
  NAND4X1 U262 ( .A(tx_en), .B(n543), .C(n296), .D(n297), .Y(n278) );
  AOI21X1 U263 ( .B(n550), .C(n277), .A(n298), .Y(n297) );
  NAND3X1 U264 ( .A(n299), .B(n300), .C(n301), .Y(n296) );
  NAND2X1 U265 ( .A(n57), .B(n544), .Y(n494) );
  AOI22X1 U266 ( .A(N173), .B(n103), .C(N145), .D(n18), .Y(n184) );
  AOI221XL U267 ( .A(n65), .B(n545), .C(n392), .D(n71), .E(n246), .Y(n395) );
  NAND2X1 U268 ( .A(n374), .B(n127), .Y(n380) );
  AOI21X1 U269 ( .B(n105), .C(n69), .A(add_263_carry[1]), .Y(n328) );
  AOI211X1 U270 ( .C(n298), .D(n113), .A(n246), .B(n312), .Y(n313) );
  INVX1 U271 ( .A(n277), .Y(n57) );
  ENOX1 U272 ( .A(n153), .B(n151), .C(adp_tx_ui_6_), .D(n392), .Y(n400) );
  NOR2X1 U273 ( .A(n62), .B(n108), .Y(n335) );
  INVX1 U274 ( .A(n342), .Y(n69) );
  ENOX1 U275 ( .A(n332), .B(n333), .C(n107), .D(n316), .Y(n317) );
  AOI22AXL U276 ( .A(n334), .B(n122), .D(n335), .C(n336), .Y(n333) );
  AOI221XL U277 ( .A(n336), .B(n122), .C(n62), .D(n108), .E(n337), .Y(n332) );
  NAND21X1 U278 ( .B(n336), .A(n335), .Y(n334) );
  NOR2X1 U279 ( .A(n119), .B(n65), .Y(n453) );
  NOR2X1 U280 ( .A(n543), .B(n122), .Y(add_274_2_carry[6]) );
  NAND2X1 U281 ( .A(n123), .B(n121), .Y(n274) );
  INVX1 U282 ( .A(n374), .Y(n112) );
  INVX1 U283 ( .A(n312), .Y(n60) );
  NOR2X1 U284 ( .A(n142), .B(n141), .Y(add_264_carry[1]) );
  NOR32XL U285 ( .B(add_274_2_carry[8]), .C(n192), .A(n198), .Y(n203) );
  XNOR2XL U286 ( .A(adp_tx_1_4[3]), .B(n124), .Y(n430) );
  NAND2X1 U287 ( .A(n489), .B(n532), .Y(n295) );
  NOR2X1 U288 ( .A(n310), .B(n149), .Y(n539) );
  NAND2X1 U289 ( .A(n367), .B(n542), .Y(n298) );
  OAI32X1 U290 ( .A(n279), .B(n476), .C(n414), .D(n109), .E(n420), .Y(n474) );
  INVX1 U291 ( .A(n419), .Y(n109) );
  NOR3XL U292 ( .A(n417), .B(n550), .C(n301), .Y(n364) );
  OAI21X1 U293 ( .B(n360), .C(n96), .A(n418), .Y(n416) );
  INVX1 U294 ( .A(n18), .Y(n103) );
  INVX1 U295 ( .A(n150), .Y(n88) );
  INVX1 U296 ( .A(n535), .Y(n549) );
  NAND4X1 U297 ( .A(n436), .B(n437), .C(n438), .D(n439), .Y(n421) );
  XNOR2XL U298 ( .A(n142), .B(n119), .Y(n437) );
  NOR21XL U299 ( .B(n427), .A(n443), .Y(n438) );
  XNOR2XL U300 ( .A(n153), .B(n122), .Y(n436) );
  NAND2X1 U301 ( .A(n339), .B(n124), .Y(n329) );
  NOR2X1 U302 ( .A(n136), .B(n137), .Y(n134) );
  XNOR2XL U303 ( .A(rx_ui_5_8[3]), .B(n124), .Y(n136) );
  XNOR2XL U304 ( .A(n138), .B(n139), .Y(n137) );
  INVX1 U305 ( .A(n299), .Y(n551) );
  NAND2X1 U306 ( .A(n121), .B(n217), .Y(n210) );
  INVX1 U307 ( .A(n227), .Y(n128) );
  XNOR2XL U308 ( .A(n143), .B(n118), .Y(n132) );
  OR2X1 U309 ( .A(n139), .B(n144), .Y(n143) );
  INVX1 U310 ( .A(n417), .Y(n97) );
  INVX1 U311 ( .A(n354), .Y(n94) );
  OAI22X1 U312 ( .A(n110), .B(n287), .C(n473), .D(n273), .Y(n419) );
  INVX1 U313 ( .A(ff_chg), .Y(n75) );
  XNOR2XL U314 ( .A(adp_tx_1_4[0]), .B(n104), .Y(n435) );
  XNOR2XL U315 ( .A(adp_tx_1_4[1]), .B(n105), .Y(n434) );
  OAI32X1 U316 ( .A(n113), .B(n490), .C(n151), .D(n287), .E(n491), .Y(n475) );
  NAND2X1 U317 ( .A(n112), .B(n538), .Y(n491) );
  NAND4X1 U318 ( .A(n403), .B(n129), .C(n123), .D(n111), .Y(n538) );
  AOI31X1 U319 ( .A(n519), .B(n57), .C(n114), .D(n299), .Y(n484) );
  NOR3XL U320 ( .A(n144), .B(n153), .C(n339), .Y(n316) );
  INVX1 U321 ( .A(n490), .Y(n117) );
  INVX1 U322 ( .A(n217), .Y(n120) );
  NOR2X1 U323 ( .A(n378), .B(n127), .Y(n519) );
  NOR3XL U324 ( .A(n76), .B(n476), .C(n279), .Y(n413) );
  NOR2X1 U325 ( .A(n300), .B(n149), .Y(n497) );
  NAND2X1 U326 ( .A(ff_chg), .B(n545), .Y(n275) );
  INVX1 U327 ( .A(n279), .Y(n552) );
  NAND2X1 U328 ( .A(n96), .B(n57), .Y(n483) );
  INVX1 U329 ( .A(n360), .Y(n554) );
  XNOR2XL U330 ( .A(n140), .B(n141), .Y(n133) );
  XNOR2XL U331 ( .A(n142), .B(n104), .Y(n140) );
  NOR3XL U332 ( .A(n349), .B(n299), .C(n126), .Y(n496) );
  NAND2X1 U333 ( .A(n288), .B(n222), .Y(n245) );
  INVX1 U334 ( .A(n273), .Y(n555) );
  NAND2X1 U335 ( .A(n349), .B(n405), .Y(N1043) );
  OAI21X1 U336 ( .B(n406), .C(n300), .A(n299), .Y(n405) );
  OAI21X1 U337 ( .B(n90), .C(n89), .A(n295), .Y(n289) );
  AOI21X1 U338 ( .B(n89), .C(n90), .A(n289), .Y(n506) );
  NOR2X1 U339 ( .A(n75), .B(n279), .Y(n540) );
  NAND3X1 U340 ( .A(n532), .B(fcp_state[0]), .C(fcp_state[3]), .Y(n299) );
  NAND3X1 U341 ( .A(n492), .B(n557), .C(fcp_state[2]), .Y(n360) );
  NAND3X1 U342 ( .A(fcp_state[0]), .B(n493), .C(fcp_state[3]), .Y(n535) );
  NOR2X1 U343 ( .A(n557), .B(fcp_state[2]), .Y(n493) );
  NOR2X1 U344 ( .A(n556), .B(fcp_state[0]), .Y(n492) );
  NOR2X1 U345 ( .A(fcp_state[2]), .B(fcp_state[1]), .Y(n532) );
  INVX1 U346 ( .A(fcp_state[1]), .Y(n557) );
  INVX1 U347 ( .A(fcp_state[3]), .Y(n556) );
  AOI22X1 U348 ( .A(n34), .B(n79), .C(r_dat[7]), .D(n40), .Y(n264) );
  AOI22X1 U349 ( .A(n21), .B(n79), .C(r_dat[2]), .D(n40), .Y(n255) );
  AOI22X1 U350 ( .A(r_wdat[1]), .B(n79), .C(r_dat[1]), .D(n40), .Y(n256) );
  AOI22X1 U351 ( .A(r_wdat[0]), .B(n79), .C(r_dat[0]), .D(n40), .Y(n259) );
  ENOX1 U352 ( .A(n33), .B(n269), .C(r_dat[6]), .D(n40), .Y(n252) );
  ENOX1 U353 ( .A(n23), .B(n269), .C(r_dat[3]), .D(n40), .Y(n253) );
  ENOX1 U354 ( .A(n24), .B(n269), .C(r_dat[4]), .D(n40), .Y(n250) );
  ENOX1 U355 ( .A(n25), .B(n269), .C(r_dat[5]), .D(n40), .Y(n249) );
  AOI211X1 U356 ( .C(n269), .D(n344), .A(n43), .B(n345), .Y(n251) );
  OAI21BBX1 U357 ( .A(n346), .B(n347), .C(r_ctl[0]), .Y(n345) );
  OAI32X1 U358 ( .A(n72), .B(n513), .C(n269), .D(n514), .E(n494), .Y(n495) );
  INVX1 U359 ( .A(r_ctl[4]), .Y(n72) );
  AOI22X1 U360 ( .A(n549), .B(n515), .C(n96), .D(n554), .Y(n514) );
  NAND31X1 U361 ( .C(n498), .A(n481), .B(n499), .Y(N1007) );
  AOI32X1 U362 ( .A(n552), .B(ff_idn), .C(n476), .D(n500), .E(n44), .Y(n499)
         );
  OAI21X1 U363 ( .B(r_ctl[0]), .C(n73), .A(n261), .Y(n500) );
  INVX1 U364 ( .A(n501), .Y(n44) );
  AO33X1 U365 ( .A(n43), .B(n548), .C(r_ctl[5]), .D(n262), .E(n261), .F(n251), 
        .Y(trans_buf[0]) );
  NAND41X1 U366 ( .D(n413), .A(n418), .B(n505), .C(n508), .Y(N1006) );
  AOI31X1 U367 ( .A(r_ctl[4]), .B(n553), .C(n513), .D(n484), .Y(n505) );
  AOI221XL U368 ( .A(n510), .B(n73), .C(n549), .D(n277), .E(n498), .Y(n508) );
  GEN2XL U369 ( .D(n497), .E(n57), .C(n496), .B(n544), .A(n495), .Y(n510) );
  AO2222XL U370 ( .A(n43), .B(rxtx_buf[5]), .C(n251), .D(n249), .E(n38), .F(
        n74), .G(n254), .H(n250), .Y(trans_buf[6]) );
  AO2222XL U371 ( .A(n43), .B(rxtx_buf[4]), .C(n251), .D(n250), .E(n36), .F(
        n74), .G(n254), .H(n253), .Y(trans_buf[5]) );
  AO2222XL U372 ( .A(n43), .B(rxtx_buf[7]), .C(n250), .D(n74), .E(n251), .F(
        n39), .G(n42), .H(n252), .Y(trans_buf[8]) );
  AO2222XL U373 ( .A(n43), .B(rxtx_buf[6]), .C(n253), .D(n74), .E(n251), .F(
        n252), .G(n254), .H(n249), .Y(trans_buf[7]) );
  AO2222XL U374 ( .A(rxtx_buf[9]), .B(n43), .C(n252), .D(n74), .E(n251), .F(
        n39), .G(n42), .H(n264), .Y(trans_buf[10]) );
  AO2222XL U375 ( .A(n43), .B(rxtx_buf[3]), .C(n251), .D(n253), .E(n37), .F(
        n74), .G(n254), .H(n38), .Y(trans_buf[4]) );
  NAND4X1 U376 ( .A(n290), .B(n291), .C(n292), .D(n293), .Y(intr) );
  AOI22X1 U377 ( .A(r_msk[2]), .B(r_irq[2]), .C(r_msk[3]), .D(r_irq[3]), .Y(
        n292) );
  AOI22X1 U378 ( .A(r_msk[4]), .B(r_irq[4]), .C(r_msk[5]), .D(r_irq[5]), .Y(
        n291) );
  AOI22X1 U379 ( .A(r_msk[6]), .B(r_irq[6]), .C(r_msk[7]), .D(r_irq[7]), .Y(
        n290) );
  OAI21BBX1 U380 ( .A(n483), .B(n554), .C(n486), .Y(N1008) );
  AOI32X1 U381 ( .A(r_ctl[0]), .B(n487), .C(r_ctl[1]), .D(ff_idn), .E(n488), 
        .Y(n486) );
  OR2X1 U382 ( .A(n475), .B(n555), .Y(n488) );
  OAI21X1 U383 ( .B(n485), .C(n494), .A(n46), .Y(n487) );
  OAI21BBX1 U384 ( .A(N363), .B(n8), .C(n41), .Y(N261) );
  NAND2X1 U385 ( .A(n263), .B(n248), .Y(trans_buf[11]) );
  AOI22X1 U386 ( .A(n39), .B(n74), .C(rxtx_buf[10]), .D(n43), .Y(n263) );
  NAND2X1 U387 ( .A(n247), .B(n248), .Y(trans_buf[9]) );
  AOI22X1 U388 ( .A(n249), .B(n74), .C(rxtx_buf[8]), .D(n43), .Y(n247) );
  OAI22X1 U389 ( .A(n20), .B(n81), .C(n155), .D(n163), .Y(tui_wdat[1]) );
  XNOR2XL U390 ( .A(n164), .B(n165), .Y(n163) );
  NAND2X1 U391 ( .A(n10), .B(N142), .Y(n165) );
  OAI22X1 U392 ( .A(n19), .B(n81), .C(n166), .D(n155), .Y(tui_wdat[0]) );
  XNOR2XL U393 ( .A(N142), .B(n10), .Y(n166) );
  ENOX1 U394 ( .A(n78), .B(n23), .C(n78), .D(rxtx_buf[3]), .Y(upd_dbuf[3]) );
  ENOX1 U395 ( .A(n14), .B(n24), .C(n78), .D(rxtx_buf[4]), .Y(upd_dbuf[4]) );
  ENOX1 U396 ( .A(n14), .B(n25), .C(n78), .D(rxtx_buf[5]), .Y(upd_dbuf[5]) );
  ENOX1 U397 ( .A(n14), .B(n33), .C(n78), .D(rxtx_buf[6]), .Y(upd_dbuf[6]) );
  AO22AXL U398 ( .A(n78), .B(rxtx_buf[7]), .C(r_wdat[7]), .D(n78), .Y(
        upd_dbuf[7]) );
  BUFX3 U399 ( .A(ff_idn), .Y(r_ctl[5]) );
  OAI22X1 U400 ( .A(r_tui[7]), .B(r_tui[3]), .C(catch_sync[1]), .D(n70), .Y(
        n142) );
  OAI22X1 U401 ( .A(r_tui[7]), .B(r_tui[4]), .C(catch_sync[2]), .D(n70), .Y(
        n331) );
  OAI22X1 U402 ( .A(r_tui[7]), .B(r_tui[2]), .C(catch_sync[0]), .D(n70), .Y(
        n342) );
  AO22X1 U403 ( .A(n409), .B(n12), .C(n29), .D(n408), .Y(N1013) );
  INVX1 U404 ( .A(r_tui[7]), .Y(n70) );
  OAI21X1 U405 ( .B(ui_intv_cnt[5]), .C(n461), .A(n462), .Y(n460) );
  AOI33X1 U406 ( .A(n458), .B(n108), .C(rx_ui_3_8[4]), .D(n63), .E(n107), .F(
        add_263_carry[5]), .Y(n462) );
  OAI32X1 U407 ( .A(n117), .B(new_rx_sync_cnt[1]), .C(new_rx_sync_cnt[0]), .D(
        n444), .E(n445), .Y(n410) );
  NOR4XL U408 ( .A(n446), .B(n447), .C(n75), .D(n87), .Y(n445) );
  OAI31XL U409 ( .A(n448), .B(ui_intv_cnt[6]), .C(ui_intv_cnt[5]), .D(n349), 
        .Y(n447) );
  AOI32X1 U410 ( .A(n457), .B(n458), .C(n459), .D(n58), .E(n460), .Y(n446) );
  ENOX1 U411 ( .A(n407), .B(n111), .C(n26), .D(n408), .Y(N1016) );
  ENOX1 U412 ( .A(n407), .B(n543), .C(n32), .D(n408), .Y(N1010) );
  NAND2X1 U413 ( .A(n461), .B(ui_intv_cnt[5]), .Y(n458) );
  OAI22X1 U414 ( .A(catch_sync[4]), .B(n70), .C(r_tui[7]), .D(adp_tx_ui_6_), 
        .Y(n153) );
  OAI22X1 U415 ( .A(r_tui[7]), .B(n71), .C(catch_sync[3]), .D(n70), .Y(n339)
         );
  NOR21XL U416 ( .B(n211), .A(n212), .Y(n170) );
  OAI31XL U417 ( .A(n213), .B(n103), .C(n214), .D(n111), .Y(n212) );
  AOI33X1 U418 ( .A(n103), .B(n120), .C(symb_cnt[4]), .D(n214), .E(n18), .F(
        n213), .Y(n211) );
  NAND2X1 U419 ( .A(n215), .B(n216), .Y(n214) );
  GEN2XL U420 ( .D(n64), .E(n124), .C(rx_ui_3_8[3]), .B(n465), .A(n466), .Y(
        n457) );
  INVX1 U421 ( .A(n470), .Y(n64) );
  NAND2X1 U422 ( .A(N141), .B(n470), .Y(n465) );
  AOI211X1 U423 ( .C(N141), .D(n59), .A(n467), .B(n468), .Y(n466) );
  INVX1 U424 ( .A(N159), .Y(n543) );
  AOI21X1 U425 ( .B(n241), .C(symb_cnt[3]), .A(n242), .Y(n232) );
  OAI21X1 U426 ( .B(r_tui[6]), .C(n71), .A(adp_tx_ui_7_), .Y(adp_tx_ui_6_) );
  INVX1 U427 ( .A(symb_cnt[2]), .Y(n127) );
  INVX1 U428 ( .A(N160), .Y(n542) );
  OAI2B11X1 U429 ( .D(n410), .C(n310), .A(n411), .B(n412), .Y(n408) );
  AOI31X1 U430 ( .A(ff_idn), .B(n419), .C(n420), .D(n364), .Y(n411) );
  AOI22X1 U431 ( .A(n413), .B(n414), .C(n57), .D(n415), .Y(n412) );
  AO222X1 U432 ( .A(n126), .B(n551), .C(n416), .D(n417), .E(n129), .F(n547), 
        .Y(n415) );
  INVX1 U433 ( .A(r_tui[5]), .Y(n71) );
  NAND2X1 U434 ( .A(r_tui[6]), .B(n71), .Y(adp_tx_ui_7_) );
  NOR2X1 U435 ( .A(n241), .B(symb_cnt[3]), .Y(n242) );
  NAND2X1 U436 ( .A(n7), .B(n404), .Y(n403) );
  XNOR2XL U437 ( .A(N159), .B(n235), .Y(N108) );
  OAI22X1 U438 ( .A(catch_sync[5]), .B(n70), .C(r_tui[7]), .D(adp_tx_ui_7_), 
        .Y(n144) );
  XNOR2XL U439 ( .A(N363), .B(n4), .Y(n371) );
  NAND3X1 U440 ( .A(n349), .B(n368), .C(n369), .Y(n361) );
  NAND42X1 U441 ( .C(n359), .D(n112), .A(n370), .B(n357), .Y(n369) );
  OAI22X1 U442 ( .A(N362), .B(N159), .C(N160), .D(n371), .Y(n370) );
  XOR2X1 U443 ( .A(n215), .B(n229), .Y(n208) );
  OAI21X1 U444 ( .B(n230), .C(symb_cnt[5]), .A(n216), .Y(n229) );
  OAI32X1 U445 ( .A(n218), .B(n103), .C(n213), .D(n219), .E(n18), .Y(n171) );
  AOI31X1 U446 ( .A(n202), .B(n210), .C(n203), .D(symb_cnt[5]), .Y(n219) );
  NAND2X1 U447 ( .A(n118), .B(n464), .Y(n463) );
  OAI21BBX1 U448 ( .A(n63), .B(add_263_carry[5]), .C(ui_intv_cnt[6]), .Y(n464)
         );
  OAI211X1 U449 ( .C(n372), .D(n129), .A(n373), .B(n374), .Y(n354) );
  NOR2X1 U450 ( .A(n95), .B(n375), .Y(n372) );
  NAND3X1 U451 ( .A(symb_cnt[2]), .B(n375), .C(n95), .Y(n373) );
  OAI211X1 U452 ( .C(n376), .D(n371), .A(n377), .B(n378), .Y(n375) );
  NAND2X1 U453 ( .A(ui_intv_cnt[0]), .B(n142), .Y(n454) );
  NAND2X1 U454 ( .A(N160), .B(N159), .Y(n378) );
  OAI21X1 U455 ( .B(n63), .C(n108), .A(n449), .Y(n448) );
  OAI22X1 U456 ( .A(N142), .B(n144), .C(n450), .D(n451), .Y(n449) );
  AOI22AXL U457 ( .A(n452), .B(n124), .D(n453), .C(n61), .Y(n451) );
  AOI211X1 U458 ( .C(n66), .D(n454), .A(n455), .B(n456), .Y(n450) );
  OAI22X1 U459 ( .A(N141), .B(n153), .C(ui_intv_cnt[2]), .D(n339), .Y(n455) );
  OAI21X1 U460 ( .B(N160), .C(symb_cnt[2]), .A(n379), .Y(n377) );
  AOI21X1 U461 ( .B(n68), .C(n331), .A(ui_intv_cnt[1]), .Y(n456) );
  XNOR2XL U462 ( .A(N159), .B(n127), .Y(N161) );
  NOR32XL U463 ( .B(r_ctl[7]), .C(n276), .A(n277), .Y(setsta[0]) );
  NOR2X1 U464 ( .A(N159), .B(n122), .Y(add_274_carry[6]) );
  AND4X1 U465 ( .A(n383), .B(n384), .C(n385), .D(n386), .Y(n382) );
  XNOR2XL U466 ( .A(n401), .B(n104), .Y(n383) );
  XNOR2XL U467 ( .A(ui_intv_cnt[6]), .B(n400), .Y(n384) );
  NOR2X1 U468 ( .A(n396), .B(n397), .Y(n385) );
  NOR21XL U469 ( .B(n230), .A(symb_cnt[5]), .Y(n218) );
  NAND31X1 U470 ( .C(n380), .A(N362), .B(N363), .Y(n368) );
  OAI21X1 U471 ( .B(n228), .C(n221), .A(n222), .Y(n227) );
  NOR2X1 U472 ( .A(N160), .B(symb_cnt[3]), .Y(n228) );
  INVX1 U473 ( .A(n517), .Y(n96) );
  OAI211X1 U474 ( .C(n518), .D(n380), .A(n368), .B(n444), .Y(n517) );
  AOI22X1 U475 ( .A(N363), .B(n378), .C(N362), .D(n542), .Y(n518) );
  INVX1 U476 ( .A(N141), .Y(n124) );
  XNOR2XL U477 ( .A(n105), .B(r_tui[1]), .Y(n526) );
  XNOR2XL U478 ( .A(n391), .B(n119), .Y(n390) );
  ENOX1 U479 ( .A(n151), .B(n342), .C(r_tui[2]), .D(n392), .Y(n391) );
  XNOR2XL U480 ( .A(n108), .B(r_tui[4]), .Y(n527) );
  XNOR2XL U481 ( .A(n399), .B(n108), .Y(n396) );
  ENOX1 U482 ( .A(n151), .B(n331), .C(r_tui[4]), .D(n392), .Y(n399) );
  NOR2X1 U483 ( .A(n274), .B(symb_cnt[6]), .Y(n374) );
  AOI21X1 U484 ( .B(symb_cnt[3]), .C(symb_cnt[2]), .A(n112), .Y(n288) );
  INVX1 U485 ( .A(ui_intv_cnt[5]), .Y(n122) );
  NAND4X1 U486 ( .A(n520), .B(n88), .C(n521), .D(n522), .Y(n277) );
  XNOR2XL U487 ( .A(ui_intv_cnt[2]), .B(r_tui[2]), .Y(n520) );
  NOR4XL U488 ( .A(n523), .B(n524), .C(n526), .D(n527), .Y(n522) );
  NOR3XL U489 ( .A(n528), .B(n529), .C(n530), .Y(n521) );
  OAI21X1 U490 ( .B(n221), .C(n222), .A(n223), .Y(n192) );
  AOI32X1 U491 ( .A(n221), .B(n542), .C(symb_cnt[3]), .D(n224), .E(n129), .Y(
        n223) );
  XNOR2XL U492 ( .A(N160), .B(n221), .Y(n224) );
  INVX1 U493 ( .A(N142), .Y(n108) );
  NAND3X1 U494 ( .A(n493), .B(n556), .C(fcp_state[0]), .Y(n151) );
  INVX1 U495 ( .A(ui_intv_cnt[2]), .Y(n119) );
  OAI22X1 U496 ( .A(n128), .B(n127), .C(n226), .D(n121), .Y(n225) );
  NOR2X1 U497 ( .A(symb_cnt[2]), .B(n227), .Y(n226) );
  INVX1 U498 ( .A(ui_intv_cnt[1]), .Y(n105) );
  INVX1 U499 ( .A(ui_intv_cnt[0]), .Y(n104) );
  INVX1 U500 ( .A(N362), .Y(n106) );
  INVX1 U501 ( .A(symb_cnt[4]), .Y(n121) );
  OAI22X1 U502 ( .A(n322), .B(n323), .C(ui_intv_cnt[5]), .D(n321), .Y(n319) );
  NOR2X1 U503 ( .A(n324), .B(n325), .Y(n323) );
  AOI21X1 U504 ( .B(n324), .C(n325), .A(n5), .Y(n322) );
  AND2X1 U505 ( .A(n326), .B(n327), .Y(n324) );
  INVX1 U506 ( .A(symb_cnt[5]), .Y(n123) );
  AOI22X1 U507 ( .A(r_msk[0]), .B(r_irq[0]), .C(r_msk[1]), .D(r_irq[1]), .Y(
        n293) );
  OAI32X1 U508 ( .A(n84), .B(new_rx_sync_cnt[1]), .C(n60), .D(n311), .E(n85), 
        .Y(N349) );
  AOI21X1 U509 ( .B(n312), .C(n84), .A(n313), .Y(n311) );
  INVX1 U510 ( .A(new_rx_sync_cnt[0]), .Y(n84) );
  XNOR2XL U511 ( .A(ui_intv_cnt[7]), .B(n398), .Y(n397) );
  AOI221XL U512 ( .A(n545), .B(n63), .C(n392), .D(adp_tx_ui_7_), .E(n246), .Y(
        n398) );
  AOI21X1 U513 ( .B(N362), .C(N363), .A(n127), .Y(n359) );
  NAND4X1 U514 ( .A(n426), .B(n427), .C(n428), .D(n429), .Y(n301) );
  NOR2X1 U515 ( .A(n434), .B(n435), .Y(n428) );
  XNOR2XL U516 ( .A(ui_intv_cnt[2]), .B(adp_tx_1_4[2]), .Y(n426) );
  NOR4XL U517 ( .A(n430), .B(n431), .C(n432), .D(n433), .Y(n429) );
  ENOX1 U518 ( .A(n141), .B(n151), .C(r_tui[1]), .D(n392), .Y(n394) );
  ENOX1 U519 ( .A(n142), .B(n151), .C(r_tui[3]), .D(n392), .Y(n393) );
  NOR2X1 U520 ( .A(fcp_state[3]), .B(fcp_state[0]), .Y(n489) );
  NOR4XL U521 ( .A(n387), .B(n388), .C(n389), .D(n390), .Y(n386) );
  XNOR2XL U522 ( .A(ui_intv_cnt[5]), .B(n395), .Y(n387) );
  XNOR2XL U523 ( .A(n394), .B(n105), .Y(n388) );
  XNOR2XL U524 ( .A(n393), .B(n124), .Y(n389) );
  NAND2X1 U525 ( .A(symb_cnt[2]), .B(N159), .Y(n221) );
  AOI22X1 U526 ( .A(n338), .B(n329), .C(n65), .D(N141), .Y(n337) );
  OAI21X1 U527 ( .B(n66), .C(n340), .A(n341), .Y(n338) );
  OAI21BBX1 U528 ( .A(n340), .B(n66), .C(ui_intv_cnt[2]), .Y(n341) );
  OAI221X1 U529 ( .A(ui_intv_cnt[1]), .B(n68), .C(ui_intv_cnt[0]), .D(n142), 
        .E(n328), .Y(n340) );
  OAI211X1 U530 ( .C(ui_intv_cnt[0]), .D(n328), .A(n329), .B(n330), .Y(n327)
         );
  AOI22X1 U531 ( .A(n66), .B(n119), .C(n67), .D(n105), .Y(n330) );
  NAND2X1 U532 ( .A(n371), .B(N160), .Y(n357) );
  ENOX1 U533 ( .A(new_rx_sync_cnt[0]), .B(n60), .C(new_rx_sync_cnt[0]), .D(
        n313), .Y(N348) );
  OAI211X1 U534 ( .C(n545), .D(n552), .A(ff_chg), .B(n115), .Y(n315) );
  OAI211X1 U535 ( .C(n316), .D(n107), .A(n317), .B(n318), .Y(n314) );
  AOI31X1 U536 ( .A(n319), .B(n107), .C(n320), .D(ui_intv_cnt[7]), .Y(n318) );
  BUFX3 U537 ( .A(n188), .Y(n18) );
  GEN2XL U538 ( .D(N142), .E(n243), .C(ui_intv_cnt[5]), .B(ui_intv_cnt[6]), 
        .A(ui_intv_cnt[7]), .Y(n188) );
  NAND4X1 U539 ( .A(n124), .B(n104), .C(n105), .D(n119), .Y(n243) );
  NOR2X1 U540 ( .A(N159), .B(N362), .Y(n376) );
  NOR43XL U541 ( .B(n119), .C(n122), .D(n477), .A(N141), .Y(n420) );
  NOR2X1 U542 ( .A(n107), .B(n478), .Y(n477) );
  AOI21X1 U543 ( .B(n367), .C(n471), .A(n115), .Y(n472) );
  NAND2X1 U544 ( .A(N159), .B(n106), .Y(n471) );
  XNOR2XL U545 ( .A(n220), .B(n128), .Y(n198) );
  XNOR2XL U546 ( .A(symb_cnt[4]), .B(symb_cnt[2]), .Y(n220) );
  XNOR2XL U547 ( .A(ui_intv_cnt[6]), .B(n144), .Y(n138) );
  XNOR2XL U548 ( .A(n152), .B(n153), .Y(n145) );
  XNOR2XL U549 ( .A(n13), .B(add_264_carry[5]), .Y(n152) );
  INVX1 U550 ( .A(symb_cnt[3]), .Y(n129) );
  XNOR2XL U551 ( .A(n104), .B(r_tui[0]), .Y(n524) );
  XNOR2XL U552 ( .A(n124), .B(r_tui[3]), .Y(n523) );
  NAND4X1 U553 ( .A(n295), .B(n91), .C(us_cnt_0_), .D(n531), .Y(n150) );
  NOR2X1 U554 ( .A(n89), .B(n92), .Y(n531) );
  XNOR2XL U555 ( .A(ui_intv_cnt[5]), .B(r_tui[5]), .Y(n529) );
  INVX1 U556 ( .A(ui_intv_cnt[6]), .Y(n107) );
  INVX1 U557 ( .A(ui_intv_cnt[7]), .Y(n118) );
  NAND2X1 U558 ( .A(symb_cnt[3]), .B(n225), .Y(n217) );
  OAI31XL U559 ( .A(n380), .B(n366), .C(n381), .D(n349), .Y(n351) );
  AOI21X1 U560 ( .B(N362), .C(n543), .A(n542), .Y(n381) );
  NOR2X1 U561 ( .A(n349), .B(symb_cnt[2]), .Y(n367) );
  NOR2X1 U562 ( .A(n150), .B(ui_intv_cnt[7]), .Y(n427) );
  NOR4XL U563 ( .A(n440), .B(n441), .C(n442), .D(n138), .Y(n439) );
  XNOR2XL U564 ( .A(n141), .B(ui_intv_cnt[0]), .Y(n441) );
  XNOR2XL U565 ( .A(ui_intv_cnt[1]), .B(n342), .Y(n440) );
  XNOR2XL U566 ( .A(N142), .B(n339), .Y(n442) );
  AOI21X1 U567 ( .B(n541), .C(N362), .A(N363), .Y(n366) );
  NAND2X1 U568 ( .A(r_tui[1]), .B(n70), .Y(n141) );
  AOI31X1 U569 ( .A(n57), .B(n362), .C(n363), .D(n364), .Y(n350) );
  AO21X1 U570 ( .B(n298), .C(n365), .A(n366), .Y(n363) );
  AO222X1 U571 ( .A(n546), .B(n351), .C(n94), .D(n551), .E(n554), .F(n361), 
        .Y(n362) );
  NAND3X1 U572 ( .A(N362), .B(n543), .C(n367), .Y(n365) );
  AOI32X1 U573 ( .A(n331), .B(n329), .C(ui_intv_cnt[2]), .D(n65), .E(N141), 
        .Y(n326) );
  NAND21X1 U574 ( .B(n402), .A(r_tui[0]), .Y(n401) );
  AOI21X1 U575 ( .B(n70), .C(n545), .A(n392), .Y(n402) );
  NAND2X1 U576 ( .A(N160), .B(symb_cnt[3]), .Y(n222) );
  NAND4X1 U577 ( .A(n427), .B(N142), .C(n104), .D(n105), .Y(n478) );
  INVX1 U578 ( .A(us_cnt_1_), .Y(n89) );
  INVX1 U579 ( .A(test_so), .Y(n92) );
  NAND2X1 U580 ( .A(ui_intv_cnt[5]), .B(n321), .Y(n320) );
  XNOR2XL U581 ( .A(N141), .B(n331), .Y(n443) );
  XNOR2XL U582 ( .A(rx_ui_5_8[4]), .B(N142), .Y(n146) );
  NOR4XL U583 ( .A(n543), .B(n129), .C(n380), .D(N160), .Y(n490) );
  NOR4XL U584 ( .A(n286), .B(n287), .C(n288), .D(n110), .Y(n525) );
  NAND2X1 U585 ( .A(ff_idn), .B(ff_chg), .Y(n286) );
  AOI31X1 U586 ( .A(fcp_state[2]), .B(fcp_state[1]), .C(n492), .D(n246), .Y(
        n287) );
  NOR42XL U587 ( .C(n479), .D(n107), .A(n119), .B(n478), .Y(n414) );
  XNOR2XL U588 ( .A(ui_intv_cnt[5]), .B(N141), .Y(n479) );
  NOR3XL U589 ( .A(n75), .B(n15), .C(n298), .Y(n513) );
  INVX1 U590 ( .A(us_cnt_2_), .Y(n91) );
  NOR32XL U591 ( .B(symb_cnt[5]), .C(n480), .A(n111), .Y(n473) );
  NAND3X1 U592 ( .A(n129), .B(n121), .C(n127), .Y(n480) );
  NOR21XL U593 ( .B(n539), .A(n302), .Y(N356) );
  XNOR2XL U594 ( .A(rxtx_buf[0]), .B(n303), .Y(n302) );
  XNOR2XL U595 ( .A(n304), .B(n305), .Y(n303) );
  XNOR2XL U596 ( .A(n306), .B(n307), .Y(n305) );
  AND4X1 U597 ( .A(n502), .B(n503), .C(n504), .D(n418), .Y(n481) );
  OAI21BBX1 U598 ( .A(n349), .B(n406), .C(n547), .Y(n503) );
  NAND4X1 U599 ( .A(ff_idn), .B(n444), .C(n9), .D(n117), .Y(n504) );
  NAND2X1 U600 ( .A(n277), .B(n546), .Y(n502) );
  XNOR2XL U601 ( .A(ui_intv_cnt[2]), .B(rx_ui_5_8[2]), .Y(n147) );
  INVX1 U602 ( .A(ff_idn), .Y(n76) );
  AND3X1 U603 ( .A(n11), .B(n367), .C(n543), .Y(n476) );
  NOR3XL U604 ( .A(n85), .B(new_rx_sync_cnt[0]), .C(n275), .Y(setsta[3]) );
  NAND3X1 U605 ( .A(fcp_state[0]), .B(n556), .C(n532), .Y(n279) );
  NAND3X1 U606 ( .A(n489), .B(n557), .C(fcp_state[2]), .Y(n273) );
  INVX1 U607 ( .A(symb_cnt[6]), .Y(n111) );
  NAND2X1 U608 ( .A(symb_cnt[3]), .B(n406), .Y(n149) );
  INVX1 U609 ( .A(r_ctl[7]), .Y(n544) );
  NAND2X1 U610 ( .A(n511), .B(n512), .Y(n498) );
  NAND4X1 U611 ( .A(n552), .B(n115), .C(n15), .D(n76), .Y(n512) );
  OAI21X1 U612 ( .B(n490), .C(n113), .A(n545), .Y(n511) );
  INVX1 U613 ( .A(rx_trans_8_chg), .Y(n87) );
  NOR3XL U614 ( .A(n272), .B(n76), .C(n273), .Y(setsta[6]) );
  NAND3X1 U615 ( .A(symb_cnt[6]), .B(n274), .C(ff_chg), .Y(n272) );
  XNOR2XL U616 ( .A(ui_intv_cnt[1]), .B(rx_ui_5_8[1]), .Y(n135) );
  XNOR2XL U617 ( .A(r_dat[7]), .B(n76), .Y(n344) );
  AND3X1 U618 ( .A(n545), .B(n245), .C(ff_idn), .Y(n284) );
  INVX1 U619 ( .A(new_rx_sync_cnt[1]), .Y(n85) );
  NAND42X1 U620 ( .C(n536), .D(n9), .A(n548), .B(n537), .Y(N1005) );
  AOI21BX1 U621 ( .C(n492), .B(fcp_state[2]), .A(n110), .Y(n537) );
  OAI211X1 U622 ( .C(n75), .D(n288), .A(ff_idn), .B(fcp_state[1]), .Y(n536) );
  XNOR2XL U623 ( .A(rxtx_buf[5]), .B(rxtx_buf[4]), .Y(n306) );
  XNOR2XL U624 ( .A(n308), .B(n309), .Y(n304) );
  XNOR2XL U625 ( .A(rxtx_buf[3]), .B(rxtx_buf[2]), .Y(n309) );
  XNOR2XL U626 ( .A(rxtx_buf[1]), .B(ff_idn), .Y(n308) );
  XNOR2XL U627 ( .A(rxtx_buf[7]), .B(rxtx_buf[6]), .Y(n307) );
  OAI32X1 U628 ( .A(n275), .B(rx_trans_8_chg), .C(n149), .D(ff_chg), .E(n87), 
        .Y(n516) );
  OAI32X1 U629 ( .A(n91), .B(test_so), .C(n294), .D(n92), .E(n289), .Y(N88) );
  OAI22X1 U630 ( .A(n289), .B(n91), .C(us_cnt_2_), .D(n294), .Y(N87) );
  INVX1 U631 ( .A(r_ctl[1]), .Y(n73) );
  NAND2X1 U632 ( .A(r_ctl[0]), .B(n73), .Y(n261) );
  NAND4X1 U633 ( .A(us_cnt_1_), .B(us_cnt_0_), .C(n150), .D(n295), .Y(n294) );
  INVX1 U634 ( .A(r_ctl[0]), .Y(n74) );
  INVX1 U635 ( .A(us_cnt_0_), .Y(n90) );
  INVX1 U636 ( .A(rxtx_buf[1]), .Y(n82) );
  INVX1 U637 ( .A(rxtx_buf[2]), .Y(n83) );
  NOR2X1 U638 ( .A(us_cnt_0_), .B(n553), .Y(N85) );
  INVX1 U639 ( .A(rxtx_buf[0]), .Y(n86) );
  BUFX3 U640 ( .A(tx_en), .Y(r_ctl[6]) );
  NAND3X1 U641 ( .A(n299), .B(n300), .C(n550), .Y(tx_en) );
endmodule


module fcpegn_a0_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module fcpegn_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(SUM[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
endmodule


module fcpegn_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9555;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9555), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9555), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9555), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9555), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9555), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9555), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9555), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9555), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9555), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9573;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9573), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9573), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9573), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9573), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9573), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9573), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9573), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9573), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9573), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9591;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9591), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9591), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9591), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9591), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9591), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9591), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9591), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9591), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9591), 
        .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_0 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_0 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[1]), .Y(n9) );
  INVX1 U4 ( .A(set2[4]), .Y(n11) );
  NAND3X1 U5 ( .A(n15), .B(n12), .C(n16), .Y(n21) );
  INVX1 U6 ( .A(set2[0]), .Y(n10) );
  INVX1 U7 ( .A(set2[2]), .Y(n14) );
  INVX1 U8 ( .A(set2[3]), .Y(n13) );
  INVX1 U9 ( .A(set2[7]), .Y(n12) );
  NOR2X1 U10 ( .A(rdat[6]), .B(n15), .Y(irq[6]) );
  NOR2X1 U11 ( .A(rdat[7]), .B(n12), .Y(irq[7]) );
  AOI211X1 U12 ( .C(n10), .D(n8), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U13 ( .A(rdat[0]), .Y(n8) );
  AOI211X1 U14 ( .C(n9), .D(n7), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U15 ( .A(rdat[1]), .Y(n7) );
  AOI211X1 U16 ( .C(n14), .D(n6), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U17 ( .A(rdat[2]), .Y(n6) );
  AOI211X1 U18 ( .C(n13), .D(n5), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U19 ( .A(rdat[3]), .Y(n5) );
  AOI211X1 U20 ( .C(n11), .D(n4), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U21 ( .A(rdat[4]), .Y(n4) );
  AOI211X1 U22 ( .C(n16), .D(n3), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U23 ( .A(rdat[5]), .Y(n3) );
  AOI211X1 U24 ( .C(n15), .D(n2), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U25 ( .A(rdat[6]), .Y(n2) );
  AOI211X1 U26 ( .C(n12), .D(n1), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U27 ( .A(rdat[7]), .Y(n1) );
  NAND4X1 U28 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U29 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U30 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U31 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR2X1 U32 ( .A(rdat[0]), .B(n10), .Y(irq[0]) );
  NOR2X1 U33 ( .A(rdat[1]), .B(n9), .Y(irq[1]) );
  NOR2X1 U34 ( .A(rdat[4]), .B(n11), .Y(irq[4]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n14), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[3]), .B(n13), .Y(irq[3]) );
  INVX1 U37 ( .A(set2[6]), .Y(n15) );
  INVX1 U38 ( .A(set2[5]), .Y(n16) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9609;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9609), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9609), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9609), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9609), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9609), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9609), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9609), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9609), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9609), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000000 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9627;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9627), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9627), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9627), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9627), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9627), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9627), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9627), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9627), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9627), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dpdmacc_a0 ( dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, r_wdat, r_acc, 
        r_dpdmsta, r_dm, r_dmchg, r_int, clk, rstz, test_si, test_se );
  input [7:0] r_wdat;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, clk, rstz, test_si, test_se;
  output r_dm, r_dmchg, r_int;
  wire   dp_chg, dp_rise, dm_fall, dp_active_acc, dp_inacti_acc, dm_active_acc,
         dm_inacti_acc, upd00, n3, n4, n5, n6, n28, n29, n30, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n31,
         n32, n33, n34, n35, n36, n37, n38, n2, n7, n8, n9, n10, n11, n39;
  wire   [7:0] wd00;

  INVX1 U4 ( .A(n6), .Y(n4) );
  INVX1 U5 ( .A(n6), .Y(n3) );
  INVX1 U6 ( .A(n6), .Y(n5) );
  INVX1 U7 ( .A(rstz), .Y(n6) );
  ff_sync_2 u0_dpsync ( .i_org(dp_comp), .o_dbc(r_dpdmsta[6]), .o_chg(dp_chg), 
        .clk(clk), .rstz(n4), .test_si(n28), .test_se(test_se) );
  ff_sync_1 u0_dmsync ( .i_org(dm_comp), .o_dbc(r_dm), .o_chg(r_dmchg), .clk(
        clk), .rstz(n4), .test_si(n30), .test_so(n29), .test_se(test_se) );
  ff_sync_0 u0_idsync ( .i_org(id_comp), .o_dbc(r_dpdmsta[5]), .o_chg(), .clk(
        clk), .rstz(n5), .test_si(r_dpdmsta[6]), .test_se(test_se) );
  filter150us_a0_1 u0_dpfltr ( .active_hit(dp_active_acc), .inacti_hit(
        dp_inacti_acc), .start_edge(dp_rise), .any_edge(dp_chg), .clk(clk), 
        .rstz(n5), .test_si(r_dpdmsta[4]), .test_so(n28), .test_se(test_se) );
  filter150us_a0_0 u0_dmfltr ( .active_hit(dm_active_acc), .inacti_hit(
        dm_inacti_acc), .start_edge(dm_fall), .any_edge(r_dmchg), .clk(clk), 
        .rstz(n5), .test_si(r_acc[7]), .test_so(n30), .test_se(test_se) );
  glreg_a0_5 u0_accmltr ( .clk(clk), .arstz(n3), .we(upd00), .wdat(wd00), 
        .rdat(r_acc), .test_si(test_si), .test_se(test_se) );
  glreg_WIDTH5_0 u0_dpdmsta ( .clk(clk), .arstz(n4), .we(r_wr_1), .wdat(
        r_wdat[4:0]), .rdat(r_dpdmsta[4:0]), .test_si(n29), .test_se(test_se)
         );
  INVX1 U3 ( .A(r_re_0), .Y(n39) );
  NAND2X1 U8 ( .A(n33), .B(n39), .Y(upd00) );
  NOR2X1 U9 ( .A(n2), .B(n8), .Y(n33) );
  OAI22X1 U10 ( .A(n39), .B(n27), .C(r_re_0), .D(n31), .Y(wd00[0]) );
  XNOR2XL U11 ( .A(n26), .B(n11), .Y(n31) );
  OAI22X1 U12 ( .A(n18), .B(n39), .C(r_re_0), .D(n19), .Y(wd00[4]) );
  XNOR2XL U13 ( .A(n17), .B(n10), .Y(n19) );
  INVX1 U14 ( .A(n27), .Y(n8) );
  INVX1 U15 ( .A(n18), .Y(n2) );
  NOR2X1 U16 ( .A(n17), .B(n10), .Y(n15) );
  NOR2X1 U17 ( .A(n26), .B(n11), .Y(n24) );
  OAI21X1 U18 ( .B(n33), .C(n39), .A(n34), .Y(r_int) );
  AOI33X1 U19 ( .A(n8), .B(n11), .C(n35), .D(n2), .E(n10), .F(n36), .Y(n34) );
  NOR3XL U20 ( .A(r_acc[5]), .B(r_acc[7]), .C(r_acc[6]), .Y(n36) );
  AOI21BX1 U21 ( .C(r_acc[3]), .B(n21), .A(r_re_0), .Y(wd00[3]) );
  NAND21X1 U22 ( .B(n22), .A(r_acc[2]), .Y(n21) );
  AOI21BX1 U23 ( .C(r_acc[7]), .B(n12), .A(r_re_0), .Y(wd00[7]) );
  NAND21X1 U24 ( .B(n13), .A(r_acc[6]), .Y(n12) );
  NOR2X1 U25 ( .A(r_re_0), .B(n25), .Y(wd00[1]) );
  XNOR2XL U26 ( .A(r_acc[1]), .B(n24), .Y(n25) );
  NOR2X1 U27 ( .A(r_re_0), .B(n23), .Y(wd00[2]) );
  XOR2X1 U28 ( .A(n22), .B(r_acc[2]), .Y(n23) );
  NOR2X1 U29 ( .A(r_re_0), .B(n16), .Y(wd00[5]) );
  XNOR2XL U30 ( .A(r_acc[5]), .B(n15), .Y(n16) );
  NOR2X1 U31 ( .A(r_re_0), .B(n14), .Y(wd00[6]) );
  XOR2X1 U32 ( .A(n13), .B(r_acc[6]), .Y(n14) );
  OAI21X1 U33 ( .B(dm_inacti_acc), .C(n7), .A(n38), .Y(n18) );
  OAI21BX1 U34 ( .C(dm_active_acc), .B(r_dm), .A(n7), .Y(n38) );
  INVX1 U35 ( .A(r_dpdmsta[1]), .Y(n7) );
  OAI21X1 U36 ( .B(dp_inacti_acc), .C(n9), .A(n37), .Y(n27) );
  OAI21BBX1 U37 ( .A(r_dpdmsta[6]), .B(dp_active_acc), .C(n9), .Y(n37) );
  INVX1 U38 ( .A(r_dpdmsta[0]), .Y(n9) );
  AND2X1 U39 ( .A(r_dmchg), .B(r_dm), .Y(dm_fall) );
  NOR21XL U40 ( .B(dp_chg), .A(r_dpdmsta[6]), .Y(dp_rise) );
  NAND2X1 U41 ( .A(n2), .B(n20), .Y(n17) );
  NAND4X1 U42 ( .A(r_acc[6]), .B(r_acc[5]), .C(r_acc[4]), .D(r_acc[7]), .Y(n20) );
  NAND2X1 U43 ( .A(n15), .B(r_acc[5]), .Y(n13) );
  INVX1 U44 ( .A(r_acc[0]), .Y(n11) );
  NOR3XL U45 ( .A(r_acc[1]), .B(r_acc[3]), .C(r_acc[2]), .Y(n35) );
  NAND2X1 U46 ( .A(n8), .B(n32), .Y(n26) );
  NAND4X1 U47 ( .A(r_acc[2]), .B(r_acc[1]), .C(r_acc[0]), .D(r_acc[3]), .Y(n32) );
  NAND2X1 U48 ( .A(n24), .B(r_acc[1]), .Y(n22) );
  INVX1 U49 ( .A(r_acc[4]), .Y(n10) );
  BUFX3 U50 ( .A(r_dm), .Y(r_dpdmsta[7]) );
endmodule


module glreg_WIDTH5_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9645;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9645), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9645), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9645), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9645), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9645), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9645), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9663;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9663), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9663), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9663), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9663), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9663), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9663), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9663), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9663), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9663), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_0 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz, test_si, test_so, test_se );
  input start_edge, any_edge, clk, rstz, test_si, test_se;
  output active_hit, inacti_hit, test_so;
  wire   dbcnt_10_, dbcnt_9_, dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_,
         dbcnt_3_, dbcnt_2_, dbcnt_1_, dbcnt_0_, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, net9681, n2, n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n4, n14;

  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9681), .TE(test_se) );
  filter150us_a0_0_DW01_inc_0 add_76 ( .A({test_so, dbcnt_10_, dbcnt_9_, 
        dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_, dbcnt_3_, dbcnt_2_, 
        dbcnt_1_, dbcnt_0_}), .SUM({N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12}) );
  SDFFRQX1 dbcnt_reg_4_ ( .D(N29), .SIN(dbcnt_3_), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_4_) );
  SDFFRQX1 dbcnt_reg_3_ ( .D(N28), .SIN(dbcnt_2_), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_3_) );
  SDFFRQX1 dbcnt_reg_11_ ( .D(N36), .SIN(dbcnt_10_), .SMC(test_se), .C(net9681), .XR(n2), .Q(test_so) );
  SDFFRQX1 dbcnt_reg_2_ ( .D(N27), .SIN(dbcnt_1_), .SMC(test_se), .C(net9681), 
        .XR(rstz), .Q(dbcnt_2_) );
  SDFFRQX1 dbcnt_reg_1_ ( .D(N26), .SIN(dbcnt_0_), .SMC(test_se), .C(net9681), 
        .XR(rstz), .Q(dbcnt_1_) );
  SDFFRQX1 dbcnt_reg_0_ ( .D(N25), .SIN(test_si), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_0_) );
  SDFFRQX1 dbcnt_reg_7_ ( .D(N32), .SIN(dbcnt_6_), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_7_) );
  SDFFRQX1 dbcnt_reg_5_ ( .D(N30), .SIN(dbcnt_4_), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_5_) );
  SDFFRQX1 dbcnt_reg_6_ ( .D(N31), .SIN(dbcnt_5_), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_6_) );
  SDFFRQX1 dbcnt_reg_9_ ( .D(N34), .SIN(dbcnt_8_), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_9_) );
  SDFFRQX1 dbcnt_reg_8_ ( .D(N33), .SIN(dbcnt_7_), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_8_) );
  SDFFRQX1 dbcnt_reg_10_ ( .D(N35), .SIN(dbcnt_9_), .SMC(test_se), .C(net9681), 
        .XR(n2), .Q(dbcnt_10_) );
  BUFX3 U3 ( .A(n9), .Y(n1) );
  INVX1 U6 ( .A(any_edge), .Y(n14) );
  AND2X1 U7 ( .A(N22), .B(n9), .Y(N35) );
  AND2X1 U8 ( .A(N20), .B(n9), .Y(N33) );
  AND2X1 U9 ( .A(N21), .B(n9), .Y(N34) );
  NOR3XL U10 ( .A(n11), .B(any_edge), .C(n4), .Y(n9) );
  AND2X1 U11 ( .A(N16), .B(n9), .Y(N29) );
  AND2X1 U12 ( .A(N15), .B(n9), .Y(N28) );
  AND2X1 U13 ( .A(N19), .B(n9), .Y(N32) );
  AND2X1 U14 ( .A(N17), .B(n9), .Y(N30) );
  AND2X1 U15 ( .A(N18), .B(n9), .Y(N31) );
  AND2X1 U16 ( .A(N14), .B(n1), .Y(N27) );
  AND2X1 U17 ( .A(N13), .B(n1), .Y(N26) );
  INVX1 U18 ( .A(n5), .Y(n4) );
  OR2X1 U19 ( .A(n1), .B(any_edge), .Y(N24) );
  AOI211X1 U20 ( .C(n5), .D(n6), .A(n14), .B(start_edge), .Y(inacti_hit) );
  AOI21X1 U21 ( .B(n7), .C(n8), .A(test_so), .Y(n5) );
  NAND32X1 U22 ( .B(dbcnt_4_), .C(dbcnt_3_), .A(n13), .Y(n7) );
  NOR3XL U23 ( .A(dbcnt_5_), .B(dbcnt_7_), .C(dbcnt_6_), .Y(n13) );
  AND3X1 U24 ( .A(dbcnt_8_), .B(dbcnt_10_), .C(dbcnt_9_), .Y(n8) );
  NOR3XL U25 ( .A(n6), .B(test_so), .C(n7), .Y(active_hit) );
  NAND4X1 U26 ( .A(dbcnt_2_), .B(dbcnt_1_), .C(dbcnt_0_), .D(n8), .Y(n6) );
  AND2X1 U27 ( .A(N23), .B(n1), .Y(N36) );
  NOR4XL U28 ( .A(dbcnt_0_), .B(dbcnt_10_), .C(n7), .D(n12), .Y(n11) );
  OR4X1 U29 ( .A(dbcnt_9_), .B(dbcnt_8_), .C(dbcnt_2_), .D(dbcnt_1_), .Y(n12)
         );
  OAI21BBX1 U30 ( .A(N12), .B(n9), .C(n10), .Y(N25) );
  OAI21X1 U31 ( .B(n11), .C(n4), .A(any_edge), .Y(n10) );
endmodule


module filter150us_a0_0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_1 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz, test_si, test_so, test_se );
  input start_edge, any_edge, clk, rstz, test_si, test_se;
  output active_hit, inacti_hit, test_so;
  wire   dbcnt_10_, dbcnt_9_, dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_,
         dbcnt_3_, dbcnt_2_, dbcnt_1_, dbcnt_0_, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, net9699, n2, n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n1, n4, n14;

  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9699), .TE(test_se) );
  filter150us_a0_1_DW01_inc_0 add_76 ( .A({test_so, dbcnt_10_, dbcnt_9_, 
        dbcnt_8_, dbcnt_7_, dbcnt_6_, dbcnt_5_, dbcnt_4_, dbcnt_3_, dbcnt_2_, 
        dbcnt_1_, dbcnt_0_}), .SUM({N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12}) );
  SDFFRQX1 dbcnt_reg_4_ ( .D(N29), .SIN(dbcnt_3_), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_4_) );
  SDFFRQX1 dbcnt_reg_3_ ( .D(N28), .SIN(dbcnt_2_), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_3_) );
  SDFFRQX1 dbcnt_reg_11_ ( .D(N36), .SIN(dbcnt_10_), .SMC(test_se), .C(net9699), .XR(n2), .Q(test_so) );
  SDFFRQX1 dbcnt_reg_2_ ( .D(N27), .SIN(dbcnt_1_), .SMC(test_se), .C(net9699), 
        .XR(rstz), .Q(dbcnt_2_) );
  SDFFRQX1 dbcnt_reg_1_ ( .D(N26), .SIN(dbcnt_0_), .SMC(test_se), .C(net9699), 
        .XR(rstz), .Q(dbcnt_1_) );
  SDFFRQX1 dbcnt_reg_0_ ( .D(N25), .SIN(test_si), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_0_) );
  SDFFRQX1 dbcnt_reg_7_ ( .D(N32), .SIN(dbcnt_6_), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_7_) );
  SDFFRQX1 dbcnt_reg_5_ ( .D(N30), .SIN(dbcnt_4_), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_5_) );
  SDFFRQX1 dbcnt_reg_6_ ( .D(N31), .SIN(dbcnt_5_), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_6_) );
  SDFFRQX1 dbcnt_reg_9_ ( .D(N34), .SIN(dbcnt_8_), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_9_) );
  SDFFRQX1 dbcnt_reg_8_ ( .D(N33), .SIN(dbcnt_7_), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_8_) );
  SDFFRQX1 dbcnt_reg_10_ ( .D(N35), .SIN(dbcnt_9_), .SMC(test_se), .C(net9699), 
        .XR(n2), .Q(dbcnt_10_) );
  BUFX3 U3 ( .A(n9), .Y(n1) );
  INVX1 U6 ( .A(any_edge), .Y(n14) );
  AND2X1 U7 ( .A(N22), .B(n9), .Y(N35) );
  AND2X1 U8 ( .A(N20), .B(n9), .Y(N33) );
  AND2X1 U9 ( .A(N21), .B(n9), .Y(N34) );
  NOR3XL U10 ( .A(n11), .B(any_edge), .C(n4), .Y(n9) );
  AND2X1 U11 ( .A(N15), .B(n9), .Y(N28) );
  AND2X1 U12 ( .A(N19), .B(n9), .Y(N32) );
  AND2X1 U13 ( .A(N17), .B(n9), .Y(N30) );
  AND2X1 U14 ( .A(N18), .B(n9), .Y(N31) );
  AND2X1 U15 ( .A(N14), .B(n9), .Y(N27) );
  AND2X1 U16 ( .A(N13), .B(n1), .Y(N26) );
  AND2X1 U17 ( .A(N16), .B(n1), .Y(N29) );
  INVX1 U18 ( .A(n5), .Y(n4) );
  OR2X1 U19 ( .A(n1), .B(any_edge), .Y(N24) );
  AOI211X1 U20 ( .C(n5), .D(n6), .A(n14), .B(start_edge), .Y(inacti_hit) );
  AOI21X1 U21 ( .B(n7), .C(n8), .A(test_so), .Y(n5) );
  NAND32X1 U22 ( .B(dbcnt_4_), .C(dbcnt_3_), .A(n13), .Y(n7) );
  NOR3XL U23 ( .A(dbcnt_5_), .B(dbcnt_7_), .C(dbcnt_6_), .Y(n13) );
  AND3X1 U24 ( .A(dbcnt_8_), .B(dbcnt_10_), .C(dbcnt_9_), .Y(n8) );
  NOR3XL U25 ( .A(n6), .B(test_so), .C(n7), .Y(active_hit) );
  NAND4X1 U26 ( .A(dbcnt_2_), .B(dbcnt_1_), .C(dbcnt_0_), .D(n8), .Y(n6) );
  AND2X1 U27 ( .A(N23), .B(n1), .Y(N36) );
  NOR4XL U28 ( .A(dbcnt_0_), .B(dbcnt_10_), .C(n7), .D(n12), .Y(n11) );
  OR4X1 U29 ( .A(dbcnt_9_), .B(dbcnt_8_), .C(dbcnt_2_), .D(dbcnt_1_), .Y(n12)
         );
  OAI21BBX1 U30 ( .A(N12), .B(n9), .C(n10), .Y(N25) );
  OAI21X1 U31 ( .B(n11), .C(n4), .A(any_edge), .Y(n10) );
endmodule


module filter150us_a0_1_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ff_sync_0 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg;
  wire   d_org_0_;

  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_1 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  INVX1 U3 ( .A(test_so), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(o_dbc) );
  XOR2X1 U5 ( .A(d_org_0_), .B(test_so), .Y(o_chg) );
endmodule


module ff_sync_2 ( i_org, o_dbc, o_chg, clk, rstz, test_si, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg;
  wire   d_org_0_;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module dacmux_a0 ( clk, srstz, i_comp, r_comp_opt, r_wdat, r_adofs, r_isofs, 
        r_wr, dacv_wr, o_dacv, o_shrst, o_hold, o_dac1, o_daci_sel, o_dat, 
        r_dac_en, r_sar_en, o_dactl, o_cmpsta, x_daclsb, o_intr, o_smpl, 
        test_si2, test_si1, test_so1, test_se );
  input [2:0] r_comp_opt;
  input [7:0] r_wdat;
  output [7:0] r_adofs;
  output [7:0] r_isofs;
  input [10:0] r_wr;
  input [17:0] dacv_wr;
  output [143:0] o_dacv;
  output [9:0] o_dac1;
  output [17:0] o_daci_sel;
  output [17:0] o_dat;
  output [17:0] r_dac_en;
  output [17:0] r_sar_en;
  output [7:0] o_dactl;
  output [7:0] o_cmpsta;
  output [5:0] x_daclsb;
  output [4:0] o_smpl;
  input clk, srstz, i_comp, test_si2, test_si1, test_se;
  output o_shrst, o_hold, o_intr, test_so1;
  wire   n570, n578, dacyc_done, updcmp, semi_start, sacyc_done, sar_ini,
         sar_nxt, ps_sample, sampl_begn, sampl_done, ps_md4ch, updlsb, N1239,
         N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1250, N1251,
         N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1261, N1262, N1263,
         N1264, N1265, N1266, N1267, N1268, N1269, N1272, N1273, N1274, N1275,
         N1276, N1277, N1278, N1279, N1280, N1283, N1284, N1285, N1286, N1287,
         N1288, N1289, N1290, N1291, N1294, N1295, N1296, N1297, N1298, N1299,
         N1300, N1301, N1302, N1305, N1306, N1307, N1308, N1309, N1310, N1311,
         N1312, N1313, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323,
         N1324, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335,
         N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1349,
         N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1360, N1361,
         N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1371, N1372, N1373,
         N1374, N1375, N1376, N1377, N1378, N1379, N1382, N1383, N1384, N1385,
         N1386, N1387, N1388, N1389, N1390, N1393, N1394, N1395, N1396, N1397,
         N1398, N1399, N1400, N1401, N1404, N1405, N1406, N1407, N1408, N1409,
         N1410, N1411, N1412, N1415, N1416, N1417, N1418, N1419, N1420, N1421,
         N1422, N1423, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433,
         N1434, n569, n577, n572, n576, n573, n571, n568, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n204, n205, n206, n574, n575, n64, n90, n91, n92, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n199, n200, n203, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n303, n304, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n457, n458, n459, n460, n461,
         n462, n463, n464, n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13,
         n15, n16, n17, n18, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n107, n110, n112, n113, n114, n115, n116, n117, n118, n120, n121,
         n122, n123, n124, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n201, n202, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n456,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567;
  wire   [1:0] syn_comp;
  wire   [4:0] cs_ptr;
  wire   [17:0] datcmp;
  wire   [4:0] ps_ptr;
  wire   [9:0] r_dac1v;
  wire   [9:0] r_rpt_v;
  wire   [17:0] app_dacis;
  wire   [17:0] pos_dacis;
  wire   [5:0] wdlsb;
  wire   [17:0] upd;
  wire   [7:6] wda;
  wire   [143:0] r_dacvs;
  wire   [7:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;

  INVX1 U196 ( .A(n204), .Y(n198) );
  INVX1 U200 ( .A(n204), .Y(n192) );
  INVX1 U201 ( .A(n204), .Y(n191) );
  INVX1 U202 ( .A(n205), .Y(n190) );
  INVX1 U203 ( .A(n206), .Y(n189) );
  INVX1 U204 ( .A(n206), .Y(n188) );
  INVX1 U205 ( .A(n205), .Y(n187) );
  INVX1 U206 ( .A(n204), .Y(n186) );
  INVX1 U207 ( .A(n205), .Y(n184) );
  INVX1 U208 ( .A(n205), .Y(n183) );
  INVX1 U209 ( .A(n206), .Y(n182) );
  INVX1 U210 ( .A(n204), .Y(n181) );
  INVX1 U211 ( .A(n205), .Y(n180) );
  INVX1 U212 ( .A(n206), .Y(n179) );
  INVX1 U213 ( .A(n205), .Y(n178) );
  INVX1 U214 ( .A(n205), .Y(n177) );
  INVX1 U215 ( .A(n206), .Y(n176) );
  INVX1 U216 ( .A(n206), .Y(n175) );
  INVX1 U217 ( .A(n206), .Y(n185) );
  INVX1 U218 ( .A(n206), .Y(n174) );
  INVX1 U219 ( .A(n205), .Y(n196) );
  INVX1 U220 ( .A(n205), .Y(n195) );
  INVX1 U221 ( .A(n205), .Y(n194) );
  INVX1 U222 ( .A(n204), .Y(n193) );
  INVX1 U223 ( .A(n206), .Y(n173) );
  INVX1 U224 ( .A(n204), .Y(n197) );
  INVX1 U225 ( .A(srstz), .Y(n204) );
  INVX1 U245 ( .A(n206), .Y(n172) );
  INVX1 U246 ( .A(srstz), .Y(n206) );
  INVX1 U247 ( .A(srstz), .Y(n205) );
  glreg_00000012 u0_compi ( .clk(clk), .arstz(n198), .we(updcmp), .wdat(datcmp), .rdat(o_dat), .test_si(o_cmpsta[7]), .test_se(test_se) );
  dac2sar_a0 u0_dac2sar ( .r_dac_t(o_dactl[3:2]), .r_dacyc(o_dactl[7]), 
        .r_sar10(n64), .sar_ini(sar_ini), .sar_nxt(sar_nxt), .semi_nxt(n90), 
        .auto_sar(n462), .busy(o_dactl[0]), .stop(n464), .sync_i(syn_comp[1]), 
        .ps_sample(ps_sample), .sampl_begn(sampl_begn), .sampl_done(sampl_done), .sh_rst(o_shrst), .dacyc_done(dacyc_done), .sacyc_done(sacyc_done), .dac_v(
        r_dac1v), .rpt_v(r_rpt_v), .clk(clk), .srstz(n198), .test_si2(
        o_dat[17]), .test_si1(test_si1), .test_so1(n575), .test_se(test_se) );
  shmux_00000005_00000012_00000012 u0_shmux ( .ps_md4ch(ps_md4ch), 
        .r_comp_swtch(r_comp_opt[2]), .r_semi(n92), .r_loop(o_dactl[1]), 
        .r_dac_en({r_dac_en[17:16], n9, r_dac_en[14:0]}), .wr_dacv(dacv_wr), 
        .busy(o_dactl[0]), .sh_hold(o_hold), .stop(n464), .semi_start(
        semi_start), .auto_start(n463), .mxcyc_done(n95), .sampl_begn(
        sampl_begn), .sampl_done(sampl_done), .app_dacis(app_dacis), 
        .pos_dacis(pos_dacis), .cs_ptr(cs_ptr), .ps_ptr(ps_ptr), .clk(clk), 
        .srstz(n198), .test_si2(r_sar_en[7]), .test_si1(o_shrst), .test_so1(
        test_so1), .test_se(test_se) );
  glreg_WIDTH7_1 u0_dactl ( .clk(clk), .arstz(n197), .we(n91), .wdat({
        r_wdat[7:5], n50, r_wdat[3:1]}), .rdat(o_dactl[7:1]), .test_si(
        x_daclsb[5]), .test_se(test_se) );
  glreg_a0_49 u0_dacen ( .clk(clk), .arstz(n172), .we(r_wr[1]), .wdat({
        r_wdat[7:1], n103}), .rdat(r_dac_en[7:0]), .test_si(n575), .test_se(
        test_se) );
  glreg_a0_48 u0_saren ( .clk(clk), .arstz(n173), .we(r_wr[2]), .wdat({
        r_wdat[7:2], n11, n104}), .rdat(r_sar_en[7:0]), .test_si(r_isofs[7]), 
        .test_se(test_se) );
  glreg_WIDTH6_2 u0_daclsb ( .clk(clk), .arstz(n198), .we(updlsb), .wdat(wdlsb), .rdat(x_daclsb), .test_si(r_dac_en[7]), .test_se(test_se) );
  glreg_a0_47 dacvs_0__u0 ( .clk(clk), .arstz(n174), .we(upd[0]), .wdat({n54, 
        n58, n461, n75, n459, n458, n457, n84}), .rdat(r_dacvs[7:0]), 
        .test_si(test_si2), .test_se(test_se) );
  glreg_a0_46 dacvs_1__u0 ( .clk(clk), .arstz(n185), .we(upd[1]), .wdat({wda, 
        n60, n75, n459, n458, n457, n84}), .rdat(r_dacvs[15:8]), .test_si(
        r_dacvs[7]), .test_se(test_se) );
  glreg_a0_45 dacvs_2__u0 ( .clk(clk), .arstz(n175), .we(upd[2]), .wdat({n54, 
        n58, n60, n75, n459, n458, n457, n85}), .rdat(r_dacvs[23:16]), 
        .test_si(r_dacvs[15]), .test_se(test_se) );
  glreg_a0_44 dacvs_3__u0 ( .clk(clk), .arstz(n176), .we(upd[3]), .wdat({wda, 
        n461, n75, n459, n458, n457, n85}), .rdat(r_dacvs[31:24]), .test_si(
        r_dacvs[23]), .test_se(test_se) );
  glreg_a0_43 dacvs_4__u0 ( .clk(clk), .arstz(n177), .we(upd[4]), .wdat({wda, 
        n461, n75, n65, n72, n80, n84}), .rdat(r_dacvs[39:32]), .test_si(
        r_dacvs[31]), .test_se(test_se) );
  glreg_a0_42 dacvs_5__u0 ( .clk(clk), .arstz(n178), .we(upd[5]), .wdat({wda, 
        n461, n74, n459, n458, n457, n84}), .rdat(r_dacvs[47:40]), .test_si(
        r_dacvs[39]), .test_se(test_se) );
  glreg_a0_41 dacvs_6__u0 ( .clk(clk), .arstz(n179), .we(upd[6]), .wdat({wda, 
        n461, n74, n459, n458, n457, n85}), .rdat(r_dacvs[55:48]), .test_si(
        r_dacvs[47]), .test_se(test_se) );
  glreg_a0_40 dacvs_7__u0 ( .clk(clk), .arstz(n180), .we(upd[7]), .wdat({wda, 
        n461, n75, n459, n458, n457, n85}), .rdat(r_dacvs[63:56]), .test_si(
        r_dacvs[55]), .test_se(test_se) );
  glreg_a0_39 dacvs_8__u0 ( .clk(clk), .arstz(n181), .we(upd[8]), .wdat({n54, 
        n58, n60, n74, n65, n72, n80, n84}), .rdat(r_dacvs[71:64]), .test_si(
        r_dacvs[63]), .test_se(test_se) );
  glreg_a0_38 dacvs_9__u0 ( .clk(clk), .arstz(n182), .we(upd[9]), .wdat({wda, 
        n461, n74, n65, n72, n80, n85}), .rdat(r_dacvs[79:72]), .test_si(
        r_dacvs[71]), .test_se(test_se) );
  glreg_a0_37 dacvs_10__u0 ( .clk(clk), .arstz(n183), .we(upd[10]), .wdat({wda, 
        n461, n75, n65, n72, n80, n85}), .rdat(r_dacvs[87:80]), .test_si(
        r_dacvs[79]), .test_se(test_se) );
  glreg_a0_36 dacvs_11__u0 ( .clk(clk), .arstz(n184), .we(upd[11]), .wdat({n54, 
        n58, n60, n74, n459, n458, n457, n84}), .rdat(r_dacvs[95:88]), 
        .test_si(r_dacvs[87]), .test_se(test_se) );
  glreg_a0_35 dacvs_12__u0 ( .clk(clk), .arstz(n186), .we(upd[12]), .wdat({wda, 
        n60, n75, n459, n458, n457, n85}), .rdat(r_dacvs[103:96]), .test_si(
        r_dacvs[95]), .test_se(test_se) );
  glreg_a0_34 dacvs_13__u0 ( .clk(clk), .arstz(n187), .we(upd[13]), .wdat({n54, 
        n58, n461, n75, n65, n72, n80, n85}), .rdat(r_dacvs[111:104]), 
        .test_si(r_dacvs[103]), .test_se(test_se) );
  glreg_a0_33 dacvs_14__u0 ( .clk(clk), .arstz(n188), .we(upd[14]), .wdat({n54, 
        n58, n60, n74, n65, n72, n80, n84}), .rdat(r_dacvs[119:112]), 
        .test_si(r_dacvs[111]), .test_se(test_se) );
  glreg_a0_32 dacvs_15__u0 ( .clk(clk), .arstz(n189), .we(upd[15]), .wdat({n54, 
        n58, n60, n74, n65, n72, n80, n84}), .rdat(r_dacvs[127:120]), 
        .test_si(r_dacvs[119]), .test_se(test_se) );
  glreg_a0_31 dacvs_16__u0 ( .clk(clk), .arstz(n190), .we(upd[16]), .wdat({n54, 
        n58, n60, n74, n65, n72, n80, n85}), .rdat(r_dacvs[135:128]), 
        .test_si(r_dacvs[127]), .test_se(test_se) );
  glreg_a0_30 dacvs_17__u0 ( .clk(clk), .arstz(n191), .we(upd[17]), .wdat({n54, 
        n58, n60, n74, n65, n72, n80, n84}), .rdat(r_dacvs[143:136]), 
        .test_si(r_dacvs[135]), .test_se(test_se) );
  glsta_a0_1 u0_cmpsta ( .clk(clk), .arstz(n192), .rst0(1'b0), .set2(setsta), 
        .clr1(clrsta), .rdat(o_cmpsta), .irq(r_irq), .test_si(r_adofs[7]), 
        .test_se(test_se) );
  glreg_a0_29 u0_adofs ( .clk(clk), .arstz(n193), .we(r_wr[5]), .wdat({
        r_wdat[7:2], n11, n104}), .rdat({n568, n569, n570, n571, n572, n573, 
        n576, n577}), .test_si(syn_comp[1]), .test_se(test_se) );
  glreg_a0_28 u0_isofs ( .clk(clk), .arstz(n194), .we(r_wr[6]), .wdat({
        r_wdat[7:1], n103}), .rdat(r_isofs), .test_si(o_dactl[7]), .test_se(
        test_se) );
  glreg_a0_27 u1_dacen ( .clk(clk), .arstz(n195), .we(r_wr[7]), .wdat({
        r_wdat[7:1], n104}), .rdat({n578, r_dac_en[14:8]}), .test_si(
        pos_dacis[17]), .test_se(test_se) );
  glreg_a0_26 u1_saren ( .clk(clk), .arstz(n196), .we(r_wr[8]), .wdat({
        r_wdat[7:1], n103}), .rdat(r_sar_en[15:8]), .test_si(n9), .test_se(
        test_se) );
  glreg_WIDTH2_1 u2_dacen ( .clk(clk), .arstz(n186), .we(r_wr[9]), .wdat({n11, 
        n103}), .rdat(r_dac_en[17:16]), .test_si(r_sar_en[15]), .test_so(n574), 
        .test_se(test_se) );
  glreg_WIDTH2_0 u2_saren ( .clk(clk), .arstz(n197), .we(r_wr[10]), .wdat({
        r_wdat[1], n104}), .rdat(r_sar_en[17:16]), .test_si(n574), .test_se(
        test_se) );
  dacmux_a0_DW01_add_0 add_235_I18 ( .A({1'b0, r_dacvs[143:136]}), .B({n124, 
        n121, r_adofs[6:5], n110, n18, r_adofs[2:1], n78}), .CI(1'b0), .SUM({
        N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426}), .CO()
         );
  dacmux_a0_DW01_add_3 add_235_I15 ( .A({1'b0, r_dacvs[119:112]}), .B({n123, 
        n121, n15, n13, r_adofs[4:1], n78}), .CI(1'b0), .SUM({N1401, N1400, 
        N1399, N1398, N1397, N1396, N1395, N1394, N1393}), .CO() );
  dacmux_a0_DW01_add_4 add_235_I14 ( .A({1'b0, r_dacvs[111:104]}), .B({n123, 
        n121, n569, n570, n110, n17, r_adofs[2:0]}), .CI(1'b0), .SUM({N1390, 
        N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382}), .CO() );
  dacmux_a0_DW01_add_5 add_235_I13 ( .A({1'b0, r_dacvs[103:96]}), .B({n123, 
        n121, r_adofs[6], n570, r_adofs[4:0]}), .CI(1'b0), .SUM({N1379, N1378, 
        N1377, N1376, N1375, N1374, N1373, N1372, N1371}), .CO() );
  dacmux_a0_DW01_add_6 add_235_I12 ( .A({1'b0, r_dacvs[95:88]}), .B({n124, 
        n121, n569, r_adofs[5], n110, r_adofs[3:1], n118}), .CI(1'b0), .SUM({
        N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360}), .CO()
         );
  dacmux_a0_DW01_add_7 add_235_I11 ( .A({1'b0, r_dacvs[87:80]}), .B({n123, 
        n121, n15, n13, r_adofs[4:0]}), .CI(1'b0), .SUM({N1357, N1356, N1355, 
        N1354, N1353, N1352, N1351, N1350, N1349}), .CO() );
  dacmux_a0_DW01_add_8 add_235_I10 ( .A({1'b0, r_dacvs[79:72]}), .B({n123, 
        n121, r_adofs[6], n570, n110, n17, r_adofs[2], n576, n117}), .CI(1'b0), 
        .SUM({N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338}), 
        .CO() );
  dacmux_a0_DW01_add_9 add_235_I9 ( .A({1'b0, r_dacvs[71:64]}), .B({n123, n121, 
        n15, r_adofs[5:1], n118}), .CI(1'b0), .SUM({N1335, N1334, N1333, N1332, 
        N1331, N1330, N1329, N1328, N1327}), .CO() );
  dacmux_a0_DW01_add_10 add_235_I8 ( .A({1'b0, r_dacvs[63:56]}), .B({n122, 
        n122, n15, n13, n110, n18, r_adofs[2:1], n117}), .CI(1'b0), .SUM({
        N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316}), .CO()
         );
  dacmux_a0_DW01_add_11 add_235_I7 ( .A({1'b0, r_dacvs[55:48]}), .B({n122, 
        n122, r_adofs[6], n13, r_adofs[4:3], n3, r_adofs[1], n117}), .CI(1'b0), 
        .SUM({N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305}), 
        .CO() );
  dacmux_a0_DW01_add_12 add_235_I6 ( .A({1'b0, r_dacvs[47:40]}), .B({n122, 
        n122, n15, n13, n110, n17, n3, n69, n118}), .CI(1'b0), .SUM({N1302, 
        N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294}), .CO() );
  dacmux_a0_DW01_add_13 add_235_I5 ( .A({1'b0, r_dacvs[39:32]}), .B({n123, 
        n122, n15, n13, r_adofs[4:3], n2, n69, n78}), .CI(1'b0), .SUM({N1291, 
        N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283}), .CO() );
  dacmux_a0_DW01_add_14 add_235_I4 ( .A({1'b0, r_dacvs[31:24]}), .B({n123, 
        n122, n569, r_adofs[5], n110, n18, n2, n69, n118}), .CI(1'b0), .SUM({
        N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272}), .CO()
         );
  dacmux_a0_DW01_add_15 add_235_I3 ( .A({1'b0, r_dacvs[23:16]}), .B({
        r_isofs[7], r_isofs}), .CI(1'b0), .SUM({N1269, N1268, N1267, N1266, 
        N1265, N1264, N1263, N1262, N1261}), .CO() );
  dacmux_a0_DW01_add_16 add_235_I2 ( .A({1'b0, r_dacvs[15:8]}), .B({n123, n122, 
        r_adofs[6], n13, r_adofs[4:3], n2, n69, r_adofs[0]}), .CI(1'b0), .SUM(
        {N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250}), 
        .CO() );
  dacmux_a0_DW01_add_17 add_235 ( .A({1'b0, r_dacvs[7:0]}), .B({n123, n122, 
        n569, r_adofs[5], n110, n18, n3, n69, n118}), .CI(1'b0), .SUM({N1247, 
        N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239}), .CO() );
  dacmux_a0_DW01_add_18 add_235_I16 ( .A({1'b0, r_dacvs[127:120]}), .B({n124, 
        n121, n569, n570, r_adofs[4:3], n1, n576, n78}), .CI(1'b0), .SUM({
        N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404}), .CO()
         );
  dacmux_a0_DW01_add_19 add_235_I17 ( .A({1'b0, r_dacvs[135:128]}), .B({n124, 
        n121, n569, r_adofs[5], n110, n18, n2, n68, n117}), .CI(1'b0), .SUM({
        N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415}), .CO()
         );
  SDFFQX1 syn_comp_reg_1_ ( .D(syn_comp[0]), .SIN(syn_comp[0]), .SMC(test_se), 
        .C(clk), .Q(syn_comp[1]) );
  SDFFQX1 syn_comp_reg_0_ ( .D(i_comp), .SIN(r_dacvs[143]), .SMC(test_se), .C(
        clk), .Q(syn_comp[0]) );
  BUFX6 U21 ( .A(n107), .Y(n1) );
  BUFXL U22 ( .A(n107), .Y(n2) );
  BUFXL U23 ( .A(n107), .Y(n3) );
  BUFX6 U24 ( .A(n573), .Y(n107) );
  AO21X1 U25 ( .B(N1416), .C(n48), .A(n45), .Y(o_dacv[129]) );
  NOR21X1 U26 ( .B(n126), .A(n524), .Y(n45) );
  INVX4 U27 ( .A(r_wdat[4]), .Y(n238) );
  INVX4 U28 ( .A(n577), .Y(n120) );
  INVX1 U29 ( .A(n127), .Y(n121) );
  INVX1 U30 ( .A(n568), .Y(n127) );
  INVX1 U31 ( .A(n488), .Y(n489) );
  BUFX3 U32 ( .A(n571), .Y(r_adofs[4]) );
  NOR21X2 U33 ( .B(n126), .A(n509), .Y(n6) );
  INVX1 U34 ( .A(o_dactl[4]), .Y(n46) );
  AO21X1 U35 ( .B(N1411), .C(n523), .A(n522), .Y(o_dacv[127]) );
  INVX2 U36 ( .A(N1346), .Y(n509) );
  INVX1 U37 ( .A(N1434), .Y(n527) );
  MUX2X1 U38 ( .D0(n256), .D1(n255), .S(ps_ptr[3]), .Y(n257) );
  GEN2XL U39 ( .D(n425), .E(n424), .C(n423), .B(n432), .A(n422), .Y(n471) );
  INVXL U40 ( .A(N1357), .Y(n4) );
  AO21X1 U41 ( .B(N1396), .C(n520), .A(n519), .Y(o_dacv[115]) );
  INVX1 U42 ( .A(N1401), .Y(n520) );
  INVX3 U43 ( .A(N1379), .Y(n514) );
  NAND21X1 U44 ( .B(n124), .A(N1434), .Y(n525) );
  INVX3 U45 ( .A(N1423), .Y(n524) );
  NAND21X1 U46 ( .B(r_adofs[7]), .A(N1390), .Y(n515) );
  INVX2 U47 ( .A(N1390), .Y(n517) );
  AO21X1 U48 ( .B(N1327), .C(n508), .A(n507), .Y(o_dacv[64]) );
  INVX1 U49 ( .A(n576), .Y(n105) );
  BUFX3 U50 ( .A(n572), .Y(r_adofs[3]) );
  AND3X1 U51 ( .A(n549), .B(n550), .C(n556), .Y(n5) );
  INVXL U52 ( .A(n578), .Y(n7) );
  INVXL U53 ( .A(n7), .Y(r_dac_en[15]) );
  INVXL U54 ( .A(n7), .Y(n9) );
  INVXL U55 ( .A(r_wdat[1]), .Y(n10) );
  INVXL U56 ( .A(n10), .Y(n11) );
  INVXL U57 ( .A(n570), .Y(n12) );
  INVXL U58 ( .A(n12), .Y(n13) );
  INVXL U59 ( .A(n38), .Y(r_adofs[6]) );
  INVXL U60 ( .A(n38), .Y(n15) );
  INVXL U61 ( .A(n572), .Y(n16) );
  INVXL U62 ( .A(n16), .Y(n17) );
  INVXL U63 ( .A(n16), .Y(n18) );
  INVXL U64 ( .A(n12), .Y(r_adofs[5]) );
  INVXL U65 ( .A(n569), .Y(n38) );
  INVXL U66 ( .A(n414), .Y(n39) );
  INVXL U67 ( .A(n414), .Y(n40) );
  AO21XL U68 ( .B(N1400), .C(n520), .A(n519), .Y(o_dacv[119]) );
  NAND21XL U69 ( .B(n481), .A(n480), .Y(o_smpl[4]) );
  NAND4XL U70 ( .A(n321), .B(n312), .C(n311), .D(n421), .Y(n98) );
  AO21X1 U71 ( .B(N1377), .C(n514), .A(n43), .Y(o_dacv[102]) );
  AO21X1 U72 ( .B(N1366), .C(n513), .A(n512), .Y(o_dacv[94]) );
  INVX1 U73 ( .A(N1368), .Y(n513) );
  AO21X1 U74 ( .B(N1364), .C(n513), .A(n512), .Y(o_dacv[92]) );
  INVX2 U75 ( .A(n511), .Y(n512) );
  NOR21X1 U76 ( .B(n126), .A(n524), .Y(n44) );
  NOR21X2 U77 ( .B(n126), .A(n514), .Y(n43) );
  NOR21X4 U78 ( .B(n126), .A(n510), .Y(n41) );
  INVX2 U79 ( .A(N1357), .Y(n510) );
  NOR21XL U80 ( .B(n126), .A(n514), .Y(n42) );
  AO21XL U81 ( .B(N1399), .C(n520), .A(n519), .Y(o_dacv[118]) );
  AO21XL U82 ( .B(N1397), .C(n520), .A(n519), .Y(o_dacv[116]) );
  AO21XL U83 ( .B(N1393), .C(n520), .A(n519), .Y(o_dacv[112]) );
  AO21XL U84 ( .B(N1331), .C(n508), .A(n507), .Y(o_dacv[68]) );
  NAND21XL U85 ( .B(r_adofs[7]), .A(N1368), .Y(n511) );
  NAND21X2 U86 ( .B(r_adofs[7]), .A(N1335), .Y(n506) );
  INVX2 U87 ( .A(N1335), .Y(n508) );
  INVX2 U88 ( .A(n515), .Y(n516) );
  AO21X1 U89 ( .B(N1330), .C(n508), .A(n507), .Y(o_dacv[67]) );
  MUX2IX2 U90 ( .D0(n238), .D1(n46), .S(n250), .Y(ps_sample) );
  AO21X1 U91 ( .B(N1333), .C(n508), .A(n507), .Y(o_dacv[70]) );
  INVXL U92 ( .A(n524), .Y(n47) );
  INVXL U93 ( .A(n47), .Y(n48) );
  INVX3 U94 ( .A(n506), .Y(n507) );
  INVX4 U95 ( .A(n120), .Y(n78) );
  INVX3 U96 ( .A(n518), .Y(n519) );
  INVX3 U97 ( .A(n120), .Y(r_adofs[0]) );
  INVX3 U98 ( .A(n120), .Y(n117) );
  INVX3 U99 ( .A(n120), .Y(n118) );
  OAI21BBXL U100 ( .A(n104), .B(o_dactl[0]), .C(r_wr[0]), .Y(n49) );
  AND2XL U101 ( .A(r_wdat[4]), .B(r_wr[4]), .Y(clrsta[4]) );
  INVXL U102 ( .A(n49), .Y(n91) );
  INVX1 U103 ( .A(n238), .Y(n50) );
  INVXL U104 ( .A(dacv_wr[14]), .Y(n535) );
  AOI21X1 U105 ( .B(n92), .C(dacyc_done), .A(sacyc_done), .Y(n545) );
  INVX1 U106 ( .A(n545), .Y(n51) );
  INVX1 U107 ( .A(n545), .Y(n52) );
  INVX1 U108 ( .A(wda[7]), .Y(n53) );
  INVX1 U109 ( .A(n53), .Y(n54) );
  BUFX3 U110 ( .A(n338), .Y(n55) );
  BUFX3 U111 ( .A(n335), .Y(n56) );
  INVX1 U112 ( .A(wda[6]), .Y(n57) );
  INVX1 U113 ( .A(n57), .Y(n58) );
  INVX1 U114 ( .A(n461), .Y(n59) );
  INVX1 U115 ( .A(n59), .Y(n60) );
  BUFX3 U116 ( .A(n333), .Y(n61) );
  BUFX3 U117 ( .A(n337), .Y(n62) );
  INVX1 U118 ( .A(n459), .Y(n63) );
  INVX1 U119 ( .A(n63), .Y(n65) );
  NOR2X1 U120 ( .A(n155), .B(n565), .Y(n66) );
  INVX1 U121 ( .A(r_wr[3]), .Y(n67) );
  INVXL U122 ( .A(n105), .Y(n68) );
  INVX1 U123 ( .A(n105), .Y(n69) );
  NOR2X1 U124 ( .A(n155), .B(cs_ptr[1]), .Y(n70) );
  INVX1 U125 ( .A(n458), .Y(n71) );
  INVX1 U126 ( .A(n71), .Y(n72) );
  BUFX3 U127 ( .A(n334), .Y(n73) );
  BUFX3 U128 ( .A(n202), .Y(n460) );
  INVX1 U129 ( .A(n460), .Y(n74) );
  INVX1 U130 ( .A(n460), .Y(n75) );
  INVX1 U131 ( .A(n199), .Y(n76) );
  AO21X1 U132 ( .B(n274), .C(n273), .A(n272), .Y(sar_ini) );
  NOR2X1 U133 ( .A(n150), .B(cs_ptr[1]), .Y(n77) );
  INVX1 U134 ( .A(n457), .Y(n79) );
  INVX1 U135 ( .A(n79), .Y(n80) );
  NOR2X1 U136 ( .A(n147), .B(n565), .Y(n81) );
  NOR2X1 U137 ( .A(o_dactl[0]), .B(semi_start), .Y(n141) );
  INVX1 U138 ( .A(n141), .Y(n82) );
  INVX1 U139 ( .A(n141), .Y(n83) );
  MUX2IX1 U140 ( .D0(r_rpt_v[2]), .D1(n104), .S(n136), .Y(n88) );
  INVX1 U141 ( .A(n88), .Y(n84) );
  INVX1 U142 ( .A(n88), .Y(n85) );
  BUFX12 U143 ( .A(n573), .Y(r_adofs[2]) );
  BUFX6 U144 ( .A(n576), .Y(r_adofs[1]) );
  MUX2BXL U145 ( .D0(n294), .D1(n291), .S(pos_dacis[7]), .Y(n320) );
  AO2222XL U146 ( .A(r_dac_en[4]), .B(n267), .C(r_dac_en[0]), .D(n265), .E(
        r_dac_en[2]), .F(n266), .G(n89), .H(r_dac_en[6]), .Y(n256) );
  INVX1 U147 ( .A(pos_dacis[3]), .Y(n280) );
  AND2X1 U148 ( .A(ps_ptr[2]), .B(ps_ptr[1]), .Y(n89) );
  NAND21XL U149 ( .B(ps_ptr[2]), .A(ps_ptr[1]), .Y(n254) );
  AO21X1 U150 ( .B(N1305), .C(n502), .A(n501), .Y(o_dacv[48]) );
  MUX2IX1 U151 ( .D0(n87), .D1(n427), .S(pos_dacis[14]), .Y(n434) );
  MUX2X1 U152 ( .D0(n435), .D1(n456), .S(pos_dacis[16]), .Y(n474) );
  AO21XL U153 ( .B(N1262), .C(n490), .A(n489), .Y(o_dacv[17]) );
  AO21XL U154 ( .B(N1263), .C(n490), .A(n489), .Y(o_dacv[18]) );
  INVXL U155 ( .A(n429), .Y(n431) );
  OAI21BXL U156 ( .C(n474), .B(pos_dacis[17]), .A(n473), .Y(o_smpl[2]) );
  AOI21XL U157 ( .B(n432), .C(n318), .A(n422), .Y(n87) );
  INVXL U158 ( .A(dacv_wr[12]), .Y(n246) );
  NAND21XL U159 ( .B(n124), .A(N1280), .Y(n491) );
  NAND21XL U160 ( .B(n124), .A(N1258), .Y(n485) );
  NAND21XL U161 ( .B(n124), .A(N1247), .Y(n482) );
  NAND21XL U162 ( .B(n124), .A(N1302), .Y(n497) );
  NAND21XL U163 ( .B(n124), .A(N1291), .Y(n494) );
  OAI21BBX1 U164 ( .A(r_wdat[0]), .B(o_dactl[0]), .C(r_wr[0]), .Y(n250) );
  AO21X1 U165 ( .B(N1239), .C(n484), .A(n483), .Y(o_dacv[0]) );
  AO21XL U166 ( .B(N1240), .C(n484), .A(n483), .Y(o_dacv[1]) );
  AO21XL U167 ( .B(N1251), .C(n487), .A(n486), .Y(o_dacv[9]) );
  AO21XL U168 ( .B(N1318), .C(n505), .A(n504), .Y(o_dacv[58]) );
  AO21XL U169 ( .B(N1274), .C(n493), .A(n492), .Y(o_dacv[26]) );
  AO21XL U170 ( .B(N1307), .C(n502), .A(n501), .Y(o_dacv[50]) );
  INVXL U171 ( .A(N1269), .Y(n490) );
  AO21XL U172 ( .B(N1296), .C(n499), .A(n498), .Y(o_dacv[42]) );
  AO21XL U173 ( .B(N1284), .C(n496), .A(n495), .Y(o_dacv[33]) );
  AO21XL U174 ( .B(N1273), .C(n493), .A(n492), .Y(o_dacv[25]) );
  OAI21BBXL U175 ( .A(ps_ptr[4]), .B(r_sar_en[17]), .C(n86), .Y(n270) );
  MUX2IX1 U176 ( .D0(n269), .D1(n268), .S(ps_ptr[3]), .Y(n86) );
  BUFX3 U177 ( .A(n571), .Y(n110) );
  AO2222XL U178 ( .A(r_dac_en[5]), .B(n267), .C(r_dac_en[1]), .D(n265), .E(
        r_dac_en[3]), .F(n266), .G(n89), .H(r_dac_en[7]), .Y(n259) );
  INVXL U179 ( .A(n568), .Y(n126) );
  OAI31XL U180 ( .A(n283), .B(pos_dacis[0]), .C(n282), .D(n322), .Y(n312) );
  OAI222XL U181 ( .A(n208), .B(n544), .C(n209), .D(n543), .E(cs_ptr[4]), .F(
        n437), .Y(n139) );
  AOI22XL U182 ( .A(r_dacvs[30]), .B(n334), .C(r_dacvs[78]), .D(n335), .Y(n352) );
  AOI22XL U183 ( .A(r_dacvs[52]), .B(n336), .C(r_dacvs[36]), .D(n337), .Y(n367) );
  AOI22XL U184 ( .A(r_dacvs[53]), .B(n81), .C(r_dacvs[37]), .D(n337), .Y(n357)
         );
  AOI22XL U185 ( .A(r_dacvs[22]), .B(n334), .C(r_dacvs[70]), .D(n335), .Y(n348) );
  AOI22XL U186 ( .A(r_dacvs[60]), .B(n336), .C(r_dacvs[44]), .D(n337), .Y(n371) );
  AOI22XL U187 ( .A(r_dacvs[61]), .B(n81), .C(r_dacvs[45]), .D(n62), .Y(n361)
         );
  AOI22XL U188 ( .A(r_dacvs[134]), .B(n338), .C(r_dacvs[6]), .D(n339), .Y(n346) );
  AOI22XL U189 ( .A(r_dacvs[142]), .B(n338), .C(r_dacvs[14]), .D(n77), .Y(n350) );
  AOI22XL U190 ( .A(r_dacvs[143]), .B(n55), .C(r_dacvs[15]), .D(n77), .Y(n340)
         );
  INVX1 U191 ( .A(dacv_wr[5]), .Y(n539) );
  INVX1 U192 ( .A(dacv_wr[4]), .Y(n538) );
  INVXL U193 ( .A(n249), .Y(n464) );
  INVX1 U194 ( .A(dacv_wr[10]), .Y(n534) );
  INVX1 U195 ( .A(dacv_wr[13]), .Y(n232) );
  INVX1 U197 ( .A(dacv_wr[6]), .Y(n540) );
  NOR2X1 U198 ( .A(n532), .B(n541), .Y(clrsta[5]) );
  NOR2X1 U199 ( .A(n10), .B(n541), .Y(clrsta[1]) );
  NOR2X1 U226 ( .A(n533), .B(n541), .Y(clrsta[2]) );
  NOR2X1 U227 ( .A(n531), .B(n541), .Y(clrsta[6]) );
  NOR2X1 U228 ( .A(n243), .B(n541), .Y(clrsta[3]) );
  AND2X1 U229 ( .A(n103), .B(r_wr[4]), .Y(clrsta[0]) );
  NOR2X1 U230 ( .A(n530), .B(n541), .Y(clrsta[7]) );
  INVX1 U231 ( .A(r_wdat[3]), .Y(n243) );
  INVXL U232 ( .A(dacv_wr[17]), .Y(n536) );
  INVX1 U233 ( .A(r_wdat[5]), .Y(n532) );
  NAND21X1 U234 ( .B(n272), .A(n251), .Y(semi_start) );
  INVX1 U235 ( .A(n251), .Y(n90) );
  INVX1 U236 ( .A(r_wdat[2]), .Y(n533) );
  INVX1 U237 ( .A(r_wdat[6]), .Y(n531) );
  INVX1 U238 ( .A(r_wdat[7]), .Y(n530) );
  NOR2X1 U239 ( .A(n115), .B(n40), .Y(n323) );
  NOR2X1 U240 ( .A(n39), .B(n114), .Y(n325) );
  INVX1 U241 ( .A(r_wr[4]), .Y(n541) );
  INVX1 U242 ( .A(r_wr[3]), .Y(n542) );
  INVX1 U243 ( .A(n51), .Y(n136) );
  INVX1 U244 ( .A(n161), .Y(n563) );
  INVX1 U248 ( .A(n162), .Y(n562) );
  NAND2X1 U249 ( .A(n563), .B(n52), .Y(n143) );
  NAND2X1 U250 ( .A(n562), .B(n52), .Y(n144) );
  NAND2X1 U251 ( .A(n73), .B(n115), .Y(n149) );
  NAND2X1 U252 ( .A(n73), .B(n114), .Y(n148) );
  NAND2X1 U253 ( .A(n331), .B(n114), .Y(n153) );
  NAND2X1 U254 ( .A(n61), .B(n115), .Y(n157) );
  NAND2X1 U255 ( .A(n66), .B(n115), .Y(n154) );
  NAND2X1 U256 ( .A(n61), .B(n114), .Y(n156) );
  INVX1 U257 ( .A(N1412), .Y(n523) );
  INVX1 U258 ( .A(n521), .Y(n522) );
  NAND21X1 U259 ( .B(r_adofs[7]), .A(N1412), .Y(n521) );
  NAND21X1 U260 ( .B(r_adofs[7]), .A(N1401), .Y(n518) );
  INVX1 U261 ( .A(n525), .Y(n526) );
  INVX1 U262 ( .A(N1313), .Y(n502) );
  INVX1 U263 ( .A(N1324), .Y(n505) );
  INVX1 U264 ( .A(N1258), .Y(n487) );
  INVX1 U265 ( .A(N1280), .Y(n493) );
  INVX1 U266 ( .A(N1247), .Y(n484) );
  INVX1 U267 ( .A(N1302), .Y(n499) );
  INVX1 U268 ( .A(N1291), .Y(n496) );
  INVX1 U269 ( .A(n500), .Y(n501) );
  NAND21X1 U270 ( .B(r_adofs[7]), .A(N1313), .Y(n500) );
  INVX1 U271 ( .A(n503), .Y(n504) );
  NAND21X1 U272 ( .B(r_adofs[7]), .A(N1324), .Y(n503) );
  INVX1 U273 ( .A(n485), .Y(n486) );
  INVX1 U274 ( .A(n491), .Y(n492) );
  INVX1 U275 ( .A(n482), .Y(n483) );
  INVX1 U276 ( .A(n497), .Y(n498) );
  INVX1 U277 ( .A(n494), .Y(n495) );
  INVX1 U278 ( .A(n248), .Y(n463) );
  INVX1 U279 ( .A(n456), .Y(n470) );
  INVX1 U280 ( .A(n253), .Y(n265) );
  NAND21X1 U281 ( .B(ps_ptr[4]), .A(n93), .Y(n253) );
  AO21X1 U282 ( .B(n465), .C(n472), .A(n97), .Y(o_smpl[0]) );
  INVX1 U283 ( .A(n254), .Y(n266) );
  INVX1 U284 ( .A(n252), .Y(n267) );
  NAND21XL U285 ( .B(ps_ptr[1]), .A(ps_ptr[2]), .Y(n252) );
  NOR2XL U286 ( .A(ps_ptr[2]), .B(ps_ptr[1]), .Y(n93) );
  INVX1 U287 ( .A(n309), .Y(n316) );
  NAND21X1 U288 ( .B(n308), .A(n307), .Y(n309) );
  INVX1 U289 ( .A(n242), .Y(n272) );
  INVX1 U290 ( .A(n244), .Y(n241) );
  OR4X1 U291 ( .A(n244), .B(n533), .C(n243), .D(n94), .Y(n251) );
  OR3XL U292 ( .A(n532), .B(r_wdat[6]), .C(n104), .Y(n94) );
  OAI22AXL U293 ( .D(dacv_wr[16]), .C(n82), .A(n136), .B(n152), .Y(upd[16]) );
  OAI22AXL U294 ( .D(dacv_wr[13]), .C(n82), .A(n143), .B(n155), .Y(upd[13]) );
  OAI22AX1 U295 ( .D(dacv_wr[7]), .C(n83), .A(n136), .B(n145), .Y(upd[7]) );
  OAI22AX1 U296 ( .D(dacv_wr[3]), .C(n83), .A(n545), .B(n148), .Y(upd[3]) );
  OAI22AX1 U297 ( .D(dacv_wr[2]), .C(n83), .A(n545), .B(n149), .Y(upd[2]) );
  OAI22AX1 U298 ( .D(dacv_wr[0]), .C(n83), .A(n144), .B(n150), .Y(upd[0]) );
  OAI22AX1 U299 ( .D(dacv_wr[1]), .C(n83), .A(n143), .B(n150), .Y(upd[1]) );
  OAI22X1 U300 ( .A(n83), .B(n245), .C(n153), .D(n136), .Y(upd[15]) );
  OAI22X1 U301 ( .A(n136), .B(n146), .C(n540), .D(n82), .Y(upd[6]) );
  OAI22X1 U302 ( .A(n83), .B(n246), .C(n144), .D(n155), .Y(upd[12]) );
  OAI22X1 U303 ( .A(n136), .B(n151), .C(n536), .D(n82), .Y(upd[17]) );
  OAI22X1 U304 ( .A(n136), .B(n154), .C(n535), .D(n82), .Y(upd[14]) );
  OAI22X1 U305 ( .A(n136), .B(n156), .C(n537), .D(n82), .Y(upd[11]) );
  OAI22X1 U306 ( .A(n136), .B(n157), .C(n534), .D(n82), .Y(upd[10]) );
  INVX1 U307 ( .A(n115), .Y(n114) );
  INVX1 U308 ( .A(cs_ptr[0]), .Y(n115) );
  NAND2X1 U309 ( .A(n114), .B(n565), .Y(n161) );
  NAND2X1 U310 ( .A(n565), .B(n115), .Y(n162) );
  NAND21X1 U311 ( .B(cs_ptr[4]), .A(n215), .Y(n155) );
  NAND21X1 U312 ( .B(cs_ptr[4]), .A(n561), .Y(n142) );
  NOR2X1 U313 ( .A(n142), .B(n565), .Y(n333) );
  NOR2X1 U314 ( .A(n155), .B(n565), .Y(n331) );
  NOR2X1 U315 ( .A(n150), .B(n565), .Y(n334) );
  INVX1 U316 ( .A(n199), .Y(n559) );
  NAND2X1 U317 ( .A(cs_ptr[4]), .B(n115), .Y(n209) );
  NAND2X1 U318 ( .A(cs_ptr[4]), .B(n114), .Y(n208) );
  NOR32XL U319 ( .B(cs_ptr[4]), .C(n565), .A(n199), .Y(n338) );
  MUX2AXL U320 ( .D0(n557), .D1(sacyc_done), .S(n462), .Y(n95) );
  INVX1 U321 ( .A(dacyc_done), .Y(n557) );
  NOR2X1 U322 ( .A(n162), .B(n164), .Y(setsta[0]) );
  NOR2X1 U323 ( .A(n161), .B(n164), .Y(setsta[1]) );
  NOR2X1 U324 ( .A(n160), .B(n164), .Y(setsta[2]) );
  NOR2X1 U325 ( .A(n158), .B(n164), .Y(setsta[3]) );
  NOR2X1 U326 ( .A(n162), .B(n159), .Y(setsta[4]) );
  NOR2X1 U327 ( .A(n160), .B(n159), .Y(setsta[6]) );
  NOR2X1 U328 ( .A(n158), .B(n159), .Y(setsta[7]) );
  NOR2X1 U329 ( .A(n161), .B(n159), .Y(setsta[5]) );
  NAND3X1 U330 ( .A(n76), .B(cs_ptr[4]), .C(n563), .Y(n151) );
  NAND3X1 U331 ( .A(n76), .B(cs_ptr[4]), .C(n562), .Y(n152) );
  NAND2X1 U332 ( .A(n336), .B(n114), .Y(n145) );
  NAND2X1 U333 ( .A(n81), .B(n115), .Y(n146) );
  AO21XL U334 ( .B(N1241), .C(n484), .A(n483), .Y(o_dacv[2]) );
  AO21X1 U335 ( .B(N1356), .C(n510), .A(n41), .Y(o_dacv[87]) );
  AO21X1 U336 ( .B(n517), .C(N1389), .A(n516), .Y(o_dacv[111]) );
  AO21XL U337 ( .B(N1355), .C(n4), .A(n41), .Y(o_dacv[86]) );
  AO21XL U338 ( .B(N1353), .C(n4), .A(n41), .Y(o_dacv[84]) );
  AO21XL U339 ( .B(N1398), .C(n520), .A(n519), .Y(o_dacv[117]) );
  AO21XL U340 ( .B(N1354), .C(n510), .A(n41), .Y(o_dacv[85]) );
  AO21XL U341 ( .B(N1352), .C(n4), .A(n41), .Y(o_dacv[83]) );
  AO21XL U342 ( .B(N1388), .C(n517), .A(n516), .Y(o_dacv[110]) );
  AO21XL U343 ( .B(N1386), .C(n517), .A(n516), .Y(o_dacv[108]) );
  AO21XL U344 ( .B(N1387), .C(n517), .A(n516), .Y(o_dacv[109]) );
  AO21XL U345 ( .B(N1385), .C(n517), .A(n516), .Y(o_dacv[107]) );
  AO21X1 U346 ( .B(N1367), .C(n513), .A(n512), .Y(o_dacv[95]) );
  AO21X1 U347 ( .B(n514), .C(N1378), .A(n42), .Y(o_dacv[103]) );
  AO21XL U348 ( .B(N1365), .C(n513), .A(n512), .Y(o_dacv[93]) );
  AO21XL U349 ( .B(N1363), .C(n513), .A(n512), .Y(o_dacv[91]) );
  AO21XL U350 ( .B(N1375), .C(n514), .A(n43), .Y(o_dacv[100]) );
  AO21XL U351 ( .B(N1376), .C(n514), .A(n43), .Y(o_dacv[101]) );
  AO21XL U352 ( .B(N1374), .C(n514), .A(n43), .Y(o_dacv[99]) );
  NAND32X1 U353 ( .B(n312), .C(n292), .A(n321), .Y(n289) );
  NAND21X1 U354 ( .B(n480), .A(n465), .Y(n456) );
  OAI211X1 U355 ( .C(n288), .D(n286), .A(n285), .B(n284), .Y(n292) );
  AO21X1 U356 ( .B(n319), .C(n320), .A(n429), .Y(n318) );
  OR2X1 U357 ( .A(n297), .B(n96), .Y(n308) );
  AOI21X1 U358 ( .B(n320), .C(n299), .A(n425), .Y(n96) );
  AO21XL U359 ( .B(N1394), .C(n520), .A(n519), .Y(o_dacv[113]) );
  AO21XL U360 ( .B(N1350), .C(n4), .A(n41), .Y(o_dacv[81]) );
  AO21XL U361 ( .B(N1383), .C(n517), .A(n516), .Y(o_dacv[105]) );
  AO21XL U362 ( .B(N1395), .C(n520), .A(n519), .Y(o_dacv[114]) );
  AO21XL U363 ( .B(N1351), .C(n4), .A(n41), .Y(o_dacv[82]) );
  AO21XL U364 ( .B(N1384), .C(n517), .A(n516), .Y(o_dacv[106]) );
  AO21XL U365 ( .B(N1361), .C(n513), .A(n512), .Y(o_dacv[89]) );
  AO21XL U366 ( .B(N1360), .C(n513), .A(n512), .Y(o_dacv[88]) );
  AO21XL U367 ( .B(N1372), .C(n514), .A(n43), .Y(o_dacv[97]) );
  AO21XL U368 ( .B(N1362), .C(n513), .A(n512), .Y(o_dacv[90]) );
  AO21XL U369 ( .B(N1371), .C(n514), .A(n43), .Y(o_dacv[96]) );
  AO21XL U370 ( .B(N1373), .C(n514), .A(n43), .Y(o_dacv[98]) );
  OAI211X1 U371 ( .C(n470), .D(n469), .A(n468), .B(n467), .Y(n479) );
  AND2X1 U372 ( .A(n473), .B(n466), .Y(n467) );
  OAI211X1 U373 ( .C(n286), .D(n284), .A(n285), .B(n288), .Y(n420) );
  OAI22X1 U374 ( .A(n317), .B(n475), .C(n432), .D(n310), .Y(n422) );
  AND2X1 U375 ( .A(n316), .B(n318), .Y(n310) );
  INVX1 U376 ( .A(n296), .Y(n314) );
  NAND32XL U377 ( .B(n308), .C(n295), .A(n320), .Y(n296) );
  AND2XL U378 ( .A(n474), .B(n470), .Y(n97) );
  INVX1 U379 ( .A(n312), .Y(n288) );
  GEN2XL U380 ( .D(n318), .E(n317), .C(n432), .B(n316), .A(n315), .Y(n433) );
  AND3X1 U381 ( .A(n314), .B(n432), .C(n313), .Y(n315) );
  AO21XL U382 ( .B(N1252), .C(n487), .A(n486), .Y(o_dacv[10]) );
  AO21X1 U383 ( .B(n472), .C(n471), .A(n479), .Y(o_smpl[1]) );
  OAI211X1 U384 ( .C(n294), .D(n421), .A(n293), .B(n311), .Y(n297) );
  INVXL U385 ( .A(n292), .Y(n293) );
  INVX1 U386 ( .A(n428), .Y(n465) );
  OAI211X1 U387 ( .C(n434), .D(n466), .A(n433), .B(n468), .Y(n428) );
  INVX1 U388 ( .A(n127), .Y(n123) );
  INVX1 U389 ( .A(n126), .Y(n124) );
  INVX1 U390 ( .A(n127), .Y(n122) );
  INVX1 U391 ( .A(n126), .Y(r_adofs[7]) );
  INVX1 U392 ( .A(n295), .Y(n425) );
  NAND6XL U393 ( .A(n92), .B(r_wdat[7]), .C(n240), .D(n239), .E(n10), .F(n238), 
        .Y(n244) );
  INVX1 U394 ( .A(o_dactl[0]), .Y(n239) );
  NAND43X1 U395 ( .B(n237), .C(n236), .D(n235), .A(n234), .Y(n240) );
  NAND2X1 U396 ( .A(n98), .B(n319), .Y(n430) );
  INVX1 U397 ( .A(n276), .Y(n319) );
  NAND21X1 U398 ( .B(n295), .A(n307), .Y(n276) );
  INVX1 U399 ( .A(n302), .Y(n307) );
  OAI221X1 U400 ( .A(n539), .B(n553), .C(n538), .D(n555), .E(n223), .Y(n236)
         );
  OA222X1 U401 ( .A(n540), .B(n552), .C(n543), .D(n222), .E(n554), .F(n221), 
        .Y(n223) );
  INVX1 U402 ( .A(dacv_wr[7]), .Y(n221) );
  INVXL U403 ( .A(dacv_wr[16]), .Y(n222) );
  AO21XL U404 ( .B(N1264), .C(n490), .A(n489), .Y(o_dacv[19]) );
  AO21XL U405 ( .B(N1253), .C(n487), .A(n486), .Y(o_dacv[11]) );
  AO21XL U406 ( .B(N1242), .C(n484), .A(n483), .Y(o_dacv[3]) );
  OAI22X1 U407 ( .A(n539), .B(n83), .C(n143), .D(n147), .Y(upd[5]) );
  OAI22X1 U408 ( .A(n538), .B(n83), .C(n144), .D(n147), .Y(upd[4]) );
  INVX1 U409 ( .A(n481), .Y(n472) );
  INVX1 U410 ( .A(n137), .Y(n64) );
  AO21XL U411 ( .B(N1265), .C(n490), .A(n489), .Y(o_dacv[20]) );
  AO21XL U412 ( .B(N1254), .C(n487), .A(n486), .Y(o_dacv[12]) );
  INVX1 U413 ( .A(cs_ptr[1]), .Y(n565) );
  AO21XL U414 ( .B(N1243), .C(n484), .A(n483), .Y(o_dacv[4]) );
  AO21XL U415 ( .B(N1266), .C(n490), .A(n489), .Y(o_dacv[21]) );
  AO21XL U416 ( .B(N1267), .C(n490), .A(n489), .Y(o_dacv[22]) );
  AO21XL U417 ( .B(N1255), .C(n487), .A(n486), .Y(o_dacv[13]) );
  AO21XL U418 ( .B(N1256), .C(n487), .A(n486), .Y(o_dacv[14]) );
  AO21XL U419 ( .B(N1257), .C(n487), .A(n486), .Y(o_dacv[15]) );
  AO21XL U420 ( .B(N1244), .C(n484), .A(n483), .Y(o_dacv[5]) );
  AO21XL U421 ( .B(N1245), .C(n484), .A(n483), .Y(o_dacv[6]) );
  AO21XL U422 ( .B(N1246), .C(n484), .A(n483), .Y(o_dacv[7]) );
  AO21XL U423 ( .B(N1268), .C(n490), .A(n489), .Y(o_dacv[23]) );
  NOR2X1 U424 ( .A(n560), .B(n564), .Y(n215) );
  NAND2X1 U425 ( .A(o_dactl[0]), .B(n139), .Y(n414) );
  NAND2X1 U426 ( .A(cs_ptr[1]), .B(n114), .Y(n158) );
  OAI22X1 U427 ( .A(n217), .B(n548), .C(n200), .D(n554), .Y(n444) );
  OAI22X1 U428 ( .A(n217), .B(n547), .C(n200), .D(n552), .Y(n445) );
  INVX1 U429 ( .A(n217), .Y(n561) );
  NOR2X1 U430 ( .A(n147), .B(n565), .Y(n336) );
  NOR2X1 U431 ( .A(n155), .B(cs_ptr[1]), .Y(n332) );
  NOR2X1 U432 ( .A(n147), .B(cs_ptr[1]), .Y(n337) );
  NOR2X1 U433 ( .A(n150), .B(cs_ptr[1]), .Y(n339) );
  NAND2X1 U434 ( .A(n564), .B(n560), .Y(n199) );
  NAND2X1 U435 ( .A(n415), .B(n564), .Y(n150) );
  NAND2X1 U436 ( .A(cs_ptr[1]), .B(n115), .Y(n160) );
  NOR2X1 U437 ( .A(n142), .B(cs_ptr[1]), .Y(n335) );
  INVX1 U438 ( .A(n203), .Y(n92) );
  NAND21X1 U439 ( .B(n436), .A(n5), .Y(n129) );
  NAND3X1 U440 ( .A(n7), .B(n546), .C(n551), .Y(n436) );
  OAI21X1 U441 ( .B(n545), .C(n137), .A(n542), .Y(updlsb) );
  INVX1 U442 ( .A(n247), .Y(n462) );
  NAND21X1 U443 ( .B(n92), .A(n139), .Y(n247) );
  NAND21X1 U444 ( .B(n147), .A(n163), .Y(n159) );
  NAND21X1 U445 ( .B(n150), .A(n163), .Y(n164) );
  NAND2X1 U446 ( .A(n303), .B(n304), .Y(o_intr) );
  NOR4XL U447 ( .A(r_irq[3]), .B(r_irq[2]), .C(r_irq[1]), .D(r_irq[0]), .Y(
        n303) );
  NOR4XL U448 ( .A(r_irq[7]), .B(r_irq[6]), .C(r_irq[5]), .D(r_irq[4]), .Y(
        n304) );
  INVX1 U449 ( .A(n200), .Y(n558) );
  AOI21X1 U450 ( .B(n203), .C(n207), .A(n557), .Y(sar_nxt) );
  NAND2X1 U451 ( .A(n140), .B(n139), .Y(n207) );
  NOR2X1 U452 ( .A(n138), .B(n557), .Y(updcmp) );
  XNOR2XL U453 ( .A(n139), .B(n140), .Y(n138) );
  OAI22X1 U454 ( .A(n150), .B(n446), .C(n452), .D(n567), .Y(datcmp[1]) );
  NOR2X1 U455 ( .A(n161), .B(n150), .Y(n452) );
  OAI22X1 U456 ( .A(n147), .B(n446), .C(n450), .D(n566), .Y(datcmp[5]) );
  NOR2X1 U457 ( .A(n161), .B(n147), .Y(n450) );
  AO21X1 U458 ( .B(N1294), .C(n499), .A(n498), .Y(o_dacv[40]) );
  AO21X1 U459 ( .B(N1317), .C(n505), .A(n504), .Y(o_dacv[57]) );
  AO21X1 U460 ( .B(N1283), .C(n496), .A(n495), .Y(o_dacv[32]) );
  AO21XL U461 ( .B(N1285), .C(n496), .A(n495), .Y(o_dacv[34]) );
  AO21X1 U462 ( .B(N1295), .C(n499), .A(n498), .Y(o_dacv[41]) );
  AO21X1 U463 ( .B(N1261), .C(n490), .A(n489), .Y(o_dacv[16]) );
  AO21X1 U464 ( .B(N1306), .C(n502), .A(n501), .Y(o_dacv[49]) );
  AO21XL U465 ( .B(N1316), .C(n505), .A(n504), .Y(o_dacv[56]) );
  AO21X1 U466 ( .B(N1345), .C(n509), .A(n6), .Y(o_dacv[79]) );
  AO21X1 U467 ( .B(N1422), .C(n524), .A(n44), .Y(o_dacv[135]) );
  AO21XL U468 ( .B(N1339), .C(n509), .A(n6), .Y(o_dacv[73]) );
  AO21XL U469 ( .B(N1338), .C(n509), .A(n6), .Y(o_dacv[72]) );
  AO21XL U470 ( .B(N1344), .C(n509), .A(n6), .Y(o_dacv[78]) );
  AO21XL U471 ( .B(N1342), .C(n509), .A(n6), .Y(o_dacv[76]) );
  AO21XL U472 ( .B(N1340), .C(n509), .A(n6), .Y(o_dacv[74]) );
  AO21XL U473 ( .B(N1343), .C(n509), .A(n6), .Y(o_dacv[77]) );
  AO21XL U474 ( .B(N1341), .C(n509), .A(n6), .Y(o_dacv[75]) );
  AO21XL U475 ( .B(N1405), .C(n523), .A(n522), .Y(o_dacv[121]) );
  AO21XL U476 ( .B(N1410), .C(n523), .A(n522), .Y(o_dacv[126]) );
  AO21XL U477 ( .B(N1404), .C(n523), .A(n522), .Y(o_dacv[120]) );
  AO21XL U478 ( .B(N1408), .C(n523), .A(n522), .Y(o_dacv[124]) );
  AO21XL U479 ( .B(N1409), .C(n523), .A(n522), .Y(o_dacv[125]) );
  AO21XL U480 ( .B(N1407), .C(n523), .A(n522), .Y(o_dacv[123]) );
  AO21XL U481 ( .B(N1415), .C(n524), .A(n45), .Y(o_dacv[128]) );
  AO21XL U482 ( .B(N1421), .C(n524), .A(n44), .Y(o_dacv[134]) );
  AO21XL U483 ( .B(N1419), .C(n524), .A(n45), .Y(o_dacv[132]) );
  AO21XL U484 ( .B(N1417), .C(n48), .A(n45), .Y(o_dacv[130]) );
  AO21XL U485 ( .B(N1420), .C(n48), .A(n45), .Y(o_dacv[133]) );
  AO21XL U486 ( .B(N1418), .C(n524), .A(n45), .Y(o_dacv[131]) );
  AO21X1 U487 ( .B(N1334), .C(n508), .A(n507), .Y(o_dacv[71]) );
  AO21X1 U488 ( .B(N1433), .C(n527), .A(n526), .Y(o_dacv[143]) );
  AO21XL U489 ( .B(N1328), .C(n508), .A(n507), .Y(o_dacv[65]) );
  AO21XL U490 ( .B(N1427), .C(n527), .A(n526), .Y(o_dacv[137]) );
  AO21XL U491 ( .B(N1432), .C(n527), .A(n526), .Y(o_dacv[142]) );
  AO21XL U492 ( .B(N1426), .C(n527), .A(n526), .Y(o_dacv[136]) );
  AO21XL U493 ( .B(N1430), .C(n527), .A(n526), .Y(o_dacv[140]) );
  AO21XL U494 ( .B(N1332), .C(n508), .A(n507), .Y(o_dacv[69]) );
  AO21XL U495 ( .B(N1431), .C(n527), .A(n526), .Y(o_dacv[141]) );
  AO21XL U496 ( .B(N1429), .C(n527), .A(n526), .Y(o_dacv[139]) );
  NAND5XL U497 ( .A(n432), .B(n431), .C(n430), .D(n468), .E(n466), .Y(n435) );
  XOR2X1 U498 ( .A(n277), .B(pos_dacis[1]), .Y(n281) );
  MUX3XL U499 ( .D0(n420), .D1(n288), .D2(n289), .S0(n321), .S1(pos_dacis[6]), 
        .Y(n294) );
  AND4X1 U500 ( .A(n426), .B(n433), .C(n476), .D(n471), .Y(n427) );
  INVX1 U501 ( .A(n430), .Y(n426) );
  AND2X1 U502 ( .A(n290), .B(n311), .Y(n291) );
  INVXL U503 ( .A(n289), .Y(n290) );
  NAND31X1 U504 ( .C(pos_dacis[6]), .A(n99), .B(n421), .Y(n424) );
  MUX2IXL U505 ( .D0(n420), .D1(n322), .S(n321), .Y(n99) );
  NAND21X1 U506 ( .B(n97), .A(pos_dacis[17]), .Y(n473) );
  MUX2IXL U507 ( .D0(n434), .D1(n100), .S(pos_dacis[15]), .Y(n480) );
  NAND3X1 U508 ( .A(n434), .B(n433), .C(n468), .Y(n100) );
  XOR2X1 U509 ( .A(n280), .B(pos_dacis[2]), .Y(n282) );
  INVXL U510 ( .A(n281), .Y(n283) );
  NAND21X1 U511 ( .B(n479), .A(n478), .Y(o_smpl[3]) );
  NAND21X1 U512 ( .B(n481), .A(n477), .Y(n478) );
  NAND21X1 U513 ( .B(n476), .A(n475), .Y(n477) );
  OAI22X1 U514 ( .A(n313), .B(n306), .C(n314), .D(n305), .Y(n429) );
  INVX1 U515 ( .A(pos_dacis[11]), .Y(n306) );
  INVX1 U516 ( .A(n423), .Y(n305) );
  AO21XL U517 ( .B(N1406), .C(n523), .A(n522), .Y(o_dacv[122]) );
  AO21XL U518 ( .B(N1329), .C(n508), .A(n507), .Y(o_dacv[66]) );
  AO21XL U519 ( .B(N1428), .C(n527), .A(n526), .Y(o_dacv[138]) );
  AO21X1 U520 ( .B(N1272), .C(n493), .A(n492), .Y(o_dacv[24]) );
  NAND32X1 U521 ( .B(pos_dacis[2]), .C(n281), .A(n280), .Y(n322) );
  AO21XL U522 ( .B(N1349), .C(n4), .A(n41), .Y(o_dacv[80]) );
  AO21XL U523 ( .B(N1382), .C(n517), .A(n516), .Y(o_dacv[104]) );
  AO21X1 U524 ( .B(N1250), .C(n487), .A(n486), .Y(o_dacv[8]) );
  INVX1 U525 ( .A(pos_dacis[0]), .Y(n277) );
  MUX2X1 U526 ( .D0(n271), .D1(n270), .S(ps_ptr[0]), .Y(n273) );
  OA21XL U527 ( .B(n463), .C(n95), .A(n261), .Y(n274) );
  AO21XL U528 ( .B(ps_ptr[4]), .C(r_sar_en[16]), .A(n264), .Y(n271) );
  NAND31X1 U529 ( .C(n302), .A(n301), .B(n300), .Y(n423) );
  NAND21X1 U530 ( .B(n299), .A(pos_dacis[9]), .Y(n300) );
  NAND21X1 U531 ( .B(n425), .A(n298), .Y(n301) );
  NAND21XL U532 ( .B(n297), .A(n320), .Y(n298) );
  MUX2IX1 U533 ( .D0(n101), .D1(n102), .S(ps_ptr[0]), .Y(n261) );
  AOI21XL U534 ( .B(ps_ptr[4]), .C(r_dac_en[16]), .A(n257), .Y(n101) );
  AOI21XL U535 ( .B(ps_ptr[4]), .C(r_dac_en[17]), .A(n260), .Y(n102) );
  MUX2X1 U536 ( .D0(n263), .D1(n262), .S(ps_ptr[3]), .Y(n264) );
  AO2222XL U537 ( .A(n89), .B(r_sar_en[14]), .C(n267), .D(r_sar_en[12]), .E(
        n93), .F(r_sar_en[8]), .G(n266), .H(r_sar_en[10]), .Y(n262) );
  AO2222XL U538 ( .A(n267), .B(r_sar_en[4]), .C(n265), .D(r_sar_en[0]), .E(
        n266), .F(r_sar_en[2]), .G(n89), .H(r_sar_en[6]), .Y(n263) );
  MUX2X1 U539 ( .D0(n259), .D1(n258), .S(ps_ptr[3]), .Y(n260) );
  AO2222XL U540 ( .A(n89), .B(r_dac_en[15]), .C(r_dac_en[13]), .D(n267), .E(
        r_dac_en[9]), .F(n93), .G(r_dac_en[11]), .H(n266), .Y(n258) );
  AO2222XL U541 ( .A(n89), .B(r_sar_en[15]), .C(n267), .D(r_sar_en[13]), .E(
        n93), .F(r_sar_en[9]), .G(n266), .H(r_sar_en[11]), .Y(n268) );
  AO2222XL U542 ( .A(n267), .B(r_sar_en[5]), .C(n265), .D(r_sar_en[1]), .E(
        n266), .F(r_sar_en[3]), .G(n89), .H(r_sar_en[7]), .Y(n269) );
  NAND21X1 U543 ( .B(r_isofs[7]), .A(N1269), .Y(n488) );
  INVX1 U544 ( .A(n279), .Y(n285) );
  OAI211XL U545 ( .C(n281), .D(n280), .A(n278), .B(n277), .Y(n279) );
  INVXL U546 ( .A(pos_dacis[2]), .Y(n278) );
  AO2222XL U547 ( .A(n89), .B(r_dac_en[14]), .C(r_dac_en[12]), .D(n267), .E(
        r_dac_en[8]), .F(n93), .G(r_dac_en[10]), .H(n266), .Y(n255) );
  NAND32XL U548 ( .B(pos_dacis[12]), .C(n320), .A(n319), .Y(n476) );
  INVX1 U549 ( .A(n287), .Y(n321) );
  NAND21X1 U550 ( .B(pos_dacis[4]), .A(n286), .Y(n287) );
  INVX1 U551 ( .A(pos_dacis[5]), .Y(n286) );
  INVX1 U552 ( .A(pos_dacis[4]), .Y(n284) );
  NAND21X1 U553 ( .B(pos_dacis[9]), .A(n299), .Y(n295) );
  INVX1 U554 ( .A(pos_dacis[7]), .Y(n421) );
  INVX1 U555 ( .A(pos_dacis[6]), .Y(n311) );
  INVX1 U556 ( .A(pos_dacis[8]), .Y(n299) );
  NAND21X1 U557 ( .B(pos_dacis[11]), .A(n313), .Y(n302) );
  INVX1 U558 ( .A(pos_dacis[10]), .Y(n313) );
  INVX1 U559 ( .A(pos_dacis[12]), .Y(n317) );
  INVX1 U560 ( .A(n275), .Y(n432) );
  NAND21X1 U561 ( .B(pos_dacis[13]), .A(n317), .Y(n275) );
  INVX1 U562 ( .A(pos_dacis[13]), .Y(n475) );
  OAI221X1 U563 ( .A(n537), .B(n548), .C(n246), .D(n229), .E(n228), .Y(n235)
         );
  INVX1 U564 ( .A(r_sar_en[12]), .Y(n229) );
  OA222X1 U565 ( .A(n534), .B(n547), .C(n227), .D(n226), .E(n225), .F(n224), 
        .Y(n228) );
  INVX1 U566 ( .A(r_sar_en[8]), .Y(n226) );
  OA2222XL U567 ( .A(n245), .B(n233), .C(n536), .D(n544), .E(n232), .F(n231), 
        .G(n535), .H(n230), .Y(n234) );
  INVX1 U568 ( .A(r_sar_en[15]), .Y(n233) );
  INVX1 U569 ( .A(r_sar_en[13]), .Y(n231) );
  INVX1 U570 ( .A(r_sar_en[14]), .Y(n230) );
  NOR21XL U571 ( .B(app_dacis[10]), .A(n113), .Y(o_daci_sel[10]) );
  NOR21XL U572 ( .B(app_dacis[11]), .A(n112), .Y(o_daci_sel[11]) );
  NOR21XL U573 ( .B(app_dacis[6]), .A(n112), .Y(o_daci_sel[6]) );
  NOR21XL U574 ( .B(app_dacis[5]), .A(n113), .Y(o_daci_sel[5]) );
  NOR21XL U575 ( .B(app_dacis[7]), .A(n113), .Y(o_daci_sel[7]) );
  NOR21XL U576 ( .B(app_dacis[4]), .A(n112), .Y(o_daci_sel[4]) );
  NOR21XL U577 ( .B(app_dacis[16]), .A(n113), .Y(o_daci_sel[16]) );
  NOR21XL U578 ( .B(app_dacis[3]), .A(n113), .Y(o_daci_sel[3]) );
  NOR21XL U579 ( .B(app_dacis[2]), .A(n112), .Y(o_daci_sel[2]) );
  NOR21XL U580 ( .B(app_dacis[1]), .A(n113), .Y(o_daci_sel[1]) );
  NOR21XL U581 ( .B(app_dacis[14]), .A(n113), .Y(o_daci_sel[14]) );
  NOR21XL U582 ( .B(app_dacis[12]), .A(n113), .Y(o_daci_sel[12]) );
  NOR21XL U583 ( .B(app_dacis[0]), .A(n112), .Y(o_daci_sel[0]) );
  NOR21XL U584 ( .B(app_dacis[17]), .A(n112), .Y(o_daci_sel[17]) );
  NOR21XL U585 ( .B(app_dacis[15]), .A(n112), .Y(o_daci_sel[15]) );
  NOR21XL U586 ( .B(app_dacis[8]), .A(n112), .Y(o_daci_sel[8]) );
  NOR21XL U587 ( .B(app_dacis[9]), .A(n113), .Y(o_daci_sel[9]) );
  INVX1 U588 ( .A(pos_dacis[14]), .Y(n468) );
  INVX1 U589 ( .A(pos_dacis[15]), .Y(n466) );
  NOR21XL U590 ( .B(app_dacis[13]), .A(n112), .Y(o_daci_sel[13]) );
  AO21XL U591 ( .B(N1297), .C(n499), .A(n498), .Y(o_dacv[43]) );
  AO21XL U592 ( .B(N1319), .C(n505), .A(n504), .Y(o_dacv[59]) );
  AO21XL U593 ( .B(N1308), .C(n502), .A(n501), .Y(o_dacv[51]) );
  AO21XL U594 ( .B(N1286), .C(n496), .A(n495), .Y(o_dacv[35]) );
  AO21XL U595 ( .B(N1275), .C(n493), .A(n492), .Y(o_dacv[27]) );
  NAND21X1 U596 ( .B(pos_dacis[17]), .A(n469), .Y(n481) );
  INVX1 U597 ( .A(pos_dacis[16]), .Y(n469) );
  MUX2BXL U598 ( .D0(o_dactl[5]), .D1(n532), .S(n91), .Y(ps_md4ch) );
  AO2222XL U599 ( .A(r_sar_en[2]), .B(dacv_wr[2]), .C(r_sar_en[3]), .D(
        dacv_wr[3]), .E(r_sar_en[0]), .F(dacv_wr[0]), .G(r_sar_en[1]), .H(
        dacv_wr[1]), .Y(n237) );
  AO21XL U600 ( .B(N1309), .C(n502), .A(n501), .Y(o_dacv[52]) );
  ENOX1 U601 ( .A(n10), .B(n52), .C(r_rpt_v[3]), .D(n51), .Y(n457) );
  ENOX1 U602 ( .A(n533), .B(n52), .C(r_rpt_v[4]), .D(n51), .Y(n458) );
  ENOX1 U603 ( .A(n532), .B(n52), .C(r_rpt_v[7]), .D(n51), .Y(n461) );
  AO21XL U604 ( .B(N1320), .C(n505), .A(n504), .Y(o_dacv[60]) );
  NAND4X1 U605 ( .A(o_dactl[6]), .B(n415), .C(n416), .D(n417), .Y(n137) );
  NOR2X1 U606 ( .A(n418), .B(n419), .Y(n417) );
  XNOR2XL U607 ( .A(x_daclsb[3]), .B(n114), .Y(n416) );
  XNOR2XL U608 ( .A(n564), .B(x_daclsb[5]), .Y(n418) );
  ENOX1 U609 ( .A(n542), .B(n532), .C(n542), .D(x_daclsb[4]), .Y(wdlsb[4]) );
  AO21XL U610 ( .B(N1310), .C(n502), .A(n501), .Y(o_dacv[53]) );
  AO21XL U611 ( .B(N1321), .C(n505), .A(n504), .Y(o_dacv[61]) );
  AO21XL U612 ( .B(N1311), .C(n502), .A(n501), .Y(o_dacv[54]) );
  AO21XL U613 ( .B(N1276), .C(n493), .A(n492), .Y(o_dacv[28]) );
  AO21XL U614 ( .B(N1277), .C(n493), .A(n492), .Y(o_dacv[29]) );
  AO21XL U615 ( .B(N1288), .C(n496), .A(n495), .Y(o_dacv[37]) );
  AO21XL U616 ( .B(N1299), .C(n499), .A(n498), .Y(o_dacv[45]) );
  AO21XL U617 ( .B(N1287), .C(n496), .A(n495), .Y(o_dacv[36]) );
  AO21XL U618 ( .B(N1298), .C(n499), .A(n498), .Y(o_dacv[44]) );
  ENOX1 U619 ( .A(n531), .B(n52), .C(r_rpt_v[8]), .D(n52), .Y(wda[6]) );
  ENOX1 U620 ( .A(n52), .B(n243), .C(r_rpt_v[5]), .D(n51), .Y(n459) );
  ENOX1 U621 ( .A(n52), .B(n530), .C(r_rpt_v[9]), .D(n52), .Y(wda[7]) );
  XNOR2XL U622 ( .A(n565), .B(x_daclsb[4]), .Y(n419) );
  INVX1 U623 ( .A(cs_ptr[2]), .Y(n564) );
  AO21XL U624 ( .B(N1322), .C(n505), .A(n504), .Y(o_dacv[62]) );
  NOR2X1 U625 ( .A(cs_ptr[3]), .B(cs_ptr[4]), .Y(n415) );
  ENOX1 U626 ( .A(n531), .B(n542), .C(n542), .D(x_daclsb[5]), .Y(wdlsb[5]) );
  ENOX1 U627 ( .A(n542), .B(n10), .C(r_rpt_v[1]), .D(n542), .Y(wdlsb[1]) );
  ENOX1 U628 ( .A(n542), .B(n533), .C(x_daclsb[2]), .D(n542), .Y(wdlsb[2]) );
  AO21XL U629 ( .B(N1312), .C(n502), .A(n501), .Y(o_dacv[55]) );
  AO21XL U630 ( .B(N1278), .C(n493), .A(n492), .Y(o_dacv[30]) );
  AO21XL U631 ( .B(N1279), .C(n493), .A(n492), .Y(o_dacv[31]) );
  AO21XL U632 ( .B(N1289), .C(n496), .A(n495), .Y(o_dacv[38]) );
  AO21XL U633 ( .B(N1300), .C(n499), .A(n498), .Y(o_dacv[46]) );
  AO21XL U634 ( .B(N1290), .C(n496), .A(n495), .Y(o_dacv[39]) );
  AO21XL U635 ( .B(N1301), .C(n499), .A(n498), .Y(o_dacv[47]) );
  AO21XL U636 ( .B(N1323), .C(n505), .A(n504), .Y(o_dacv[63]) );
  MUX2XL U637 ( .D0(r_wdat[4]), .D1(x_daclsb[3]), .S(n542), .Y(wdlsb[3]) );
  MUX2AXL U638 ( .D0(r_rpt_v[6]), .D1(n238), .S(n136), .Y(n202) );
  OA2222XL U639 ( .A(n438), .B(n160), .C(n439), .D(n158), .E(n440), .F(n161), 
        .G(n441), .H(n162), .Y(n437) );
  AOI221XL U640 ( .A(r_sar_en[2]), .B(n559), .C(r_sar_en[14]), .D(n215), .E(
        n445), .Y(n438) );
  AOI221XL U641 ( .A(r_sar_en[3]), .B(n559), .C(r_sar_en[15]), .D(n215), .E(
        n444), .Y(n439) );
  AO222X1 U642 ( .A(n323), .B(n384), .C(n325), .D(n385), .E(r_dac1v[4]), .F(
        n39), .Y(o_dac1[4]) );
  NAND4X1 U643 ( .A(n390), .B(n391), .C(n392), .D(n393), .Y(n384) );
  NAND4X1 U644 ( .A(n386), .B(n387), .C(n388), .D(n389), .Y(n385) );
  AOI22XL U645 ( .A(r_dacvs[26]), .B(n334), .C(r_dacvs[74]), .D(n335), .Y(n392) );
  AO222X1 U646 ( .A(n323), .B(n374), .C(n325), .D(n375), .E(r_dac1v[5]), .F(
        n40), .Y(o_dac1[5]) );
  NAND4X1 U647 ( .A(n380), .B(n381), .C(n382), .D(n383), .Y(n374) );
  NAND4X1 U648 ( .A(n376), .B(n377), .C(n378), .D(n379), .Y(n375) );
  AOI22XL U649 ( .A(r_dacvs[27]), .B(n73), .C(r_dacvs[75]), .D(n56), .Y(n382)
         );
  AO222X1 U650 ( .A(n323), .B(n364), .C(n325), .D(n365), .E(r_dac1v[6]), .F(
        n39), .Y(o_dac1[6]) );
  NAND4X1 U651 ( .A(n370), .B(n371), .C(n372), .D(n373), .Y(n364) );
  NAND4X1 U652 ( .A(n366), .B(n367), .C(n368), .D(n369), .Y(n365) );
  AOI22XL U653 ( .A(r_dacvs[28]), .B(n73), .C(r_dacvs[76]), .D(n56), .Y(n372)
         );
  AO222X1 U654 ( .A(n323), .B(n344), .C(n325), .D(n345), .E(r_dac1v[8]), .F(
        n40), .Y(o_dac1[8]) );
  NAND4X1 U655 ( .A(n350), .B(n351), .C(n352), .D(n353), .Y(n344) );
  NAND4X1 U656 ( .A(n346), .B(n347), .C(n348), .D(n349), .Y(n345) );
  AO222X1 U657 ( .A(n323), .B(n404), .C(n325), .D(n405), .E(r_dac1v[2]), .F(
        n39), .Y(o_dac1[2]) );
  NAND4X1 U658 ( .A(n410), .B(n411), .C(n412), .D(n413), .Y(n404) );
  NAND4X1 U659 ( .A(n406), .B(n407), .C(n408), .D(n409), .Y(n405) );
  AOI22XL U660 ( .A(r_dacvs[24]), .B(n73), .C(r_dacvs[72]), .D(n56), .Y(n412)
         );
  AO222X1 U661 ( .A(n323), .B(n394), .C(n325), .D(n395), .E(r_dac1v[3]), .F(
        n40), .Y(o_dac1[3]) );
  NAND4X1 U662 ( .A(n400), .B(n401), .C(n402), .D(n403), .Y(n394) );
  NAND4X1 U663 ( .A(n396), .B(n397), .C(n398), .D(n399), .Y(n395) );
  AOI22XL U664 ( .A(r_dacvs[25]), .B(n73), .C(r_dacvs[73]), .D(n56), .Y(n402)
         );
  AO222X1 U665 ( .A(n323), .B(n354), .C(n325), .D(n355), .E(r_dac1v[7]), .F(
        n39), .Y(o_dac1[7]) );
  NAND4X1 U666 ( .A(n360), .B(n361), .C(n362), .D(n363), .Y(n354) );
  NAND4X1 U667 ( .A(n356), .B(n357), .C(n358), .D(n359), .Y(n355) );
  AOI22XL U668 ( .A(r_dacvs[29]), .B(n73), .C(r_dacvs[77]), .D(n56), .Y(n362)
         );
  AO222X1 U669 ( .A(n323), .B(n324), .C(n325), .D(n326), .E(r_dac1v[9]), .F(
        n40), .Y(o_dac1[9]) );
  NAND4X1 U670 ( .A(n340), .B(n341), .C(n342), .D(n343), .Y(n324) );
  NAND4X1 U671 ( .A(n327), .B(n328), .C(n329), .D(n330), .Y(n326) );
  AOI22X1 U672 ( .A(r_dacvs[31]), .B(n73), .C(r_dacvs[79]), .D(n56), .Y(n342)
         );
  AO22X1 U673 ( .A(x_daclsb[0]), .B(n414), .C(r_dac1v[0]), .D(n39), .Y(
        o_dac1[0]) );
  AO22X1 U674 ( .A(x_daclsb[1]), .B(n414), .C(r_dac1v[1]), .D(n40), .Y(
        o_dac1[1]) );
  NAND2X1 U675 ( .A(cs_ptr[2]), .B(n560), .Y(n200) );
  INVX1 U676 ( .A(cs_ptr[3]), .Y(n560) );
  NAND2X1 U677 ( .A(cs_ptr[3]), .B(n564), .Y(n217) );
  AOI221XL U678 ( .A(r_sar_en[0]), .B(n559), .C(r_sar_en[12]), .D(n215), .E(
        n442), .Y(n441) );
  ENOX1 U679 ( .A(n200), .B(n555), .C(n561), .D(r_sar_en[8]), .Y(n442) );
  AOI221XL U680 ( .A(r_sar_en[1]), .B(n559), .C(r_sar_en[13]), .D(n215), .E(
        n443), .Y(n440) );
  ENOX1 U681 ( .A(n200), .B(n553), .C(n561), .D(r_sar_en[9]), .Y(n443) );
  INVX1 U682 ( .A(r_sar_en[7]), .Y(n554) );
  NAND2X1 U683 ( .A(n415), .B(cs_ptr[2]), .Y(n147) );
  AOI222XL U684 ( .A(r_dacvs[112]), .B(n331), .C(r_dacvs[96]), .D(n332), .E(
        r_dacvs[80]), .F(n333), .Y(n409) );
  AOI222XL U685 ( .A(r_dacvs[120]), .B(n331), .C(r_dacvs[104]), .D(n332), .E(
        r_dacvs[88]), .F(n61), .Y(n413) );
  AOI222XL U686 ( .A(r_dacvs[113]), .B(n66), .C(r_dacvs[97]), .D(n70), .E(
        r_dacvs[81]), .F(n333), .Y(n399) );
  AOI222XL U687 ( .A(r_dacvs[121]), .B(n66), .C(r_dacvs[105]), .D(n70), .E(
        r_dacvs[89]), .F(n61), .Y(n403) );
  AOI222XL U688 ( .A(r_dacvs[114]), .B(n331), .C(r_dacvs[98]), .D(n332), .E(
        r_dacvs[82]), .F(n333), .Y(n389) );
  AOI222XL U689 ( .A(r_dacvs[122]), .B(n331), .C(r_dacvs[106]), .D(n332), .E(
        r_dacvs[90]), .F(n333), .Y(n393) );
  AOI222XL U690 ( .A(r_dacvs[115]), .B(n66), .C(r_dacvs[99]), .D(n70), .E(
        r_dacvs[83]), .F(n333), .Y(n379) );
  AOI222XL U691 ( .A(r_dacvs[123]), .B(n66), .C(r_dacvs[107]), .D(n70), .E(
        r_dacvs[91]), .F(n61), .Y(n383) );
  AOI222XL U692 ( .A(r_dacvs[116]), .B(n331), .C(r_dacvs[100]), .D(n332), .E(
        r_dacvs[84]), .F(n333), .Y(n369) );
  AOI222XL U693 ( .A(r_dacvs[124]), .B(n331), .C(r_dacvs[108]), .D(n332), .E(
        r_dacvs[92]), .F(n61), .Y(n373) );
  AOI222XL U694 ( .A(r_dacvs[117]), .B(n331), .C(r_dacvs[101]), .D(n332), .E(
        r_dacvs[85]), .F(n333), .Y(n359) );
  AOI222XL U695 ( .A(r_dacvs[125]), .B(n331), .C(r_dacvs[109]), .D(n332), .E(
        r_dacvs[93]), .F(n61), .Y(n363) );
  AOI222XL U696 ( .A(r_dacvs[118]), .B(n66), .C(r_dacvs[102]), .D(n70), .E(
        r_dacvs[86]), .F(n333), .Y(n349) );
  AOI222XL U697 ( .A(r_dacvs[126]), .B(n66), .C(r_dacvs[110]), .D(n70), .E(
        r_dacvs[94]), .F(n61), .Y(n353) );
  AOI222XL U698 ( .A(r_dacvs[119]), .B(n66), .C(r_dacvs[103]), .D(n70), .E(
        r_dacvs[87]), .F(n333), .Y(n330) );
  AOI222XL U699 ( .A(r_dacvs[127]), .B(n66), .C(r_dacvs[111]), .D(n70), .E(
        r_dacvs[95]), .F(n61), .Y(n343) );
  AOI22XL U700 ( .A(r_dacvs[16]), .B(n334), .C(r_dacvs[64]), .D(n335), .Y(n408) );
  AOI22XL U701 ( .A(r_dacvs[17]), .B(n334), .C(r_dacvs[65]), .D(n335), .Y(n398) );
  AOI22XL U702 ( .A(r_dacvs[18]), .B(n334), .C(r_dacvs[66]), .D(n335), .Y(n388) );
  AOI22XL U703 ( .A(r_dacvs[19]), .B(n334), .C(r_dacvs[67]), .D(n335), .Y(n378) );
  AOI22XL U704 ( .A(r_dacvs[20]), .B(n334), .C(r_dacvs[68]), .D(n335), .Y(n368) );
  AOI22XL U705 ( .A(r_dacvs[21]), .B(n334), .C(r_dacvs[69]), .D(n335), .Y(n358) );
  AOI22X1 U706 ( .A(r_dacvs[23]), .B(n73), .C(r_dacvs[71]), .D(n56), .Y(n329)
         );
  AOI22XL U707 ( .A(r_dacvs[48]), .B(n336), .C(r_dacvs[32]), .D(n337), .Y(n407) );
  AOI22XL U708 ( .A(r_dacvs[56]), .B(n336), .C(r_dacvs[40]), .D(n62), .Y(n411)
         );
  AOI22XL U709 ( .A(r_dacvs[49]), .B(n81), .C(r_dacvs[33]), .D(n337), .Y(n397)
         );
  AOI22XL U710 ( .A(r_dacvs[57]), .B(n81), .C(r_dacvs[41]), .D(n62), .Y(n401)
         );
  AOI22XL U711 ( .A(r_dacvs[50]), .B(n81), .C(r_dacvs[34]), .D(n337), .Y(n387)
         );
  AOI22XL U712 ( .A(r_dacvs[58]), .B(n81), .C(r_dacvs[42]), .D(n337), .Y(n391)
         );
  AOI22XL U713 ( .A(r_dacvs[51]), .B(n336), .C(r_dacvs[35]), .D(n337), .Y(n377) );
  AOI22XL U714 ( .A(r_dacvs[59]), .B(n336), .C(r_dacvs[43]), .D(n337), .Y(n381) );
  AOI22X1 U715 ( .A(r_dacvs[54]), .B(n336), .C(r_dacvs[38]), .D(n62), .Y(n347)
         );
  AOI22X1 U716 ( .A(r_dacvs[62]), .B(n336), .C(r_dacvs[46]), .D(n62), .Y(n351)
         );
  AOI22X1 U717 ( .A(r_dacvs[55]), .B(n81), .C(r_dacvs[39]), .D(n62), .Y(n328)
         );
  AOI22X1 U718 ( .A(r_dacvs[63]), .B(n81), .C(r_dacvs[47]), .D(n62), .Y(n341)
         );
  AOI22XL U719 ( .A(r_dacvs[128]), .B(n338), .C(r_dacvs[0]), .D(n339), .Y(n406) );
  AOI22XL U720 ( .A(r_dacvs[129]), .B(n338), .C(r_dacvs[1]), .D(n77), .Y(n396)
         );
  AOI22XL U721 ( .A(r_dacvs[130]), .B(n338), .C(r_dacvs[2]), .D(n77), .Y(n386)
         );
  AOI22XL U722 ( .A(r_dacvs[131]), .B(n338), .C(r_dacvs[3]), .D(n339), .Y(n376) );
  AOI22XL U723 ( .A(r_dacvs[132]), .B(n338), .C(r_dacvs[4]), .D(n77), .Y(n366)
         );
  AOI22XL U724 ( .A(r_dacvs[133]), .B(n338), .C(r_dacvs[5]), .D(n339), .Y(n356) );
  AOI22X1 U725 ( .A(r_dacvs[135]), .B(n55), .C(r_dacvs[7]), .D(n77), .Y(n327)
         );
  INVX1 U726 ( .A(r_sar_en[5]), .Y(n553) );
  INVX1 U727 ( .A(r_sar_en[4]), .Y(n555) );
  INVX1 U728 ( .A(r_sar_en[6]), .Y(n552) );
  INVX1 U729 ( .A(r_sar_en[10]), .Y(n547) );
  INVX1 U730 ( .A(r_sar_en[11]), .Y(n548) );
  NAND42X1 U731 ( .C(r_dac_en[2]), .D(n201), .A(n135), .B(n134), .Y(n203) );
  NOR43XL U732 ( .B(n133), .C(n132), .D(n131), .A(n130), .Y(n134) );
  NAND21X1 U733 ( .B(r_dac_en[0]), .A(n128), .Y(n201) );
  NOR32XL U734 ( .B(n529), .C(n528), .A(n129), .Y(n135) );
  INVX1 U735 ( .A(r_dac_en[7]), .Y(n556) );
  INVX1 U736 ( .A(r_dac_en[9]), .Y(n550) );
  INVX1 U737 ( .A(r_dac_en[8]), .Y(n549) );
  AOI22XL U738 ( .A(r_dacvs[136]), .B(n55), .C(r_dacvs[8]), .D(n339), .Y(n410)
         );
  AOI22XL U739 ( .A(r_dacvs[137]), .B(n55), .C(r_dacvs[9]), .D(n77), .Y(n400)
         );
  AOI22XL U740 ( .A(r_dacvs[138]), .B(n338), .C(r_dacvs[10]), .D(n339), .Y(
        n390) );
  AOI22XL U741 ( .A(r_dacvs[139]), .B(n55), .C(r_dacvs[11]), .D(n77), .Y(n380)
         );
  AOI22XL U742 ( .A(r_dacvs[140]), .B(n55), .C(r_dacvs[12]), .D(n339), .Y(n370) );
  AOI22XL U743 ( .A(r_dacvs[141]), .B(n55), .C(r_dacvs[13]), .D(n339), .Y(n360) );
  INVX1 U744 ( .A(r_dac_en[14]), .Y(n551) );
  INVX1 U745 ( .A(r_dac_en[16]), .Y(n546) );
  INVX1 U746 ( .A(r_sar_en[16]), .Y(n543) );
  INVX1 U747 ( .A(r_sar_en[17]), .Y(n544) );
  OR4X1 U748 ( .A(r_dac_en[3]), .B(r_dac_en[4]), .C(r_dac_en[13]), .D(
        r_dac_en[5]), .Y(n130) );
  INVX1 U749 ( .A(r_dac_en[1]), .Y(n128) );
  INVX1 U750 ( .A(r_dac_en[6]), .Y(n528) );
  INVX1 U751 ( .A(r_dac_en[17]), .Y(n529) );
  INVX1 U752 ( .A(r_dac_en[12]), .Y(n132) );
  INVX1 U753 ( .A(r_dac_en[11]), .Y(n133) );
  INVX1 U754 ( .A(r_dac_en[10]), .Y(n131) );
  INVX1 U755 ( .A(r_sar_en[9]), .Y(n224) );
  BUFX3 U756 ( .A(r_comp_opt[0]), .Y(n112) );
  BUFX3 U757 ( .A(r_comp_opt[0]), .Y(n113) );
  NOR42XL U758 ( .C(n165), .D(o_dactl[1]), .A(n557), .B(n139), .Y(n163) );
  XNOR2XL U759 ( .A(syn_comp[1]), .B(n166), .Y(n165) );
  AOI221XL U760 ( .A(n563), .B(n167), .C(n562), .D(n168), .E(n169), .Y(n166)
         );
  OAI22X1 U761 ( .A(n199), .B(n567), .C(n200), .D(n566), .Y(n167) );
  OAI22X1 U762 ( .A(n170), .B(n158), .C(n171), .D(n160), .Y(n169) );
  AOI22X1 U763 ( .A(o_dat[7]), .B(n558), .C(o_dat[3]), .D(n559), .Y(n170) );
  AOI22X1 U764 ( .A(o_dat[6]), .B(n558), .C(o_dat[2]), .D(n559), .Y(n171) );
  AO22X1 U765 ( .A(n559), .B(o_dat[0]), .C(n558), .D(o_dat[4]), .Y(n168) );
  OAI222XL U766 ( .A(n208), .B(n529), .C(n209), .D(n546), .E(cs_ptr[4]), .F(
        n210), .Y(n140) );
  OA2222XL U767 ( .A(n211), .B(n160), .C(n212), .D(n158), .E(n213), .F(n161), 
        .G(n214), .H(n162), .Y(n210) );
  AOI221XL U768 ( .A(r_dac_en[2]), .B(n76), .C(r_dac_en[14]), .D(n215), .E(
        n220), .Y(n211) );
  AOI221XL U769 ( .A(r_dac_en[1]), .B(n559), .C(r_dac_en[13]), .D(n215), .E(
        n218), .Y(n213) );
  AOI221XL U770 ( .A(r_dac_en[0]), .B(n559), .C(r_dac_en[12]), .D(n215), .E(
        n216), .Y(n214) );
  ENOX1 U771 ( .A(n217), .B(n549), .C(n558), .D(r_dac_en[4]), .Y(n216) );
  AOI221XL U772 ( .A(r_dac_en[3]), .B(n559), .C(n9), .D(n215), .E(n219), .Y(
        n212) );
  ENOX1 U773 ( .A(n200), .B(n556), .C(n561), .D(r_dac_en[11]), .Y(n219) );
  INVX1 U774 ( .A(o_dat[5]), .Y(n566) );
  INVX1 U775 ( .A(o_dat[1]), .Y(n567) );
  ENOX1 U776 ( .A(n217), .B(n550), .C(n558), .D(r_dac_en[5]), .Y(n218) );
  ENOX1 U777 ( .A(n200), .B(n528), .C(n561), .D(r_dac_en[10]), .Y(n220) );
  ENOX1 U778 ( .A(n151), .B(n116), .C(o_dat[17]), .D(n151), .Y(datcmp[17]) );
  OAI21X1 U779 ( .B(n142), .C(n448), .A(n449), .Y(datcmp[8]) );
  OAI21X1 U780 ( .B(n162), .C(n142), .A(o_dat[8]), .Y(n449) );
  OAI21X1 U781 ( .B(n155), .C(n448), .A(n454), .Y(datcmp[12]) );
  OAI21X1 U782 ( .B(n162), .C(n155), .A(o_dat[12]), .Y(n454) );
  OAI21X1 U783 ( .B(n142), .C(n446), .A(n447), .Y(datcmp[9]) );
  OAI21X1 U784 ( .B(n161), .C(n142), .A(o_dat[9]), .Y(n447) );
  OAI21X1 U785 ( .B(n155), .C(n446), .A(n453), .Y(datcmp[13]) );
  OAI21X1 U786 ( .B(n161), .C(n155), .A(o_dat[13]), .Y(n453) );
  OAI21X1 U787 ( .B(n150), .C(n448), .A(n455), .Y(datcmp[0]) );
  OAI21X1 U788 ( .B(n162), .C(n150), .A(o_dat[0]), .Y(n455) );
  OAI21X1 U789 ( .B(n147), .C(n448), .A(n451), .Y(datcmp[4]) );
  OAI21X1 U790 ( .B(n162), .C(n147), .A(o_dat[4]), .Y(n451) );
  ENOX1 U791 ( .A(n153), .B(n116), .C(o_dat[15]), .D(n153), .Y(datcmp[15]) );
  ENOX1 U792 ( .A(n152), .B(n116), .C(o_dat[16]), .D(n152), .Y(datcmp[16]) );
  ENOX1 U793 ( .A(n157), .B(n116), .C(o_dat[10]), .D(n157), .Y(datcmp[10]) );
  ENOX1 U794 ( .A(n154), .B(n116), .C(o_dat[14]), .D(n154), .Y(datcmp[14]) );
  ENOX1 U795 ( .A(n156), .B(n116), .C(o_dat[11]), .D(n156), .Y(datcmp[11]) );
  ENOX1 U796 ( .A(n149), .B(n116), .C(n149), .D(o_dat[2]), .Y(datcmp[2]) );
  ENOX1 U797 ( .A(n148), .B(n116), .C(n148), .D(o_dat[3]), .Y(datcmp[3]) );
  ENOX1 U798 ( .A(n145), .B(n116), .C(n145), .D(o_dat[7]), .Y(datcmp[7]) );
  ENOX1 U799 ( .A(n146), .B(n116), .C(n146), .D(o_dat[6]), .Y(datcmp[6]) );
  NAND2X1 U800 ( .A(syn_comp[1]), .B(n563), .Y(n446) );
  NAND2X1 U801 ( .A(syn_comp[1]), .B(n562), .Y(n448) );
  INVX1 U802 ( .A(syn_comp[1]), .Y(n116) );
  NAND32XL U803 ( .B(n92), .C(n49), .A(n249), .Y(n248) );
  INVXL U804 ( .A(dacv_wr[11]), .Y(n537) );
  OAI22AXL U805 ( .D(dacv_wr[9]), .C(n82), .A(n142), .B(n143), .Y(upd[9]) );
  INVXL U806 ( .A(dacv_wr[9]), .Y(n225) );
  OAI22AXL U807 ( .D(dacv_wr[8]), .C(n83), .A(n142), .B(n144), .Y(upd[8]) );
  INVXL U808 ( .A(dacv_wr[8]), .Y(n227) );
  BUFXL U809 ( .A(n104), .Y(n103) );
  BUFXL U810 ( .A(r_wdat[0]), .Y(n104) );
  INVXL U811 ( .A(dacv_wr[15]), .Y(n245) );
  MUX2XL U812 ( .D0(n103), .D1(r_rpt_v[0]), .S(n67), .Y(wdlsb[0]) );
  NAND6XL U813 ( .A(r_wdat[6]), .B(n103), .C(n241), .D(n533), .E(n243), .F(
        n532), .Y(n242) );
  NAND21XL U814 ( .B(n104), .A(r_wr[0]), .Y(n249) );
endmodule


module dacmux_a0_DW01_add_19 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55;

  FAD1X1 U3 ( .A(B[6]), .B(A[6]), .CI(n4), .CO(n3), .SO(SUM[6]) );
  FAD1X1 U4 ( .A(B[5]), .B(A[5]), .CI(n5), .CO(n4), .SO(SUM[5]) );
  FAD1X1 U5 ( .A(B[4]), .B(A[4]), .CI(n6), .CO(n5), .SO(SUM[4]) );
  FAD1X1 U6 ( .A(B[3]), .B(A[3]), .CI(n7), .CO(n6), .SO(SUM[3]) );
  FAD1X1 U7 ( .A(B[2]), .B(A[2]), .CI(n8), .CO(n7), .SO(SUM[2]) );
  FAD1X1 U8 ( .A(B[1]), .B(A[1]), .CI(n11), .CO(n8), .SO(SUM[1]) );
  INVX2 U19 ( .A(n10), .Y(n11) );
  NAND3X1 U20 ( .A(n54), .B(n53), .C(n52), .Y(n2) );
  INVX1 U21 ( .A(n2), .Y(n46) );
  NAND2X1 U22 ( .A(n2), .B(n55), .Y(n48) );
  NAND2X2 U23 ( .A(n46), .B(n47), .Y(n49) );
  NAND2X2 U24 ( .A(n48), .B(n49), .Y(SUM[8]) );
  INVX1 U25 ( .A(n55), .Y(n47) );
  INVXL U26 ( .A(n55), .Y(n50) );
  INVX1 U27 ( .A(B[8]), .Y(n55) );
  XOR2XL U28 ( .A(A[7]), .B(n50), .Y(n51) );
  XOR2XL U29 ( .A(n51), .B(n3), .Y(SUM[7]) );
  NAND2XL U30 ( .A(n3), .B(B[7]), .Y(n52) );
  NAND2XL U31 ( .A(n3), .B(A[7]), .Y(n53) );
  NAND2X1 U32 ( .A(n50), .B(A[7]), .Y(n54) );
  NAND2X2 U33 ( .A(B[0]), .B(A[0]), .Y(n10) );
  NOR2XL U34 ( .A(B[0]), .B(A[0]), .Y(n9) );
  INVX1 U35 ( .A(n1), .Y(SUM[0]) );
  NAND21XL U36 ( .B(n9), .A(n10), .Y(n1) );
endmodule


module dacmux_a0_DW01_add_18 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n13, n14, n15, n16, n17, n18, n56,
         n57;

  FAD1X1 U2 ( .A(B[7]), .B(A[7]), .CI(n5), .CO(n4), .SO(SUM[7]) );
  FAD1X1 U3 ( .A(B[6]), .B(A[6]), .CI(n6), .CO(n5), .SO(SUM[6]) );
  FAD1X1 U4 ( .A(B[5]), .B(A[5]), .CI(n7), .CO(n6), .SO(SUM[5]) );
  FAD1X1 U5 ( .A(B[4]), .B(A[4]), .CI(n8), .CO(n7), .SO(SUM[4]) );
  FAD1X1 U6 ( .A(B[3]), .B(A[3]), .CI(n57), .CO(n8), .SO(SUM[3]) );
  XOR2X1 U16 ( .A(n2), .B(n18), .Y(SUM[1]) );
  OAI21X1 U17 ( .B(n15), .C(n18), .A(n16), .Y(n14) );
  NOR2X1 U25 ( .A(B[0]), .B(A[0]), .Y(n17) );
  NOR2XL U31 ( .A(B[1]), .B(A[1]), .Y(n15) );
  NAND2X1 U32 ( .A(B[0]), .B(A[0]), .Y(n18) );
  OR2X1 U33 ( .A(B[2]), .B(A[2]), .Y(n56) );
  XOR2X1 U34 ( .A(n4), .B(B[8]), .Y(SUM[8]) );
  NAND21XL U35 ( .B(n15), .A(n16), .Y(n2) );
  NAND2XL U36 ( .A(B[2]), .B(A[2]), .Y(n13) );
  NAND21XL U37 ( .B(n17), .A(n18), .Y(n3) );
  XNOR2XL U38 ( .A(n1), .B(n14), .Y(SUM[2]) );
  NAND2X1 U39 ( .A(n56), .B(n13), .Y(n1) );
  OAI21BBX1 U40 ( .A(n14), .B(n56), .C(n13), .Y(n57) );
  NAND2XL U41 ( .A(B[1]), .B(A[1]), .Y(n16) );
  INVX1 U42 ( .A(n3), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_17 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2XL U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_16 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2XL U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_15 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  XOR2X1 U3 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_14 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2XL U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_13 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2XL U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_12 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2XL U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_11 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2XL U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_10 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2XL U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_9 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  NAND2X1 U1 ( .A(B[5]), .B(A[5]), .Y(n4) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U3 ( .A(A[5]), .B(B[5]), .Y(n1) );
  XOR2XL U4 ( .A(n1), .B(carry[5]), .Y(SUM[5]) );
  NAND2X1 U5 ( .A(carry[5]), .B(B[5]), .Y(n2) );
  NAND2XL U6 ( .A(carry[5]), .B(A[5]), .Y(n3) );
  NAND3X1 U7 ( .A(n4), .B(n3), .C(n2), .Y(carry[6]) );
  XOR3XL U8 ( .A(carry[6]), .B(B[6]), .C(A[6]), .Y(SUM[6]) );
  NAND2XL U9 ( .A(carry[6]), .B(B[6]), .Y(n5) );
  NAND2XL U10 ( .A(carry[6]), .B(A[6]), .Y(n6) );
  NAND2X1 U11 ( .A(B[6]), .B(A[6]), .Y(n7) );
  NAND3X1 U12 ( .A(n7), .B(n6), .C(n5), .Y(carry[7]) );
  AND2X2 U13 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U14 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [8:2] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  NAND2XL U1 ( .A(A[1]), .B(B[1]), .Y(n3) );
  NAND3X2 U2 ( .A(n3), .B(n4), .C(n5), .Y(carry[2]) );
  NAND2XL U3 ( .A(n10), .B(carry[8]), .Y(n8) );
  NAND2X1 U4 ( .A(n6), .B(n7), .Y(n9) );
  NAND2X1 U5 ( .A(n8), .B(n9), .Y(SUM[8]) );
  INVX1 U6 ( .A(n10), .Y(n6) );
  INVX1 U7 ( .A(carry[8]), .Y(n7) );
  INVX1 U8 ( .A(B[8]), .Y(n10) );
  AND2X2 U9 ( .A(A[0]), .B(B[0]), .Y(n11) );
  NAND2X1 U10 ( .A(A[1]), .B(n11), .Y(n4) );
  NAND2X1 U11 ( .A(B[1]), .B(n11), .Y(n5) );
  XOR2XL U12 ( .A(n2), .B(n11), .Y(SUM[1]) );
  XOR2XL U13 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2XL U14 ( .A(A[1]), .B(B[1]), .Y(n2) );
endmodule


module dacmux_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4;
  wire   [8:1] carry;

  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR3XL U2 ( .A(carry[7]), .B(B[7]), .C(A[7]), .Y(SUM[7]) );
  NAND2XL U3 ( .A(carry[7]), .B(B[7]), .Y(n2) );
  NAND2XL U4 ( .A(carry[7]), .B(A[7]), .Y(n3) );
  NAND2X1 U5 ( .A(B[7]), .B(A[7]), .Y(n4) );
  NAND3X1 U6 ( .A(n4), .B(n3), .C(n2), .Y(carry[8]) );
  XOR2X1 U7 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U8 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_6 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  INVX1 U1 ( .A(A[0]), .Y(n3) );
  INVX1 U2 ( .A(B[0]), .Y(n4) );
  NOR2X4 U3 ( .A(n3), .B(n4), .Y(carry[1]) );
  XNOR2X1 U4 ( .A(n5), .B(carry[8]), .Y(SUM[8]) );
  INVXL U5 ( .A(B[8]), .Y(n5) );
  XOR2XL U6 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_5 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  INVX1 U1 ( .A(n11), .Y(n3) );
  NAND2X1 U2 ( .A(n11), .B(carry[8]), .Y(n5) );
  NAND2X2 U3 ( .A(n3), .B(n4), .Y(n6) );
  NAND2X2 U4 ( .A(n5), .B(n6), .Y(SUM[8]) );
  INVX1 U5 ( .A(carry[8]), .Y(n4) );
  XOR2X1 U6 ( .A(A[5]), .B(B[5]), .Y(n7) );
  XOR2XL U7 ( .A(n7), .B(carry[5]), .Y(SUM[5]) );
  NAND2X1 U8 ( .A(carry[5]), .B(B[5]), .Y(n8) );
  NAND2XL U9 ( .A(carry[5]), .B(A[5]), .Y(n9) );
  NAND2X1 U10 ( .A(B[5]), .B(A[5]), .Y(n10) );
  NAND3X1 U11 ( .A(n10), .B(n9), .C(n8), .Y(carry[6]) );
  AND2X2 U12 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  INVXL U13 ( .A(B[8]), .Y(n11) );
  XOR2XL U14 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[6]), .B(B[6]), .Y(n8) );
  NAND2X1 U2 ( .A(n2), .B(n3), .Y(n5) );
  INVX1 U3 ( .A(n17), .Y(n2) );
  INVX1 U4 ( .A(B[5]), .Y(n10) );
  INVX1 U5 ( .A(A[5]), .Y(n9) );
  INVX1 U6 ( .A(B[6]), .Y(n7) );
  NAND2X1 U7 ( .A(n17), .B(carry[8]), .Y(n4) );
  NAND2X2 U8 ( .A(n4), .B(n5), .Y(SUM[8]) );
  INVX1 U9 ( .A(carry[8]), .Y(n3) );
  INVXL U10 ( .A(n17), .Y(n6) );
  INVX1 U11 ( .A(B[8]), .Y(n17) );
  NAND21X1 U12 ( .B(n7), .A(carry[6]), .Y(n16) );
  NAND31X4 U13 ( .C(n8), .A(n15), .B(n16), .Y(carry[7]) );
  NAND21XL U14 ( .B(n9), .A(carry[5]), .Y(n12) );
  NAND21XL U15 ( .B(n10), .A(carry[5]), .Y(n13) );
  XOR3XL U16 ( .A(A[5]), .B(B[5]), .C(carry[5]), .Y(SUM[5]) );
  NAND2X1 U17 ( .A(A[5]), .B(B[5]), .Y(n11) );
  NAND3X4 U18 ( .A(n11), .B(n12), .C(n13), .Y(carry[6]) );
  XOR2XL U19 ( .A(A[6]), .B(B[6]), .Y(n14) );
  XOR2XL U20 ( .A(n14), .B(carry[6]), .Y(SUM[6]) );
  NAND2X1 U21 ( .A(A[6]), .B(carry[6]), .Y(n15) );
  AND2XL U22 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U23 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X2 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(n7), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  NAND2XL U1 ( .A(n12), .B(carry[8]), .Y(n5) );
  NAND3X1 U2 ( .A(n11), .B(n10), .C(n9), .Y(carry[4]) );
  NAND2X1 U3 ( .A(n5), .B(n6), .Y(SUM[8]) );
  NAND2X1 U4 ( .A(n3), .B(n4), .Y(n6) );
  INVX1 U5 ( .A(n12), .Y(n3) );
  INVX1 U6 ( .A(carry[8]), .Y(n4) );
  INVXL U7 ( .A(n12), .Y(n7) );
  XOR2X1 U8 ( .A(A[3]), .B(B[3]), .Y(n8) );
  XOR2XL U9 ( .A(n8), .B(carry[3]), .Y(SUM[3]) );
  NAND2XL U10 ( .A(carry[3]), .B(B[3]), .Y(n9) );
  NAND2XL U11 ( .A(carry[3]), .B(A[3]), .Y(n10) );
  NAND2X1 U12 ( .A(B[3]), .B(A[3]), .Y(n11) );
  AND2X1 U13 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  INVX1 U14 ( .A(B[8]), .Y(n12) );
  XOR2XL U15 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module glreg_WIDTH2_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n4, n5, n1;

  SDFFRQX1 mem_reg_0_ ( .D(n5), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(n4), .SIN(rdat[0]), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[1]) );
  AO22XL U2 ( .A(wdat[1]), .B(we), .C(rdat[1]), .D(n1), .Y(n4) );
  INVXL U3 ( .A(we), .Y(n1) );
  AO22XL U4 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(n1), .Y(n5) );
endmodule


module glreg_WIDTH2_1 ( clk, arstz, we, wdat, rdat, test_si, test_so, test_se
 );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  output test_so;
  wire   n8, n9;

  SDFFRQX1 mem_reg_0_ ( .D(n9), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(n8), .SIN(rdat[0]), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[1]) );
  AO22AXL U2 ( .A(wdat[1]), .B(we), .C(rdat[1]), .D(we), .Y(n8) );
  BUFX3 U3 ( .A(rdat[1]), .Y(test_so) );
  AO22AXL U4 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n9) );
endmodule


module glreg_a0_26 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9717;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_26 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9717), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9717), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9717), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9717), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9717), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9717), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9717), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9717), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9717), 
        .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_27 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n11, n12, n13, n14, n15, net9735, n1, n3, n5, n7, n9;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_27 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9735), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9735), 
        .XR(arstz), .Q(n15) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9735), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9735), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(n15), .SMC(test_se), .C(net9735), 
        .XR(arstz), .Q(n14) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(n12), .SMC(test_se), .C(net9735), 
        .XR(arstz), .Q(n11) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(n13), .SMC(test_se), .C(net9735), 
        .XR(arstz), .Q(n12) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(n14), .SMC(test_se), .C(net9735), 
        .XR(arstz), .Q(n13) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(n11), .SMC(test_se), .C(net9735), 
        .XR(arstz), .Q(rdat[7]) );
  INVXL U2 ( .A(n13), .Y(n1) );
  INVXL U3 ( .A(n1), .Y(rdat[4]) );
  INVXL U4 ( .A(n12), .Y(n3) );
  INVXL U5 ( .A(n3), .Y(rdat[5]) );
  INVXL U6 ( .A(n15), .Y(n5) );
  INVXL U7 ( .A(n5), .Y(rdat[2]) );
  INVXL U8 ( .A(n14), .Y(n7) );
  INVXL U9 ( .A(n7), .Y(rdat[3]) );
  INVX1 U10 ( .A(n11), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_28 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9753;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_28 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9753), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9753), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9753), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9753), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9753), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9753), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9753), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9753), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9753), 
        .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_29 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9771;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_29 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9771), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9771), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9771), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9771), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9771), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQXX2 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9771), .XR(arstz), .Q(rdat[0]), .XQ() );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9771), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9771), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX2 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9771), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_1 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_1 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[0]), .Y(n9) );
  INVX1 U4 ( .A(set2[1]), .Y(n10) );
  INVX1 U5 ( .A(set2[2]), .Y(n11) );
  INVX1 U6 ( .A(set2[3]), .Y(n12) );
  INVX1 U7 ( .A(set2[4]), .Y(n13) );
  NAND3X1 U8 ( .A(n15), .B(n16), .C(n14), .Y(n21) );
  INVX1 U9 ( .A(set2[6]), .Y(n15) );
  INVX1 U10 ( .A(set2[7]), .Y(n16) );
  INVX1 U11 ( .A(set2[5]), .Y(n14) );
  AOI211X1 U12 ( .C(n10), .D(n8), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U13 ( .A(rdat[1]), .Y(n8) );
  AOI211X1 U14 ( .C(n14), .D(n3), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U15 ( .A(rdat[5]), .Y(n3) );
  NAND4X1 U16 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U17 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U18 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U19 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U20 ( .C(n11), .D(n7), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U21 ( .A(rdat[2]), .Y(n7) );
  AOI211X1 U22 ( .C(n12), .D(n5), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U23 ( .A(rdat[3]), .Y(n5) );
  AOI211X1 U24 ( .C(n15), .D(n2), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U25 ( .A(rdat[6]), .Y(n2) );
  AOI211X1 U26 ( .C(n16), .D(n1), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U27 ( .A(rdat[7]), .Y(n1) );
  AOI211X1 U28 ( .C(n9), .D(n6), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U29 ( .A(rdat[0]), .Y(n6) );
  AOI211X1 U30 ( .C(n13), .D(n4), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U31 ( .A(rdat[4]), .Y(n4) );
  NOR2X1 U32 ( .A(rdat[5]), .B(n14), .Y(irq[5]) );
  NOR2X1 U33 ( .A(rdat[1]), .B(n10), .Y(irq[1]) );
  NOR2X1 U34 ( .A(rdat[0]), .B(n9), .Y(irq[0]) );
  NOR2X1 U35 ( .A(rdat[4]), .B(n13), .Y(irq[4]) );
  NOR2X1 U36 ( .A(rdat[6]), .B(n15), .Y(irq[6]) );
  NOR2X1 U37 ( .A(rdat[2]), .B(n11), .Y(irq[2]) );
  NOR2X1 U38 ( .A(rdat[7]), .B(n16), .Y(irq[7]) );
  NOR2X1 U39 ( .A(rdat[3]), .B(n12), .Y(irq[3]) );
endmodule


module glreg_WIDTH8_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9789;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9789), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9789), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9789), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9789), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9789), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9789), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9789), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9789), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9789), 
        .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_30 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9807;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_30 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9807), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9807), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9807), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9807), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9807), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9807), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9807), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9807), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9807), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_31 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9825;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_31 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9825), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9825), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9825), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9825), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9825), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9825), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9825), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9825), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9825), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_32 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9843;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_32 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9843), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9843), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9843), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9843), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9843), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9843), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9843), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9843), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9843), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_33 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9861;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_33 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9861), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9861), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9861), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9861), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9861), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9861), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9861), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9861), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9861), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_34 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9879;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_34 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9879), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9879), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9879), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9879), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9879), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9879), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9879), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9879), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9879), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_35 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9897;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_35 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9897), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9897), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9897), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9897), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9897), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9897), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9897), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9897), 
        .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9897), 
        .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_36 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9915;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_36 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9915), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9915), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9915), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9915), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9915), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9915), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9915), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9915), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9915), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_37 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9933;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_37 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9933), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9933), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9933), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9933), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9933), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9933), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9933), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9933), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9933), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_38 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9951;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_38 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9951), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9951), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9951), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9951), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9951), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9951), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9951), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9951), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9951), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_39 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9969;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_39 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9969), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9969), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9969), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9969), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9969), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9969), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9969), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9969), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9969), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_40 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net9987;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_40 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9987), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net9987), 
        .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net9987), 
        .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net9987), 
        .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net9987), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net9987), 
        .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net9987), 
        .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net9987), 
        .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net9987), 
        .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_41 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10005;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_41 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10005), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10005), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10005), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10005), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10005), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10005), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10005), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10005), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10005), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_42 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10023;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_42 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10023), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10023), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10023), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10023), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10023), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10023), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10023), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10023), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10023), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_43 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10041;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_43 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10041), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10041), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10041), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10041), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10041), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10041), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10041), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10041), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10041), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_44 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10059;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_44 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10059), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10059), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10059), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10059), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10059), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10059), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10059), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10059), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10059), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_45 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10077;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_45 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10077), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10077), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10077), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10077), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10077), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10077), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10077), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10077), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10077), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_46 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10095;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_46 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10095), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10095), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10095), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10095), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10095), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10095), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10095), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10095), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10095), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_47 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10113;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_47 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10113), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10113), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10113), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10113), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10113), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10113), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10113), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10113), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10113), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10131;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10131), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10131), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10131), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10131), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10131), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10131), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10131), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_48 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10149;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_48 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10149), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10149), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10149), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10149), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10149), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10149), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10149), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10149), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10149), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_49 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n7, n8, n9, net10167, n1, n3, n5;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_49 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10167), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(n7), .SMC(test_se), .C(net10167), 
        .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10167), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10167), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10167), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(n8), .SMC(test_se), .C(net10167), 
        .XR(arstz), .Q(n7) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10167), .XR(arstz), .Q(n8) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10167), .XR(arstz), .Q(n9) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(n9), .SMC(test_se), .C(net10167), 
        .XR(arstz), .Q(rdat[1]) );
  INVXL U2 ( .A(n9), .Y(n1) );
  INVXL U3 ( .A(n1), .Y(rdat[0]) );
  INVXL U4 ( .A(n8), .Y(n3) );
  INVXL U5 ( .A(n3), .Y(rdat[2]) );
  INVXL U6 ( .A(n7), .Y(n5) );
  INVXL U7 ( .A(n5), .Y(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH7_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10185;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10185), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10185), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10185), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10185), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10185), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10185), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10185), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10185), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module shmux_00000005_00000012_00000012 ( ps_md4ch, r_comp_swtch, r_semi, 
        r_loop, r_dac_en, wr_dacv, busy, sh_hold, stop, semi_start, auto_start, 
        mxcyc_done, sampl_begn, sampl_done, app_dacis, pos_dacis, cs_ptr, 
        ps_ptr, clk, srstz, test_si2, test_si1, test_so1, test_se );
  input [17:0] r_dac_en;
  input [17:0] wr_dacv;
  output [17:0] app_dacis;
  output [17:0] pos_dacis;
  output [4:0] cs_ptr;
  output [4:0] ps_ptr;
  input ps_md4ch, r_comp_swtch, r_semi, r_loop, stop, semi_start, auto_start,
         mxcyc_done, sampl_begn, sampl_done, clk, srstz, test_si2, test_si1,
         test_se;
  output busy, sh_hold, test_so1;
  wire   cs_mux_5_, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958,
         N959, N960, N961, N962, N963, N964, N965, N966, N967, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N994, N995, N996, N997, N998,
         N999, N1139, N1148, N1230, N1262, N1271, N1312, N1394, net10203,
         net10221, net10226, n671, n1, n37, n38, n39, n43, n47, n51, n54, n56,
         n79, n80, n82, n736, n735, n734, n820, n821, n822, n823, n824, n825,
         n192, n193, n195, n197, n198, n200, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n238, n239, n240, n241, n242, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n255, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n301, n304, n305, n306, n308, n309, n310, n311, n312, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n375, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n458, n459, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n502, n503, n505, n506, n507, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n592, n593, n594,
         n595, n649, n652, n654, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n41, n44, n45, n46, n48,
         n49, n52, n53, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n81, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n194, n196, n199, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n243, n253, n254, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n302, n303, n307, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n374, n376, n392,
         n412, n439, n457, n460, n472, n501, n504, n508, n520, n553, n574,
         n591, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n650,
         n651, n653, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733;
  wire   [16:4] neg_dacis;
  wire   [5:4] sub_398_S2_I7_aco_carry;
  wire   [5:4] sub_398_S2_I5_aco_carry;
  wire   [5:4] sub_398_S2_I4_aco_carry;
  wire   [5:4] sub_398_S2_I3_aco_carry;
  wire   [5:4] sub_398_S2_aco_carry;

  FAD1X1 sub_398_S2_I7_aco_U2_4 ( .A(n722), .B(n80), .CI(
        sub_398_S2_I7_aco_carry[4]), .CO(sub_398_S2_I7_aco_carry[5]), .SO(
        N1394) );
  FAD1X1 sub_398_S2_I5_aco_U2_4 ( .A(n721), .B(n708), .CI(
        sub_398_S2_I5_aco_carry[4]), .CO(sub_398_S2_I5_aco_carry[5]), .SO(
        N1312) );
  FAD1X1 sub_398_S2_I4_aco_U2_4 ( .A(N1262), .B(n1), .CI(
        sub_398_S2_I4_aco_carry[4]), .CO(sub_398_S2_I4_aco_carry[5]), .SO(
        N1271) );
  FAD1X1 sub_398_S2_I3_aco_U2_4 ( .A(n720), .B(n82), .CI(
        sub_398_S2_I3_aco_carry[4]), .CO(sub_398_S2_I3_aco_carry[5]), .SO(
        N1230) );
  FAD1X1 sub_398_S2_aco_U2_4 ( .A(N1139), .B(n79), .CI(sub_398_S2_aco_carry[4]), .CO(sub_398_S2_aco_carry[5]), .SO(N1148) );
  SNPS_CLOCK_GATE_LOW_shmux_00000005_00000012_00000012 clk_gate_neg_dacis_reg ( 
        .CLK(clk), .EN(N949), .ENCLK(net10203), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 clk_gate_r_dacis_reg ( 
        .CLK(clk), .EN(N971), .ENCLK(net10221), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 clk_gate_cs_mux_reg ( 
        .CLK(clk), .EN(N994), .ENCLK(net10226), .TE(test_se) );
  SDFFQX1 cs_mux_reg_3_ ( .D(N998), .SIN(n18), .SMC(test_se), .C(net10226), 
        .Q(cs_ptr[3]) );
  SDFFQX1 cs_mux_reg_1_ ( .D(N996), .SIN(n45), .SMC(test_se), .C(net10226), 
        .Q(n735) );
  SDFFQX1 cs_mux_reg_4_ ( .D(N999), .SIN(n19), .SMC(test_se), .C(net10226), 
        .Q(n734) );
  SDFFQX1 cs_mux_reg_2_ ( .D(N997), .SIN(n735), .SMC(test_se), .C(net10226), 
        .Q(cs_ptr[2]) );
  SDFFQX1 cs_mux_reg_0_ ( .D(N995), .SIN(test_si2), .SMC(test_se), .C(net10226), .Q(n736) );
  SDFFQX1 r_dacis_reg_17_ ( .D(N989), .SIN(pos_dacis[16]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[17]) );
  SDFFQX1 r_dacis_reg_16_ ( .D(N988), .SIN(pos_dacis[15]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[16]) );
  SDFFQX1 r_dacis_reg_15_ ( .D(N987), .SIN(pos_dacis[14]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[15]) );
  SDFFQX1 r_dacis_reg_14_ ( .D(N986), .SIN(pos_dacis[13]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[14]) );
  SDFFQX1 cs_mux_reg_5_ ( .D(n671), .SIN(n53), .SMC(test_se), .C(clk), .Q(
        cs_mux_5_) );
  SDFFQX1 r_dacis_reg_12_ ( .D(N984), .SIN(pos_dacis[11]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[12]) );
  SDFFQX1 r_dacis_reg_13_ ( .D(N985), .SIN(pos_dacis[12]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[13]) );
  SDFFQX1 r_dacis_reg_10_ ( .D(N982), .SIN(pos_dacis[9]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[10]) );
  SDFFQX1 r_dacis_reg_11_ ( .D(N983), .SIN(pos_dacis[10]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[11]) );
  SDFFQX1 r_dacis_reg_9_ ( .D(N981), .SIN(pos_dacis[8]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[9]) );
  SDFFQX1 r_dacis_reg_8_ ( .D(N980), .SIN(pos_dacis[7]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[8]) );
  SDFFQX1 r_dacis_reg_7_ ( .D(N979), .SIN(pos_dacis[6]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[7]) );
  SDFFQX1 r_dacis_reg_5_ ( .D(N977), .SIN(pos_dacis[4]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[5]) );
  SDFFQX1 r_dacis_reg_4_ ( .D(N976), .SIN(pos_dacis[3]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[4]) );
  SDFFQX1 r_dacis_reg_6_ ( .D(N978), .SIN(pos_dacis[5]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[6]) );
  SDFFQX1 r_dacis_reg_2_ ( .D(N974), .SIN(pos_dacis[1]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[2]) );
  SDFFQX1 r_dacis_reg_1_ ( .D(N973), .SIN(pos_dacis[0]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[1]) );
  SDFFQX1 r_dacis_reg_0_ ( .D(N972), .SIN(cs_mux_5_), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[0]) );
  SDFFQX1 r_dacis_reg_3_ ( .D(N975), .SIN(pos_dacis[2]), .SMC(test_se), .C(
        net10221), .Q(pos_dacis[3]) );
  SDFFNQX4 neg_dacis_reg_12_ ( .D(N962), .SIN(n825), .SMC(test_se), .XC(
        net10203), .Q(neg_dacis[12]) );
  SDFFNQX4 neg_dacis_reg_4_ ( .D(N954), .SIN(n822), .SMC(test_se), .XC(
        net10203), .Q(neg_dacis[4]) );
  SDFFNQX4 neg_dacis_reg_9_ ( .D(N959), .SIN(n608), .SMC(test_se), .XC(
        net10203), .Q(neg_dacis[9]) );
  SDFFNQX4 neg_dacis_reg_16_ ( .D(N966), .SIN(n605), .SMC(test_se), .XC(
        net10203), .Q(neg_dacis[16]) );
  SDFFNQXX4 neg_dacis_reg_6_ ( .D(N956), .SIN(n604), .SMC(test_se), .XC(
        net10203), .Q(n607), .XQ(n43) );
  SDFFNQXX4 neg_dacis_reg_17_ ( .D(N967), .SIN(neg_dacis[16]), .SMC(test_se), 
        .XC(net10203), .Q(test_so1), .XQ(n37) );
  SDFFNQXX4 neg_dacis_reg_2_ ( .D(N952), .SIN(n821), .SMC(test_se), .XC(
        net10203), .Q(n823), .XQ(n7) );
  SDFFNQXX4 neg_dacis_reg_14_ ( .D(N964), .SIN(neg_dacis[13]), .SMC(test_se), 
        .XC(net10203), .Q(n606), .XQ(n51) );
  SDFFNQXX4 neg_dacis_reg_15_ ( .D(N965), .SIN(n606), .SMC(test_se), .XC(
        net10203), .Q(n605), .XQ(n56) );
  SDFFNQXX4 neg_dacis_reg_7_ ( .D(N957), .SIN(n607), .SMC(test_se), .XC(
        net10203), .Q(n38), .XQ(n39) );
  SDFFNQXX4 neg_dacis_reg_11_ ( .D(N961), .SIN(n820), .SMC(test_se), .XC(
        net10203), .Q(n825), .XQ(n4) );
  SDFFNQXX4 neg_dacis_reg_0_ ( .D(N950), .SIN(test_si1), .SMC(test_se), .XC(
        net10203), .Q(n824), .XQ(n5) );
  SDFFNQXX4 neg_dacis_reg_1_ ( .D(N951), .SIN(n824), .SMC(test_se), .XC(
        net10203), .Q(n821), .XQ(n3) );
  SDFFNQXX4 neg_dacis_reg_10_ ( .D(N960), .SIN(neg_dacis[9]), .SMC(test_se), 
        .XC(net10203), .Q(n820), .XQ(n2) );
  SDFFNQXX4 neg_dacis_reg_8_ ( .D(N958), .SIN(n38), .SMC(test_se), .XC(
        net10203), .Q(n608), .XQ(n47) );
  SDFFNQXX4 neg_dacis_reg_5_ ( .D(N955), .SIN(neg_dacis[4]), .SMC(test_se), 
        .XC(net10203), .Q(n604), .XQ(n54) );
  SDFFNQXX4 neg_dacis_reg_3_ ( .D(N953), .SIN(n823), .SMC(test_se), .XC(
        net10203), .Q(n822), .XQ(n6) );
  SDFFNQX4 neg_dacis_reg_13_ ( .D(N963), .SIN(neg_dacis[12]), .SMC(test_se), 
        .XC(net10203), .Q(neg_dacis[13]) );
  OR3XL U3 ( .A(n357), .B(n189), .C(n165), .Y(n259) );
  NOR43XL U4 ( .B(n199), .C(n196), .D(n356), .A(n10), .Y(n201) );
  MUX2X1 U5 ( .D0(n640), .D1(n456), .S(cs_ptr[0]), .Y(n60) );
  MUX2X1 U6 ( .D0(n77), .D1(n76), .S(n263), .Y(n78) );
  OR3XL U7 ( .A(n187), .B(n253), .C(n259), .Y(n286) );
  OAI221X1 U8 ( .A(n263), .B(n349), .C(n22), .D(n350), .E(n262), .Y(ps_ptr[2])
         );
  OAI221X1 U9 ( .A(n206), .B(n349), .C(n205), .D(n350), .E(n204), .Y(ps_ptr[1]) );
  AOI221XL U10 ( .A(n203), .B(n351), .C(n599), .D(n202), .E(n201), .Y(n204) );
  INVX1 U11 ( .A(pos_dacis[16]), .Y(n14) );
  AOI21AX1 U12 ( .B(n313), .C(n646), .A(n307), .Y(n8) );
  INVX1 U13 ( .A(pos_dacis[13]), .Y(n15) );
  INVX3 U14 ( .A(n612), .Y(n9) );
  INVX3 U15 ( .A(n612), .Y(n21) );
  BUFXL U16 ( .A(r_dac_en[1]), .Y(n10) );
  INVXL U17 ( .A(n116), .Y(n11) );
  OR2X1 U18 ( .A(n617), .B(n13), .Y(N949) );
  NOR21XL U19 ( .B(n21), .A(n15), .Y(N963) );
  INVXL U20 ( .A(sampl_done), .Y(n12) );
  INVXL U21 ( .A(n12), .Y(n13) );
  NOR21XL U22 ( .B(n9), .A(n14), .Y(N966) );
  INVX1 U23 ( .A(n735), .Y(n16) );
  INVX1 U24 ( .A(n19), .Y(n17) );
  INVX1 U25 ( .A(n640), .Y(n18) );
  AO21X1 U26 ( .B(ps_md4ch), .C(n636), .A(n18), .Y(n665) );
  BUFX3 U27 ( .A(cs_ptr[3]), .Y(n19) );
  BUFX3 U28 ( .A(n732), .Y(n20) );
  NAND21X4 U29 ( .B(n617), .A(sampl_done), .Y(n612) );
  INVXL U30 ( .A(n111), .Y(n128) );
  NAND2X1 U31 ( .A(n129), .B(n128), .Y(n360) );
  OA222X1 U32 ( .A(n24), .B(n360), .C(n261), .D(n353), .E(n260), .F(n259), .Y(
        n262) );
  NAND21XL U33 ( .B(n25), .A(n113), .Y(n349) );
  INVXL U34 ( .A(wr_dacv[12]), .Y(n153) );
  AND2XL U35 ( .A(n350), .B(n349), .Y(n169) );
  XNOR2XL U36 ( .A(n529), .B(n695), .Y(n527) );
  OAI211X1 U37 ( .C(n317), .D(n360), .A(n316), .B(n315), .Y(ps_ptr[3]) );
  AOI32XL U38 ( .A(n303), .B(n302), .C(n300), .D(n599), .E(n299), .Y(n316) );
  NAND32X1 U39 ( .B(n130), .C(n129), .A(n128), .Y(n353) );
  INVXL U40 ( .A(n286), .Y(n303) );
  AND2XL U41 ( .A(ps_ptr[4]), .B(n318), .Y(N999) );
  OAI222XL U42 ( .A(n524), .B(n693), .C(n240), .D(n380), .E(n523), .F(n301), 
        .Y(n372) );
  AOI221XL U43 ( .A(n52), .B(n729), .C(n442), .D(n637), .E(n647), .Y(n567) );
  XNOR2XL U44 ( .A(n497), .B(n498), .Y(n244) );
  NAND32XL U45 ( .B(n188), .C(n243), .A(n287), .Y(n132) );
  INVXL U46 ( .A(n182), .Y(n183) );
  AND3XL U47 ( .A(n153), .B(n152), .C(n151), .Y(n156) );
  OAI211XL U48 ( .C(n150), .D(n180), .A(n149), .B(n148), .Y(n151) );
  AOI31XL U49 ( .A(n147), .B(n146), .C(n145), .D(n181), .Y(n150) );
  OAI211XL U50 ( .C(n17), .D(n289), .A(n288), .B(n287), .Y(n300) );
  INVXL U51 ( .A(n349), .Y(n457) );
  AOI221XL U52 ( .A(n647), .B(n729), .C(n57), .D(n442), .E(n637), .Y(n440) );
  AOI221XL U53 ( .A(n57), .B(n731), .C(n476), .D(n647), .E(n637), .Y(n479) );
  AOI221XL U54 ( .A(n647), .B(n730), .C(n57), .D(n537), .E(n637), .Y(n492) );
  XNOR2XL U55 ( .A(n537), .B(n638), .Y(n490) );
  INVXL U56 ( .A(n115), .Y(n194) );
  NAND21XL U57 ( .B(n19), .A(ps_ptr[3]), .Y(n348) );
  NOR42XL U58 ( .C(n193), .D(n192), .A(pos_dacis[2]), .B(pos_dacis[0]), .Y(
        n634) );
  INVX1 U59 ( .A(wr_dacv[1]), .Y(n196) );
  INVX1 U60 ( .A(wr_dacv[2]), .Y(n168) );
  INVX1 U61 ( .A(n462), .Y(n703) );
  INVX1 U62 ( .A(n313), .Y(n102) );
  INVX1 U63 ( .A(n95), .Y(n113) );
  INVX1 U64 ( .A(n360), .Y(n203) );
  INVX1 U65 ( .A(wr_dacv[10]), .Y(n154) );
  NOR2X1 U66 ( .A(n704), .B(n661), .Y(n465) );
  INVX1 U67 ( .A(n228), .Y(n600) );
  NOR2X1 U68 ( .A(n659), .B(n592), .Y(n583) );
  NOR2X1 U69 ( .A(n592), .B(n593), .Y(n580) );
  INVX1 U70 ( .A(n593), .Y(n659) );
  INVX1 U71 ( .A(n428), .Y(n711) );
  INVX1 U72 ( .A(n488), .Y(n690) );
  AOI21X1 U73 ( .B(n704), .C(n661), .A(n465), .Y(n462) );
  NOR2X1 U74 ( .A(n310), .B(n346), .Y(n386) );
  INVX1 U75 ( .A(n483), .Y(n691) );
  INVX1 U76 ( .A(n527), .Y(n692) );
  INVX1 U77 ( .A(n480), .Y(n687) );
  INVX1 U78 ( .A(n519), .Y(n264) );
  INVX1 U79 ( .A(n205), .Y(n392) );
  INVX1 U80 ( .A(n81), .Y(n99) );
  NAND21X1 U81 ( .B(n661), .A(n20), .Y(n81) );
  INVX1 U82 ( .A(n526), .Y(n694) );
  NAND21X1 U83 ( .B(n100), .A(n99), .Y(n313) );
  INVX1 U84 ( .A(n542), .Y(n657) );
  NAND21X1 U85 ( .B(auto_start), .A(n596), .Y(n95) );
  NAND21XL U86 ( .B(n95), .A(n25), .Y(n111) );
  INVX1 U87 ( .A(n353), .Y(n599) );
  INVX1 U88 ( .A(wr_dacv[16]), .Y(n147) );
  AO21X1 U89 ( .B(n355), .C(n354), .A(n353), .Y(n359) );
  AOI221XL U90 ( .A(n352), .B(n643), .C(n338), .D(n600), .E(n335), .Y(n354) );
  AND2X1 U91 ( .A(ps_ptr[3]), .B(n318), .Y(N998) );
  AND2X1 U92 ( .A(n331), .B(n332), .Y(N974) );
  AND2X1 U93 ( .A(n331), .B(n328), .Y(N978) );
  INVX1 U94 ( .A(N1312), .Y(n707) );
  NOR2X1 U95 ( .A(n435), .B(n655), .Y(n436) );
  INVX1 U96 ( .A(n653), .Y(n732) );
  AO22X1 U97 ( .A(n338), .B(n600), .C(n352), .D(n643), .Y(n179) );
  INVX1 U98 ( .A(n473), .Y(n704) );
  OA2222XL U99 ( .A(n178), .B(n290), .C(n177), .D(n295), .E(n700), .F(n294), 
        .G(n293), .H(n176), .Y(n355) );
  INVX1 U100 ( .A(n334), .Y(n178) );
  INVX1 U101 ( .A(n339), .Y(n177) );
  INVX1 U102 ( .A(n644), .Y(n176) );
  NAND21X1 U103 ( .B(n125), .A(n375), .Y(n228) );
  OA2222XL U104 ( .A(n295), .B(n717), .C(n542), .D(n294), .E(n564), .F(n293), 
        .G(n511), .H(n290), .Y(n127) );
  AOI21X1 U105 ( .B(n699), .C(n590), .A(n587), .Y(n593) );
  NAND21X1 U106 ( .B(n732), .A(n655), .Y(n393) );
  AOI21X1 U107 ( .B(n435), .C(n655), .A(n436), .Y(n428) );
  NAND2X1 U108 ( .A(n125), .B(n375), .Y(n295) );
  INVX1 U109 ( .A(N1148), .Y(n706) );
  INVX1 U110 ( .A(n589), .Y(n698) );
  NOR2X1 U111 ( .A(n653), .B(n82), .Y(n488) );
  INVX1 U112 ( .A(n643), .Y(n592) );
  INVX1 U113 ( .A(n347), .Y(n709) );
  NOR2X1 U114 ( .A(n393), .B(n79), .Y(n390) );
  NOR2X1 U115 ( .A(n659), .B(n643), .Y(n582) );
  NOR2X1 U116 ( .A(n690), .B(n478), .Y(n489) );
  NOR2X1 U117 ( .A(n643), .B(n593), .Y(n577) );
  INVX1 U118 ( .A(n478), .Y(n661) );
  NOR2X1 U119 ( .A(n590), .B(n699), .Y(n587) );
  INVX1 U120 ( .A(n255), .Y(n697) );
  INVX1 U121 ( .A(n466), .Y(n705) );
  INVX1 U122 ( .A(n281), .Y(n688) );
  AOI32X1 U123 ( .A(n567), .B(n568), .C(n569), .D(n723), .E(n716), .Y(n564) );
  INVX1 U124 ( .A(n567), .Y(n723) );
  AOI21X1 U125 ( .B(n653), .C(n82), .A(n488), .Y(n483) );
  INVX1 U126 ( .A(n568), .Y(n716) );
  OAI21X1 U127 ( .B(n417), .C(n699), .A(sub_398_S2_I4_aco_carry[4]), .Y(n278)
         );
  NAND2X1 U128 ( .A(n417), .B(n699), .Y(sub_398_S2_I4_aco_carry[4]) );
  NAND21X1 U129 ( .B(n390), .A(n635), .Y(n310) );
  XOR2X1 U130 ( .A(n653), .B(n716), .Y(n644) );
  AOI21X1 U131 ( .B(n478), .C(n690), .A(n489), .Y(n480) );
  NAND21X1 U132 ( .B(n529), .A(n530), .Y(n240) );
  XNOR2XL U133 ( .A(n531), .B(n532), .Y(n530) );
  NOR2X1 U134 ( .A(n645), .B(n393), .Y(n519) );
  NOR2X1 U135 ( .A(n535), .B(n478), .Y(n529) );
  NAND2X1 U136 ( .A(n732), .B(n532), .Y(n535) );
  NOR2X1 U137 ( .A(n732), .B(n79), .Y(n346) );
  OR2X1 U138 ( .A(n100), .B(n85), .Y(n307) );
  XOR2X1 U139 ( .A(n101), .B(n20), .Y(n205) );
  OAI21X1 U140 ( .B(n20), .C(n532), .A(n535), .Y(n526) );
  AOI21X1 U141 ( .B(n478), .C(n535), .A(n529), .Y(n301) );
  INVX1 U142 ( .A(n314), .Y(n70) );
  INVX1 U143 ( .A(n101), .Y(n100) );
  INVX1 U144 ( .A(n136), .Y(n110) );
  INVX1 U145 ( .A(n398), .Y(n684) );
  NAND21X1 U146 ( .B(n26), .A(n67), .Y(n137) );
  XOR2X1 U147 ( .A(n20), .B(n67), .Y(n69) );
  NAND2X1 U148 ( .A(n546), .B(n547), .Y(n542) );
  XNOR2XL U149 ( .A(n543), .B(n548), .Y(n546) );
  NOR2X1 U150 ( .A(n102), .B(n23), .Y(n22) );
  AOI21X1 U151 ( .B(n101), .C(n20), .A(n478), .Y(n23) );
  INVX1 U152 ( .A(n394), .Y(n727) );
  INVX1 U153 ( .A(n90), .Y(n175) );
  XNOR2XL U154 ( .A(n90), .B(n641), .Y(n24) );
  INVX1 U155 ( .A(n273), .Y(n296) );
  INVX1 U156 ( .A(n326), .Y(n615) );
  NAND32XL U157 ( .B(n129), .C(n111), .A(n130), .Y(n350) );
  OA22XL U158 ( .A(n314), .B(n349), .C(n8), .D(n350), .Y(n315) );
  INVX1 U159 ( .A(n254), .Y(n287) );
  NAND21X1 U160 ( .B(n44), .A(ps_ptr[0]), .Y(n460) );
  INVX1 U161 ( .A(n237), .Y(n258) );
  AND2XL U162 ( .A(ps_ptr[2]), .B(n318), .Y(N997) );
  AND2XL U163 ( .A(ps_ptr[1]), .B(n318), .Y(N996) );
  AND2X1 U164 ( .A(ps_ptr[0]), .B(n318), .Y(N995) );
  AND2X1 U165 ( .A(n614), .B(n29), .Y(N981) );
  AND2X1 U166 ( .A(n615), .B(n29), .Y(N980) );
  INVX1 U167 ( .A(n197), .Y(n318) );
  INVX1 U168 ( .A(n329), .Y(n332) );
  AND2X1 U169 ( .A(n616), .B(n615), .Y(N988) );
  AND2X1 U170 ( .A(n332), .B(n614), .Y(N973) );
  AND2X1 U171 ( .A(n324), .B(n614), .Y(N985) );
  AND2X1 U172 ( .A(n324), .B(n615), .Y(N984) );
  AND2X1 U173 ( .A(n324), .B(n331), .Y(N986) );
  AND2X1 U174 ( .A(n324), .B(n330), .Y(N987) );
  AND2X1 U175 ( .A(n330), .B(n332), .Y(N975) );
  AND2X1 U176 ( .A(n330), .B(n328), .Y(N979) );
  NOR21XL U177 ( .B(n330), .A(n649), .Y(N983) );
  AND2X1 U178 ( .A(n614), .B(n616), .Y(N989) );
  INVX1 U179 ( .A(n652), .Y(n328) );
  INVX1 U180 ( .A(n195), .Y(n708) );
  NAND2X1 U181 ( .A(n653), .B(n195), .Y(n435) );
  INVX1 U182 ( .A(n440), .Y(n721) );
  XOR2X1 U183 ( .A(n642), .B(n44), .Y(n653) );
  NOR21XL U184 ( .B(n362), .A(n363), .Y(n214) );
  OAI21X1 U185 ( .B(n653), .C(n195), .A(n435), .Y(n347) );
  OAI221X1 U186 ( .A(n458), .B(n703), .C(n380), .D(n702), .E(n459), .Y(n217)
         );
  GEN2XL U187 ( .D(n648), .E(n650), .C(n705), .B(n461), .A(n462), .Y(n459) );
  INVX1 U188 ( .A(N1394), .Y(n702) );
  AOI22X1 U189 ( .A(n466), .B(n467), .C(n468), .D(n705), .Y(n458) );
  AND3X1 U190 ( .A(n363), .B(n367), .C(n362), .Y(n250) );
  INVX1 U191 ( .A(n73), .Y(n655) );
  NOR2X1 U192 ( .A(n653), .B(n80), .Y(n473) );
  INVX1 U193 ( .A(n476), .Y(n731) );
  AOI22AXL U194 ( .A(n250), .B(n684), .D(n251), .C(n252), .Y(n247) );
  AOI22X1 U195 ( .A(n249), .B(n53), .C(n219), .D(N1271), .Y(n248) );
  NOR2X1 U196 ( .A(n217), .B(n378), .Y(n365) );
  AOI22X1 U197 ( .A(n214), .B(N1230), .C(n223), .D(N1148), .Y(n246) );
  INVX1 U198 ( .A(n211), .Y(n667) );
  AOI221XL U199 ( .A(n255), .B(n352), .C(n242), .D(n600), .E(n238), .Y(n126)
         );
  OAI22X1 U200 ( .A(n656), .B(n239), .C(n240), .D(n241), .Y(n238) );
  NAND4X1 U201 ( .A(n245), .B(n246), .C(n247), .D(n248), .Y(n242) );
  AOI22X1 U202 ( .A(n667), .B(N1312), .C(N1394), .D(n217), .Y(n245) );
  AOI22X1 U203 ( .A(n214), .B(n687), .C(n223), .D(n310), .Y(n305) );
  NAND2X1 U204 ( .A(n465), .B(n646), .Y(sub_398_S2_I7_aco_carry[4]) );
  NAND4X1 U205 ( .A(n340), .B(n341), .C(n342), .D(n343), .Y(n338) );
  AOI22X1 U206 ( .A(n667), .B(n347), .C(n217), .D(n705), .Y(n340) );
  AOI22X1 U207 ( .A(n250), .B(n344), .C(n252), .D(n345), .Y(n342) );
  AOI22X1 U208 ( .A(n214), .B(n691), .C(n346), .D(n223), .Y(n341) );
  INVX1 U209 ( .A(n479), .Y(n722) );
  INVX1 U210 ( .A(n442), .Y(n729) );
  OAI21X1 U211 ( .B(n522), .C(n477), .A(n224), .Y(N1139) );
  NOR21XL U212 ( .B(n594), .A(n595), .Y(n589) );
  OAI21X1 U213 ( .B(n699), .C(n420), .A(n588), .Y(n594) );
  NOR21XL U214 ( .B(n378), .A(n217), .Y(n252) );
  XOR2X1 U215 ( .A(n642), .B(n698), .Y(n643) );
  OA222X1 U216 ( .A(n480), .B(n481), .C(n482), .D(n687), .E(n380), .F(n689), 
        .Y(n363) );
  INVX1 U217 ( .A(N1230), .Y(n689) );
  AOI21X1 U218 ( .B(n486), .C(n691), .A(n487), .Y(n481) );
  AOI22X1 U219 ( .A(n483), .B(n484), .C(n485), .D(n691), .Y(n482) );
  NAND21X1 U220 ( .B(n420), .A(n698), .Y(n590) );
  OAI21X1 U221 ( .B(n489), .C(n490), .A(sub_398_S2_I3_aco_carry[4]), .Y(n281)
         );
  OAI32X1 U222 ( .A(n587), .B(n588), .C(n589), .D(n698), .E(n715), .Y(n255) );
  INVX1 U223 ( .A(n588), .Y(n715) );
  AOI21X1 U224 ( .B(n653), .C(n80), .A(n473), .Y(n466) );
  NOR41XL U225 ( .D(n369), .A(n371), .B(n372), .C(n370), .Y(n375) );
  NAND2X1 U226 ( .A(n537), .B(n476), .Y(n478) );
  NAND32X1 U227 ( .B(n270), .C(n298), .A(n297), .Y(n299) );
  OAI22X1 U228 ( .A(n656), .B(n271), .C(n692), .D(n241), .Y(n270) );
  OA2222XL U229 ( .A(n296), .B(n295), .C(n294), .D(n696), .E(n293), .F(n292), 
        .G(n291), .H(n290), .Y(n297) );
  AO22X1 U230 ( .A(n272), .B(n600), .C(n352), .D(n659), .Y(n298) );
  NOR3XL U231 ( .A(n728), .B(n393), .C(n224), .Y(n79) );
  INVX1 U232 ( .A(n477), .Y(n714) );
  AOI21X1 U233 ( .B(n442), .C(n53), .A(n714), .Y(n225) );
  OAI21X1 U234 ( .B(n465), .C(n646), .A(sub_398_S2_I7_aco_carry[4]), .Y(n284)
         );
  INVX1 U235 ( .A(n490), .Y(n695) );
  NOR2X1 U236 ( .A(n477), .B(n733), .Y(n595) );
  INVX1 U237 ( .A(n421), .Y(n699) );
  AOI211X1 U238 ( .C(n720), .D(n695), .A(n491), .B(n222), .Y(n82) );
  AOI21X1 U239 ( .B(n732), .C(n661), .A(n492), .Y(n491) );
  NAND2X1 U240 ( .A(n455), .B(n448), .Y(n447) );
  NAND2X1 U241 ( .A(n489), .B(n490), .Y(sub_398_S2_I3_aco_carry[4]) );
  INVX1 U242 ( .A(n492), .Y(n720) );
  INVX1 U243 ( .A(n283), .Y(n710) );
  INVX1 U244 ( .A(n280), .Y(n726) );
  INVX1 U245 ( .A(n537), .Y(n730) );
  OAI21X1 U246 ( .B(n567), .C(n573), .A(n477), .Y(n568) );
  NAND43X1 U247 ( .B(n371), .C(n124), .D(n372), .A(n369), .Y(n290) );
  INVX1 U248 ( .A(n370), .Y(n124) );
  NOR32XL U249 ( .B(n239), .C(n660), .A(n712), .Y(n555) );
  NAND32X1 U250 ( .B(n121), .C(n120), .A(n119), .Y(n294) );
  INVX1 U251 ( .A(n371), .Y(n121) );
  INVX1 U252 ( .A(n372), .Y(n119) );
  INVX1 U253 ( .A(n369), .Y(n120) );
  AOI221XL U254 ( .A(N1262), .B(n421), .C(n420), .D(N1262), .E(n220), .Y(n1)
         );
  NAND31X1 U255 ( .C(n732), .A(n568), .B(n73), .Y(n572) );
  OAI21X1 U256 ( .B(n564), .C(n380), .A(n63), .Y(n368) );
  MUX2X1 U257 ( .D0(n562), .D1(n563), .S(n227), .Y(n63) );
  AOI22AXL U258 ( .A(n644), .B(n570), .D(n644), .C(n571), .Y(n562) );
  AOI221XL U259 ( .A(n644), .B(n565), .C(n669), .D(n268), .E(n566), .Y(n563)
         );
  OAI221X1 U260 ( .A(n413), .B(n308), .C(n397), .D(n686), .E(n414), .Y(n379)
         );
  OAI31XL U261 ( .A(n415), .B(n674), .C(n408), .D(n308), .Y(n414) );
  INVX1 U262 ( .A(N1271), .Y(n686) );
  AOI22X1 U263 ( .A(n416), .B(n418), .C(n685), .D(n419), .Y(n413) );
  ENOX1 U264 ( .A(n694), .B(n241), .C(n336), .D(n337), .Y(n335) );
  OAI22X1 U265 ( .A(n292), .B(n648), .C(n650), .D(n268), .Y(n571) );
  NOR2X1 U266 ( .A(n420), .B(n1), .Y(n417) );
  NAND2X1 U267 ( .A(n369), .B(n372), .Y(n241) );
  INVX1 U268 ( .A(n448), .Y(n725) );
  NAND2X1 U269 ( .A(n573), .B(n568), .Y(n569) );
  OAI22X1 U270 ( .A(n503), .B(n498), .C(n502), .D(n267), .Y(n273) );
  AND2X1 U271 ( .A(n266), .B(n641), .Y(n267) );
  OAI21X1 U272 ( .B(n550), .C(n548), .A(n477), .Y(n543) );
  INVX1 U273 ( .A(n301), .Y(n693) );
  AOI221XL U274 ( .A(n525), .B(n526), .C(n527), .D(n669), .E(n528), .Y(n524)
         );
  AOI22X1 U275 ( .A(n694), .B(n533), .C(n534), .D(n526), .Y(n523) );
  AO21X1 U276 ( .B(n642), .C(n641), .A(n417), .Y(n308) );
  NAND21X1 U277 ( .B(n653), .A(n73), .Y(n635) );
  NOR21XL U278 ( .B(n572), .A(n62), .Y(n227) );
  NOR21XL U279 ( .B(n655), .A(n61), .Y(n62) );
  NOR21XL U280 ( .B(n653), .A(n716), .Y(n61) );
  OAI21X1 U281 ( .B(n511), .C(n380), .A(n123), .Y(n370) );
  MUX2X1 U282 ( .D0(n509), .D1(n510), .S(n230), .Y(n123) );
  AOI22AXL U283 ( .A(n334), .B(n512), .D(n334), .C(n513), .Y(n510) );
  AOI222XL U284 ( .A(n334), .B(n517), .C(n291), .D(n518), .E(n269), .F(n673), 
        .Y(n509) );
  AOI32X1 U285 ( .A(n718), .B(n514), .C(n515), .D(n516), .E(n645), .Y(n511) );
  INVX1 U286 ( .A(n516), .Y(n718) );
  NAND21X1 U287 ( .B(n336), .A(n368), .Y(n293) );
  OAI21X1 U288 ( .B(n717), .C(n397), .A(n118), .Y(n125) );
  INVX1 U289 ( .A(n244), .Y(n717) );
  MUX2X1 U290 ( .D0(n493), .D1(n494), .S(n27), .Y(n118) );
  AOI221XL U291 ( .A(n339), .B(n495), .C(n670), .D(n273), .E(n496), .Y(n494)
         );
  OAI211X1 U292 ( .C(n531), .D(n695), .A(n536), .B(n477), .Y(n532) );
  AO21X1 U293 ( .B(n732), .C(n661), .A(n531), .Y(n536) );
  AOI21X1 U294 ( .B(n497), .C(n503), .A(n53), .Y(n498) );
  AND4X1 U295 ( .A(n295), .B(n656), .C(n294), .D(n139), .Y(n140) );
  AOI21X1 U296 ( .B(n373), .C(n600), .A(n352), .Y(n139) );
  OR4X1 U297 ( .A(n249), .B(n219), .C(n250), .D(n252), .Y(n373) );
  AOI221XL U298 ( .A(n537), .B(n637), .C(n53), .D(n730), .E(n647), .Y(n531) );
  INVX1 U299 ( .A(n505), .Y(n641) );
  AND3X1 U300 ( .A(n241), .B(n293), .C(n138), .Y(n141) );
  OA21X1 U301 ( .B(n361), .C(n228), .A(n290), .Y(n138) );
  NOR4XL U302 ( .A(n223), .B(n667), .C(n214), .D(n217), .Y(n361) );
  NAND2X1 U303 ( .A(n519), .B(n728), .Y(n515) );
  INVX1 U304 ( .A(n231), .Y(n352) );
  INVX1 U305 ( .A(n271), .Y(n712) );
  OAI22X1 U306 ( .A(n648), .B(n692), .C(n650), .D(n527), .Y(n533) );
  INVX1 U307 ( .A(n514), .Y(n645) );
  OAI211X1 U308 ( .C(n538), .D(n700), .A(n539), .B(n540), .Y(n371) );
  AOI22X1 U309 ( .A(n675), .B(n285), .C(n696), .D(n682), .Y(n538) );
  AOI32X1 U310 ( .A(n660), .B(n542), .C(n696), .D(n670), .E(n285), .Y(n539) );
  AOI22X1 U311 ( .A(n541), .B(n311), .C(n657), .D(n668), .Y(n540) );
  INVX1 U312 ( .A(n416), .Y(n685) );
  AOI21X1 U313 ( .B(n648), .C(n650), .A(n691), .Y(n487) );
  INVX1 U314 ( .A(n173), .Y(n266) );
  NOR2X1 U315 ( .A(n647), .B(n637), .Y(n548) );
  INVX1 U316 ( .A(n556), .Y(n713) );
  INVX1 U317 ( .A(n285), .Y(n696) );
  MUX4X1 U318 ( .D0(n98), .D1(n96), .D2(n518), .D3(n673), .S0(n70), .S1(n69), 
        .Y(n77) );
  AO21X1 U319 ( .B(n85), .C(n83), .A(n714), .Y(n101) );
  AO21X1 U320 ( .B(n498), .C(n642), .A(n266), .Y(n339) );
  XOR2X1 U321 ( .A(n514), .B(n20), .Y(n334) );
  XOR2X1 U322 ( .A(n74), .B(n728), .Y(n314) );
  NAND21X1 U323 ( .B(n86), .A(n307), .Y(n136) );
  XOR2X1 U324 ( .A(n101), .B(n84), .Y(n86) );
  INVX1 U325 ( .A(n83), .Y(n84) );
  NAND21X1 U326 ( .B(n646), .A(n99), .Y(n85) );
  OAI21X1 U327 ( .B(n53), .C(n403), .A(n404), .Y(n398) );
  XOR2X1 U328 ( .A(n642), .B(n543), .Y(n700) );
  NAND21X1 U329 ( .B(n393), .A(n174), .Y(n74) );
  AO21X1 U330 ( .B(n392), .C(n97), .A(n669), .Y(n106) );
  AO21X1 U331 ( .B(n392), .C(n96), .A(n673), .Y(n107) );
  AND2X1 U332 ( .A(n636), .B(n733), .Y(n403) );
  AOI21BX1 U333 ( .C(n137), .B(n109), .A(n78), .Y(n25) );
  AOI21X1 U334 ( .B(n94), .C(n45), .A(n53), .Y(n26) );
  NAND2X1 U335 ( .A(n550), .B(n543), .Y(n547) );
  INVX1 U336 ( .A(n134), .Y(n94) );
  INVX1 U337 ( .A(n336), .Y(n656) );
  INVX1 U338 ( .A(n122), .Y(n230) );
  OAI211X1 U339 ( .C(n514), .D(n655), .A(n635), .B(n264), .Y(n122) );
  INVX1 U340 ( .A(n279), .Y(n683) );
  NOR2X1 U341 ( .A(n639), .B(n410), .Y(n394) );
  INVX1 U342 ( .A(n651), .Y(n669) );
  INVX1 U343 ( .A(n174), .Y(n67) );
  XNOR2XL U344 ( .A(n173), .B(n641), .Y(n27) );
  INVX1 U345 ( .A(n408), .Y(n680) );
  INVX1 U346 ( .A(n545), .Y(n678) );
  INVX1 U347 ( .A(n75), .Y(n263) );
  OAI211X1 U348 ( .C(n655), .D(n174), .A(n74), .B(n635), .Y(n75) );
  AO21X1 U349 ( .B(n94), .C(n668), .A(n93), .Y(n129) );
  MUX2X1 U350 ( .D0(n92), .D1(n91), .S(n24), .Y(n93) );
  MUX4X1 U351 ( .D0(n545), .D1(n676), .D2(n408), .D3(n674), .S0(n88), .S1(n87), 
        .Y(n92) );
  MUX4X1 U352 ( .D0(n682), .D1(n675), .D2(n89), .D3(n670), .S0(n88), .S1(n87), 
        .Y(n91) );
  NAND21X1 U353 ( .B(n642), .A(n52), .Y(n90) );
  INVX1 U354 ( .A(n648), .Y(n673) );
  INVX1 U355 ( .A(n650), .Y(n518) );
  INVX1 U356 ( .A(n317), .Y(n88) );
  AND2X1 U357 ( .A(n134), .B(n660), .Y(n89) );
  INVX1 U358 ( .A(n397), .Y(n668) );
  INVX1 U359 ( .A(n269), .Y(n291) );
  INVX1 U360 ( .A(n268), .Y(n292) );
  XOR2X1 U361 ( .A(n174), .B(n20), .Y(n439) );
  INVX1 U362 ( .A(n380), .Y(n109) );
  INVX1 U363 ( .A(r_semi), .Y(n596) );
  OAI221X1 U364 ( .A(n210), .B(n211), .C(n212), .D(n666), .E(n213), .Y(n200)
         );
  XOR2X1 U365 ( .A(sub_398_S2_aco_carry[5]), .B(n224), .Y(n212) );
  XNOR2XL U366 ( .A(sub_398_S2_I5_aco_carry[5]), .B(n225), .Y(n210) );
  INVX1 U367 ( .A(n223), .Y(n666) );
  AOI222XL U368 ( .A(n214), .B(n215), .C(n216), .D(n217), .E(n218), .F(n219), 
        .Y(n213) );
  XNOR2XL U369 ( .A(sub_398_S2_I4_aco_carry[5]), .B(n220), .Y(n218) );
  XNOR2XL U370 ( .A(sub_398_S2_I3_aco_carry[5]), .B(n222), .Y(n215) );
  XNOR2XL U371 ( .A(sub_398_S2_I7_aco_carry[5]), .B(n221), .Y(n216) );
  INVX1 U372 ( .A(n351), .Y(n374) );
  NAND32X1 U373 ( .B(n44), .C(n323), .A(n16), .Y(n326) );
  INVX1 U374 ( .A(n325), .Y(n331) );
  OAI221X1 U375 ( .A(n137), .B(n349), .C(n136), .D(n350), .E(n135), .Y(
        ps_ptr[4]) );
  OA222X1 U376 ( .A(n134), .B(n360), .C(n133), .D(n132), .E(n131), .F(n353), 
        .Y(n135) );
  AND2X1 U377 ( .A(n127), .B(n126), .Y(n131) );
  AO21X1 U378 ( .B(n256), .C(n55), .A(n286), .Y(n133) );
  INVX1 U379 ( .A(n439), .Y(n206) );
  NAND32X1 U380 ( .B(n335), .C(n179), .A(n355), .Y(n202) );
  AND2X1 U381 ( .A(n236), .B(n235), .Y(n261) );
  NOR21XL U382 ( .B(n258), .A(n257), .Y(n260) );
  OR2X1 U383 ( .A(n181), .B(n180), .Y(n184) );
  OR3XL U384 ( .A(n180), .B(n182), .C(n181), .Y(n254) );
  OAI221XL U385 ( .A(n172), .B(n353), .C(n171), .D(n357), .E(n170), .Y(
        ps_ptr[0]) );
  MUX2X1 U386 ( .D0(n141), .D1(n140), .S(n44), .Y(n172) );
  AOI31X1 U387 ( .A(n168), .B(n167), .C(n166), .D(n165), .Y(n171) );
  MUX2XL U388 ( .D0(n169), .D1(n360), .S(n44), .Y(n170) );
  INVX1 U389 ( .A(n289), .Y(n256) );
  INVXL U390 ( .A(wr_dacv[13]), .Y(n149) );
  INVX1 U391 ( .A(n243), .Y(n288) );
  NAND32XL U392 ( .B(n44), .C(wr_dacv[17]), .A(n144), .Y(n145) );
  NAND2X1 U393 ( .A(n28), .B(n348), .Y(n553) );
  OAI22XL U394 ( .A(n640), .B(ps_ptr[2]), .C(n17), .D(ps_ptr[3]), .Y(n28) );
  NAND21X1 U395 ( .B(n603), .A(n602), .Y(n671) );
  INVX1 U396 ( .A(n198), .Y(n603) );
  MUX2X1 U397 ( .D0(n601), .D1(busy), .S(n197), .Y(n602) );
  AOI32XL U398 ( .A(n200), .B(n600), .C(n599), .D(n598), .E(busy), .Y(n601) );
  OAI22X1 U399 ( .A(n52), .B(n508), .C(n504), .D(n501), .Y(n520) );
  INVXL U400 ( .A(ps_ptr[4]), .Y(n508) );
  INVX1 U401 ( .A(n553), .Y(n504) );
  OR2X1 U402 ( .A(n188), .B(n187), .Y(n237) );
  NAND32X1 U403 ( .B(wr_dacv[2]), .C(n162), .A(n167), .Y(n189) );
  AOI221XL U404 ( .A(n457), .B(n439), .C(n412), .D(n392), .E(n376), .Y(n472)
         );
  INVXL U405 ( .A(n350), .Y(n412) );
  OAI211XL U406 ( .C(n374), .D(n360), .A(n359), .B(n358), .Y(n376) );
  INVX1 U407 ( .A(n188), .Y(n302) );
  OAI31XL U408 ( .A(auto_start), .B(semi_start), .C(mxcyc_done), .D(n198), .Y(
        n197) );
  OAI21X1 U409 ( .B(n662), .C(n652), .A(n649), .Y(n29) );
  NAND2X1 U410 ( .A(n636), .B(n665), .Y(n652) );
  NAND21X1 U411 ( .B(n665), .A(n637), .Y(n649) );
  NAND21X1 U412 ( .B(n665), .A(n636), .Y(n329) );
  INVX1 U413 ( .A(n320), .Y(n324) );
  NAND21X1 U414 ( .B(n507), .A(n665), .Y(n320) );
  INVX1 U415 ( .A(n613), .Y(n616) );
  NAND21X1 U416 ( .B(n665), .A(n647), .Y(n613) );
  AND3X1 U417 ( .A(n614), .B(n662), .C(n328), .Y(N977) );
  OAI32X1 U418 ( .A(n329), .B(n662), .C(n326), .D(n649), .E(n325), .Y(N982) );
  AND2X1 U419 ( .A(n333), .B(n332), .Y(N972) );
  AND2X1 U420 ( .A(n333), .B(n328), .Y(N976) );
  INVX1 U421 ( .A(n48), .Y(cs_ptr[0]) );
  NOR32XL U422 ( .B(n365), .C(n364), .A(n379), .Y(n362) );
  NOR42XL U423 ( .C(n363), .D(n362), .A(n367), .B(n366), .Y(n249) );
  OA2222XL U424 ( .A(n230), .B(n290), .C(n27), .D(n295), .E(n229), .F(n228), 
        .G(n227), .H(n293), .Y(n236) );
  AND4X1 U425 ( .A(n305), .B(n306), .C(n304), .D(n226), .Y(n229) );
  AOI22X1 U426 ( .A(n667), .B(n711), .C(n217), .D(n703), .Y(n304) );
  AOI22X1 U427 ( .A(n250), .B(n727), .C(n252), .D(n309), .Y(n306) );
  OAI211X1 U428 ( .C(n440), .D(n438), .A(n441), .B(n225), .Y(n195) );
  OAI21X1 U429 ( .B(n655), .C(n732), .A(n721), .Y(n441) );
  INVX1 U430 ( .A(n507), .Y(n637) );
  INVX1 U431 ( .A(n55), .Y(n52) );
  INVX1 U432 ( .A(n55), .Y(cs_ptr[4]) );
  NAND2X1 U433 ( .A(n436), .B(n438), .Y(sub_398_S2_I5_aco_carry[4]) );
  AOI22AXL U434 ( .A(n219), .B(n308), .D(n640), .C(n249), .Y(n226) );
  NOR43XL U435 ( .B(n363), .C(n366), .D(n362), .A(n367), .Y(n223) );
  AO21X1 U436 ( .B(n642), .C(n49), .A(n640), .Y(n476) );
  AND3X1 U437 ( .A(n379), .B(n364), .C(n365), .Y(n219) );
  NAND21X1 U438 ( .B(n364), .A(n365), .Y(n211) );
  OAI21X1 U439 ( .B(n642), .C(n49), .A(n640), .Y(n442) );
  NAND2X1 U440 ( .A(n453), .B(n60), .Y(n73) );
  INVX1 U441 ( .A(cs_ptr[1]), .Y(n642) );
  INVX1 U442 ( .A(n719), .Y(n647) );
  INVX1 U443 ( .A(n48), .Y(n44) );
  AOI22X1 U444 ( .A(n249), .B(n735), .C(n219), .D(n685), .Y(n343) );
  OAI31XL U445 ( .A(n284), .B(N1394), .C(n471), .D(n651), .Y(n467) );
  AOI211X1 U446 ( .C(n722), .D(n474), .A(n475), .B(n221), .Y(n80) );
  AOI21X1 U447 ( .B(n478), .C(n732), .A(n479), .Y(n475) );
  NAND21X1 U448 ( .B(n638), .A(n52), .Y(n477) );
  NAND2X1 U449 ( .A(n456), .B(n453), .Y(n505) );
  OAI21X1 U450 ( .B(n455), .C(n449), .A(n57), .Y(n448) );
  OAI21X1 U451 ( .B(n436), .C(n438), .A(sub_398_S2_I5_aco_carry[4]), .Y(n283)
         );
  AOI211X1 U452 ( .C(n57), .D(n733), .A(n636), .B(n595), .Y(n588) );
  OAI21BBX1 U453 ( .A(n453), .B(n454), .C(n447), .Y(n280) );
  AOI21X1 U454 ( .B(n638), .C(n411), .A(n550), .Y(n421) );
  NOR3XL U455 ( .A(n377), .B(n368), .C(n336), .Y(n369) );
  OAI222XL U456 ( .A(n724), .B(n443), .C(n444), .D(n309), .E(n397), .F(n251), 
        .Y(n378) );
  INVX1 U457 ( .A(n309), .Y(n724) );
  AOI22AXL U458 ( .A(n345), .B(n450), .D(n345), .C(n451), .Y(n443) );
  AOI222XL U459 ( .A(n345), .B(n445), .C(n251), .D(n660), .E(n280), .F(n670), 
        .Y(n444) );
  NAND2X1 U460 ( .A(n733), .B(n46), .Y(n537) );
  INVX1 U461 ( .A(n411), .Y(n733) );
  OAI21X1 U462 ( .B(n476), .C(n57), .A(n477), .Y(n221) );
  INVX1 U463 ( .A(n319), .Y(n636) );
  NAND21X1 U464 ( .B(n52), .A(n638), .Y(n319) );
  INVX1 U465 ( .A(n55), .Y(n53) );
  OAI21X1 U466 ( .B(n406), .C(n726), .A(n405), .Y(n445) );
  OAI22X1 U467 ( .A(n469), .B(n688), .C(n470), .D(n281), .Y(n485) );
  OAI21X1 U468 ( .B(n464), .C(n688), .A(n463), .Y(n486) );
  NOR2X1 U469 ( .A(n411), .B(n638), .Y(n550) );
  OAI31XL U470 ( .A(n281), .B(N1230), .C(n471), .D(n651), .Y(n484) );
  NAND2X1 U471 ( .A(n41), .B(n505), .Y(n420) );
  NAND2X1 U472 ( .A(n390), .B(n391), .Y(sub_398_S2_aco_carry[4]) );
  NAND4X1 U473 ( .A(n274), .B(n275), .C(n276), .D(n277), .Y(n272) );
  AOI22X1 U474 ( .A(n667), .B(n283), .C(n217), .D(n284), .Y(n274) );
  AOI22X1 U475 ( .A(n250), .B(n279), .C(n252), .D(n280), .Y(n276) );
  AOI22X1 U476 ( .A(n214), .B(n281), .C(n223), .D(n282), .Y(n275) );
  OAI21BBX1 U477 ( .A(n463), .B(n464), .C(n705), .Y(n461) );
  OAI21BBX1 U478 ( .A(n572), .B(n438), .C(n569), .Y(n268) );
  AOI21X1 U479 ( .B(n559), .C(n557), .A(n714), .Y(n556) );
  OAI21X1 U480 ( .B(n239), .C(n397), .A(n59), .Y(n336) );
  MUX2X1 U481 ( .D0(n551), .D1(n552), .S(n234), .Y(n59) );
  AOI221XL U482 ( .A(n337), .B(n554), .C(n712), .D(n670), .E(n555), .Y(n552)
         );
  AOI222XL U483 ( .A(n337), .B(n560), .C(n712), .D(n674), .E(n271), .F(n408), 
        .Y(n551) );
  OA2222XL U484 ( .A(n234), .B(n656), .C(n301), .D(n241), .E(n233), .F(n294), 
        .G(n232), .H(n231), .Y(n235) );
  INVX1 U485 ( .A(n311), .Y(n233) );
  INVX1 U486 ( .A(n312), .Y(n232) );
  XNOR2XL U487 ( .A(n41), .B(n725), .Y(n345) );
  NAND21X1 U488 ( .B(n48), .A(n639), .Y(n522) );
  OAI221X1 U489 ( .A(n411), .B(n719), .C(n53), .D(n733), .E(n507), .Y(N1262)
         );
  INVX1 U490 ( .A(n506), .Y(n639) );
  INVX1 U491 ( .A(n391), .Y(n728) );
  OAI21X1 U492 ( .B(n522), .C(n638), .A(n57), .Y(n224) );
  OAI21X1 U493 ( .B(n556), .C(n557), .A(n558), .Y(n239) );
  XNOR2XL U494 ( .A(n556), .B(n559), .Y(n558) );
  OAI21X1 U495 ( .B(n730), .C(n55), .A(n477), .Y(n222) );
  INVX1 U496 ( .A(n474), .Y(n646) );
  AOI21X1 U497 ( .B(n638), .C(n733), .A(n57), .Y(n220) );
  NOR3XL U498 ( .A(n438), .B(n655), .C(n732), .Y(n573) );
  OAI22X1 U499 ( .A(n678), .B(n712), .C(n409), .D(n271), .Y(n560) );
  OAI22X1 U500 ( .A(n292), .B(n469), .C(n470), .D(n268), .Y(n565) );
  OAI21BBX1 U501 ( .A(n713), .B(n455), .C(n561), .Y(n271) );
  OAI21X1 U502 ( .B(n556), .C(n453), .A(n454), .Y(n561) );
  OAI22X1 U503 ( .A(n292), .B(n464), .C(n463), .D(n268), .Y(n570) );
  NOR2X1 U504 ( .A(n453), .B(n454), .Y(n455) );
  OAI21X1 U505 ( .B(n409), .C(n726), .A(n678), .Y(n450) );
  OAI31XL U506 ( .A(n278), .B(N1271), .C(n401), .D(n402), .Y(n418) );
  NOR3XL U507 ( .A(n268), .B(n471), .C(n658), .Y(n566) );
  INVX1 U508 ( .A(n564), .Y(n658) );
  NAND2X1 U509 ( .A(n446), .B(n447), .Y(n251) );
  XNOR2XL U510 ( .A(n448), .B(n449), .Y(n446) );
  OAI21BBX1 U511 ( .A(n391), .B(n264), .C(n515), .Y(n269) );
  NAND21X1 U512 ( .B(n52), .A(n521), .Y(n514) );
  OAI21X1 U513 ( .B(n393), .C(n391), .A(n516), .Y(n521) );
  NAND21X1 U514 ( .B(n209), .A(n208), .Y(n312) );
  NAND21X1 U515 ( .B(n505), .A(n207), .Y(n208) );
  INVX1 U516 ( .A(n590), .Y(n209) );
  NAND21X1 U517 ( .B(n589), .A(n41), .Y(n207) );
  NAND21X1 U518 ( .B(n498), .A(n41), .Y(n173) );
  XNOR2XL U519 ( .A(n41), .B(n1), .Y(n416) );
  NAND32X1 U520 ( .B(n368), .C(n336), .A(n377), .Y(n231) );
  OAI211X1 U521 ( .C(n52), .D(n522), .A(n507), .B(n719), .Y(n516) );
  NOR32XL U522 ( .B(n692), .C(n240), .A(n471), .Y(n528) );
  XNOR2XL U523 ( .A(n41), .B(n556), .Y(n337) );
  NAND21X1 U524 ( .B(n453), .A(n454), .Y(n557) );
  OAI21X1 U525 ( .B(n390), .C(n391), .A(sub_398_S2_aco_carry[4]), .Y(n282) );
  NAND2X1 U526 ( .A(n549), .B(n547), .Y(n285) );
  OAI21X1 U527 ( .B(n701), .C(n411), .A(n638), .Y(n549) );
  INVX1 U528 ( .A(n543), .Y(n701) );
  OAI211X1 U529 ( .C(n52), .D(n506), .A(n507), .B(n719), .Y(n497) );
  OAI222XL U530 ( .A(n680), .B(n285), .C(n696), .D(n452), .E(n544), .F(n700), 
        .Y(n541) );
  AOI22X1 U531 ( .A(n676), .B(n285), .C(n696), .D(n545), .Y(n544) );
  INVX1 U532 ( .A(n265), .Y(n502) );
  OAI22X1 U533 ( .A(n469), .B(n692), .C(n470), .D(n527), .Y(n525) );
  OAI22X1 U534 ( .A(n405), .B(n712), .C(n406), .D(n271), .Y(n554) );
  OAI21X1 U535 ( .B(n464), .C(n291), .A(n463), .Y(n517) );
  OAI21X1 U536 ( .B(n296), .C(n406), .A(n405), .Y(n495) );
  OAI22X1 U537 ( .A(n464), .B(n692), .C(n463), .D(n527), .Y(n534) );
  OAI22AX1 U538 ( .D(n511), .C(n471), .A(n651), .B(n291), .Y(n513) );
  OAI21X1 U539 ( .B(n469), .C(n291), .A(n470), .Y(n512) );
  AOI22AXL U540 ( .A(n339), .B(n499), .D(n339), .C(n500), .Y(n493) );
  OAI21X1 U541 ( .B(n296), .C(n409), .A(n678), .Y(n499) );
  OAI22X1 U542 ( .A(n680), .B(n273), .C(n296), .D(n452), .Y(n500) );
  AOI21X1 U543 ( .B(n678), .C(n409), .A(n416), .Y(n415) );
  NOR3XL U544 ( .A(n273), .B(n401), .C(n244), .Y(n496) );
  NAND3X1 U545 ( .A(n41), .B(n502), .C(n641), .Y(n503) );
  NAND21X1 U546 ( .B(n714), .A(n66), .Y(n174) );
  NAND21X1 U547 ( .B(n26), .A(n65), .Y(n66) );
  NAND21X1 U548 ( .B(n393), .A(n391), .Y(n65) );
  MUX2X1 U549 ( .D0(n143), .D1(n114), .S(n44), .Y(n651) );
  MUX4X1 U550 ( .D0(n72), .D1(n97), .D2(n71), .D3(n669), .S0(n70), .S1(n69), 
        .Y(n76) );
  INVX1 U551 ( .A(n470), .Y(n72) );
  AND2X1 U552 ( .A(n137), .B(n68), .Y(n71) );
  INVX1 U553 ( .A(n471), .Y(n68) );
  NAND21X1 U554 ( .B(n507), .A(n639), .Y(n134) );
  OAI21X1 U555 ( .B(n410), .C(n638), .A(n404), .Y(n279) );
  OR2X1 U556 ( .A(n647), .B(n30), .Y(n83) );
  MUX2IX1 U557 ( .D0(n55), .D1(n507), .S(n731), .Y(n30) );
  AO21X1 U558 ( .B(n110), .C(n109), .A(n108), .Y(n130) );
  MUX4X1 U559 ( .D0(n107), .D1(n106), .D2(n105), .D3(n104), .S0(n22), .S1(n103), .Y(n108) );
  OA21X1 U560 ( .B(n474), .C(n102), .A(n307), .Y(n103) );
  AO21X1 U561 ( .B(n392), .C(n98), .A(n518), .Y(n105) );
  OAI222XL U562 ( .A(n394), .B(n395), .C(n396), .D(n727), .E(n397), .F(n398), 
        .Y(n367) );
  AOI211X1 U563 ( .C(n344), .D(n407), .A(n674), .B(n408), .Y(n395) );
  AOI22AXL U564 ( .A(n344), .B(n399), .D(n344), .C(n400), .Y(n396) );
  OAI21X1 U565 ( .B(n683), .C(n409), .A(n678), .Y(n407) );
  NOR2X1 U566 ( .A(n411), .B(n403), .Y(n410) );
  INVX1 U567 ( .A(n48), .Y(n45) );
  OAI22X1 U568 ( .A(n470), .B(n205), .C(n471), .D(n110), .Y(n104) );
  OAI22X1 U569 ( .A(n405), .B(n279), .C(n683), .D(n406), .Y(n399) );
  OAI21X1 U570 ( .B(n401), .C(n684), .A(n402), .Y(n400) );
  INVX1 U571 ( .A(n401), .Y(n660) );
  INVX1 U572 ( .A(n402), .Y(n670) );
  NAND2X1 U573 ( .A(n410), .B(n638), .Y(n404) );
  NAND2X1 U574 ( .A(n469), .B(n470), .Y(n468) );
  NAND2X1 U575 ( .A(n680), .B(n452), .Y(n451) );
  MUX2X1 U576 ( .D0(n144), .D1(n146), .S(cs_ptr[0]), .Y(n380) );
  MUX2X1 U577 ( .D0(n146), .D1(n144), .S(cs_ptr[0]), .Y(n397) );
  MUX2X1 U578 ( .D0(n148), .D1(n152), .S(n44), .Y(n648) );
  MUX2X1 U579 ( .D0(n663), .D1(n664), .S(cs_ptr[0]), .Y(n650) );
  OAI21X1 U580 ( .B(n49), .C(n663), .A(n664), .Y(n408) );
  OAI21X1 U581 ( .B(n49), .C(n681), .A(n679), .Y(n545) );
  OR2X1 U582 ( .A(n639), .B(n31), .Y(n311) );
  MUX2IX1 U583 ( .D0(n640), .D1(n411), .S(n543), .Y(n31) );
  NOR2X1 U584 ( .A(n41), .B(n403), .Y(n344) );
  INVX1 U585 ( .A(n452), .Y(n674) );
  INVX1 U586 ( .A(n409), .Y(n676) );
  NAND2X1 U587 ( .A(n405), .B(n406), .Y(n419) );
  XNOR2XL U588 ( .A(n265), .B(n32), .Y(n317) );
  NAND2X1 U589 ( .A(n175), .B(n641), .Y(n32) );
  OA21X1 U590 ( .B(n53), .C(n735), .A(n90), .Y(n87) );
  INVX1 U591 ( .A(n406), .Y(n675) );
  INVX1 U592 ( .A(n469), .Y(n97) );
  INVX1 U593 ( .A(n405), .Y(n682) );
  INVX1 U594 ( .A(n463), .Y(n98) );
  INVX1 U595 ( .A(n464), .Y(n96) );
  NOR41XL U596 ( .D(n634), .A(n33), .B(n34), .C(n35), .Y(sh_hold) );
  NAND4X1 U597 ( .A(n626), .B(n625), .C(n624), .D(n623), .Y(n33) );
  NAND4X1 U598 ( .A(n630), .B(n629), .C(n628), .D(n627), .Y(n34) );
  NAND4X1 U599 ( .A(n15), .B(n633), .C(n632), .D(n631), .Y(n35) );
  AO21X1 U600 ( .B(n16), .C(n57), .A(n175), .Y(n351) );
  NAND32X1 U601 ( .B(n16), .C(n323), .A(n46), .Y(n325) );
  INVX1 U602 ( .A(n654), .Y(n323) );
  INVX1 U603 ( .A(n321), .Y(n330) );
  NAND32X1 U604 ( .B(n48), .C(n16), .A(n654), .Y(n321) );
  INVX1 U605 ( .A(n322), .Y(n614) );
  NAND32X1 U606 ( .B(n48), .C(n323), .A(n16), .Y(n322) );
  AND2XL U607 ( .A(n9), .B(pos_dacis[9]), .Y(N959) );
  AND2XL U608 ( .A(n21), .B(pos_dacis[6]), .Y(N956) );
  AND2XL U609 ( .A(n9), .B(pos_dacis[2]), .Y(N952) );
  AND2XL U610 ( .A(n21), .B(pos_dacis[15]), .Y(N965) );
  AND2XL U611 ( .A(n9), .B(pos_dacis[7]), .Y(N957) );
  AND2XL U612 ( .A(n9), .B(pos_dacis[14]), .Y(N964) );
  AND2XL U613 ( .A(n9), .B(pos_dacis[4]), .Y(N954) );
  AND2XL U614 ( .A(n21), .B(pos_dacis[11]), .Y(N961) );
  AND2XL U615 ( .A(n21), .B(pos_dacis[12]), .Y(N962) );
  AND2XL U616 ( .A(n9), .B(pos_dacis[0]), .Y(N950) );
  AND2XL U617 ( .A(n9), .B(pos_dacis[10]), .Y(N960) );
  AND2XL U618 ( .A(n9), .B(pos_dacis[3]), .Y(N953) );
  AND2XL U619 ( .A(n21), .B(pos_dacis[5]), .Y(N955) );
  AND2XL U620 ( .A(n21), .B(pos_dacis[17]), .Y(N967) );
  AND2XL U621 ( .A(n21), .B(pos_dacis[8]), .Y(N958) );
  AND2XL U622 ( .A(n21), .B(pos_dacis[1]), .Y(N951) );
  NAND32X1 U623 ( .B(wr_dacv[0]), .C(n113), .A(n112), .Y(n357) );
  INVX1 U624 ( .A(r_dac_en[0]), .Y(n112) );
  OR2XL U625 ( .A(wr_dacv[14]), .B(r_dac_en[14]), .Y(n180) );
  GEN2XL U626 ( .D(n194), .E(n191), .C(n237), .B(n190), .A(n189), .Y(n356) );
  INVX1 U627 ( .A(n253), .Y(n190) );
  GEN2XL U628 ( .D(n256), .E(n735), .C(n184), .B(n183), .A(n11), .Y(n186) );
  INVXL U629 ( .A(n357), .Y(n199) );
  GEN2XL U630 ( .D(n256), .E(n18), .C(n254), .B(n288), .A(n253), .Y(n257) );
  NAND43X1 U631 ( .B(r_dac_en[13]), .C(r_dac_en[12]), .D(wr_dacv[13]), .A(n153), .Y(n182) );
  NAND43X1 U632 ( .B(r_dac_en[17]), .C(r_dac_en[16]), .D(wr_dacv[17]), .A(n147), .Y(n289) );
  OR2XL U633 ( .A(wr_dacv[15]), .B(r_dac_en[15]), .Y(n181) );
  GEN2XL U634 ( .D(n159), .E(n158), .C(n157), .B(n302), .A(n187), .Y(n160) );
  AND2X1 U635 ( .A(n143), .B(n142), .Y(n159) );
  AND2X1 U636 ( .A(n154), .B(n185), .Y(n155) );
  NAND5XL U637 ( .A(n117), .B(n185), .C(n116), .D(n194), .E(n154), .Y(n243) );
  INVX1 U638 ( .A(r_dac_en[11]), .Y(n116) );
  OAI31XL U639 ( .A(n164), .B(wr_dacv[4]), .C(r_dac_en[4]), .D(n163), .Y(n166)
         );
  INVX1 U640 ( .A(n162), .Y(n163) );
  AND3X1 U641 ( .A(n663), .B(n161), .C(n160), .Y(n164) );
  INVX1 U642 ( .A(wr_dacv[5]), .Y(n161) );
  NAND32X1 U643 ( .B(r_dac_en[9]), .C(n157), .A(n142), .Y(n115) );
  INVX1 U644 ( .A(cs_mux_5_), .Y(busy) );
  OAI21X1 U645 ( .B(r_loop), .C(n597), .A(n596), .Y(n598) );
  OA21XL U646 ( .B(n55), .C(ps_ptr[4]), .A(n591), .Y(n597) );
  GEN2XL U647 ( .D(ps_ptr[2]), .E(n640), .C(n574), .B(n553), .A(n520), .Y(n591) );
  INVX1 U648 ( .A(n348), .Y(n574) );
  NAND21X1 U649 ( .B(pos_dacis[10]), .A(n2), .Y(app_dacis[10]) );
  NAND43X1 U650 ( .B(wr_dacv[4]), .C(wr_dacv[5]), .D(r_dac_en[4]), .A(n663), 
        .Y(n253) );
  OR2X1 U651 ( .A(wr_dacv[7]), .B(r_dac_en[7]), .Y(n188) );
  OR2X1 U652 ( .A(wr_dacv[6]), .B(r_dac_en[6]), .Y(n187) );
  NAND21X1 U653 ( .B(pos_dacis[11]), .A(n4), .Y(app_dacis[11]) );
  NAND21X1 U654 ( .B(pos_dacis[6]), .A(n43), .Y(app_dacis[6]) );
  NAND21XL U655 ( .B(pos_dacis[5]), .A(n54), .Y(app_dacis[5]) );
  NAND21X1 U656 ( .B(pos_dacis[7]), .A(n39), .Y(app_dacis[7]) );
  NAND21XL U657 ( .B(pos_dacis[4]), .A(n618), .Y(app_dacis[4]) );
  NAND21X1 U658 ( .B(pos_dacis[16]), .A(n622), .Y(app_dacis[16]) );
  NAND21XL U659 ( .B(pos_dacis[3]), .A(n6), .Y(app_dacis[3]) );
  NAND21XL U660 ( .B(pos_dacis[2]), .A(n7), .Y(app_dacis[2]) );
  NAND21XL U661 ( .B(pos_dacis[1]), .A(n3), .Y(app_dacis[1]) );
  NAND21X1 U662 ( .B(pos_dacis[14]), .A(n51), .Y(app_dacis[14]) );
  NAND21X1 U663 ( .B(pos_dacis[12]), .A(n620), .Y(app_dacis[12]) );
  NAND21XL U664 ( .B(pos_dacis[0]), .A(n5), .Y(app_dacis[0]) );
  NAND21X1 U665 ( .B(pos_dacis[17]), .A(n37), .Y(app_dacis[17]) );
  NAND21X1 U666 ( .B(pos_dacis[15]), .A(n56), .Y(app_dacis[15]) );
  NAND21X1 U667 ( .B(pos_dacis[8]), .A(n47), .Y(app_dacis[8]) );
  NAND21X1 U668 ( .B(pos_dacis[9]), .A(n619), .Y(app_dacis[9]) );
  OR2X1 U669 ( .A(wr_dacv[3]), .B(r_dac_en[3]), .Y(n162) );
  NAND43X1 U670 ( .B(wr_dacv[1]), .C(n357), .D(n10), .A(n356), .Y(n358) );
  INVX1 U671 ( .A(neg_dacis[9]), .Y(n619) );
  INVX1 U672 ( .A(neg_dacis[12]), .Y(n620) );
  INVX1 U673 ( .A(neg_dacis[4]), .Y(n618) );
  INVX1 U674 ( .A(neg_dacis[16]), .Y(n622) );
  NAND21X1 U675 ( .B(pos_dacis[13]), .A(n621), .Y(app_dacis[13]) );
  INVX1 U676 ( .A(neg_dacis[13]), .Y(n621) );
  NAND21X1 U677 ( .B(n10), .A(n196), .Y(n165) );
  OAI21X1 U678 ( .B(stop), .C(srstz), .A(n197), .Y(N994) );
  NOR21XL U679 ( .B(srstz), .A(stop), .Y(n198) );
  INVX1 U680 ( .A(n736), .Y(n48) );
  NAND21X1 U681 ( .B(n52), .A(cs_ptr[3]), .Y(n507) );
  BUFX3 U682 ( .A(n735), .Y(cs_ptr[1]) );
  OAI22X1 U683 ( .A(n422), .B(n423), .C(n49), .D(n424), .Y(n364) );
  OAI21BBX1 U684 ( .A(r_dac_en[17]), .B(N1312), .C(n432), .Y(n423) );
  GEN2XL U685 ( .D(n709), .E(n672), .C(n434), .B(n428), .A(n736), .Y(n422) );
  OAI21BBX1 U686 ( .A(r_dac_en[16]), .B(N1312), .C(n425), .Y(n424) );
  OAI32X1 U687 ( .A(n426), .B(r_dac_en[8]), .C(n710), .D(n283), .E(n427), .Y(
        n425) );
  ENOX1 U688 ( .A(n428), .B(n431), .C(n347), .D(r_dac_en[10]), .Y(n426) );
  OAI22X1 U689 ( .A(n428), .B(n429), .C(n430), .D(n711), .Y(n427) );
  AOI21X1 U690 ( .B(r_dac_en[14]), .C(n347), .A(r_dac_en[12]), .Y(n431) );
  AOI32X1 U691 ( .A(r_dac_en[0]), .B(n707), .C(n709), .D(r_dac_en[2]), .E(n347), .Y(n430) );
  INVX1 U692 ( .A(n734), .Y(n55) );
  NAND21X1 U693 ( .B(n41), .A(cs_ptr[2]), .Y(n453) );
  NAND21X1 U694 ( .B(cs_ptr[3]), .A(n52), .Y(n719) );
  NAND21X1 U695 ( .B(cs_ptr[2]), .A(n41), .Y(n456) );
  XNOR2XL U696 ( .A(cs_ptr[3]), .B(n729), .Y(n438) );
  BUFX3 U697 ( .A(n735), .Y(n41) );
  INVX1 U698 ( .A(cs_ptr[2]), .Y(n640) );
  NAND6XL U699 ( .A(n620), .B(n618), .C(n622), .D(n619), .E(n611), .F(n610), 
        .Y(n617) );
  NOR5X1 U700 ( .A(neg_dacis[13]), .B(n825), .C(n824), .D(n823), .E(n822), .Y(
        n611) );
  NOR6XL U701 ( .A(n609), .B(n608), .C(n607), .D(n606), .E(n605), .F(n604), 
        .Y(n610) );
  NAND5XL U702 ( .A(n39), .B(n37), .C(srstz), .D(n2), .E(n3), .Y(n609) );
  INVX1 U703 ( .A(n736), .Y(n49) );
  INVX1 U704 ( .A(n437), .Y(n672) );
  AOI31X1 U705 ( .A(n710), .B(n707), .C(n10), .D(r_dac_en[9]), .Y(n437) );
  NAND21X1 U706 ( .B(cs_ptr[2]), .A(n642), .Y(n411) );
  XOR2X1 U707 ( .A(n476), .B(cs_ptr[3]), .Y(n474) );
  AO2222XL U708 ( .A(n577), .B(r_dac_en[12]), .C(n582), .D(r_dac_en[4]), .E(
        n580), .F(r_dac_en[14]), .G(n583), .H(r_dac_en[6]), .Y(n578) );
  AO2222XL U709 ( .A(n577), .B(r_dac_en[13]), .C(n582), .D(r_dac_en[5]), .E(
        n580), .F(r_dac_en[15]), .G(n583), .H(r_dac_en[7]), .Y(n584) );
  INVX1 U710 ( .A(cs_ptr[3]), .Y(n638) );
  OAI21X1 U711 ( .B(n697), .C(n397), .A(n64), .Y(n377) );
  MUX2X1 U712 ( .D0(n576), .D1(n575), .S(cs_ptr[0]), .Y(n64) );
  AOI221XL U713 ( .A(n577), .B(r_dac_en[9]), .C(n584), .D(n312), .E(n585), .Y(
        n575) );
  AOI221XL U714 ( .A(n577), .B(r_dac_en[8]), .C(n578), .D(n312), .E(n579), .Y(
        n576) );
  AOI221XL U715 ( .A(n640), .B(n647), .C(n55), .D(cs_ptr[2]), .E(n637), .Y(
        n449) );
  AOI22X1 U716 ( .A(n249), .B(n19), .C(n219), .D(n278), .Y(n277) );
  OAI211X1 U717 ( .C(n380), .D(n706), .A(n381), .B(n382), .Y(n366) );
  OAI31XL U718 ( .A(n387), .B(r_dac_en[10]), .C(n388), .D(n44), .Y(n381) );
  OAI31XL U719 ( .A(n383), .B(r_dac_en[11]), .C(n384), .D(n48), .Y(n382) );
  OR3XL U720 ( .A(r_dac_en[14]), .B(r_dac_en[8]), .C(r_dac_en[12]), .Y(n387)
         );
  INVX1 U721 ( .A(n736), .Y(n46) );
  OAI21BBX1 U722 ( .A(r_dac_en[10]), .B(n580), .C(n581), .Y(n579) );
  AOI32X1 U723 ( .A(n697), .B(r_dac_en[0]), .C(n582), .D(n583), .E(r_dac_en[2]), .Y(n581) );
  OAI21BBX1 U724 ( .A(r_dac_en[11]), .B(n580), .C(n586), .Y(n585) );
  AOI32X1 U725 ( .A(n697), .B(n10), .C(n582), .D(n583), .E(r_dac_en[3]), .Y(
        n586) );
  AOI21X1 U726 ( .B(r_dac_en[6]), .C(n347), .A(r_dac_en[4]), .Y(n429) );
  AOI31X1 U727 ( .A(n663), .B(n681), .C(n385), .D(n282), .Y(n384) );
  AOI31X1 U728 ( .A(n10), .B(n706), .C(n386), .D(r_dac_en[3]), .Y(n385) );
  INVX1 U729 ( .A(n734), .Y(n57) );
  XOR2X1 U730 ( .A(n522), .B(n19), .Y(n391) );
  NAND21X1 U731 ( .B(n642), .A(cs_ptr[2]), .Y(n506) );
  XNOR2XL U732 ( .A(cs_ptr[3]), .B(cs_ptr[2]), .Y(n454) );
  GEN2XL U733 ( .D(n677), .E(n681), .C(n709), .B(n433), .A(n428), .Y(n432) );
  INVX1 U734 ( .A(r_dac_en[15]), .Y(n677) );
  OAI21X1 U735 ( .B(r_dac_en[5]), .C(r_dac_en[13]), .A(n709), .Y(n433) );
  AOI21BBXL U736 ( .B(r_dac_en[11]), .C(r_dac_en[3]), .A(n709), .Y(n434) );
  OAI221X1 U737 ( .A(n640), .B(n507), .C(n18), .D(n57), .E(n719), .Y(n559) );
  AOI31X1 U738 ( .A(n664), .B(n679), .C(n389), .D(n282), .Y(n388) );
  AOI31X1 U739 ( .A(r_dac_en[0]), .B(n706), .C(n386), .D(r_dac_en[2]), .Y(n389) );
  XOR2X1 U740 ( .A(n506), .B(n19), .Y(n265) );
  OAI221X1 U741 ( .A(n18), .B(n448), .C(n725), .D(n453), .E(n456), .Y(n309) );
  AOI22X1 U742 ( .A(n45), .B(r_dac_en[0]), .C(n46), .D(n10), .Y(n471) );
  AOI22X1 U743 ( .A(n45), .B(r_dac_en[2]), .C(n46), .D(r_dac_en[3]), .Y(n470)
         );
  AOI21X1 U744 ( .B(n45), .C(r_dac_en[11]), .A(r_dac_en[10]), .Y(n406) );
  AOI22X1 U745 ( .A(n45), .B(r_dac_en[3]), .C(n46), .D(r_dac_en[2]), .Y(n405)
         );
  AOI22X1 U746 ( .A(n45), .B(r_dac_en[10]), .C(n46), .D(r_dac_en[11]), .Y(n469) );
  AOI21X1 U747 ( .B(n45), .C(r_dac_en[15]), .A(r_dac_en[14]), .Y(n409) );
  AOI22X1 U748 ( .A(n45), .B(r_dac_en[6]), .C(n49), .D(r_dac_en[7]), .Y(n463)
         );
  AOI22X1 U749 ( .A(n736), .B(r_dac_en[14]), .C(n49), .D(r_dac_en[15]), .Y(
        n464) );
  AOI21X1 U750 ( .B(n44), .C(r_dac_en[13]), .A(r_dac_en[12]), .Y(n452) );
  AOI22X1 U751 ( .A(n45), .B(n10), .C(n46), .D(r_dac_en[0]), .Y(n401) );
  AOI22X1 U752 ( .A(n736), .B(r_dac_en[9]), .C(n49), .D(r_dac_en[8]), .Y(n402)
         );
  INVX1 U753 ( .A(n58), .Y(n234) );
  OAI221X1 U754 ( .A(n556), .B(n453), .C(n713), .D(n18), .E(n456), .Y(n58) );
  INVX1 U755 ( .A(r_dac_en[5]), .Y(n663) );
  INVX1 U756 ( .A(r_dac_en[7]), .Y(n681) );
  INVX1 U757 ( .A(r_dac_en[6]), .Y(n679) );
  INVX1 U758 ( .A(r_dac_en[12]), .Y(n152) );
  INVX1 U759 ( .A(r_dac_en[9]), .Y(n143) );
  INVX1 U760 ( .A(r_dac_en[13]), .Y(n148) );
  INVX1 U761 ( .A(r_dac_en[8]), .Y(n114) );
  INVX1 U762 ( .A(r_dac_en[4]), .Y(n664) );
  INVX1 U763 ( .A(r_dac_en[17]), .Y(n144) );
  INVX1 U764 ( .A(r_dac_en[16]), .Y(n146) );
  OR3XL U765 ( .A(r_dac_en[13]), .B(r_dac_en[9]), .C(r_dac_en[15]), .Y(n383)
         );
  NOR2X1 U766 ( .A(pos_dacis[9]), .B(pos_dacis[8]), .Y(n193) );
  INVX1 U767 ( .A(pos_dacis[6]), .Y(n629) );
  INVX1 U768 ( .A(pos_dacis[14]), .Y(n631) );
  INVX1 U769 ( .A(pos_dacis[15]), .Y(n632) );
  INVX1 U770 ( .A(pos_dacis[7]), .Y(n630) );
  INVXL U771 ( .A(pos_dacis[4]), .Y(n623) );
  INVX1 U772 ( .A(pos_dacis[11]), .Y(n628) );
  INVX1 U773 ( .A(pos_dacis[12]), .Y(n633) );
  INVX1 U774 ( .A(pos_dacis[10]), .Y(n627) );
  INVXL U775 ( .A(pos_dacis[5]), .Y(n624) );
  INVXL U776 ( .A(pos_dacis[3]), .Y(n626) );
  NOR2X1 U777 ( .A(pos_dacis[17]), .B(pos_dacis[16]), .Y(n192) );
  INVXL U778 ( .A(pos_dacis[1]), .Y(n625) );
  INVX1 U779 ( .A(r_dac_en[10]), .Y(n185) );
  INVX1 U780 ( .A(r_dac_en[2]), .Y(n167) );
  AND2X1 U781 ( .A(sampl_begn), .B(srstz), .Y(n654) );
  INVX1 U782 ( .A(n327), .Y(n333) );
  NAND21X1 U783 ( .B(r_comp_swtch), .A(n615), .Y(n327) );
  INVX1 U784 ( .A(r_comp_swtch), .Y(n662) );
  NAND32XL U785 ( .B(sampl_begn), .C(n13), .A(n198), .Y(N971) );
  OAI31XL U786 ( .A(n156), .B(n11), .C(wr_dacv[11]), .D(n155), .Y(n158) );
  INVXL U787 ( .A(wr_dacv[11]), .Y(n117) );
  NAND43X1 U788 ( .B(wr_dacv[11]), .C(wr_dacv[10]), .D(n186), .A(n185), .Y(
        n191) );
  INVXL U789 ( .A(wr_dacv[9]), .Y(n142) );
  NAND21XL U790 ( .B(wr_dacv[8]), .A(n114), .Y(n157) );
  MAJ3X1 U791 ( .A(n472), .B(n735), .C(n460), .Y(n501) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_LOW_shmux_00000005_00000012_00000012 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLNXL latch ( .CKN(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dac2sar_a0 ( r_dac_t, r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, 
        auto_sar, busy, stop, sync_i, ps_sample, sampl_begn, sampl_done, 
        sh_rst, dacyc_done, sacyc_done, dac_v, rpt_v, clk, srstz, test_si2, 
        test_si1, test_so1, test_se );
  input [1:0] r_dac_t;
  output [9:0] dac_v;
  output [9:0] rpt_v;
  input r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, auto_sar, busy, stop,
         sync_i, ps_sample, clk, srstz, test_si2, test_si1, test_se;
  output sampl_begn, sampl_done, sh_rst, dacyc_done, sacyc_done, test_so1;
  wire   N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N71, N72, N73, N74, N75, N79, updlo, updup, upd1v, r_lt_up_8_,
         r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, r_lt_up_3_,
         r_lt_up_2_, r_lt_up_1_, r_lt_up_0_, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102,
         net10243, net10249, n136, n45, n46, n47, n48, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n64, n66, n67, n71, n72, n73, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n1, n3, n7, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n68,
         n69, n70, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3;
  wire   [3:0] sarcyc;
  wire   [6:0] dacnt;
  wire   [9:0] r_lt_lo;
  wire   [9:0] r_avg00;
  wire   [9:0] r_avgup;
  wire   [9:0] r_dacvo;

  INVX1 U55 ( .A(n48), .Y(n46) );
  INVX1 U56 ( .A(n48), .Y(n47) );
  INVX1 U57 ( .A(srstz), .Y(n48) );
  INVX1 U58 ( .A(n48), .Y(n45) );
  glreg_WIDTH10_2 u0_dac1v ( .clk(clk), .arstz(n47), .we(upd1v), .wdat(r_dacvo), .rdat({dac_v[9:1], n136}), .test_si(sarcyc[3]), .test_se(test_se) );
  glreg_WIDTH10_1 u0_lt_lo ( .clk(clk), .arstz(n46), .we(updlo), .wdat({n40, 
        n39, n38, n37, n36, n35, n31, n33, n32, n34}), .rdat(r_lt_lo), 
        .test_si(dac_v[9]), .test_se(test_se) );
  glreg_WIDTH10_0 u0_lt_up ( .clk(clk), .arstz(n45), .we(updup), .wdat(r_avgup), .rdat({test_so1, r_lt_up_8_, r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, 
        r_lt_up_3_, r_lt_up_2_, r_lt_up_1_, r_lt_up_0_}), .test_si(r_lt_lo[9]), 
        .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 clk_gate_dacnt_reg ( .CLK(clk), .EN(N54), 
        .ENCLK(net10243), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 clk_gate_sarcyc_reg ( .CLK(clk), .EN(N71), 
        .ENCLK(net10249), .TE(test_se) );
  dac2sar_a0_DW01_add_0 add_312 ( .A({1'b0, n9, n11, n13, n15, n17, n19, n21, 
        n23, n25, n27}), .B({1'b0, n8, n10, n12, n14, n16, n18, n20, n22, n24, 
        n26}), .CI(1'b0), .SUM({N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, SYNOPSYS_UNCONNECTED_1}), .CO() );
  dac2sar_a0_DW01_add_1 add_310 ( .A({1'b0, n40, n39, n38, n37, n36, n35, n31, 
        n33, n32, n34}), .B({1'b0, r_avgup}), .CI(1'b0), .SUM({N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, SYNOPSYS_UNCONNECTED_2}), .CO() );
  dac2sar_a0_DW01_add_2 add_305 ( .A({1'b0, r_lt_lo}), .B({1'b0, test_so1, 
        r_lt_up_8_, r_lt_up_7_, r_lt_up_6_, r_lt_up_5_, r_lt_up_4_, r_lt_up_3_, 
        r_lt_up_2_, r_lt_up_1_, r_lt_up_0_}), .CI(1'b0), .SUM({r_avg00, 
        SYNOPSYS_UNCONNECTED_3}), .CO() );
  dac2sar_a0_DW01_inc_0 add_285 ( .A(dacnt), .SUM({N53, N52, N51, N50, N49, 
        N48, N47}) );
  SDFFQX1 dacnt_reg_1_ ( .D(N56), .SIN(dacnt[0]), .SMC(test_se), .C(net10243), 
        .Q(dacnt[1]) );
  SDFFQX1 dacnt_reg_0_ ( .D(N55), .SIN(test_si2), .SMC(test_se), .C(net10243), 
        .Q(dacnt[0]) );
  SDFFQX1 sarcyc_reg_3_ ( .D(N75), .SIN(sarcyc[2]), .SMC(test_se), .C(net10249), .Q(sarcyc[3]) );
  SDFFQX1 sarcyc_reg_1_ ( .D(N73), .SIN(sarcyc[0]), .SMC(test_se), .C(net10249), .Q(sarcyc[1]) );
  SDFFQX1 dacnt_reg_2_ ( .D(N57), .SIN(dacnt[1]), .SMC(test_se), .C(net10243), 
        .Q(dacnt[2]) );
  SDFFQX1 sarcyc_reg_2_ ( .D(N74), .SIN(sarcyc[1]), .SMC(test_se), .C(net10249), .Q(sarcyc[2]) );
  SDFFQX1 dacnt_reg_3_ ( .D(N58), .SIN(dacnt[2]), .SMC(test_se), .C(net10243), 
        .Q(dacnt[3]) );
  SDFFQX1 sarcyc_reg_0_ ( .D(N72), .SIN(dacnt[6]), .SMC(test_se), .C(net10249), 
        .Q(sarcyc[0]) );
  SDFFQX1 dacnt_reg_5_ ( .D(N60), .SIN(dacnt[4]), .SMC(test_se), .C(net10243), 
        .Q(dacnt[5]) );
  SDFFQX1 dacnt_reg_6_ ( .D(N61), .SIN(dacnt[5]), .SMC(test_se), .C(net10243), 
        .Q(dacnt[6]) );
  SDFFQX1 dacnt_reg_4_ ( .D(N59), .SIN(dacnt[3]), .SMC(test_se), .C(net10243), 
        .Q(dacnt[4]) );
  SDFFNQX1 sh_rst_n_reg ( .D(N79), .SIN(test_si1), .SMC(test_se), .XC(clk), 
        .Q(sh_rst) );
  INVX1 U6 ( .A(dacnt[0]), .Y(n42) );
  INVXL U7 ( .A(n136), .Y(n1) );
  INVXL U8 ( .A(n1), .Y(dac_v[0]) );
  INVXL U9 ( .A(n1), .Y(n3) );
  MUX2IX2 U10 ( .D0(n29), .D1(n30), .S(ps_sample), .Y(n43) );
  BUFX3 U11 ( .A(semi_nxt), .Y(n7) );
  BUFX3 U12 ( .A(sar_ini), .Y(n28) );
  INVX1 U13 ( .A(sar_ini), .Y(n51) );
  INVX1 U14 ( .A(n77), .Y(n30) );
  INVX1 U15 ( .A(n78), .Y(n29) );
  INVX1 U16 ( .A(n96), .Y(n129) );
  NAND2X1 U17 ( .A(n100), .B(n96), .Y(N71) );
  INVX1 U18 ( .A(n113), .Y(n132) );
  INVX1 U19 ( .A(n106), .Y(n62) );
  NAND2X1 U20 ( .A(n81), .B(n51), .Y(r_avgup[1]) );
  MUX2X1 U21 ( .D0(N91), .D1(r_avg00[9]), .S(semi_nxt), .Y(r_dacvo[9]) );
  MUX2X1 U22 ( .D0(N90), .D1(r_avg00[8]), .S(semi_nxt), .Y(r_dacvo[8]) );
  NAND2X1 U23 ( .A(n80), .B(n51), .Y(r_avgup[0]) );
  NOR2XL U24 ( .A(sar_ini), .B(n90), .Y(n31) );
  NAND2XL U25 ( .A(n82), .B(n51), .Y(r_avgup[2]) );
  NAND2XL U26 ( .A(n83), .B(n51), .Y(r_avgup[3]) );
  NAND2XL U27 ( .A(n120), .B(n51), .Y(r_avgup[4]) );
  MUX2X1 U28 ( .D0(N89), .D1(r_avg00[7]), .S(n7), .Y(r_dacvo[7]) );
  MUX2X1 U29 ( .D0(N88), .D1(r_avg00[6]), .S(n7), .Y(r_dacvo[6]) );
  MUX2X1 U30 ( .D0(N87), .D1(r_avg00[5]), .S(semi_nxt), .Y(r_dacvo[5]) );
  NOR2XL U31 ( .A(sar_ini), .B(n92), .Y(n32) );
  NOR2XL U32 ( .A(sar_ini), .B(n91), .Y(n33) );
  NOR2XL U33 ( .A(sar_ini), .B(n93), .Y(n34) );
  NOR2XL U34 ( .A(sar_ini), .B(n89), .Y(n35) );
  NOR2XL U35 ( .A(sar_ini), .B(n88), .Y(n36) );
  NAND2XL U36 ( .A(n121), .B(n51), .Y(r_avgup[5]) );
  MUX2X1 U37 ( .D0(N85), .D1(r_avg00[3]), .S(semi_nxt), .Y(r_dacvo[3]) );
  MUX2X1 U38 ( .D0(N86), .D1(r_avg00[4]), .S(semi_nxt), .Y(r_dacvo[4]) );
  NOR2XL U39 ( .A(sar_ini), .B(n87), .Y(n37) );
  NOR2XL U40 ( .A(sar_ini), .B(n86), .Y(n38) );
  NAND2XL U41 ( .A(n122), .B(n51), .Y(r_avgup[6]) );
  NAND2XL U42 ( .A(n123), .B(n51), .Y(r_avgup[7]) );
  MUX2X1 U43 ( .D0(N84), .D1(r_avg00[2]), .S(semi_nxt), .Y(r_dacvo[2]) );
  NOR2XL U44 ( .A(n28), .B(n85), .Y(n39) );
  NOR2XL U45 ( .A(n28), .B(n84), .Y(n40) );
  NAND2XL U46 ( .A(n124), .B(n51), .Y(r_avgup[8]) );
  MUX2X1 U47 ( .D0(N82), .D1(r_avg00[0]), .S(semi_nxt), .Y(r_dacvo[0]) );
  MUX2X1 U48 ( .D0(N83), .D1(r_avg00[1]), .S(semi_nxt), .Y(r_dacvo[1]) );
  NAND2XL U49 ( .A(n125), .B(n51), .Y(r_avgup[9]) );
  AO21XL U50 ( .B(sar_nxt), .C(sync_i), .A(n28), .Y(updlo) );
  OR3XL U51 ( .A(sar_nxt), .B(n28), .C(semi_nxt), .Y(upd1v) );
  NOR21XL U52 ( .B(n102), .A(sacyc_done), .Y(n100) );
  NAND3X1 U53 ( .A(n100), .B(dacyc_done), .C(auto_sar), .Y(n96) );
  XNOR2XL U54 ( .A(n135), .B(r_sar10), .Y(n104) );
  NAND2X1 U59 ( .A(n129), .B(n97), .Y(n98) );
  NOR2X1 U60 ( .A(n99), .B(n98), .Y(N73) );
  NOR21XL U61 ( .B(n116), .A(n115), .Y(n113) );
  NOR21XL U62 ( .B(n79), .A(n65), .Y(n68) );
  NAND3X1 U63 ( .A(busy), .B(n101), .C(n102), .Y(n106) );
  NOR21XL U64 ( .B(N52), .A(n106), .Y(N60) );
  NOR21XL U65 ( .B(N51), .A(n106), .Y(N59) );
  NOR21XL U66 ( .B(N49), .A(n106), .Y(N57) );
  NOR21XL U67 ( .B(N50), .A(n106), .Y(N58) );
  AND2X1 U68 ( .A(N48), .B(n62), .Y(N56) );
  NAND3X1 U69 ( .A(n106), .B(n101), .C(n102), .Y(N54) );
  XOR2X1 U70 ( .A(n133), .B(n116), .Y(n65) );
  INVX1 U71 ( .A(n117), .Y(n131) );
  INVX1 U72 ( .A(n110), .Y(n134) );
  NOR2X1 U73 ( .A(n101), .B(n64), .Y(sacyc_done) );
  INVX1 U74 ( .A(n101), .Y(dacyc_done) );
  INVX1 U75 ( .A(n89), .Y(n19) );
  INVX1 U76 ( .A(n120), .Y(n18) );
  INVX1 U77 ( .A(n88), .Y(n17) );
  INVX1 U78 ( .A(n121), .Y(n16) );
  INVX1 U79 ( .A(n87), .Y(n15) );
  INVX1 U80 ( .A(n122), .Y(n14) );
  INVX1 U81 ( .A(n91), .Y(n23) );
  INVX1 U82 ( .A(n82), .Y(n22) );
  INVX1 U83 ( .A(n123), .Y(n12) );
  INVX1 U84 ( .A(n86), .Y(n13) );
  INVX1 U85 ( .A(n90), .Y(n21) );
  INVX1 U86 ( .A(n83), .Y(n20) );
  INVX1 U87 ( .A(n124), .Y(n10) );
  INVX1 U88 ( .A(n85), .Y(n11) );
  INVX1 U89 ( .A(n92), .Y(n25) );
  INVX1 U90 ( .A(n81), .Y(n24) );
  INVX1 U91 ( .A(n84), .Y(n9) );
  INVX1 U92 ( .A(n125), .Y(n8) );
  INVX1 U93 ( .A(r_avg00[4]), .Y(n57) );
  INVX1 U94 ( .A(r_avg00[0]), .Y(n61) );
  INVX1 U95 ( .A(r_avg00[5]), .Y(n56) );
  INVX1 U96 ( .A(r_avg00[1]), .Y(n60) );
  INVX1 U97 ( .A(r_avg00[6]), .Y(n55) );
  INVX1 U98 ( .A(r_avg00[2]), .Y(n59) );
  INVX1 U99 ( .A(r_avg00[7]), .Y(n54) );
  INVX1 U100 ( .A(r_avg00[3]), .Y(n58) );
  INVX1 U101 ( .A(r_avg00[8]), .Y(n53) );
  INVX1 U102 ( .A(n80), .Y(n26) );
  INVX1 U103 ( .A(n93), .Y(n27) );
  INVX1 U104 ( .A(r_avg00[9]), .Y(n52) );
  INVX1 U105 ( .A(n50), .Y(n49) );
  INVX1 U106 ( .A(n50), .Y(n44) );
  NOR32X4 U107 ( .B(n42), .C(dacnt[1]), .A(n43), .Y(sampl_done) );
  AO21XL U108 ( .B(sar_nxt), .C(n50), .A(n28), .Y(updup) );
  ENOX1 U109 ( .A(dac_v[0]), .B(n83), .C(N96), .D(n3), .Y(rpt_v[3]) );
  ENOX1 U110 ( .A(n3), .B(n120), .C(N97), .D(dac_v[0]), .Y(rpt_v[4]) );
  ENOX1 U111 ( .A(dac_v[0]), .B(n123), .C(N100), .D(n3), .Y(rpt_v[7]) );
  NOR21XL U112 ( .B(n47), .A(stop), .Y(n102) );
  NAND42X1 U113 ( .C(n64), .D(n76), .A(n75), .B(n74), .Y(n77) );
  XOR2X1 U114 ( .A(n70), .B(r_dacyc), .Y(n75) );
  XOR2X1 U115 ( .A(n130), .B(dacnt[2]), .Y(n74) );
  NAND31X1 U116 ( .C(dacnt[6]), .A(n126), .B(n66), .Y(n76) );
  GEN2XL U117 ( .D(n129), .E(n135), .C(n128), .B(sarcyc[3]), .A(n95), .Y(N75)
         );
  NOR4XL U118 ( .A(sarcyc[3]), .B(n135), .C(n96), .D(n97), .Y(n95) );
  INVX1 U119 ( .A(n98), .Y(n128) );
  NAND41X1 U120 ( .D(n63), .A(n105), .B(n103), .C(n104), .Y(n64) );
  INVX1 U121 ( .A(sarcyc[0]), .Y(n63) );
  XOR2X1 U122 ( .A(sarcyc[1]), .B(r_sar10), .Y(n105) );
  XNOR2XL U123 ( .A(sarcyc[3]), .B(r_sar10), .Y(n103) );
  OAI32X1 U124 ( .A(n97), .B(sarcyc[2]), .C(n96), .D(n135), .E(n98), .Y(N74)
         );
  NOR2X1 U125 ( .A(sarcyc[0]), .B(n96), .Y(N72) );
  ENOX1 U126 ( .A(n136), .B(n124), .C(N101), .D(dac_v[0]), .Y(rpt_v[8]) );
  ENOX1 U127 ( .A(n3), .B(n121), .C(N98), .D(n3), .Y(rpt_v[5]) );
  ENOX1 U128 ( .A(n3), .B(n125), .C(n3), .D(N102), .Y(rpt_v[9]) );
  NAND42X1 U129 ( .C(n72), .D(n71), .A(n69), .B(n68), .Y(n78) );
  XNOR2XL U130 ( .A(n131), .B(dacnt[2]), .Y(n72) );
  XOR2X1 U131 ( .A(dacnt[5]), .B(n113), .Y(n69) );
  XNOR2XL U132 ( .A(n132), .B(dacnt[6]), .Y(n71) );
  ENOX1 U133 ( .A(dac_v[0]), .B(n82), .C(N95), .D(n3), .Y(rpt_v[2]) );
  AOI21BBXL U134 ( .B(r_dac_t[0]), .C(n115), .A(n117), .Y(n116) );
  NOR21XL U135 ( .B(N53), .A(n106), .Y(N61) );
  NOR2X1 U136 ( .A(r_dac_t[1]), .B(n115), .Y(n117) );
  NOR2X1 U137 ( .A(r_dac_t[0]), .B(r_dac_t[1]), .Y(n115) );
  XOR2X1 U138 ( .A(n70), .B(n114), .Y(n79) );
  OAI21X1 U139 ( .B(r_dac_t[0]), .C(n115), .A(n132), .Y(n114) );
  AND2X1 U140 ( .A(N47), .B(n62), .Y(N55) );
  ENOX1 U141 ( .A(n3), .B(n81), .C(N94), .D(dac_v[0]), .Y(rpt_v[1]) );
  ENOX1 U142 ( .A(n136), .B(n80), .C(N93), .D(n136), .Y(rpt_v[0]) );
  ENOX1 U143 ( .A(dac_v[0]), .B(n122), .C(N99), .D(n3), .Y(rpt_v[6]) );
  XNOR2XL U144 ( .A(n130), .B(dacnt[3]), .Y(n66) );
  INVX1 U145 ( .A(dacnt[4]), .Y(n70) );
  INVX1 U146 ( .A(r_dacyc), .Y(n130) );
  INVX1 U147 ( .A(sarcyc[2]), .Y(n135) );
  INVX1 U148 ( .A(dacnt[3]), .Y(n133) );
  NAND32X1 U149 ( .B(sarcyc[2]), .C(sarcyc[3]), .A(n99), .Y(n110) );
  NAND42X1 U150 ( .C(dacnt[1]), .D(dacnt[2]), .A(n134), .B(n94), .Y(n73) );
  NOR4XL U151 ( .A(dacnt[6]), .B(dacnt[5]), .C(dacnt[4]), .D(dacnt[3]), .Y(n94) );
  NOR2X1 U152 ( .A(sarcyc[1]), .B(sarcyc[0]), .Y(n99) );
  NOR31X1 U153 ( .C(busy), .A(dacnt[0]), .B(n73), .Y(N79) );
  INVX1 U154 ( .A(dacnt[5]), .Y(n126) );
  NAND4X1 U155 ( .A(dacnt[0]), .B(dacnt[1]), .C(n107), .D(n108), .Y(n101) );
  XNOR2XL U156 ( .A(dacnt[2]), .B(n119), .Y(n107) );
  AOI221XL U157 ( .A(dacnt[6]), .B(dacnt[5]), .C(n109), .D(n110), .E(n111), 
        .Y(n108) );
  AOI22X1 U158 ( .A(n134), .B(n131), .C(n110), .D(n130), .Y(n119) );
  AOI31X1 U159 ( .A(n67), .B(n79), .C(n112), .D(n110), .Y(n111) );
  INVX1 U160 ( .A(n65), .Y(n67) );
  AOI22X1 U161 ( .A(n113), .B(n127), .C(n132), .D(n126), .Y(n112) );
  INVX1 U162 ( .A(dacnt[6]), .Y(n127) );
  OAI221X1 U163 ( .A(n70), .B(n133), .C(dacnt[4]), .D(n130), .E(n118), .Y(n109) );
  AOI211X1 U164 ( .C(n133), .D(n130), .A(dacnt[6]), .B(dacnt[5]), .Y(n118) );
  MUX2BXL U165 ( .D0(n59), .D1(r_lt_up_2_), .S(n49), .Y(n82) );
  MUX2BXL U166 ( .D0(n55), .D1(r_lt_up_6_), .S(n49), .Y(n122) );
  MUX2BXL U167 ( .D0(n58), .D1(r_lt_up_3_), .S(n49), .Y(n83) );
  MUX2BXL U168 ( .D0(n57), .D1(r_lt_up_4_), .S(n49), .Y(n120) );
  MUX2BXL U169 ( .D0(n56), .D1(r_lt_up_5_), .S(n49), .Y(n121) );
  MUX2BXL U170 ( .D0(n54), .D1(r_lt_up_7_), .S(n49), .Y(n123) );
  MUX2BXL U171 ( .D0(n53), .D1(r_lt_up_8_), .S(n49), .Y(n124) );
  MUX2BXL U172 ( .D0(n61), .D1(r_lt_up_0_), .S(n49), .Y(n80) );
  MUX2BXL U173 ( .D0(n60), .D1(r_lt_up_1_), .S(n49), .Y(n81) );
  MUX2AXL U174 ( .D0(r_lt_lo[4]), .D1(n57), .S(n44), .Y(n89) );
  MUX2AXL U175 ( .D0(r_lt_lo[0]), .D1(n61), .S(n49), .Y(n93) );
  MUX2AXL U176 ( .D0(r_lt_lo[5]), .D1(n56), .S(n44), .Y(n88) );
  MUX2AXL U177 ( .D0(r_lt_lo[1]), .D1(n60), .S(n44), .Y(n92) );
  MUX2AXL U178 ( .D0(r_lt_lo[6]), .D1(n55), .S(n44), .Y(n87) );
  MUX2AXL U179 ( .D0(r_lt_lo[2]), .D1(n59), .S(n44), .Y(n91) );
  MUX2AXL U180 ( .D0(r_lt_lo[7]), .D1(n54), .S(n44), .Y(n86) );
  MUX2AXL U181 ( .D0(r_lt_lo[3]), .D1(n58), .S(n44), .Y(n90) );
  MUX2AXL U182 ( .D0(r_lt_lo[8]), .D1(n53), .S(n44), .Y(n85) );
  MUX2BXL U183 ( .D0(n52), .D1(test_so1), .S(n44), .Y(n125) );
  MUX2AXL U184 ( .D0(r_lt_lo[9]), .D1(n52), .S(n44), .Y(n84) );
  INVX1 U185 ( .A(sync_i), .Y(n50) );
  NOR21XL U186 ( .B(dacnt[0]), .A(n73), .Y(sampl_begn) );
  NAND2X1 U187 ( .A(sarcyc[0]), .B(sarcyc[1]), .Y(n97) );
endmodule


module dac2sar_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module dac2sar_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module dac2sar_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module dac2sar_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10266;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10266), .TE(test_se) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10266), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10284;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10284), .TE(test_se) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10284), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10302;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10302), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[1]) );
  SDFFRQXL mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[9]) );
  SDFFRQXL mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[8]) );
  SDFFRQXL mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[7]) );
  SDFFRQXL mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10302), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_00000012 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [17:0] wdat;
  output [17:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10320, n1, n2, n3;

  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(arstz), .Y(n3) );
  SNPS_CLOCK_GATE_HIGH_glreg_00000012 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10320), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10320), .XR(n2), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10320), .XR(n2), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10320), .XR(n2), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10320), .XR(n2), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10320), .XR(n2), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_10_ ( .D(wdat[10]), .SIN(rdat[9]), .SMC(test_se), .C(
        net10320), .XR(n1), .Q(rdat[10]) );
  SDFFRQX1 mem_reg_16_ ( .D(wdat[16]), .SIN(rdat[15]), .SMC(test_se), .C(
        net10320), .XR(n1), .Q(rdat[16]) );
  SDFFRQX1 mem_reg_17_ ( .D(wdat[17]), .SIN(rdat[16]), .SMC(test_se), .C(
        net10320), .XR(n1), .Q(rdat[17]) );
  SDFFRQX1 mem_reg_9_ ( .D(wdat[9]), .SIN(rdat[8]), .SMC(test_se), .C(net10320), .XR(n1), .Q(rdat[9]) );
  SDFFRQX1 mem_reg_12_ ( .D(wdat[12]), .SIN(rdat[11]), .SMC(test_se), .C(
        net10320), .XR(n1), .Q(rdat[12]) );
  SDFFRQX1 mem_reg_8_ ( .D(wdat[8]), .SIN(rdat[7]), .SMC(test_se), .C(net10320), .XR(n1), .Q(rdat[8]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10320), .XR(n2), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10320), .XR(n2), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10320), .XR(n2), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_11_ ( .D(wdat[11]), .SIN(rdat[10]), .SMC(test_se), .C(
        net10320), .XR(n1), .Q(rdat[11]) );
  SDFFRQX1 mem_reg_14_ ( .D(wdat[14]), .SIN(rdat[13]), .SMC(test_se), .C(
        net10320), .XR(n1), .Q(rdat[14]) );
  SDFFRQX1 mem_reg_15_ ( .D(wdat[15]), .SIN(rdat[14]), .SMC(test_se), .C(
        net10320), .XR(n1), .Q(rdat[15]) );
  SDFFRQX1 mem_reg_13_ ( .D(wdat[13]), .SIN(rdat[12]), .SMC(test_se), .C(
        net10320), .XR(n1), .Q(rdat[13]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_00000012 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( i_cc, i_cc_49, i_sqlch, r_sqlch, 
        r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, 
        r_fiforst, r_unlock, r_first, r_last, r_set_cpmsgid, r_rdy, r_wdat, 
        r_rdat, r_txnumk, r_txendk, r_txshrt, r_auto_discard, r_txauto, 
        r_rxords_ena, r_spec, r_dat_spec, r_auto_gdcrc, r_rxdb_opt, r_pshords, 
        r_dat_portrole, r_dat_datarole, r_discard, pid_goidle, pid_gobusy, 
        pff_ack, pff_rdat, pff_rxpart, prx_rcvinf, pff_obsd, pff_ptr, 
        pff_empty, pff_full, ptx_ack, ptx_cc, ptx_oe, prx_setsta, prx_rst, 
        prl_c0set, prl_cany0, prl_cany0r, prl_cany0w, prl_discard, 
        prl_GCTxDone, prl_cany0adr, prl_cpmsgid, prx_fifowdat, ptx_fsm, 
        prl_fsm, prx_fsm, prx_adpn, dbgpo, clk, srstz, test_si, test_so, 
        test_se );
  input [1:0] r_sqlch;
  input [7:0] r_wdat;
  input [7:0] r_rdat;
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [6:0] r_rxords_ena;
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [1:0] r_auto_gdcrc;
  input [1:0] r_rxdb_opt;
  output [1:0] pff_ack;
  output [7:0] pff_rdat;
  output [15:0] pff_rxpart;
  output [4:0] prx_rcvinf;
  output [5:0] pff_ptr;
  output [6:0] prx_setsta;
  output [1:0] prx_rst;
  output [7:0] prl_cany0adr;
  output [2:0] prl_cpmsgid;
  output [7:0] prx_fifowdat;
  output [2:0] ptx_fsm;
  output [3:0] prl_fsm;
  output [3:0] prx_fsm;
  output [5:0] prx_adpn;
  output [31:0] dbgpo;
  input i_cc, i_cc_49, i_sqlch, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4,
         r_fifopsh, r_fifopop, r_fiforst, r_unlock, r_first, r_last,
         r_set_cpmsgid, r_rdy, r_txendk, r_txshrt, r_auto_discard, r_pshords,
         r_dat_portrole, r_dat_datarole, r_discard, clk, srstz, test_si,
         test_se;
  output pid_goidle, pid_gobusy, pff_obsd, pff_empty, pff_full, ptx_ack,
         ptx_cc, ptx_oe, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_discard, prl_GCTxDone, test_so;
  wire   n116, rx_pshords, auto_rx_gdcrc, prx_trans, prx_fiforst, pcc_rxgood,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd, x_trans, ptx_goidle,
         c0_txendk, mux_one, ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4,
         crcstart, crcshfi4, crcshfo4, prl_idle, lockena, fifosrstz,
         fifopop_pff, fifopsh_pff, pff_txreq, pff_one, obsd, prl_last,
         prl_txreq, fifopop_prl, fifopsh_prl, prx_gdmsgrcvd, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, d_sqlch, net10338, n114, n117, n68, n69,
         n70, n71, n55, n56, n57, n58, n64, n65, n66, n67, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n5, n7, n9, n11, n12, n15, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n59, n60, n61, n62, n63, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4;
  wire   [1:0] prx_cccnt;
  wire   [3:0] prx_crcsidat;
  wire   [4:0] c0_txnumk;
  wire   [6:0] c0_txauto;
  wire   [7:0] mux_rdat;
  wire   [3:0] ptx_crcsidat;
  wire   [3:0] crc32_3_0;
  wire   [3:0] crcsidat;
  wire   [55:0] pff_dat_7_1;
  wire   [47:16] pff_c0dat;
  wire   [7:0] prl_rdat;
  wire   [4:0] prl_txauto;
  wire   [1:0] d_cc;
  wire   [8:0] cclow_cnt;

  phyrx_a0 u0_phyrx ( .i_cc(i_cc), .ptx_txact(ptx_oe), .r_adprx_en(r_adprx_en), 
        .r_adp2nd(r_adp2nd), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), 
        .r_rxdb_opt(r_rxdb_opt), .r_ords_ena(r_rxords_ena), .r_pshords(
        rx_pshords), .r_rgdcrc(auto_rx_gdcrc), .prx_cccnt(prx_cccnt), 
        .prx_rst(prx_rst), .prx_setsta({prx_setsta[6:1], 
        SYNOPSYS_UNCONNECTED_1}), .prx_idle(), .prx_d_cc(dbgpo[17]), .prx_bmc(
        dbgpo[18]), .prx_trans(prx_trans), .prx_fiforst(prx_fiforst), 
        .prx_fifopsh(n117), .prx_fifowdat(prx_fifowdat), .pff_txreq(n15), 
        .pid_gobusy(pid_gobusy), .pid_goidle(pid_goidle), .pid_ccidle(
        prx_rcvinf[4]), .pcc_rxgood(pcc_rxgood), .prx_crcstart(prx_crcstart), 
        .prx_crcshfi4(prx_crcshfi4), .prx_crcsidat(prx_crcsidat), .prx_rxcode(
        dbgpo[28:24]), .prx_adpn(prx_adpn), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_eoprcvd(prx_eoprcvd), .prx_fsm(prx_fsm), .clk(clk), .srstz(n41), 
        .test_si(n70), .test_so(n69), .test_se(test_se) );
  phyidd_a0 u0_phyidd ( .i_trans(x_trans), .i_goidle(ptx_goidle), .o_ccidle(
        prx_rcvinf[4]), .o_goidle(pid_goidle), .o_gobusy(pid_gobusy), .clk(clk), .srstz(n41), .test_si(pff_ptr[5]), .test_so(n70), .test_se(test_se) );
  phytx_a0 u0_phytx ( .r_txnumk(c0_txnumk), .r_txendk(c0_txendk), .r_txshrt(
        r_txshrt), .r_txauto(c0_txauto), .prx_cccnt(prx_cccnt), .ptx_txact(
        n114), .ptx_cc(ptx_cc), .ptx_goidle(ptx_goidle), .ptx_fifopop(n116), 
        .ptx_pspyld(), .i_rdat(mux_rdat), .i_txreq(n15), .i_one(mux_one), 
        .ptx_crcstart(ptx_crcstart), .ptx_crcshfi4(ptx_crcshfi4), 
        .ptx_crcshfo4(ptx_crcshfo4), .ptx_crcsidat(ptx_crcsidat), .ptx_fsm(
        ptx_fsm), .pcc_crc30(crc32_3_0), .clk(clk), .srstz(n41), .test_si(n69), 
        .test_se(test_se) );
  phycrc_a0 u0_phycrc ( .crc32_3_0(crc32_3_0), .rx_good(pcc_rxgood), 
        .i_shfidat(crcsidat), .i_start(crcstart), .i_shfi4(crcshfi4), 
        .i_shfo4(crcshfo4), .clk(clk), .test_si(d_cc[1]), .test_so(n71), 
        .test_se(test_se) );
  phyff_DEPTH_NUM34_DEPTH_NBT6 u0_phyff ( .r_psh(r_fifopsh), .r_pop(r_fifopop), 
        .prx_psh(fifopsh_pff), .ptx_pop(fifopop_pff), .r_last(r_last), 
        .r_unlock(r_unlock), .i_lockena(lockena), .r_fiforst(r_fiforst), 
        .i_ccidle(prx_rcvinf[4]), .r_wdat(r_wdat), .prx_wdat(prx_fifowdat), 
        .txreq(pff_txreq), .ffack(pff_ack), .rdat0(pff_rdat), .full(pff_full), 
        .empty(pff_empty), .one(pff_one), .half(), .obsd(obsd), .dat_7_1(
        pff_dat_7_1), .ptr(pff_ptr), .fifowdat(dbgpo[7:0]), .fifopsh(dbgpo[16]), .clk(clk), .srstz(fifosrstz), .test_si(n71), .test_se(test_se) );
  updprl_a0 u0_updprl ( .r_spec(r_spec), .r_dat_spec(r_dat_spec), 
        .r_auto_txgdcrc(r_auto_gdcrc[0]), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_auto_discard(r_auto_discard), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_dat_cpmsgid(r_wdat[2:0]), .r_rdat(
        r_rdat), .r_rdy(r_rdy), .pid_ccidle(prx_rcvinf[4]), .r_discard(
        r_discard), .ptx_ack(ptx_goidle), .ptx_txact(n7), .ptx_fifopop(
        fifopop_prl), .prx_fifopsh(fifopsh_prl), .prx_gdmsgrcvd(prx_gdmsgrcvd), 
        .prx_eoprcvd(prx_eoprcvd), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_fifowdat(prx_fifowdat), .pff_c0dat({pff_c0dat, pff_rxpart}), 
        .prl_rdat(prl_rdat), .prl_txauto({SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, prl_txauto[4], SYNOPSYS_UNCONNECTED_4, 
        prl_txauto[2:0]}), .prl_last(prl_last), .prl_txreq(prl_txreq), 
        .prl_c0set(prl_c0set), .prl_cany0(prl_cany0), .prl_cany0r(prl_cany0r), 
        .prl_cany0w(prl_cany0w), .prl_idle(prl_idle), .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_fsm(prl_fsm), .prl_cpmsgid(prl_cpmsgid), 
        .prl_cany0adr(prl_cany0adr), .clk(clk), .srstz(n40), .test_si(n68), 
        .test_so(test_so), .test_se(test_se) );
  dbnc_WIDTH3 u0_sqlch_db ( .o_dbc(d_sqlch), .o_chg(), .i_org(i_sqlch), .clk(
        clk), .rstz(n40), .test_si(ptx_cc), .test_so(n68), .test_se(test_se)
         );
  SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 clk_gate_cclow_cnt_reg ( 
        .CLK(clk), .EN(N34), .ENCLK(net10338), .TE(test_se) );
  SDFFSQX1 d_cc_reg_0_ ( .D(i_cc_49), .SIN(cclow_cnt[8]), .SMC(test_se), .C(
        clk), .XS(n41), .Q(d_cc[0]) );
  SDFFSQX1 d_cc_reg_1_ ( .D(d_cc[0]), .SIN(d_cc[0]), .SMC(test_se), .C(clk), 
        .XS(n41), .Q(d_cc[1]) );
  SDFFQX1 cclow_cnt_reg_1_ ( .D(N36), .SIN(cclow_cnt[0]), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[1]) );
  SDFFQX1 cclow_cnt_reg_3_ ( .D(N38), .SIN(cclow_cnt[2]), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[3]) );
  SDFFQX1 cclow_cnt_reg_8_ ( .D(n108), .SIN(cclow_cnt[7]), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[8]) );
  SDFFQX1 cclow_cnt_reg_4_ ( .D(N39), .SIN(cclow_cnt[3]), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[4]) );
  SDFFQX1 cclow_cnt_reg_5_ ( .D(N40), .SIN(cclow_cnt[4]), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[5]) );
  SDFFQX1 cclow_cnt_reg_6_ ( .D(N41), .SIN(cclow_cnt[5]), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[6]) );
  SDFFQX1 cclow_cnt_reg_2_ ( .D(N37), .SIN(cclow_cnt[1]), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[2]) );
  SDFFQX1 cclow_cnt_reg_7_ ( .D(N42), .SIN(cclow_cnt[6]), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[7]) );
  SDFFQX1 cclow_cnt_reg_0_ ( .D(N35), .SIN(test_si), .SMC(test_se), .C(
        net10338), .Q(cclow_cnt[0]) );
  INVX1 U3 ( .A(1'b1), .Y(dbgpo[31]) );
  INVXL U5 ( .A(n38), .Y(n35) );
  AND2X1 U6 ( .A(r_txnumk[2]), .B(n36), .Y(c0_txnumk[2]) );
  NAND2X2 U7 ( .A(n11), .B(n12), .Y(mux_rdat[6]) );
  AND2X2 U8 ( .A(r_txnumk[1]), .B(n36), .Y(c0_txnumk[1]) );
  INVX4 U9 ( .A(n38), .Y(n36) );
  INVX3 U10 ( .A(prl_idle), .Y(n38) );
  INVX1 U11 ( .A(n49), .Y(n46) );
  OAI21X1 U12 ( .B(n7), .C(prx_fsm[3]), .A(r_sqlch[1]), .Y(n55) );
  MUX2IX1 U13 ( .D0(n51), .D1(n106), .S(n44), .Y(pff_rxpart[7]) );
  MUX2IX1 U14 ( .D0(n50), .D1(n85), .S(n43), .Y(pff_rxpart[6]) );
  INVXL U15 ( .A(n114), .Y(n5) );
  INVXL U16 ( .A(n5), .Y(ptx_oe) );
  INVXL U17 ( .A(n5), .Y(n7) );
  INVX2 U18 ( .A(n38), .Y(n37) );
  MUX2X1 U19 ( .D0(prl_rdat[1]), .D1(pff_rdat[1]), .S(n37), .Y(mux_rdat[1]) );
  MUX2X1 U20 ( .D0(prl_rdat[3]), .D1(pff_rdat[3]), .S(n37), .Y(mux_rdat[3]) );
  NAND2X1 U21 ( .A(prl_rdat[6]), .B(n9), .Y(n11) );
  NAND2XL U22 ( .A(pff_rdat[6]), .B(n36), .Y(n12) );
  INVXL U23 ( .A(n36), .Y(n9) );
  MUX2X2 U24 ( .D0(prl_rdat[7]), .D1(pff_rdat[7]), .S(n37), .Y(mux_rdat[7]) );
  MUX2X2 U25 ( .D0(prl_rdat[5]), .D1(pff_rdat[5]), .S(n37), .Y(mux_rdat[5]) );
  BUFXL U26 ( .A(n116), .Y(dbgpo[30]) );
  BUFXL U27 ( .A(n117), .Y(dbgpo[29]) );
  MUX2X2 U28 ( .D0(prl_rdat[2]), .D1(pff_rdat[2]), .S(n36), .Y(mux_rdat[2]) );
  AO22XL U29 ( .A(ptx_crcshfi4), .B(n7), .C(prx_crcshfi4), .D(n5), .Y(crcshfi4) );
  AO22XL U30 ( .A(ptx_crcstart), .B(n7), .C(prx_crcstart), .D(n5), .Y(crcstart) );
  BUFXL U31 ( .A(prx_fsm[3]), .Y(dbgpo[23]) );
  BUFX3 U32 ( .A(prx_rcvinf[4]), .Y(dbgpo[19]) );
  BUFXL U33 ( .A(prx_fsm[0]), .Y(dbgpo[20]) );
  BUFXL U34 ( .A(pff_rdat[6]), .Y(dbgpo[14]) );
  BUFXL U35 ( .A(pff_rdat[0]), .Y(dbgpo[8]) );
  BUFXL U36 ( .A(pff_rdat[3]), .Y(dbgpo[11]) );
  BUFXL U37 ( .A(pff_rdat[4]), .Y(dbgpo[12]) );
  BUFXL U38 ( .A(pff_rdat[7]), .Y(dbgpo[15]) );
  BUFXL U39 ( .A(pff_rdat[2]), .Y(dbgpo[10]) );
  BUFXL U40 ( .A(pff_rdat[5]), .Y(dbgpo[13]) );
  BUFXL U41 ( .A(pff_rdat[1]), .Y(dbgpo[9]) );
  BUFXL U42 ( .A(prx_fsm[2]), .Y(dbgpo[22]) );
  BUFXL U43 ( .A(prx_fsm[1]), .Y(dbgpo[21]) );
  AND2XL U44 ( .A(r_txnumk[3]), .B(n36), .Y(c0_txnumk[3]) );
  INVXL U45 ( .A(prl_idle), .Y(n39) );
  INVXL U46 ( .A(n49), .Y(n44) );
  INVXL U47 ( .A(n49), .Y(n45) );
  MUX2X2 U48 ( .D0(prl_last), .D1(pff_one), .S(n35), .Y(mux_one) );
  AND2X2 U49 ( .A(n117), .B(n39), .Y(fifopsh_prl) );
  MUX2XL U50 ( .D0(prl_txreq), .D1(pff_txreq), .S(n35), .Y(n15) );
  AND2XL U51 ( .A(r_txnumk[0]), .B(n36), .Y(c0_txnumk[0]) );
  MUX2XL U52 ( .D0(pff_rdat[0]), .D1(pff_dat_7_1[8]), .S(n43), .Y(
        pff_rxpart[0]) );
  AND2XL U53 ( .A(n37), .B(n46), .Y(rx_pshords) );
  AND2X1 U54 ( .A(prx_setsta[3]), .B(n58), .Y(prx_gdmsgrcvd) );
  NOR2X1 U55 ( .A(prx_fiforst), .B(n42), .Y(fifosrstz) );
  NOR21XL U56 ( .B(ptx_crcshfo4), .A(n5), .Y(crcshfo4) );
  AND2XL U57 ( .A(dbgpo[30]), .B(n35), .Y(fifopop_pff) );
  MUX2X1 U58 ( .D0(pff_dat_7_1[18]), .D1(pff_dat_7_1[34]), .S(n45), .Y(
        pff_c0dat[26]) );
  MUX2X1 U59 ( .D0(pff_dat_7_1[17]), .D1(pff_dat_7_1[33]), .S(n45), .Y(
        pff_c0dat[25]) );
  MUX2X1 U60 ( .D0(pff_dat_7_1[15]), .D1(pff_dat_7_1[31]), .S(n45), .Y(
        pff_c0dat[23]) );
  INVX1 U61 ( .A(n49), .Y(n47) );
  INVX1 U62 ( .A(n49), .Y(n48) );
  INVX1 U63 ( .A(n42), .Y(n41) );
  INVX1 U64 ( .A(n42), .Y(n40) );
  INVX1 U65 ( .A(r_pshords), .Y(n49) );
  MUX2X1 U66 ( .D0(pff_dat_7_1[11]), .D1(pff_dat_7_1[27]), .S(n44), .Y(
        pff_c0dat[19]) );
  NOR21XL U67 ( .B(obsd), .A(prx_setsta[6]), .Y(pff_obsd) );
  NAND42X1 U68 ( .C(pff_rxpart[14]), .D(pff_rxpart[13]), .A(n83), .B(n63), .Y(
        n58) );
  AND3X1 U69 ( .A(n62), .B(pff_rxpart[0]), .C(n61), .Y(n63) );
  NOR32XL U70 ( .B(n60), .C(n59), .A(n54), .Y(n83) );
  NAND21X1 U71 ( .B(pff_rxpart[4]), .A(n53), .Y(n54) );
  INVX1 U72 ( .A(n49), .Y(n43) );
  INVX1 U73 ( .A(pff_rxpart[2]), .Y(n59) );
  INVX1 U74 ( .A(pff_rxpart[3]), .Y(n60) );
  INVX1 U75 ( .A(pff_rxpart[12]), .Y(n53) );
  MUX2IX1 U76 ( .D0(n85), .D1(n89), .S(n45), .Y(pff_c0dat[22]) );
  MUX2BXL U77 ( .D0(pff_dat_7_1[12]), .D1(n93), .S(n45), .Y(pff_c0dat[20]) );
  MUX2IX1 U78 ( .D0(n105), .D1(n100), .S(n45), .Y(pff_c0dat[24]) );
  MUX2IX1 U79 ( .D0(n107), .D1(n91), .S(n45), .Y(pff_c0dat[21]) );
  MUX2BXL U80 ( .D0(pff_dat_7_1[21]), .D1(n90), .S(n45), .Y(pff_c0dat[29]) );
  MUX2X1 U81 ( .D0(pff_dat_7_1[20]), .D1(pff_dat_7_1[36]), .S(n45), .Y(
        pff_c0dat[28]) );
  MUX2X1 U82 ( .D0(pff_dat_7_1[19]), .D1(pff_dat_7_1[35]), .S(n45), .Y(
        pff_c0dat[27]) );
  INVX1 U83 ( .A(n61), .Y(pff_rxpart[1]) );
  INVX1 U84 ( .A(n62), .Y(pff_rxpart[15]) );
  INVX1 U85 ( .A(srstz), .Y(n42) );
  INVX1 U86 ( .A(n72), .Y(n110) );
  INVX1 U87 ( .A(n76), .Y(n112) );
  INVX1 U88 ( .A(n74), .Y(n111) );
  MUX2X2 U89 ( .D0(prl_rdat[4]), .D1(pff_rdat[4]), .S(n36), .Y(mux_rdat[4]) );
  AND2XL U90 ( .A(r_txendk), .B(n37), .Y(c0_txendk) );
  AND2XL U91 ( .A(r_txnumk[4]), .B(n36), .Y(c0_txnumk[4]) );
  AND2XL U92 ( .A(r_txauto[6]), .B(n35), .Y(c0_txauto[6]) );
  BUFXL U93 ( .A(dbgpo[17]), .Y(prx_rcvinf[3]) );
  AOI21AXL U94 ( .B(n7), .C(n37), .A(r_first), .Y(lockena) );
  NAND21XL U95 ( .B(r_txauto[5]), .A(n35), .Y(c0_txauto[5]) );
  AO22XL U96 ( .A(ptx_crcsidat[1]), .B(ptx_oe), .C(prx_crcsidat[1]), .D(n5), 
        .Y(crcsidat[1]) );
  AO22XL U97 ( .A(ptx_crcsidat[0]), .B(ptx_oe), .C(prx_crcsidat[0]), .D(n5), 
        .Y(crcsidat[0]) );
  AO22XL U98 ( .A(ptx_crcsidat[2]), .B(n7), .C(prx_crcsidat[2]), .D(n5), .Y(
        crcsidat[2]) );
  AO22XL U99 ( .A(ptx_crcsidat[3]), .B(n7), .C(prx_crcsidat[3]), .D(n5), .Y(
        crcsidat[3]) );
  MUX2BXL U100 ( .D0(pff_rdat[5]), .D1(n107), .S(n44), .Y(pff_rxpart[5]) );
  INVX1 U101 ( .A(n52), .Y(pff_rxpart[8]) );
  MUX2AXL U102 ( .D0(pff_dat_7_1[0]), .D1(n105), .S(n43), .Y(n52) );
  NOR21XL U103 ( .B(r_auto_gdcrc[1]), .A(n58), .Y(auto_rx_gdcrc) );
  MUX2XL U104 ( .D0(pff_rdat[2]), .D1(pff_dat_7_1[10]), .S(n43), .Y(
        pff_rxpart[2]) );
  MUX2XL U105 ( .D0(pff_rdat[3]), .D1(pff_dat_7_1[11]), .S(n44), .Y(
        pff_rxpart[3]) );
  MUX2X1 U106 ( .D0(pff_dat_7_1[4]), .D1(pff_dat_7_1[20]), .S(n44), .Y(
        pff_rxpart[12]) );
  MUX2IXL U107 ( .D0(pff_rdat[1]), .D1(pff_dat_7_1[9]), .S(n43), .Y(n61) );
  MUX2IX1 U108 ( .D0(pff_dat_7_1[7]), .D1(pff_dat_7_1[23]), .S(n43), .Y(n62)
         );
  MUX2X1 U109 ( .D0(pff_dat_7_1[5]), .D1(pff_dat_7_1[21]), .S(n44), .Y(
        pff_rxpart[13]) );
  MUX2X1 U110 ( .D0(pff_dat_7_1[6]), .D1(pff_dat_7_1[22]), .S(n44), .Y(
        pff_rxpart[14]) );
  MUX2XL U111 ( .D0(pff_rdat[4]), .D1(pff_dat_7_1[12]), .S(n43), .Y(
        pff_rxpart[4]) );
  MUX2BXL U112 ( .D0(pff_dat_7_1[9]), .D1(n99), .S(n44), .Y(pff_c0dat[17]) );
  MUX2BXL U113 ( .D0(pff_dat_7_1[23]), .D1(n86), .S(n46), .Y(pff_c0dat[31]) );
  ENOX1 U114 ( .A(n47), .B(n98), .C(pff_dat_7_1[49]), .D(n48), .Y(
        pff_c0dat[41]) );
  ENOX1 U115 ( .A(n47), .B(n87), .C(pff_dat_7_1[47]), .D(n48), .Y(
        pff_c0dat[39]) );
  ENOXL U116 ( .A(n46), .B(n89), .C(pff_dat_7_1[46]), .D(n48), .Y(
        pff_c0dat[38]) );
  ENOXL U117 ( .A(n46), .B(n93), .C(pff_dat_7_1[44]), .D(n48), .Y(
        pff_c0dat[36]) );
  ENOXL U118 ( .A(n46), .B(n97), .C(pff_dat_7_1[42]), .D(n48), .Y(
        pff_c0dat[34]) );
  MUX2X1 U119 ( .D0(pff_dat_7_1[8]), .D1(pff_dat_7_1[24]), .S(n44), .Y(
        pff_c0dat[16]) );
  MUX2X1 U120 ( .D0(pff_dat_7_1[10]), .D1(pff_dat_7_1[26]), .S(n44), .Y(
        pff_c0dat[18]) );
  ENOX1 U121 ( .A(n47), .B(n86), .C(pff_dat_7_1[55]), .D(r_pshords), .Y(
        pff_c0dat[47]) );
  ENOX1 U122 ( .A(n47), .B(n90), .C(pff_dat_7_1[53]), .D(r_pshords), .Y(
        pff_c0dat[45]) );
  ENOX1 U123 ( .A(n47), .B(n88), .C(pff_dat_7_1[54]), .D(r_pshords), .Y(
        pff_c0dat[46]) );
  ENOX1 U124 ( .A(n47), .B(n100), .C(pff_dat_7_1[48]), .D(n48), .Y(
        pff_c0dat[40]) );
  ENOX1 U125 ( .A(n47), .B(n94), .C(pff_dat_7_1[51]), .D(r_pshords), .Y(
        pff_c0dat[43]) );
  ENOX1 U126 ( .A(n47), .B(n96), .C(pff_dat_7_1[50]), .D(n48), .Y(
        pff_c0dat[42]) );
  ENOX1 U127 ( .A(n47), .B(n92), .C(pff_dat_7_1[52]), .D(r_pshords), .Y(
        pff_c0dat[44]) );
  ENOXL U128 ( .A(n46), .B(n101), .C(pff_dat_7_1[40]), .D(n47), .Y(
        pff_c0dat[32]) );
  ENOXL U129 ( .A(n46), .B(n99), .C(pff_dat_7_1[41]), .D(n48), .Y(
        pff_c0dat[33]) );
  MUX2XL U130 ( .D0(pff_dat_7_1[22]), .D1(pff_dat_7_1[38]), .S(n46), .Y(
        pff_c0dat[30]) );
  ENOXL U131 ( .A(n46), .B(n91), .C(pff_dat_7_1[45]), .D(n48), .Y(
        pff_c0dat[37]) );
  ENOXL U132 ( .A(n46), .B(n95), .C(pff_dat_7_1[43]), .D(n48), .Y(
        pff_c0dat[35]) );
  MUX2XL U133 ( .D0(prl_txauto[2]), .D1(r_txauto[2]), .S(n35), .Y(c0_txauto[2]) );
  MUX2XL U134 ( .D0(prl_txauto[0]), .D1(r_txauto[0]), .S(n35), .Y(c0_txauto[0]) );
  MUX2XL U135 ( .D0(prl_txauto[1]), .D1(r_txauto[1]), .S(n35), .Y(c0_txauto[1]) );
  INVX1 U136 ( .A(pff_dat_7_1[26]), .Y(n97) );
  INVX1 U137 ( .A(pff_dat_7_1[24]), .Y(n101) );
  INVX1 U138 ( .A(pff_dat_7_1[29]), .Y(n91) );
  INVX1 U139 ( .A(pff_dat_7_1[32]), .Y(n100) );
  INVX1 U140 ( .A(pff_dat_7_1[35]), .Y(n94) );
  INVX1 U141 ( .A(pff_dat_7_1[36]), .Y(n92) );
  INVX1 U142 ( .A(pff_dat_7_1[34]), .Y(n96) );
  INVX1 U143 ( .A(pff_dat_7_1[25]), .Y(n99) );
  INVX1 U144 ( .A(pff_dat_7_1[37]), .Y(n90) );
  INVX1 U145 ( .A(pff_dat_7_1[39]), .Y(n86) );
  INVX1 U146 ( .A(pff_dat_7_1[30]), .Y(n89) );
  INVX1 U147 ( .A(pff_dat_7_1[16]), .Y(n105) );
  INVX1 U148 ( .A(pff_dat_7_1[13]), .Y(n107) );
  INVX1 U149 ( .A(pff_dat_7_1[38]), .Y(n88) );
  INVX1 U150 ( .A(pff_dat_7_1[27]), .Y(n95) );
  INVX1 U151 ( .A(pff_dat_7_1[31]), .Y(n87) );
  INVX1 U152 ( .A(pff_dat_7_1[33]), .Y(n98) );
  INVX1 U153 ( .A(pff_dat_7_1[28]), .Y(n93) );
  INVX1 U154 ( .A(pff_dat_7_1[19]), .Y(n102) );
  INVX1 U155 ( .A(pff_dat_7_1[17]), .Y(n104) );
  INVX1 U156 ( .A(pff_dat_7_1[18]), .Y(n103) );
  INVX1 U157 ( .A(pff_dat_7_1[14]), .Y(n85) );
  INVX1 U158 ( .A(pff_dat_7_1[15]), .Y(n106) );
  MUX2XL U159 ( .D0(prl_txauto[4]), .D1(r_txauto[4]), .S(n35), .Y(c0_txauto[4]) );
  NAND21XL U160 ( .B(r_txauto[3]), .A(n35), .Y(c0_txauto[3]) );
  NOR21XL U161 ( .B(ptx_goidle), .A(prl_cany0), .Y(ptx_ack) );
  AOI31X1 U162 ( .A(d_sqlch), .B(n55), .C(r_sqlch[0]), .D(n84), .Y(x_trans) );
  INVX1 U163 ( .A(prx_trans), .Y(n84) );
  OAI211X1 U164 ( .C(cclow_cnt[8]), .D(n65), .A(n41), .B(n82), .Y(n72) );
  XNOR2XL U165 ( .A(d_cc[1]), .B(d_cc[0]), .Y(n82) );
  GEN2XL U166 ( .D(cclow_cnt[1]), .E(cclow_cnt[0]), .C(n80), .B(n110), .A(n66), 
        .Y(N36) );
  GEN2XL U167 ( .D(cclow_cnt[4]), .E(n75), .C(n76), .B(n110), .A(n66), .Y(N39)
         );
  GEN2XL U168 ( .D(cclow_cnt[6]), .E(n111), .C(n73), .B(n110), .A(n66), .Y(N41) );
  GEN2XL U169 ( .D(cclow_cnt[5]), .E(n112), .C(n74), .B(n110), .A(n66), .Y(N40) );
  NOR4XL U170 ( .A(n56), .B(n57), .C(cclow_cnt[5]), .D(cclow_cnt[4]), .Y(
        prx_setsta[0]) );
  OR3XL U171 ( .A(cclow_cnt[7]), .B(cclow_cnt[6]), .C(cclow_cnt[8]), .Y(n57)
         );
  NAND43X1 U172 ( .B(cclow_cnt[3]), .C(cclow_cnt[1]), .D(cclow_cnt[2]), .A(
        cclow_cnt[0]), .Y(n56) );
  NAND21X1 U173 ( .B(cclow_cnt[2]), .A(n80), .Y(n78) );
  NAND21X1 U174 ( .B(cclow_cnt[7]), .A(n73), .Y(n65) );
  NOR2X1 U175 ( .A(n75), .B(cclow_cnt[4]), .Y(n76) );
  NOR2X1 U176 ( .A(n112), .B(cclow_cnt[5]), .Y(n74) );
  NOR2X1 U178 ( .A(n111), .B(cclow_cnt[6]), .Y(n73) );
  NOR2X1 U179 ( .A(cclow_cnt[1]), .B(cclow_cnt[0]), .Y(n80) );
  AOI21X1 U180 ( .B(n65), .C(n67), .A(n72), .Y(N42) );
  NAND21X1 U181 ( .B(n73), .A(cclow_cnt[7]), .Y(n67) );
  AOI21X1 U182 ( .B(n78), .C(n79), .A(n72), .Y(N37) );
  NAND21X1 U183 ( .B(n80), .A(cclow_cnt[2]), .Y(n79) );
  AOI21X1 U184 ( .B(n75), .C(n77), .A(n72), .Y(N38) );
  NAND2X1 U185 ( .A(cclow_cnt[3]), .B(n78), .Y(n77) );
  MUX2BXL U186 ( .D0(pff_dat_7_1[3]), .D1(n102), .S(n43), .Y(pff_rxpart[11])
         );
  MUX2BXL U187 ( .D0(pff_dat_7_1[1]), .D1(n104), .S(n43), .Y(pff_rxpart[9]) );
  MUX2BXL U188 ( .D0(pff_dat_7_1[2]), .D1(n103), .S(n43), .Y(pff_rxpart[10])
         );
  OR2X1 U189 ( .A(n78), .B(cclow_cnt[3]), .Y(n75) );
  NOR2X1 U190 ( .A(cclow_cnt[0]), .B(n72), .Y(N35) );
  INVX1 U191 ( .A(n64), .Y(n108) );
  AOI31X1 U192 ( .A(n110), .B(n65), .C(cclow_cnt[8]), .D(n66), .Y(n64) );
  NAND31X1 U193 ( .C(n66), .A(n72), .B(n81), .Y(N34) );
  AOI21X1 U194 ( .B(d_cc[0]), .C(n109), .A(n42), .Y(n81) );
  NOR3XL U195 ( .A(n42), .B(d_cc[0]), .C(n109), .Y(n66) );
  INVX1 U196 ( .A(d_cc[1]), .Y(n109) );
  INVXL U197 ( .A(pff_rdat[6]), .Y(n50) );
  INVXL U198 ( .A(pff_rdat[7]), .Y(n51) );
  AND2XL U199 ( .A(dbgpo[29]), .B(n37), .Y(fifopsh_pff) );
  MUX2X2 U200 ( .D0(prl_rdat[0]), .D1(pff_rdat[0]), .S(n36), .Y(mux_rdat[0])
         );
  AND2X2 U201 ( .A(n116), .B(n39), .Y(fifopop_prl) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, test_se
 );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_1_, db_cnt_0_, N14, N15, N16, N17, net10356, n8, n1,
         n2, n3, n4, n5;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N14), 
        .ENCLK(net10356), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N17), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net10356), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N16), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net10356), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N15), .SIN(o_dbc), .SMC(test_se), .C(net10356), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n8), .SIN(d_org_0_), .SMC(test_se), .C(net10356), 
        .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n2), .A(n1), .Y(n4) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U5 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n8) );
  NOR2X1 U6 ( .A(n1), .B(n2), .Y(o_chg) );
  NAND3X1 U7 ( .A(db_cnt_1_), .B(db_cnt_0_), .C(test_so), .Y(n1) );
  NOR2X1 U8 ( .A(n5), .B(n4), .Y(N16) );
  XNOR2XL U9 ( .A(db_cnt_1_), .B(db_cnt_0_), .Y(n5) );
  NOR2X1 U10 ( .A(db_cnt_0_), .B(n4), .Y(N15) );
  NOR2X1 U11 ( .A(n3), .B(n4), .Y(N17) );
  AOI21X1 U12 ( .B(db_cnt_1_), .C(db_cnt_0_), .A(test_so), .Y(n3) );
  NAND43X1 U13 ( .B(test_so), .C(db_cnt_0_), .D(db_cnt_1_), .A(n2), .Y(N14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updprl_a0 ( r_spec, r_dat_spec, r_auto_txgdcrc, r_dat_portrole, 
        r_dat_datarole, r_auto_discard, r_set_cpmsgid, r_dat_cpmsgid, r_rdat, 
        r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact, ptx_fifopop, 
        prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, prx_rcvdords, prx_fifowdat, 
        pff_c0dat, prl_rdat, prl_txauto, prl_last, prl_txreq, prl_c0set, 
        prl_cany0, prl_cany0r, prl_cany0w, prl_idle, prl_discard, prl_GCTxDone, 
        prl_fsm, prl_cpmsgid, prl_cany0adr, clk, srstz, test_si, test_so, 
        test_se );
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [2:0] r_dat_cpmsgid;
  input [7:0] r_rdat;
  input [2:0] prx_rcvdords;
  input [7:0] prx_fifowdat;
  input [47:0] pff_c0dat;
  output [7:0] prl_rdat;
  output [6:0] prl_txauto;
  output [3:0] prl_fsm;
  output [2:0] prl_cpmsgid;
  output [7:0] prl_cany0adr;
  input r_auto_txgdcrc, r_dat_portrole, r_dat_datarole, r_auto_discard,
         r_set_cpmsgid, r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact,
         ptx_fifopop, prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, clk, srstz,
         test_si, test_se;
  output prl_last, prl_txreq, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_idle, prl_discard, prl_GCTxDone, test_so;
  wire   n170, sendgdcrc, stoptimer, N41, c0_iop, N113, N114, N115, N116, N117,
         N118, N119, N120, N151, N152, N153, N154, N155, N156, N157, N158,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N189, N190,
         N192, N193, N194, N196, N203, N204, N205, N206, net10379, net10385,
         net10390, net10395, net10400, n99, n100, n52, n37, n49, n54, n57, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n98, n7, n8, n9, n10, n12, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n27, n28, n29, n30, n31, n35, n36, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n50, n51, n53, n55, n56, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n95, n96, n97, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166;
  wire   [1:0] PrlTo;
  wire   [8:0] c0_cnt;
  wire   [7:0] txbuf;

  PrlTimer_1112a0 u0_PrlTimer ( .to(PrlTo), .restart(sendgdcrc), .stop(
        stoptimer), .clk(clk), .srstz(srstz), .test_si(txbuf[7]), .test_so(
        test_so), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_0 clk_gate_txbuf_reg ( .CLK(clk), .EN(N41), 
        .ENCLK(net10379), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_4 clk_gate_c0_adr_reg ( .CLK(clk), .EN(N194), 
        .ENCLK(net10385), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_3 clk_gate_cs_prcl_reg ( .CLK(clk), .EN(N189), 
        .ENCLK(net10390), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_2 clk_gate_c0_cnt_reg ( .CLK(clk), .EN(N196), 
        .ENCLK(net10395), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_1 clk_gate_CpMsgId_reg ( .CLK(clk), .EN(N203), 
        .ENCLK(net10400), .TE(test_se) );
  updprl_a0_DW01_inc_0 r328 ( .A(prl_cany0adr), .SUM({N120, N119, N118, N117, 
        N116, N115, N114, N113}) );
  SDFFQX1 c0_iop_reg ( .D(n99), .SIN(c0_cnt[8]), .SMC(test_se), .C(net10390), 
        .Q(c0_iop) );
  SDFFQX1 canyon_m0_reg ( .D(n100), .SIN(c0_iop), .SMC(test_se), .C(clk), .Q(
        n170) );
  SDFFQX1 c0_adr_reg_1_ ( .D(N152), .SIN(prl_cany0adr[0]), .SMC(test_se), .C(
        net10385), .Q(prl_cany0adr[1]) );
  SDFFQX1 c0_adr_reg_5_ ( .D(N156), .SIN(prl_cany0adr[4]), .SMC(test_se), .C(
        net10385), .Q(prl_cany0adr[5]) );
  SDFFQX1 c0_adr_reg_2_ ( .D(N153), .SIN(prl_cany0adr[1]), .SMC(test_se), .C(
        net10385), .Q(prl_cany0adr[2]) );
  SDFFQX1 c0_adr_reg_0_ ( .D(N151), .SIN(prl_cpmsgid[2]), .SMC(test_se), .C(
        net10385), .Q(prl_cany0adr[0]) );
  SDFFQX1 c0_adr_reg_3_ ( .D(N154), .SIN(prl_cany0adr[2]), .SMC(test_se), .C(
        net10385), .Q(prl_cany0adr[3]) );
  SDFFQX1 c0_adr_reg_6_ ( .D(N157), .SIN(prl_cany0adr[5]), .SMC(test_se), .C(
        net10385), .Q(prl_cany0adr[6]) );
  SDFFQX1 c0_adr_reg_4_ ( .D(N155), .SIN(prl_cany0adr[3]), .SMC(test_se), .C(
        net10385), .Q(prl_cany0adr[4]) );
  SDFFQX1 c0_adr_reg_7_ ( .D(N158), .SIN(prl_cany0adr[6]), .SMC(test_se), .C(
        net10385), .Q(prl_cany0adr[7]) );
  SDFFQXL txbuf_reg_5_ ( .D(r_rdat[5]), .SIN(txbuf[4]), .SMC(test_se), .C(
        net10379), .Q(txbuf[5]) );
  SDFFQX1 txbuf_reg_7_ ( .D(r_rdat[7]), .SIN(txbuf[6]), .SMC(test_se), .C(
        net10379), .Q(txbuf[7]) );
  SDFFQX1 txbuf_reg_4_ ( .D(r_rdat[4]), .SIN(txbuf[3]), .SMC(test_se), .C(
        net10379), .Q(txbuf[4]) );
  SDFFQX1 c0_cnt_reg_7_ ( .D(N172), .SIN(c0_cnt[6]), .SMC(test_se), .C(
        net10395), .Q(c0_cnt[7]) );
  SDFFQX1 c0_cnt_reg_8_ ( .D(N173), .SIN(c0_cnt[7]), .SMC(test_se), .C(
        net10395), .Q(c0_cnt[8]) );
  SDFFQX1 txbuf_reg_0_ ( .D(r_rdat[0]), .SIN(prl_fsm[3]), .SMC(test_se), .C(
        net10379), .Q(txbuf[0]) );
  SDFFQX1 txbuf_reg_1_ ( .D(r_rdat[1]), .SIN(txbuf[0]), .SMC(test_se), .C(
        net10379), .Q(txbuf[1]) );
  SDFFQX1 txbuf_reg_3_ ( .D(r_rdat[3]), .SIN(txbuf[2]), .SMC(test_se), .C(
        net10379), .Q(txbuf[3]) );
  SDFFQX1 CpMsgId_reg_2_ ( .D(N206), .SIN(prl_cpmsgid[1]), .SMC(test_se), .C(
        net10400), .Q(prl_cpmsgid[2]) );
  SDFFQX1 c0_cnt_reg_2_ ( .D(N167), .SIN(n52), .SMC(test_se), .C(net10395), 
        .Q(c0_cnt[2]) );
  SDFFQX1 c0_cnt_reg_3_ ( .D(N168), .SIN(c0_cnt[2]), .SMC(test_se), .C(
        net10395), .Q(c0_cnt[3]) );
  SDFFQX1 c0_cnt_reg_6_ ( .D(N171), .SIN(c0_cnt[5]), .SMC(test_se), .C(
        net10395), .Q(c0_cnt[6]) );
  SDFFQX1 c0_cnt_reg_5_ ( .D(N170), .SIN(c0_cnt[4]), .SMC(test_se), .C(
        net10395), .Q(c0_cnt[5]) );
  SDFFQXL txbuf_reg_2_ ( .D(r_rdat[2]), .SIN(txbuf[1]), .SMC(test_se), .C(
        net10379), .Q(txbuf[2]) );
  SDFFQXL txbuf_reg_6_ ( .D(r_rdat[6]), .SIN(txbuf[5]), .SMC(test_se), .C(
        net10379), .Q(txbuf[6]) );
  SDFFQX1 c0_cnt_reg_4_ ( .D(N169), .SIN(c0_cnt[3]), .SMC(test_se), .C(
        net10395), .Q(c0_cnt[4]) );
  SDFFQXL CpMsgId_reg_1_ ( .D(N205), .SIN(prl_cpmsgid[0]), .SMC(test_se), .C(
        net10400), .Q(prl_cpmsgid[1]) );
  SDFFQXL CpMsgId_reg_0_ ( .D(N204), .SIN(test_si), .SMC(test_se), .C(net10400), .Q(prl_cpmsgid[0]) );
  SDFFQX2 cs_prcl_reg_3_ ( .D(N193), .SIN(prl_fsm[2]), .SMC(test_se), .C(
        net10390), .Q(n21) );
  SDFFQX2 cs_prcl_reg_0_ ( .D(N190), .SIN(n170), .SMC(test_se), .C(net10390), 
        .Q(n19) );
  SDFFQX4 cs_prcl_reg_1_ ( .D(n166), .SIN(prl_fsm[0]), .SMC(test_se), .C(
        net10390), .Q(prl_fsm[1]) );
  SDFFQX2 cs_prcl_reg_2_ ( .D(N192), .SIN(prl_fsm[1]), .SMC(test_se), .C(
        net10390), .Q(prl_fsm[2]) );
  SDFFQX1 c0_cnt_reg_1_ ( .D(N166), .SIN(c0_cnt[0]), .SMC(test_se), .C(
        net10395), .Q(n52) );
  SDFFQX4 c0_cnt_reg_0_ ( .D(N165), .SIN(prl_cany0adr[7]), .SMC(test_se), .C(
        net10395), .Q(c0_cnt[0]) );
  INVX1 U3 ( .A(1'b0), .Y(prl_txauto[3]) );
  INVX1 U5 ( .A(1'b0), .Y(prl_txauto[5]) );
  INVX1 U7 ( .A(1'b1), .Y(prl_txauto[6]) );
  INVX3 U9 ( .A(n39), .Y(n45) );
  NAND21X2 U10 ( .B(n21), .A(n19), .Y(n55) );
  INVX2 U11 ( .A(n22), .Y(prl_fsm[3]) );
  NAND21X2 U12 ( .B(c0_cnt[2]), .A(n61), .Y(n65) );
  INVX2 U13 ( .A(n63), .Y(n61) );
  NAND21X2 U14 ( .B(c0_cnt[7]), .A(n96), .Y(n104) );
  INVX3 U15 ( .A(n101), .Y(n96) );
  NAND21X2 U16 ( .B(c0_cnt[8]), .A(n102), .Y(n103) );
  INVXL U17 ( .A(c0_cnt[4]), .Y(n73) );
  NAND21X1 U18 ( .B(n20), .A(n105), .Y(prl_txauto[4]) );
  NAND32X1 U19 ( .B(prl_fsm[3]), .C(n106), .A(n20), .Y(n141) );
  INVX2 U20 ( .A(n141), .Y(prl_idle) );
  NOR21XL U21 ( .B(prx_rcvdords[0]), .A(prx_rcvdords[1]), .Y(n155) );
  INVX1 U22 ( .A(prx_rcvdords[2]), .Y(n154) );
  OAI21X1 U23 ( .B(prx_eoprcvd), .C(pid_ccidle), .A(n14), .Y(n38) );
  INVX1 U24 ( .A(c0_cnt[5]), .Y(n75) );
  INVX1 U25 ( .A(c0_cnt[3]), .Y(n74) );
  OAI21X1 U26 ( .B(ptx_txact), .C(prl_txauto[4]), .A(n142), .Y(prl_txreq) );
  NOR21X1 U27 ( .B(txbuf[7]), .A(n161), .Y(n164) );
  OAI22X1 U28 ( .A(n161), .B(n152), .C(n151), .D(n150), .Y(prl_rdat[3]) );
  NAND31X1 U29 ( .C(n9), .A(n162), .B(r_spec[1]), .Y(n163) );
  NOR21XL U30 ( .B(txbuf[6]), .A(n161), .Y(n160) );
  OR2X2 U31 ( .A(n52), .B(c0_cnt[0]), .Y(n63) );
  INVX2 U32 ( .A(prx_fifopsh), .Y(n129) );
  INVX2 U33 ( .A(n10), .Y(prl_cany0w) );
  NAND21XL U34 ( .B(n106), .A(prl_fsm[3]), .Y(n130) );
  INVXL U35 ( .A(n103), .Y(n144) );
  INVX1 U36 ( .A(n19), .Y(n20) );
  INVX1 U37 ( .A(n20), .Y(prl_fsm[0]) );
  INVX1 U38 ( .A(n130), .Y(n105) );
  INVX1 U39 ( .A(n130), .Y(n14) );
  INVXL U40 ( .A(n9), .Y(n17) );
  AND2X1 U41 ( .A(txbuf[4]), .B(n153), .Y(prl_rdat[4]) );
  BUFX3 U42 ( .A(n151), .Y(n7) );
  BUFX3 U43 ( .A(n12), .Y(n9) );
  INVXL U44 ( .A(n7), .Y(n8) );
  NAND21X1 U45 ( .B(prl_fsm[1]), .A(n42), .Y(n106) );
  NAND21X1 U46 ( .B(prl_fsm[2]), .A(prl_fsm[1]), .Y(n39) );
  NAND21X2 U47 ( .B(n46), .A(n45), .Y(n12) );
  INVX1 U48 ( .A(n21), .Y(n22) );
  OR2X2 U49 ( .A(n19), .B(n21), .Y(n46) );
  INVXL U50 ( .A(n8), .Y(n16) );
  NAND32X1 U51 ( .B(n130), .C(prl_fsm[0]), .A(prx_fifopsh), .Y(n10) );
  OAI22AXL U52 ( .D(n103), .C(n18), .A(n24), .B(n112), .Y(n15) );
  OAI21X1 U53 ( .B(n103), .C(prl_txauto[4]), .A(n16), .Y(prl_last) );
  INVXL U54 ( .A(prl_txauto[4]), .Y(n143) );
  INVX2 U55 ( .A(n65), .Y(n77) );
  INVX2 U56 ( .A(n104), .Y(n102) );
  NAND2X2 U57 ( .A(n12), .B(n151), .Y(n161) );
  INVX2 U58 ( .A(prl_fsm[2]), .Y(n42) );
  BUFXL U59 ( .A(n132), .Y(n18) );
  OAI22AX1 U60 ( .D(n103), .C(n132), .A(n129), .B(n112), .Y(prl_cany0r) );
  NAND5X2 U61 ( .A(n77), .B(n76), .C(n75), .D(n74), .E(n73), .Y(n101) );
  INVX1 U62 ( .A(n24), .Y(n23) );
  BUFXL U63 ( .A(n129), .Y(n24) );
  NAND31XL U64 ( .C(n12), .A(n158), .B(r_spec[0]), .Y(n159) );
  NAND42XL U65 ( .C(r_dat_datarole), .D(n12), .A(n155), .B(n154), .Y(n156) );
  OAI221X1 U66 ( .A(n161), .B(n145), .C(n7), .D(r_dat_portrole), .E(n9), .Y(
        prl_rdat[0]) );
  OAI22X1 U67 ( .A(n161), .B(n149), .C(n7), .D(n148), .Y(prl_rdat[2]) );
  INVX1 U68 ( .A(n165), .Y(prl_cany0) );
  OAI211XL U69 ( .C(n35), .D(n7), .A(n108), .B(n134), .Y(N192) );
  INVXL U70 ( .A(n112), .Y(n120) );
  NAND21XL U71 ( .B(n14), .A(n112), .Y(n59) );
  INVXL U72 ( .A(c0_cnt[6]), .Y(n76) );
  INVX1 U73 ( .A(r_discard), .Y(n115) );
  NOR21XL U74 ( .B(prx_gdmsgrcvd), .A(r_set_cpmsgid), .Y(n57) );
  OR3XL U75 ( .A(r_set_cpmsgid), .B(prx_gdmsgrcvd), .C(n35), .Y(N203) );
  INVXL U76 ( .A(ptx_fifopop), .Y(n123) );
  INVX1 U77 ( .A(srstz), .Y(n35) );
  INVX1 U78 ( .A(n49), .Y(prl_c0set) );
  INVX1 U79 ( .A(n117), .Y(n37) );
  NAND32X1 U80 ( .B(n116), .C(prl_discard), .A(n115), .Y(n117) );
  OR3XL U81 ( .A(pff_c0dat[26]), .B(pff_c0dat[25]), .C(pff_c0dat[23]), .Y(n87)
         );
  NAND21X1 U82 ( .B(n118), .A(n116), .Y(n142) );
  INVX1 U83 ( .A(n125), .Y(n58) );
  NAND21X2 U84 ( .B(n55), .A(n45), .Y(n151) );
  NAND21XL U85 ( .B(n55), .A(n53), .Y(n112) );
  INVX1 U86 ( .A(n51), .Y(n53) );
  NAND4X1 U87 ( .A(n79), .B(n80), .C(n81), .D(n82), .Y(n49) );
  NOR4XL U88 ( .A(n86), .B(n87), .C(pff_c0dat[22]), .D(pff_c0dat[20]), .Y(n81)
         );
  NOR4XL U89 ( .A(n83), .B(n84), .C(pff_c0dat[36]), .D(pff_c0dat[34]), .Y(n82)
         );
  NOR42XL U90 ( .C(pff_c0dat[46]), .D(pff_c0dat[40]), .A(n92), .B(n93), .Y(n79) );
  NOR42XL U91 ( .C(pff_c0dat[1]), .D(pff_c0dat[19]), .A(n89), .B(n90), .Y(n80)
         );
  NAND3X1 U92 ( .A(pff_c0dat[12]), .B(pff_c0dat[0]), .C(pff_c0dat[17]), .Y(n90) );
  NAND42X1 U93 ( .C(pff_c0dat[14]), .D(pff_c0dat[13]), .A(prx_gdmsgrcvd), .B(
        n91), .Y(n89) );
  OAI221XL U94 ( .A(n153), .B(n123), .C(n141), .D(n122), .E(n133), .Y(n127) );
  OAI22X1 U95 ( .A(n119), .B(n139), .C(n37), .D(n118), .Y(n128) );
  OAI211X1 U96 ( .C(n35), .D(n50), .A(n48), .B(n134), .Y(n166) );
  AOI31XL U97 ( .A(n114), .B(n115), .C(n47), .D(n17), .Y(n50) );
  INVX1 U98 ( .A(n142), .Y(n47) );
  OAI21BBX1 U99 ( .A(r_dat_cpmsgid[2]), .B(r_set_cpmsgid), .C(n27), .Y(N206)
         );
  AOI21X1 U100 ( .B(pff_c0dat[11]), .C(n57), .A(n35), .Y(n27) );
  OAI21BBX1 U101 ( .A(r_dat_cpmsgid[0]), .B(r_set_cpmsgid), .C(n28), .Y(N204)
         );
  AOI21X1 U102 ( .B(pff_c0dat[9]), .C(n57), .A(n35), .Y(n28) );
  OAI21BBX1 U103 ( .A(r_dat_cpmsgid[1]), .B(r_set_cpmsgid), .C(n29), .Y(N205)
         );
  AOI21X1 U104 ( .B(pff_c0dat[10]), .C(n57), .A(n35), .Y(n29) );
  INVX1 U105 ( .A(n131), .Y(n113) );
  INVX1 U106 ( .A(sendgdcrc), .Y(n122) );
  INVX1 U107 ( .A(n40), .Y(n108) );
  OAI31XL U108 ( .A(n139), .B(n35), .C(n165), .D(n48), .Y(n40) );
  NOR3XL U109 ( .A(prx_fifowdat[5]), .B(prx_fifowdat[7]), .C(prx_fifowdat[6]), 
        .Y(n98) );
  NAND32X1 U110 ( .B(pff_c0dat[28]), .C(pff_c0dat[27]), .A(n88), .Y(n86) );
  NOR3XL U111 ( .A(pff_c0dat[29]), .B(pff_c0dat[32]), .C(pff_c0dat[31]), .Y(
        n88) );
  INVX1 U112 ( .A(n54), .Y(n109) );
  AO22X1 U113 ( .A(N117), .B(n59), .C(n58), .D(prx_fifowdat[4]), .Y(N155) );
  AO22X1 U114 ( .A(N119), .B(n59), .C(prx_fifowdat[6]), .D(n58), .Y(N157) );
  AO22X1 U115 ( .A(N118), .B(n59), .C(prx_fifowdat[5]), .D(n58), .Y(N156) );
  INVX1 U116 ( .A(n44), .Y(n116) );
  NAND21X1 U117 ( .B(n121), .A(PrlTo[0]), .Y(n44) );
  OR2XL U118 ( .A(n55), .B(n106), .Y(n118) );
  AND3X1 U119 ( .A(ptx_ack), .B(n165), .C(n140), .Y(prl_GCTxDone) );
  INVX1 U120 ( .A(n139), .Y(n140) );
  INVX1 U121 ( .A(n114), .Y(prl_discard) );
  INVX1 U122 ( .A(n124), .Y(n110) );
  NAND32XL U123 ( .B(n55), .C(n42), .A(n41), .Y(n125) );
  NAND21X1 U124 ( .B(n121), .A(n120), .Y(n133) );
  INVX1 U125 ( .A(n72), .Y(n69) );
  INVX1 U126 ( .A(n68), .Y(n66) );
  INVX1 U127 ( .A(ptx_ack), .Y(n119) );
  AO22X1 U128 ( .A(N116), .B(n59), .C(n58), .D(prx_fifowdat[3]), .Y(N154) );
  NAND21X1 U129 ( .B(n157), .A(n156), .Y(prl_rdat[5]) );
  INVXL U130 ( .A(txbuf[1]), .Y(n147) );
  INVXL U131 ( .A(prl_cpmsgid[0]), .Y(n146) );
  INVXL U132 ( .A(txbuf[2]), .Y(n149) );
  INVXL U133 ( .A(prl_cpmsgid[1]), .Y(n148) );
  NAND21X1 U134 ( .B(n164), .A(n163), .Y(prl_rdat[7]) );
  INVXL U135 ( .A(txbuf[0]), .Y(n145) );
  INVXL U136 ( .A(txbuf[3]), .Y(n152) );
  NAND21X1 U137 ( .B(r_dat_spec[0]), .A(r_spec[1]), .Y(n158) );
  NAND21X1 U138 ( .B(r_dat_spec[1]), .A(r_spec[0]), .Y(n162) );
  INVXL U139 ( .A(prl_cpmsgid[2]), .Y(n150) );
  NAND21XL U140 ( .B(n41), .A(prl_fsm[2]), .Y(n51) );
  INVXL U141 ( .A(prl_fsm[1]), .Y(n41) );
  OAI21BX1 U142 ( .C(PrlTo[0]), .B(r_auto_discard), .A(n37), .Y(stoptimer) );
  NAND21X1 U143 ( .B(r_rdy), .A(n138), .Y(N41) );
  OAI21BBX1 U144 ( .A(r_auto_txgdcrc), .B(prx_gdmsgrcvd), .C(n49), .Y(
        sendgdcrc) );
  NAND43X1 U145 ( .B(prx_fifowdat[0]), .C(n54), .D(n124), .A(n113), .Y(n48) );
  MUX2X1 U146 ( .D0(prx_fifowdat[1]), .D1(c0_iop), .S(n30), .Y(n99) );
  NAND4XL U147 ( .A(n113), .B(n53), .C(n20), .D(n109), .Y(n30) );
  INVX1 U148 ( .A(c0_iop), .Y(n136) );
  INVX1 U149 ( .A(n134), .Y(n135) );
  OA21X1 U150 ( .B(n120), .C(n111), .A(n113), .Y(N193) );
  AND3X1 U151 ( .A(prx_fifowdat[0]), .B(n110), .C(n109), .Y(n111) );
  OA21X1 U152 ( .B(n170), .C(prl_c0set), .A(n113), .Y(n100) );
  NAND43X1 U153 ( .B(prx_fifowdat[3]), .C(prx_fifowdat[4]), .D(prx_fifowdat[2]), .A(n98), .Y(n54) );
  OR3XL U154 ( .A(pff_c0dat[41]), .B(pff_c0dat[39]), .C(pff_c0dat[38]), .Y(n84) );
  NOR3XL U155 ( .A(pff_c0dat[15]), .B(pff_c0dat[18]), .C(pff_c0dat[16]), .Y(
        n91) );
  NAND42X1 U156 ( .C(pff_c0dat[47]), .D(pff_c0dat[45]), .A(n165), .B(n85), .Y(
        n83) );
  NOR3XL U157 ( .A(pff_c0dat[42]), .B(pff_c0dat[44]), .C(pff_c0dat[43]), .Y(
        n85) );
  NAND4X1 U158 ( .A(pff_c0dat[33]), .B(pff_c0dat[30]), .C(n94), .D(
        pff_c0dat[2]), .Y(n92) );
  AND2X1 U162 ( .A(pff_c0dat[24]), .B(pff_c0dat[21]), .Y(n94) );
  NAND3X1 U163 ( .A(pff_c0dat[37]), .B(pff_c0dat[35]), .C(pff_c0dat[3]), .Y(
        n93) );
  BUFXL U164 ( .A(prx_rcvdords[2]), .Y(prl_txauto[2]) );
  BUFXL U165 ( .A(prx_rcvdords[0]), .Y(prl_txauto[0]) );
  BUFXL U166 ( .A(prx_rcvdords[1]), .Y(prl_txauto[1]) );
  GEN2XL U167 ( .D(c0_cnt[7]), .E(n101), .C(n102), .B(n14), .A(n97), .Y(N172)
         );
  AND2X1 U168 ( .A(prx_fifowdat[7]), .B(n120), .Y(n97) );
  GEN2XL U169 ( .D(c0_cnt[6]), .E(n95), .C(n96), .B(n14), .A(n78), .Y(N171) );
  AND2X1 U170 ( .A(prx_fifowdat[6]), .B(n120), .Y(n78) );
  GEN2XL U171 ( .D(c0_cnt[4]), .E(n68), .C(n69), .B(n14), .A(n67), .Y(N169) );
  AND2X1 U172 ( .A(n120), .B(prx_fifowdat[4]), .Y(n67) );
  AO22X1 U173 ( .A(N120), .B(n59), .C(prx_fifowdat[7]), .D(n58), .Y(N158) );
  GEN2XL U174 ( .D(c0_cnt[5]), .E(n72), .C(n71), .B(n14), .A(n70), .Y(N170) );
  INVX1 U175 ( .A(n95), .Y(n71) );
  AND2X1 U176 ( .A(prx_fifowdat[5]), .B(n120), .Y(n70) );
  INVX1 U177 ( .A(n170), .Y(n165) );
  INVX1 U178 ( .A(pid_ccidle), .Y(n121) );
  NAND32XL U179 ( .B(prl_fsm[3]), .C(n51), .A(n20), .Y(n124) );
  NAND32X1 U180 ( .B(n43), .C(n118), .A(PrlTo[1]), .Y(n114) );
  INVX1 U181 ( .A(r_auto_discard), .Y(n43) );
  OR3XL U182 ( .A(prl_fsm[1]), .B(n42), .C(n46), .Y(n139) );
  AND2X1 U183 ( .A(n120), .B(prx_fifowdat[3]), .Y(n64) );
  NAND21XL U184 ( .B(c0_cnt[4]), .A(n66), .Y(n72) );
  NAND21XL U185 ( .B(c0_cnt[5]), .A(n69), .Y(n95) );
  NAND21XL U186 ( .B(c0_cnt[3]), .A(n77), .Y(n68) );
  GEN2XL U187 ( .D(c0_cnt[2]), .E(n63), .C(n77), .B(n14), .A(n62), .Y(N167) );
  AND2X1 U188 ( .A(n120), .B(prx_fifowdat[2]), .Y(n62) );
  GEN2XL U189 ( .D(n52), .E(c0_cnt[0]), .C(n61), .B(n14), .A(n60), .Y(N166) );
  AND2X1 U190 ( .A(prx_fifowdat[1]), .B(n120), .Y(n60) );
  NOR21XL U191 ( .B(n105), .A(n31), .Y(N173) );
  AOI21XL U192 ( .B(c0_cnt[8]), .C(n104), .A(n144), .Y(n31) );
  AO22X1 U193 ( .A(N113), .B(n59), .C(prx_fifowdat[0]), .D(n58), .Y(N151) );
  AO22X1 U194 ( .A(N114), .B(n59), .C(prx_fifowdat[1]), .D(n58), .Y(N152) );
  AO22X1 U195 ( .A(N115), .B(n59), .C(n58), .D(prx_fifowdat[2]), .Y(N153) );
  OAI22XL U196 ( .A(n112), .B(n56), .C(c0_cnt[0]), .D(n130), .Y(N165) );
  INVX1 U197 ( .A(prx_fifowdat[0]), .Y(n56) );
  AND2XL U198 ( .A(n113), .B(n15), .Y(N196) );
  GEN2XL U199 ( .D(c0_cnt[3]), .E(n65), .C(n66), .B(n14), .A(n64), .Y(N168) );
  OAI22XL U200 ( .A(n161), .B(n147), .C(n151), .D(n146), .Y(prl_rdat[1]) );
  NOR21XL U201 ( .B(txbuf[5]), .A(n161), .Y(n157) );
  INVXL U202 ( .A(n161), .Y(n153) );
  INVXL U203 ( .A(n15), .Y(n138) );
  AO21XL U204 ( .B(n125), .C(n124), .A(n24), .Y(n126) );
  NAND43X1 U205 ( .B(n131), .C(n128), .D(n127), .A(n126), .Y(N189) );
  OAI211XL U206 ( .C(n112), .D(n131), .A(n108), .B(n107), .Y(N190) );
  NAND21X1 U207 ( .B(n131), .A(n58), .Y(n134) );
  NAND21X1 U208 ( .B(n160), .A(n159), .Y(prl_rdat[6]) );
  AOI31XL U209 ( .A(n133), .B(n10), .C(n18), .D(n131), .Y(n137) );
  AO21XL U210 ( .B(n141), .C(n9), .A(n35), .Y(n107) );
  OAI211XL U211 ( .C(prl_fsm[0]), .D(n38), .A(srstz), .B(n36), .Y(n131) );
  NAND21X2 U212 ( .B(prl_txauto[4]), .A(ptx_fifopop), .Y(n132) );
  AO22XL U213 ( .A(n137), .B(n136), .C(n135), .D(n23), .Y(N194) );
  AOI32XL U214 ( .A(n54), .B(n23), .C(n110), .D(ptx_ack), .E(n143), .Y(n36) );
endmodule


module updprl_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1XL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1XL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  HAD1XL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  XOR2XL U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVXL U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module PrlTimer_1112a0 ( to, restart, stop, clk, srstz, test_si, test_so, 
        test_se );
  output [1:0] to;
  input restart, stop, clk, srstz, test_si, test_se;
  output test_so;
  wire   timer_10_, timer_9_, timer_8_, timer_7_, timer_6_, timer_5_, timer_4_,
         timer_3_, timer_2_, timer_1_, timer_0_, ena, N4, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, net10417, n7, n8, n9, n10, n11, n12, n13, n1,
         n2, n3, n4;

  SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 clk_gate_timer_reg ( .CLK(clk), .EN(N18), .ENCLK(net10417), .TE(test_se) );
  PrlTimer_1112a0_DW01_inc_0 add_25 ( .A({test_so, timer_10_, timer_9_, 
        timer_8_, timer_7_, timer_6_, timer_5_, timer_4_, timer_3_, timer_2_, 
        timer_1_, timer_0_}), .SUM({N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, N4}) );
  SDFFQX1 ena_reg ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .Q(ena) );
  SDFFQX1 timer_reg_1_ ( .D(N20), .SIN(timer_0_), .SMC(test_se), .C(net10417), 
        .Q(timer_1_) );
  SDFFQX1 timer_reg_2_ ( .D(N21), .SIN(timer_1_), .SMC(test_se), .C(net10417), 
        .Q(timer_2_) );
  SDFFQX1 timer_reg_0_ ( .D(N19), .SIN(ena), .SMC(test_se), .C(net10417), .Q(
        timer_0_) );
  SDFFQX1 timer_reg_11_ ( .D(N30), .SIN(timer_10_), .SMC(test_se), .C(net10417), .Q(test_so) );
  SDFFQX1 timer_reg_9_ ( .D(N28), .SIN(timer_8_), .SMC(test_se), .C(net10417), 
        .Q(timer_9_) );
  SDFFQX1 timer_reg_10_ ( .D(N29), .SIN(timer_9_), .SMC(test_se), .C(net10417), 
        .Q(timer_10_) );
  SDFFQX1 timer_reg_7_ ( .D(N26), .SIN(timer_6_), .SMC(test_se), .C(net10417), 
        .Q(timer_7_) );
  SDFFQX1 timer_reg_6_ ( .D(N25), .SIN(timer_5_), .SMC(test_se), .C(net10417), 
        .Q(timer_6_) );
  SDFFQX1 timer_reg_8_ ( .D(N27), .SIN(timer_7_), .SMC(test_se), .C(net10417), 
        .Q(timer_8_) );
  SDFFQX1 timer_reg_3_ ( .D(N22), .SIN(timer_2_), .SMC(test_se), .C(net10417), 
        .Q(timer_3_) );
  SDFFQX1 timer_reg_4_ ( .D(N23), .SIN(timer_3_), .SMC(test_se), .C(net10417), 
        .Q(timer_4_) );
  SDFFQX1 timer_reg_5_ ( .D(N24), .SIN(timer_4_), .SMC(test_se), .C(net10417), 
        .Q(timer_5_) );
  BUFX3 U3 ( .A(n11), .Y(n1) );
  OAI31XL U4 ( .A(timer_10_), .B(timer_9_), .C(timer_8_), .D(test_so), .Y(n13)
         );
  NOR21XL U5 ( .B(N7), .A(n11), .Y(N22) );
  NOR21XL U6 ( .B(N8), .A(n11), .Y(N23) );
  NOR21XL U7 ( .B(N12), .A(n11), .Y(N27) );
  NOR21XL U8 ( .B(N11), .A(n11), .Y(N26) );
  NOR21XL U9 ( .B(N10), .A(n11), .Y(N25) );
  NOR21XL U10 ( .B(N9), .A(n11), .Y(N24) );
  NOR21XL U11 ( .B(N14), .A(n11), .Y(N29) );
  NOR21XL U12 ( .B(N13), .A(n11), .Y(N28) );
  NOR21XL U13 ( .B(N6), .A(n11), .Y(N21) );
  NOR21XL U14 ( .B(N5), .A(n1), .Y(N20) );
  NAND31X1 U15 ( .C(restart), .A(n1), .B(srstz), .Y(N18) );
  NAND3X1 U16 ( .A(srstz), .B(ena), .C(n12), .Y(n11) );
  NOR3XL U17 ( .A(to[1]), .B(stop), .C(restart), .Y(n12) );
  NOR21XL U18 ( .B(N15), .A(n1), .Y(N30) );
  NOR21XL U19 ( .B(N4), .A(n1), .Y(N19) );
  INVX1 U20 ( .A(n10), .Y(n2) );
  AOI31X1 U21 ( .A(srstz), .B(n3), .C(ena), .D(restart), .Y(n10) );
  INVX1 U22 ( .A(stop), .Y(n3) );
  AO21X1 U23 ( .B(timer_4_), .C(timer_3_), .A(timer_5_), .Y(n9) );
  INVX1 U24 ( .A(n7), .Y(to[0]) );
  AOI211X1 U25 ( .C(n4), .D(timer_9_), .A(timer_10_), .B(test_so), .Y(n7) );
  INVX1 U26 ( .A(n8), .Y(n4) );
  AOI211X1 U27 ( .C(timer_6_), .D(n9), .A(timer_8_), .B(timer_7_), .Y(n8) );
  INVX1 U28 ( .A(n13), .Y(to[1]) );
endmodule


module PrlTimer_1112a0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyff_DEPTH_NUM34_DEPTH_NBT6 ( r_psh, r_pop, prx_psh, ptx_pop, r_last, 
        r_unlock, i_lockena, r_fiforst, i_ccidle, r_wdat, prx_wdat, txreq, 
        ffack, rdat0, full, empty, one, half, obsd, dat_7_1, ptr, fifowdat, 
        fifopsh, clk, srstz, test_si, test_se );
  input [7:0] r_wdat;
  input [7:0] prx_wdat;
  output [1:0] ffack;
  output [7:0] rdat0;
  output [55:0] dat_7_1;
  output [5:0] ptr;
  output [7:0] fifowdat;
  input r_psh, r_pop, prx_psh, ptx_pop, r_last, r_unlock, i_lockena, r_fiforst,
         i_ccidle, clk, srstz, test_si, test_se;
  output txreq, full, empty, one, half, obsd, fifopsh;
  wire   ps_locked, locked, mem_8__7_, mem_8__6_, mem_8__5_, mem_8__4_,
         mem_8__3_, mem_8__2_, mem_8__1_, mem_8__0_, mem_9__7_, mem_9__6_,
         mem_9__5_, mem_9__4_, mem_9__3_, mem_9__2_, mem_9__1_, mem_9__0_,
         mem_10__7_, mem_10__6_, mem_10__5_, mem_10__4_, mem_10__3_,
         mem_10__2_, mem_10__1_, mem_10__0_, mem_11__7_, mem_11__6_,
         mem_11__5_, mem_11__4_, mem_11__3_, mem_11__2_, mem_11__1_,
         mem_11__0_, mem_12__7_, mem_12__6_, mem_12__5_, mem_12__4_,
         mem_12__3_, mem_12__2_, mem_12__1_, mem_12__0_, mem_13__7_,
         mem_13__6_, mem_13__5_, mem_13__4_, mem_13__3_, mem_13__2_,
         mem_13__1_, mem_13__0_, mem_14__7_, mem_14__6_, mem_14__5_,
         mem_14__4_, mem_14__3_, mem_14__2_, mem_14__1_, mem_14__0_,
         mem_15__7_, mem_15__6_, mem_15__5_, mem_15__4_, mem_15__3_,
         mem_15__2_, mem_15__1_, mem_15__0_, mem_16__7_, mem_16__6_,
         mem_16__5_, mem_16__4_, mem_16__3_, mem_16__2_, mem_16__1_,
         mem_16__0_, mem_17__7_, mem_17__6_, mem_17__5_, mem_17__4_,
         mem_17__3_, mem_17__2_, mem_17__1_, mem_17__0_, mem_18__7_,
         mem_18__6_, mem_18__5_, mem_18__4_, mem_18__3_, mem_18__2_,
         mem_18__1_, mem_18__0_, mem_19__7_, mem_19__6_, mem_19__5_,
         mem_19__4_, mem_19__3_, mem_19__2_, mem_19__1_, mem_19__0_,
         mem_20__7_, mem_20__6_, mem_20__5_, mem_20__4_, mem_20__3_,
         mem_20__2_, mem_20__1_, mem_20__0_, mem_21__7_, mem_21__6_,
         mem_21__5_, mem_21__4_, mem_21__3_, mem_21__2_, mem_21__1_,
         mem_21__0_, mem_22__7_, mem_22__6_, mem_22__5_, mem_22__4_,
         mem_22__3_, mem_22__2_, mem_22__1_, mem_22__0_, mem_23__7_,
         mem_23__6_, mem_23__5_, mem_23__4_, mem_23__3_, mem_23__2_,
         mem_23__1_, mem_23__0_, mem_24__7_, mem_24__6_, mem_24__5_,
         mem_24__4_, mem_24__3_, mem_24__2_, mem_24__1_, mem_24__0_,
         mem_25__7_, mem_25__6_, mem_25__5_, mem_25__4_, mem_25__3_,
         mem_25__2_, mem_25__1_, mem_25__0_, mem_26__7_, mem_26__6_,
         mem_26__5_, mem_26__4_, mem_26__3_, mem_26__2_, mem_26__1_,
         mem_26__0_, mem_27__7_, mem_27__6_, mem_27__5_, mem_27__4_,
         mem_27__3_, mem_27__2_, mem_27__1_, mem_27__0_, mem_28__7_,
         mem_28__6_, mem_28__5_, mem_28__4_, mem_28__3_, mem_28__2_,
         mem_28__1_, mem_28__0_, mem_29__7_, mem_29__6_, mem_29__5_,
         mem_29__4_, mem_29__3_, mem_29__2_, mem_29__1_, mem_29__0_,
         mem_30__7_, mem_30__6_, mem_30__5_, mem_30__4_, mem_30__3_,
         mem_30__2_, mem_30__1_, mem_30__0_, mem_31__7_, mem_31__6_,
         mem_31__5_, mem_31__4_, mem_31__3_, mem_31__2_, mem_31__1_,
         mem_31__0_, mem_32__7_, mem_32__6_, mem_32__5_, mem_32__4_,
         mem_32__3_, mem_32__2_, mem_32__1_, mem_32__0_, mem_33__7_,
         mem_33__6_, mem_33__5_, mem_33__4_, mem_33__3_, mem_33__2_,
         mem_33__1_, mem_33__0_, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1053, N1054, N1055,
         N1056, N1057, N1058, N1059, net10435, net10441, net10446, net10451,
         net10456, net10461, net10466, net10471, net10476, net10481, net10486,
         net10491, net10496, net10501, net10506, net10511, net10516, net10521,
         net10526, net10531, net10536, net10541, net10546, net10551, net10556,
         net10561, net10566, net10571, net10576, net10581, net10586, net10591,
         net10596, net10601, net10606, n58, n60, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n150, n151, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n262, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n462, n463, n464, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n29,
         n30, n31, n32, n33, n34, n35, n37, n38, n39, n40, n41, n42, n43, n45,
         n46, n47, n48, n49, n50, n51, n53, n54, n55, n56, n57, n59, n61, n78,
         n99, n126, n137, n149, n152, n163, n179, n190, n191, n203, n204, n249,
         n261, n275, n286, n298, n299, n311, n356, n357, n393, n405, n406,
         n427, n428, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n465, n466, n467, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577;

  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 clk_gate_mem_reg_0_ ( 
        .CLK(clk), .EN(N1022), .ENCLK(net10435), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 clk_gate_mem_reg_1_ ( 
        .CLK(clk), .EN(N1013), .ENCLK(net10441), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 clk_gate_mem_reg_2_ ( 
        .CLK(clk), .EN(N1004), .ENCLK(net10446), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 clk_gate_mem_reg_3_ ( 
        .CLK(clk), .EN(N995), .ENCLK(net10451), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 clk_gate_mem_reg_4_ ( 
        .CLK(clk), .EN(N986), .ENCLK(net10456), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 clk_gate_mem_reg_5_ ( 
        .CLK(clk), .EN(N977), .ENCLK(net10461), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 clk_gate_mem_reg_6_ ( 
        .CLK(clk), .EN(N968), .ENCLK(net10466), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 clk_gate_mem_reg_7_ ( 
        .CLK(clk), .EN(N959), .ENCLK(net10471), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 clk_gate_mem_reg_8_ ( 
        .CLK(clk), .EN(N950), .ENCLK(net10476), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 clk_gate_mem_reg_9_ ( 
        .CLK(clk), .EN(N941), .ENCLK(net10481), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 clk_gate_mem_reg_10_ ( 
        .CLK(clk), .EN(N932), .ENCLK(net10486), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 clk_gate_mem_reg_11_ ( 
        .CLK(clk), .EN(N923), .ENCLK(net10491), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 clk_gate_mem_reg_12_ ( 
        .CLK(clk), .EN(N914), .ENCLK(net10496), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 clk_gate_mem_reg_13_ ( 
        .CLK(clk), .EN(N905), .ENCLK(net10501), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 clk_gate_mem_reg_14_ ( 
        .CLK(clk), .EN(N896), .ENCLK(net10506), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 clk_gate_mem_reg_15_ ( 
        .CLK(clk), .EN(N887), .ENCLK(net10511), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 clk_gate_mem_reg_16_ ( 
        .CLK(clk), .EN(N878), .ENCLK(net10516), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 clk_gate_mem_reg_17_ ( 
        .CLK(clk), .EN(N869), .ENCLK(net10521), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 clk_gate_mem_reg_18_ ( 
        .CLK(clk), .EN(N860), .ENCLK(net10526), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 clk_gate_mem_reg_19_ ( 
        .CLK(clk), .EN(N851), .ENCLK(net10531), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 clk_gate_mem_reg_20_ ( 
        .CLK(clk), .EN(N842), .ENCLK(net10536), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 clk_gate_mem_reg_21_ ( 
        .CLK(clk), .EN(N833), .ENCLK(net10541), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 clk_gate_mem_reg_22_ ( 
        .CLK(clk), .EN(N824), .ENCLK(net10546), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 clk_gate_mem_reg_23_ ( 
        .CLK(clk), .EN(N815), .ENCLK(net10551), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 clk_gate_mem_reg_24_ ( 
        .CLK(clk), .EN(N806), .ENCLK(net10556), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 clk_gate_mem_reg_25_ ( 
        .CLK(clk), .EN(N797), .ENCLK(net10561), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 clk_gate_mem_reg_26_ ( 
        .CLK(clk), .EN(N788), .ENCLK(net10566), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 clk_gate_mem_reg_27_ ( 
        .CLK(clk), .EN(N779), .ENCLK(net10571), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 clk_gate_mem_reg_28_ ( 
        .CLK(clk), .EN(N770), .ENCLK(net10576), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 clk_gate_mem_reg_29_ ( 
        .CLK(clk), .EN(N761), .ENCLK(net10581), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 clk_gate_mem_reg_30_ ( 
        .CLK(clk), .EN(N752), .ENCLK(net10586), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 clk_gate_mem_reg_31_ ( 
        .CLK(clk), .EN(N743), .ENCLK(net10591), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 clk_gate_mem_reg_32_ ( 
        .CLK(clk), .EN(N734), .ENCLK(net10596), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 clk_gate_mem_reg_33_ ( 
        .CLK(clk), .EN(N733), .ENCLK(net10601), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 clk_gate_pshptr_reg ( 
        .CLK(clk), .EN(N1053), .ENCLK(net10606), .TE(test_se) );
  SDFFQX1 mem_reg_33__7_ ( .D(fifowdat[7]), .SIN(mem_33__6_), .SMC(test_se), 
        .C(net10601), .Q(mem_33__7_) );
  SDFFQX1 mem_reg_32__7_ ( .D(N742), .SIN(mem_32__6_), .SMC(test_se), .C(
        net10596), .Q(mem_32__7_) );
  SDFFQX1 mem_reg_31__7_ ( .D(N751), .SIN(mem_31__6_), .SMC(test_se), .C(
        net10591), .Q(mem_31__7_) );
  SDFFQX1 mem_reg_30__7_ ( .D(N760), .SIN(mem_30__6_), .SMC(test_se), .C(
        net10586), .Q(mem_30__7_) );
  SDFFQX1 mem_reg_29__7_ ( .D(N769), .SIN(mem_29__6_), .SMC(test_se), .C(
        net10581), .Q(mem_29__7_) );
  SDFFQX1 mem_reg_28__7_ ( .D(N778), .SIN(mem_28__6_), .SMC(test_se), .C(
        net10576), .Q(mem_28__7_) );
  SDFFQX1 mem_reg_33__6_ ( .D(fifowdat[6]), .SIN(mem_33__5_), .SMC(test_se), 
        .C(net10601), .Q(mem_33__6_) );
  SDFFQX1 mem_reg_32__6_ ( .D(N741), .SIN(mem_32__5_), .SMC(test_se), .C(
        net10596), .Q(mem_32__6_) );
  SDFFQX1 mem_reg_31__6_ ( .D(N750), .SIN(mem_31__5_), .SMC(test_se), .C(
        net10591), .Q(mem_31__6_) );
  SDFFQX1 mem_reg_30__6_ ( .D(N759), .SIN(mem_30__5_), .SMC(test_se), .C(
        net10586), .Q(mem_30__6_) );
  SDFFQX1 mem_reg_29__6_ ( .D(N768), .SIN(mem_29__5_), .SMC(test_se), .C(
        net10581), .Q(mem_29__6_) );
  SDFFQX1 mem_reg_28__6_ ( .D(N777), .SIN(mem_28__5_), .SMC(test_se), .C(
        net10576), .Q(mem_28__6_) );
  SDFFQX1 mem_reg_33__5_ ( .D(fifowdat[5]), .SIN(mem_33__4_), .SMC(test_se), 
        .C(net10601), .Q(mem_33__5_) );
  SDFFQX1 mem_reg_32__5_ ( .D(N740), .SIN(mem_32__4_), .SMC(test_se), .C(
        net10596), .Q(mem_32__5_) );
  SDFFQX1 mem_reg_31__5_ ( .D(N749), .SIN(mem_31__4_), .SMC(test_se), .C(
        net10591), .Q(mem_31__5_) );
  SDFFQX1 mem_reg_30__5_ ( .D(N758), .SIN(mem_30__4_), .SMC(test_se), .C(
        net10586), .Q(mem_30__5_) );
  SDFFQX1 mem_reg_29__5_ ( .D(N767), .SIN(mem_29__4_), .SMC(test_se), .C(
        net10581), .Q(mem_29__5_) );
  SDFFQX1 mem_reg_28__5_ ( .D(N776), .SIN(mem_28__4_), .SMC(test_se), .C(
        net10576), .Q(mem_28__5_) );
  SDFFQX1 mem_reg_33__4_ ( .D(fifowdat[4]), .SIN(mem_33__3_), .SMC(test_se), 
        .C(net10601), .Q(mem_33__4_) );
  SDFFQX1 mem_reg_32__4_ ( .D(N739), .SIN(mem_32__3_), .SMC(test_se), .C(
        net10596), .Q(mem_32__4_) );
  SDFFQX1 mem_reg_31__4_ ( .D(N748), .SIN(mem_31__3_), .SMC(test_se), .C(
        net10591), .Q(mem_31__4_) );
  SDFFQX1 mem_reg_30__4_ ( .D(N757), .SIN(mem_30__3_), .SMC(test_se), .C(
        net10586), .Q(mem_30__4_) );
  SDFFQX1 mem_reg_29__4_ ( .D(N766), .SIN(mem_29__3_), .SMC(test_se), .C(
        net10581), .Q(mem_29__4_) );
  SDFFQX1 mem_reg_28__4_ ( .D(N775), .SIN(mem_28__3_), .SMC(test_se), .C(
        net10576), .Q(mem_28__4_) );
  SDFFQX1 mem_reg_33__3_ ( .D(fifowdat[3]), .SIN(mem_33__2_), .SMC(test_se), 
        .C(net10601), .Q(mem_33__3_) );
  SDFFQX1 mem_reg_32__3_ ( .D(N738), .SIN(mem_32__2_), .SMC(test_se), .C(
        net10596), .Q(mem_32__3_) );
  SDFFQX1 mem_reg_31__3_ ( .D(N747), .SIN(mem_31__2_), .SMC(test_se), .C(
        net10591), .Q(mem_31__3_) );
  SDFFQX1 mem_reg_30__3_ ( .D(N756), .SIN(mem_30__2_), .SMC(test_se), .C(
        net10586), .Q(mem_30__3_) );
  SDFFQX1 mem_reg_29__3_ ( .D(N765), .SIN(mem_29__2_), .SMC(test_se), .C(
        net10581), .Q(mem_29__3_) );
  SDFFQX1 mem_reg_28__3_ ( .D(N774), .SIN(mem_28__2_), .SMC(test_se), .C(
        net10576), .Q(mem_28__3_) );
  SDFFQX1 mem_reg_33__2_ ( .D(fifowdat[2]), .SIN(mem_33__1_), .SMC(test_se), 
        .C(net10601), .Q(mem_33__2_) );
  SDFFQX1 mem_reg_32__2_ ( .D(N737), .SIN(mem_32__1_), .SMC(test_se), .C(
        net10596), .Q(mem_32__2_) );
  SDFFQX1 mem_reg_31__2_ ( .D(N746), .SIN(mem_31__1_), .SMC(test_se), .C(
        net10591), .Q(mem_31__2_) );
  SDFFQX1 mem_reg_30__2_ ( .D(N755), .SIN(mem_30__1_), .SMC(test_se), .C(
        net10586), .Q(mem_30__2_) );
  SDFFQX1 mem_reg_29__2_ ( .D(N764), .SIN(mem_29__1_), .SMC(test_se), .C(
        net10581), .Q(mem_29__2_) );
  SDFFQX1 mem_reg_28__2_ ( .D(N773), .SIN(mem_28__1_), .SMC(test_se), .C(
        net10576), .Q(mem_28__2_) );
  SDFFQX1 mem_reg_33__1_ ( .D(fifowdat[1]), .SIN(mem_33__0_), .SMC(test_se), 
        .C(net10601), .Q(mem_33__1_) );
  SDFFQX1 mem_reg_32__1_ ( .D(N736), .SIN(mem_32__0_), .SMC(test_se), .C(
        net10596), .Q(mem_32__1_) );
  SDFFQX1 mem_reg_31__1_ ( .D(N745), .SIN(mem_31__0_), .SMC(test_se), .C(
        net10591), .Q(mem_31__1_) );
  SDFFQX1 mem_reg_30__1_ ( .D(N754), .SIN(mem_30__0_), .SMC(test_se), .C(
        net10586), .Q(mem_30__1_) );
  SDFFQX1 mem_reg_29__1_ ( .D(N763), .SIN(mem_29__0_), .SMC(test_se), .C(
        net10581), .Q(mem_29__1_) );
  SDFFQX1 mem_reg_28__1_ ( .D(N772), .SIN(mem_28__0_), .SMC(test_se), .C(
        net10576), .Q(mem_28__1_) );
  SDFFQX1 mem_reg_33__0_ ( .D(fifowdat[0]), .SIN(mem_32__7_), .SMC(test_se), 
        .C(net10601), .Q(mem_33__0_) );
  SDFFQX1 mem_reg_32__0_ ( .D(N735), .SIN(mem_31__7_), .SMC(test_se), .C(
        net10596), .Q(mem_32__0_) );
  SDFFQX1 mem_reg_31__0_ ( .D(N744), .SIN(mem_30__7_), .SMC(test_se), .C(
        net10591), .Q(mem_31__0_) );
  SDFFQX1 mem_reg_30__0_ ( .D(N753), .SIN(mem_29__7_), .SMC(test_se), .C(
        net10586), .Q(mem_30__0_) );
  SDFFQX1 mem_reg_29__0_ ( .D(N762), .SIN(mem_28__7_), .SMC(test_se), .C(
        net10581), .Q(mem_29__0_) );
  SDFFQX1 mem_reg_28__0_ ( .D(N771), .SIN(mem_27__7_), .SMC(test_se), .C(
        net10576), .Q(mem_28__0_) );
  SDFFQX1 mem_reg_27__7_ ( .D(N787), .SIN(mem_27__6_), .SMC(test_se), .C(
        net10571), .Q(mem_27__7_) );
  SDFFQX1 mem_reg_26__7_ ( .D(N796), .SIN(mem_26__6_), .SMC(test_se), .C(
        net10566), .Q(mem_26__7_) );
  SDFFQX1 mem_reg_25__7_ ( .D(N805), .SIN(mem_25__6_), .SMC(test_se), .C(
        net10561), .Q(mem_25__7_) );
  SDFFQX1 mem_reg_24__7_ ( .D(N814), .SIN(mem_24__6_), .SMC(test_se), .C(
        net10556), .Q(mem_24__7_) );
  SDFFQX1 mem_reg_23__7_ ( .D(N823), .SIN(mem_23__6_), .SMC(test_se), .C(
        net10551), .Q(mem_23__7_) );
  SDFFQX1 mem_reg_22__7_ ( .D(N832), .SIN(mem_22__6_), .SMC(test_se), .C(
        net10546), .Q(mem_22__7_) );
  SDFFQX1 mem_reg_21__7_ ( .D(N841), .SIN(mem_21__6_), .SMC(test_se), .C(
        net10541), .Q(mem_21__7_) );
  SDFFQX1 mem_reg_20__7_ ( .D(N850), .SIN(mem_20__6_), .SMC(test_se), .C(
        net10536), .Q(mem_20__7_) );
  SDFFQX1 mem_reg_19__7_ ( .D(N859), .SIN(mem_19__6_), .SMC(test_se), .C(
        net10531), .Q(mem_19__7_) );
  SDFFQX1 mem_reg_18__7_ ( .D(N868), .SIN(mem_18__6_), .SMC(test_se), .C(
        net10526), .Q(mem_18__7_) );
  SDFFQX1 mem_reg_17__7_ ( .D(N877), .SIN(mem_17__6_), .SMC(test_se), .C(
        net10521), .Q(mem_17__7_) );
  SDFFQX1 mem_reg_16__7_ ( .D(N886), .SIN(mem_16__6_), .SMC(test_se), .C(
        net10516), .Q(mem_16__7_) );
  SDFFQX1 mem_reg_15__7_ ( .D(N895), .SIN(mem_15__6_), .SMC(test_se), .C(
        net10511), .Q(mem_15__7_) );
  SDFFQX1 mem_reg_14__7_ ( .D(N904), .SIN(mem_14__6_), .SMC(test_se), .C(
        net10506), .Q(mem_14__7_) );
  SDFFQX1 mem_reg_13__7_ ( .D(N913), .SIN(mem_13__6_), .SMC(test_se), .C(
        net10501), .Q(mem_13__7_) );
  SDFFQX1 mem_reg_12__7_ ( .D(N922), .SIN(mem_12__6_), .SMC(test_se), .C(
        net10496), .Q(mem_12__7_) );
  SDFFQX1 mem_reg_11__7_ ( .D(N931), .SIN(mem_11__6_), .SMC(test_se), .C(
        net10491), .Q(mem_11__7_) );
  SDFFQX1 mem_reg_10__7_ ( .D(N940), .SIN(mem_10__6_), .SMC(test_se), .C(
        net10486), .Q(mem_10__7_) );
  SDFFQX1 mem_reg_9__7_ ( .D(N949), .SIN(mem_9__6_), .SMC(test_se), .C(
        net10481), .Q(mem_9__7_) );
  SDFFQX1 mem_reg_8__7_ ( .D(N958), .SIN(mem_8__6_), .SMC(test_se), .C(
        net10476), .Q(mem_8__7_) );
  SDFFQX1 mem_reg_27__6_ ( .D(N786), .SIN(mem_27__5_), .SMC(test_se), .C(
        net10571), .Q(mem_27__6_) );
  SDFFQX1 mem_reg_26__6_ ( .D(N795), .SIN(mem_26__5_), .SMC(test_se), .C(
        net10566), .Q(mem_26__6_) );
  SDFFQX1 mem_reg_25__6_ ( .D(N804), .SIN(mem_25__5_), .SMC(test_se), .C(
        net10561), .Q(mem_25__6_) );
  SDFFQX1 mem_reg_24__6_ ( .D(N813), .SIN(mem_24__5_), .SMC(test_se), .C(
        net10556), .Q(mem_24__6_) );
  SDFFQX1 mem_reg_23__6_ ( .D(N822), .SIN(mem_23__5_), .SMC(test_se), .C(
        net10551), .Q(mem_23__6_) );
  SDFFQX1 mem_reg_22__6_ ( .D(N831), .SIN(mem_22__5_), .SMC(test_se), .C(
        net10546), .Q(mem_22__6_) );
  SDFFQX1 mem_reg_21__6_ ( .D(N840), .SIN(mem_21__5_), .SMC(test_se), .C(
        net10541), .Q(mem_21__6_) );
  SDFFQX1 mem_reg_20__6_ ( .D(N849), .SIN(mem_20__5_), .SMC(test_se), .C(
        net10536), .Q(mem_20__6_) );
  SDFFQX1 mem_reg_19__6_ ( .D(N858), .SIN(mem_19__5_), .SMC(test_se), .C(
        net10531), .Q(mem_19__6_) );
  SDFFQX1 mem_reg_18__6_ ( .D(N867), .SIN(mem_18__5_), .SMC(test_se), .C(
        net10526), .Q(mem_18__6_) );
  SDFFQX1 mem_reg_17__6_ ( .D(N876), .SIN(mem_17__5_), .SMC(test_se), .C(
        net10521), .Q(mem_17__6_) );
  SDFFQX1 mem_reg_16__6_ ( .D(N885), .SIN(mem_16__5_), .SMC(test_se), .C(
        net10516), .Q(mem_16__6_) );
  SDFFQX1 mem_reg_15__6_ ( .D(N894), .SIN(mem_15__5_), .SMC(test_se), .C(
        net10511), .Q(mem_15__6_) );
  SDFFQX1 mem_reg_14__6_ ( .D(N903), .SIN(mem_14__5_), .SMC(test_se), .C(
        net10506), .Q(mem_14__6_) );
  SDFFQX1 mem_reg_13__6_ ( .D(N912), .SIN(mem_13__5_), .SMC(test_se), .C(
        net10501), .Q(mem_13__6_) );
  SDFFQX1 mem_reg_12__6_ ( .D(N921), .SIN(mem_12__5_), .SMC(test_se), .C(
        net10496), .Q(mem_12__6_) );
  SDFFQX1 mem_reg_11__6_ ( .D(N930), .SIN(mem_11__5_), .SMC(test_se), .C(
        net10491), .Q(mem_11__6_) );
  SDFFQX1 mem_reg_10__6_ ( .D(N939), .SIN(mem_10__5_), .SMC(test_se), .C(
        net10486), .Q(mem_10__6_) );
  SDFFQX1 mem_reg_9__6_ ( .D(N948), .SIN(mem_9__5_), .SMC(test_se), .C(
        net10481), .Q(mem_9__6_) );
  SDFFQX1 mem_reg_8__6_ ( .D(N957), .SIN(mem_8__5_), .SMC(test_se), .C(
        net10476), .Q(mem_8__6_) );
  SDFFQX1 mem_reg_27__5_ ( .D(N785), .SIN(mem_27__4_), .SMC(test_se), .C(
        net10571), .Q(mem_27__5_) );
  SDFFQX1 mem_reg_26__5_ ( .D(N794), .SIN(mem_26__4_), .SMC(test_se), .C(
        net10566), .Q(mem_26__5_) );
  SDFFQX1 mem_reg_25__5_ ( .D(N803), .SIN(mem_25__4_), .SMC(test_se), .C(
        net10561), .Q(mem_25__5_) );
  SDFFQX1 mem_reg_24__5_ ( .D(N812), .SIN(mem_24__4_), .SMC(test_se), .C(
        net10556), .Q(mem_24__5_) );
  SDFFQX1 mem_reg_23__5_ ( .D(N821), .SIN(mem_23__4_), .SMC(test_se), .C(
        net10551), .Q(mem_23__5_) );
  SDFFQX1 mem_reg_22__5_ ( .D(N830), .SIN(mem_22__4_), .SMC(test_se), .C(
        net10546), .Q(mem_22__5_) );
  SDFFQX1 mem_reg_21__5_ ( .D(N839), .SIN(mem_21__4_), .SMC(test_se), .C(
        net10541), .Q(mem_21__5_) );
  SDFFQX1 mem_reg_20__5_ ( .D(N848), .SIN(mem_20__4_), .SMC(test_se), .C(
        net10536), .Q(mem_20__5_) );
  SDFFQX1 mem_reg_19__5_ ( .D(N857), .SIN(mem_19__4_), .SMC(test_se), .C(
        net10531), .Q(mem_19__5_) );
  SDFFQX1 mem_reg_18__5_ ( .D(N866), .SIN(mem_18__4_), .SMC(test_se), .C(
        net10526), .Q(mem_18__5_) );
  SDFFQX1 mem_reg_17__5_ ( .D(N875), .SIN(mem_17__4_), .SMC(test_se), .C(
        net10521), .Q(mem_17__5_) );
  SDFFQX1 mem_reg_16__5_ ( .D(N884), .SIN(mem_16__4_), .SMC(test_se), .C(
        net10516), .Q(mem_16__5_) );
  SDFFQX1 mem_reg_15__5_ ( .D(N893), .SIN(mem_15__4_), .SMC(test_se), .C(
        net10511), .Q(mem_15__5_) );
  SDFFQX1 mem_reg_14__5_ ( .D(N902), .SIN(mem_14__4_), .SMC(test_se), .C(
        net10506), .Q(mem_14__5_) );
  SDFFQX1 mem_reg_13__5_ ( .D(N911), .SIN(mem_13__4_), .SMC(test_se), .C(
        net10501), .Q(mem_13__5_) );
  SDFFQX1 mem_reg_12__5_ ( .D(N920), .SIN(mem_12__4_), .SMC(test_se), .C(
        net10496), .Q(mem_12__5_) );
  SDFFQX1 mem_reg_11__5_ ( .D(N929), .SIN(mem_11__4_), .SMC(test_se), .C(
        net10491), .Q(mem_11__5_) );
  SDFFQX1 mem_reg_10__5_ ( .D(N938), .SIN(mem_10__4_), .SMC(test_se), .C(
        net10486), .Q(mem_10__5_) );
  SDFFQX1 mem_reg_9__5_ ( .D(N947), .SIN(mem_9__4_), .SMC(test_se), .C(
        net10481), .Q(mem_9__5_) );
  SDFFQX1 mem_reg_8__5_ ( .D(N956), .SIN(mem_8__4_), .SMC(test_se), .C(
        net10476), .Q(mem_8__5_) );
  SDFFQX1 mem_reg_27__4_ ( .D(N784), .SIN(mem_27__3_), .SMC(test_se), .C(
        net10571), .Q(mem_27__4_) );
  SDFFQX1 mem_reg_26__4_ ( .D(N793), .SIN(mem_26__3_), .SMC(test_se), .C(
        net10566), .Q(mem_26__4_) );
  SDFFQX1 mem_reg_25__4_ ( .D(N802), .SIN(mem_25__3_), .SMC(test_se), .C(
        net10561), .Q(mem_25__4_) );
  SDFFQX1 mem_reg_24__4_ ( .D(N811), .SIN(mem_24__3_), .SMC(test_se), .C(
        net10556), .Q(mem_24__4_) );
  SDFFQX1 mem_reg_23__4_ ( .D(N820), .SIN(mem_23__3_), .SMC(test_se), .C(
        net10551), .Q(mem_23__4_) );
  SDFFQX1 mem_reg_22__4_ ( .D(N829), .SIN(mem_22__3_), .SMC(test_se), .C(
        net10546), .Q(mem_22__4_) );
  SDFFQX1 mem_reg_21__4_ ( .D(N838), .SIN(mem_21__3_), .SMC(test_se), .C(
        net10541), .Q(mem_21__4_) );
  SDFFQX1 mem_reg_20__4_ ( .D(N847), .SIN(mem_20__3_), .SMC(test_se), .C(
        net10536), .Q(mem_20__4_) );
  SDFFQX1 mem_reg_19__4_ ( .D(N856), .SIN(mem_19__3_), .SMC(test_se), .C(
        net10531), .Q(mem_19__4_) );
  SDFFQX1 mem_reg_18__4_ ( .D(N865), .SIN(mem_18__3_), .SMC(test_se), .C(
        net10526), .Q(mem_18__4_) );
  SDFFQX1 mem_reg_17__4_ ( .D(N874), .SIN(mem_17__3_), .SMC(test_se), .C(
        net10521), .Q(mem_17__4_) );
  SDFFQX1 mem_reg_16__4_ ( .D(N883), .SIN(mem_16__3_), .SMC(test_se), .C(
        net10516), .Q(mem_16__4_) );
  SDFFQX1 mem_reg_15__4_ ( .D(N892), .SIN(mem_15__3_), .SMC(test_se), .C(
        net10511), .Q(mem_15__4_) );
  SDFFQX1 mem_reg_14__4_ ( .D(N901), .SIN(mem_14__3_), .SMC(test_se), .C(
        net10506), .Q(mem_14__4_) );
  SDFFQX1 mem_reg_13__4_ ( .D(N910), .SIN(mem_13__3_), .SMC(test_se), .C(
        net10501), .Q(mem_13__4_) );
  SDFFQX1 mem_reg_12__4_ ( .D(N919), .SIN(mem_12__3_), .SMC(test_se), .C(
        net10496), .Q(mem_12__4_) );
  SDFFQX1 mem_reg_11__4_ ( .D(N928), .SIN(mem_11__3_), .SMC(test_se), .C(
        net10491), .Q(mem_11__4_) );
  SDFFQX1 mem_reg_10__4_ ( .D(N937), .SIN(mem_10__3_), .SMC(test_se), .C(
        net10486), .Q(mem_10__4_) );
  SDFFQX1 mem_reg_9__4_ ( .D(N946), .SIN(mem_9__3_), .SMC(test_se), .C(
        net10481), .Q(mem_9__4_) );
  SDFFQX1 mem_reg_8__4_ ( .D(N955), .SIN(mem_8__3_), .SMC(test_se), .C(
        net10476), .Q(mem_8__4_) );
  SDFFQX1 mem_reg_27__3_ ( .D(N783), .SIN(mem_27__2_), .SMC(test_se), .C(
        net10571), .Q(mem_27__3_) );
  SDFFQX1 mem_reg_26__3_ ( .D(N792), .SIN(mem_26__2_), .SMC(test_se), .C(
        net10566), .Q(mem_26__3_) );
  SDFFQX1 mem_reg_25__3_ ( .D(N801), .SIN(mem_25__2_), .SMC(test_se), .C(
        net10561), .Q(mem_25__3_) );
  SDFFQX1 mem_reg_24__3_ ( .D(N810), .SIN(mem_24__2_), .SMC(test_se), .C(
        net10556), .Q(mem_24__3_) );
  SDFFQX1 mem_reg_23__3_ ( .D(N819), .SIN(mem_23__2_), .SMC(test_se), .C(
        net10551), .Q(mem_23__3_) );
  SDFFQX1 mem_reg_22__3_ ( .D(N828), .SIN(mem_22__2_), .SMC(test_se), .C(
        net10546), .Q(mem_22__3_) );
  SDFFQX1 mem_reg_21__3_ ( .D(N837), .SIN(mem_21__2_), .SMC(test_se), .C(
        net10541), .Q(mem_21__3_) );
  SDFFQX1 mem_reg_20__3_ ( .D(N846), .SIN(mem_20__2_), .SMC(test_se), .C(
        net10536), .Q(mem_20__3_) );
  SDFFQX1 mem_reg_19__3_ ( .D(N855), .SIN(mem_19__2_), .SMC(test_se), .C(
        net10531), .Q(mem_19__3_) );
  SDFFQX1 mem_reg_18__3_ ( .D(N864), .SIN(mem_18__2_), .SMC(test_se), .C(
        net10526), .Q(mem_18__3_) );
  SDFFQX1 mem_reg_17__3_ ( .D(N873), .SIN(mem_17__2_), .SMC(test_se), .C(
        net10521), .Q(mem_17__3_) );
  SDFFQX1 mem_reg_16__3_ ( .D(N882), .SIN(mem_16__2_), .SMC(test_se), .C(
        net10516), .Q(mem_16__3_) );
  SDFFQX1 mem_reg_15__3_ ( .D(N891), .SIN(mem_15__2_), .SMC(test_se), .C(
        net10511), .Q(mem_15__3_) );
  SDFFQX1 mem_reg_14__3_ ( .D(N900), .SIN(mem_14__2_), .SMC(test_se), .C(
        net10506), .Q(mem_14__3_) );
  SDFFQX1 mem_reg_13__3_ ( .D(N909), .SIN(mem_13__2_), .SMC(test_se), .C(
        net10501), .Q(mem_13__3_) );
  SDFFQX1 mem_reg_12__3_ ( .D(N918), .SIN(mem_12__2_), .SMC(test_se), .C(
        net10496), .Q(mem_12__3_) );
  SDFFQX1 mem_reg_11__3_ ( .D(N927), .SIN(mem_11__2_), .SMC(test_se), .C(
        net10491), .Q(mem_11__3_) );
  SDFFQX1 mem_reg_10__3_ ( .D(N936), .SIN(mem_10__2_), .SMC(test_se), .C(
        net10486), .Q(mem_10__3_) );
  SDFFQX1 mem_reg_9__3_ ( .D(N945), .SIN(mem_9__2_), .SMC(test_se), .C(
        net10481), .Q(mem_9__3_) );
  SDFFQX1 mem_reg_8__3_ ( .D(N954), .SIN(mem_8__2_), .SMC(test_se), .C(
        net10476), .Q(mem_8__3_) );
  SDFFQX1 mem_reg_27__2_ ( .D(N782), .SIN(mem_27__1_), .SMC(test_se), .C(
        net10571), .Q(mem_27__2_) );
  SDFFQX1 mem_reg_26__2_ ( .D(N791), .SIN(mem_26__1_), .SMC(test_se), .C(
        net10566), .Q(mem_26__2_) );
  SDFFQX1 mem_reg_25__2_ ( .D(N800), .SIN(mem_25__1_), .SMC(test_se), .C(
        net10561), .Q(mem_25__2_) );
  SDFFQX1 mem_reg_24__2_ ( .D(N809), .SIN(mem_24__1_), .SMC(test_se), .C(
        net10556), .Q(mem_24__2_) );
  SDFFQX1 mem_reg_23__2_ ( .D(N818), .SIN(mem_23__1_), .SMC(test_se), .C(
        net10551), .Q(mem_23__2_) );
  SDFFQX1 mem_reg_22__2_ ( .D(N827), .SIN(mem_22__1_), .SMC(test_se), .C(
        net10546), .Q(mem_22__2_) );
  SDFFQX1 mem_reg_21__2_ ( .D(N836), .SIN(mem_21__1_), .SMC(test_se), .C(
        net10541), .Q(mem_21__2_) );
  SDFFQX1 mem_reg_20__2_ ( .D(N845), .SIN(mem_20__1_), .SMC(test_se), .C(
        net10536), .Q(mem_20__2_) );
  SDFFQX1 mem_reg_19__2_ ( .D(N854), .SIN(mem_19__1_), .SMC(test_se), .C(
        net10531), .Q(mem_19__2_) );
  SDFFQX1 mem_reg_18__2_ ( .D(N863), .SIN(mem_18__1_), .SMC(test_se), .C(
        net10526), .Q(mem_18__2_) );
  SDFFQX1 mem_reg_17__2_ ( .D(N872), .SIN(mem_17__1_), .SMC(test_se), .C(
        net10521), .Q(mem_17__2_) );
  SDFFQX1 mem_reg_16__2_ ( .D(N881), .SIN(mem_16__1_), .SMC(test_se), .C(
        net10516), .Q(mem_16__2_) );
  SDFFQX1 mem_reg_15__2_ ( .D(N890), .SIN(mem_15__1_), .SMC(test_se), .C(
        net10511), .Q(mem_15__2_) );
  SDFFQX1 mem_reg_14__2_ ( .D(N899), .SIN(mem_14__1_), .SMC(test_se), .C(
        net10506), .Q(mem_14__2_) );
  SDFFQX1 mem_reg_13__2_ ( .D(N908), .SIN(mem_13__1_), .SMC(test_se), .C(
        net10501), .Q(mem_13__2_) );
  SDFFQX1 mem_reg_12__2_ ( .D(N917), .SIN(mem_12__1_), .SMC(test_se), .C(
        net10496), .Q(mem_12__2_) );
  SDFFQX1 mem_reg_11__2_ ( .D(N926), .SIN(mem_11__1_), .SMC(test_se), .C(
        net10491), .Q(mem_11__2_) );
  SDFFQX1 mem_reg_10__2_ ( .D(N935), .SIN(mem_10__1_), .SMC(test_se), .C(
        net10486), .Q(mem_10__2_) );
  SDFFQX1 mem_reg_9__2_ ( .D(N944), .SIN(mem_9__1_), .SMC(test_se), .C(
        net10481), .Q(mem_9__2_) );
  SDFFQX1 mem_reg_8__2_ ( .D(N953), .SIN(mem_8__1_), .SMC(test_se), .C(
        net10476), .Q(mem_8__2_) );
  SDFFQX1 mem_reg_27__1_ ( .D(N781), .SIN(mem_27__0_), .SMC(test_se), .C(
        net10571), .Q(mem_27__1_) );
  SDFFQX1 mem_reg_26__1_ ( .D(N790), .SIN(mem_26__0_), .SMC(test_se), .C(
        net10566), .Q(mem_26__1_) );
  SDFFQX1 mem_reg_25__1_ ( .D(N799), .SIN(mem_25__0_), .SMC(test_se), .C(
        net10561), .Q(mem_25__1_) );
  SDFFQX1 mem_reg_24__1_ ( .D(N808), .SIN(mem_24__0_), .SMC(test_se), .C(
        net10556), .Q(mem_24__1_) );
  SDFFQX1 mem_reg_23__1_ ( .D(N817), .SIN(mem_23__0_), .SMC(test_se), .C(
        net10551), .Q(mem_23__1_) );
  SDFFQX1 mem_reg_22__1_ ( .D(N826), .SIN(mem_22__0_), .SMC(test_se), .C(
        net10546), .Q(mem_22__1_) );
  SDFFQX1 mem_reg_21__1_ ( .D(N835), .SIN(mem_21__0_), .SMC(test_se), .C(
        net10541), .Q(mem_21__1_) );
  SDFFQX1 mem_reg_20__1_ ( .D(N844), .SIN(mem_20__0_), .SMC(test_se), .C(
        net10536), .Q(mem_20__1_) );
  SDFFQX1 mem_reg_19__1_ ( .D(N853), .SIN(mem_19__0_), .SMC(test_se), .C(
        net10531), .Q(mem_19__1_) );
  SDFFQX1 mem_reg_18__1_ ( .D(N862), .SIN(mem_18__0_), .SMC(test_se), .C(
        net10526), .Q(mem_18__1_) );
  SDFFQX1 mem_reg_17__1_ ( .D(N871), .SIN(mem_17__0_), .SMC(test_se), .C(
        net10521), .Q(mem_17__1_) );
  SDFFQX1 mem_reg_16__1_ ( .D(N880), .SIN(mem_16__0_), .SMC(test_se), .C(
        net10516), .Q(mem_16__1_) );
  SDFFQX1 mem_reg_15__1_ ( .D(N889), .SIN(mem_15__0_), .SMC(test_se), .C(
        net10511), .Q(mem_15__1_) );
  SDFFQX1 mem_reg_14__1_ ( .D(N898), .SIN(mem_14__0_), .SMC(test_se), .C(
        net10506), .Q(mem_14__1_) );
  SDFFQX1 mem_reg_13__1_ ( .D(N907), .SIN(mem_13__0_), .SMC(test_se), .C(
        net10501), .Q(mem_13__1_) );
  SDFFQX1 mem_reg_12__1_ ( .D(N916), .SIN(mem_12__0_), .SMC(test_se), .C(
        net10496), .Q(mem_12__1_) );
  SDFFQX1 mem_reg_11__1_ ( .D(N925), .SIN(mem_11__0_), .SMC(test_se), .C(
        net10491), .Q(mem_11__1_) );
  SDFFQX1 mem_reg_10__1_ ( .D(N934), .SIN(mem_10__0_), .SMC(test_se), .C(
        net10486), .Q(mem_10__1_) );
  SDFFQX1 mem_reg_9__1_ ( .D(N943), .SIN(mem_9__0_), .SMC(test_se), .C(
        net10481), .Q(mem_9__1_) );
  SDFFQX1 mem_reg_8__1_ ( .D(N952), .SIN(mem_8__0_), .SMC(test_se), .C(
        net10476), .Q(mem_8__1_) );
  SDFFQX1 mem_reg_27__0_ ( .D(N780), .SIN(mem_26__7_), .SMC(test_se), .C(
        net10571), .Q(mem_27__0_) );
  SDFFQX1 mem_reg_26__0_ ( .D(N789), .SIN(mem_25__7_), .SMC(test_se), .C(
        net10566), .Q(mem_26__0_) );
  SDFFQX1 mem_reg_25__0_ ( .D(N798), .SIN(mem_24__7_), .SMC(test_se), .C(
        net10561), .Q(mem_25__0_) );
  SDFFQX1 mem_reg_24__0_ ( .D(N807), .SIN(mem_23__7_), .SMC(test_se), .C(
        net10556), .Q(mem_24__0_) );
  SDFFQX1 mem_reg_23__0_ ( .D(N816), .SIN(mem_22__7_), .SMC(test_se), .C(
        net10551), .Q(mem_23__0_) );
  SDFFQX1 mem_reg_22__0_ ( .D(N825), .SIN(mem_21__7_), .SMC(test_se), .C(
        net10546), .Q(mem_22__0_) );
  SDFFQX1 mem_reg_21__0_ ( .D(N834), .SIN(mem_20__7_), .SMC(test_se), .C(
        net10541), .Q(mem_21__0_) );
  SDFFQX1 mem_reg_20__0_ ( .D(N843), .SIN(mem_19__7_), .SMC(test_se), .C(
        net10536), .Q(mem_20__0_) );
  SDFFQX1 mem_reg_19__0_ ( .D(N852), .SIN(mem_18__7_), .SMC(test_se), .C(
        net10531), .Q(mem_19__0_) );
  SDFFQX1 mem_reg_18__0_ ( .D(N861), .SIN(mem_17__7_), .SMC(test_se), .C(
        net10526), .Q(mem_18__0_) );
  SDFFQX1 mem_reg_17__0_ ( .D(N870), .SIN(mem_16__7_), .SMC(test_se), .C(
        net10521), .Q(mem_17__0_) );
  SDFFQX1 mem_reg_16__0_ ( .D(N879), .SIN(mem_15__7_), .SMC(test_se), .C(
        net10516), .Q(mem_16__0_) );
  SDFFQX1 mem_reg_15__0_ ( .D(N888), .SIN(mem_14__7_), .SMC(test_se), .C(
        net10511), .Q(mem_15__0_) );
  SDFFQX1 mem_reg_14__0_ ( .D(N897), .SIN(mem_13__7_), .SMC(test_se), .C(
        net10506), .Q(mem_14__0_) );
  SDFFQX1 mem_reg_13__0_ ( .D(N906), .SIN(mem_12__7_), .SMC(test_se), .C(
        net10501), .Q(mem_13__0_) );
  SDFFQX1 mem_reg_12__0_ ( .D(N915), .SIN(mem_11__7_), .SMC(test_se), .C(
        net10496), .Q(mem_12__0_) );
  SDFFQX1 mem_reg_11__0_ ( .D(N924), .SIN(mem_10__7_), .SMC(test_se), .C(
        net10491), .Q(mem_11__0_) );
  SDFFQX1 mem_reg_10__0_ ( .D(N933), .SIN(mem_9__7_), .SMC(test_se), .C(
        net10486), .Q(mem_10__0_) );
  SDFFQX1 mem_reg_9__0_ ( .D(N942), .SIN(mem_8__7_), .SMC(test_se), .C(
        net10481), .Q(mem_9__0_) );
  SDFFQX1 mem_reg_8__0_ ( .D(N951), .SIN(dat_7_1[55]), .SMC(test_se), .C(
        net10476), .Q(mem_8__0_) );
  SDFFQX1 mem_reg_1__0_ ( .D(N1014), .SIN(rdat0[7]), .SMC(test_se), .C(
        net10441), .Q(dat_7_1[0]) );
  SDFFQX1 mem_reg_1__3_ ( .D(N1017), .SIN(dat_7_1[2]), .SMC(test_se), .C(
        net10441), .Q(dat_7_1[3]) );
  SDFFQX1 mem_reg_1__2_ ( .D(N1016), .SIN(dat_7_1[1]), .SMC(test_se), .C(
        net10441), .Q(dat_7_1[2]) );
  SDFFQX1 mem_reg_1__1_ ( .D(N1015), .SIN(dat_7_1[0]), .SMC(test_se), .C(
        net10441), .Q(dat_7_1[1]) );
  SDFFQX1 locked_reg ( .D(ps_locked), .SIN(test_si), .SMC(test_se), .C(clk), 
        .Q(locked) );
  SDFFQX1 mem_reg_7__7_ ( .D(N967), .SIN(dat_7_1[54]), .SMC(test_se), .C(
        net10471), .Q(dat_7_1[55]) );
  SDFFQX1 mem_reg_7__5_ ( .D(N965), .SIN(dat_7_1[52]), .SMC(test_se), .C(
        net10471), .Q(dat_7_1[53]) );
  SDFFQX1 mem_reg_6__4_ ( .D(N973), .SIN(dat_7_1[43]), .SMC(test_se), .C(
        net10466), .Q(dat_7_1[44]) );
  SDFFQX1 mem_reg_6__2_ ( .D(N971), .SIN(dat_7_1[41]), .SMC(test_se), .C(
        net10466), .Q(dat_7_1[42]) );
  SDFFQX1 mem_reg_6__7_ ( .D(N976), .SIN(dat_7_1[46]), .SMC(test_se), .C(
        net10466), .Q(dat_7_1[47]) );
  SDFFQX1 mem_reg_7__6_ ( .D(N966), .SIN(dat_7_1[53]), .SMC(test_se), .C(
        net10471), .Q(dat_7_1[54]) );
  SDFFQX1 mem_reg_6__6_ ( .D(N975), .SIN(dat_7_1[45]), .SMC(test_se), .C(
        net10466), .Q(dat_7_1[46]) );
  SDFFQX1 mem_reg_6__5_ ( .D(N974), .SIN(dat_7_1[44]), .SMC(test_se), .C(
        net10466), .Q(dat_7_1[45]) );
  SDFFQX1 mem_reg_6__3_ ( .D(N972), .SIN(dat_7_1[42]), .SMC(test_se), .C(
        net10466), .Q(dat_7_1[43]) );
  SDFFQX1 mem_reg_7__1_ ( .D(N961), .SIN(dat_7_1[48]), .SMC(test_se), .C(
        net10471), .Q(dat_7_1[49]) );
  SDFFQX1 mem_reg_6__1_ ( .D(N970), .SIN(dat_7_1[40]), .SMC(test_se), .C(
        net10466), .Q(dat_7_1[41]) );
  SDFFQX1 mem_reg_7__0_ ( .D(N960), .SIN(dat_7_1[47]), .SMC(test_se), .C(
        net10471), .Q(dat_7_1[48]) );
  SDFFQX1 mem_reg_2__6_ ( .D(N1011), .SIN(dat_7_1[13]), .SMC(test_se), .C(
        net10446), .Q(dat_7_1[14]) );
  SDFFQX1 mem_reg_4__7_ ( .D(N994), .SIN(dat_7_1[30]), .SMC(test_se), .C(
        net10456), .Q(dat_7_1[31]) );
  SDFFQX1 mem_reg_5__6_ ( .D(N984), .SIN(dat_7_1[37]), .SMC(test_se), .C(
        net10461), .Q(dat_7_1[38]) );
  SDFFQX1 mem_reg_4__4_ ( .D(N991), .SIN(dat_7_1[27]), .SMC(test_se), .C(
        net10456), .Q(dat_7_1[28]) );
  SDFFQX1 mem_reg_4__3_ ( .D(N990), .SIN(dat_7_1[26]), .SMC(test_se), .C(
        net10456), .Q(dat_7_1[27]) );
  SDFFQX1 mem_reg_5__1_ ( .D(N979), .SIN(dat_7_1[32]), .SMC(test_se), .C(
        net10461), .Q(dat_7_1[33]) );
  SDFFQX1 mem_reg_3__3_ ( .D(N999), .SIN(dat_7_1[18]), .SMC(test_se), .C(
        net10451), .Q(dat_7_1[19]) );
  SDFFQX1 mem_reg_3__2_ ( .D(N998), .SIN(dat_7_1[17]), .SMC(test_se), .C(
        net10451), .Q(dat_7_1[18]) );
  SDFFQX1 mem_reg_3__1_ ( .D(N997), .SIN(dat_7_1[16]), .SMC(test_se), .C(
        net10451), .Q(dat_7_1[17]) );
  SDFFQX1 mem_reg_2__7_ ( .D(N1012), .SIN(dat_7_1[14]), .SMC(test_se), .C(
        net10446), .Q(dat_7_1[15]) );
  SDFFQX1 mem_reg_7__4_ ( .D(N964), .SIN(dat_7_1[51]), .SMC(test_se), .C(
        net10471), .Q(dat_7_1[52]) );
  SDFFQX1 mem_reg_7__3_ ( .D(N963), .SIN(dat_7_1[50]), .SMC(test_se), .C(
        net10471), .Q(dat_7_1[51]) );
  SDFFQX1 mem_reg_7__2_ ( .D(N962), .SIN(dat_7_1[49]), .SMC(test_se), .C(
        net10471), .Q(dat_7_1[50]) );
  SDFFQX1 mem_reg_6__0_ ( .D(N969), .SIN(dat_7_1[39]), .SMC(test_se), .C(
        net10466), .Q(dat_7_1[40]) );
  SDFFQX1 mem_reg_5__7_ ( .D(N985), .SIN(dat_7_1[38]), .SMC(test_se), .C(
        net10461), .Q(dat_7_1[39]) );
  SDFFQX1 mem_reg_4__6_ ( .D(N993), .SIN(dat_7_1[29]), .SMC(test_se), .C(
        net10456), .Q(dat_7_1[30]) );
  SDFFQX1 mem_reg_5__5_ ( .D(N983), .SIN(dat_7_1[36]), .SMC(test_se), .C(
        net10461), .Q(dat_7_1[37]) );
  SDFFQX1 mem_reg_4__5_ ( .D(N992), .SIN(dat_7_1[28]), .SMC(test_se), .C(
        net10456), .Q(dat_7_1[29]) );
  SDFFQX1 mem_reg_5__4_ ( .D(N982), .SIN(dat_7_1[35]), .SMC(test_se), .C(
        net10461), .Q(dat_7_1[36]) );
  SDFFQX1 mem_reg_5__3_ ( .D(N981), .SIN(dat_7_1[34]), .SMC(test_se), .C(
        net10461), .Q(dat_7_1[35]) );
  SDFFQX1 mem_reg_5__2_ ( .D(N980), .SIN(dat_7_1[33]), .SMC(test_se), .C(
        net10461), .Q(dat_7_1[34]) );
  SDFFQX1 mem_reg_4__2_ ( .D(N989), .SIN(dat_7_1[25]), .SMC(test_se), .C(
        net10456), .Q(dat_7_1[26]) );
  SDFFQX1 mem_reg_4__1_ ( .D(N988), .SIN(dat_7_1[24]), .SMC(test_se), .C(
        net10456), .Q(dat_7_1[25]) );
  SDFFQX1 mem_reg_5__0_ ( .D(N978), .SIN(dat_7_1[31]), .SMC(test_se), .C(
        net10461), .Q(dat_7_1[32]) );
  SDFFQX1 mem_reg_4__0_ ( .D(N987), .SIN(dat_7_1[23]), .SMC(test_se), .C(
        net10456), .Q(dat_7_1[24]) );
  SDFFQX1 mem_reg_3__0_ ( .D(N996), .SIN(dat_7_1[15]), .SMC(test_se), .C(
        net10451), .Q(dat_7_1[16]) );
  SDFFQX1 mem_reg_2__5_ ( .D(N1010), .SIN(dat_7_1[12]), .SMC(test_se), .C(
        net10446), .Q(dat_7_1[13]) );
  SDFFQX1 mem_reg_1__7_ ( .D(N1021), .SIN(dat_7_1[6]), .SMC(test_se), .C(
        net10441), .Q(dat_7_1[7]) );
  SDFFQX1 mem_reg_1__6_ ( .D(N1020), .SIN(dat_7_1[5]), .SMC(test_se), .C(
        net10441), .Q(dat_7_1[6]) );
  SDFFQX1 mem_reg_1__5_ ( .D(N1019), .SIN(dat_7_1[4]), .SMC(test_se), .C(
        net10441), .Q(dat_7_1[5]) );
  SDFFQX1 mem_reg_1__4_ ( .D(N1018), .SIN(dat_7_1[3]), .SMC(test_se), .C(
        net10441), .Q(dat_7_1[4]) );
  SDFFQX1 mem_reg_3__6_ ( .D(N1002), .SIN(dat_7_1[21]), .SMC(test_se), .C(
        net10451), .Q(dat_7_1[22]) );
  SDFFQX1 mem_reg_2__3_ ( .D(N1008), .SIN(dat_7_1[10]), .SMC(test_se), .C(
        net10446), .Q(dat_7_1[11]) );
  SDFFQX1 mem_reg_3__5_ ( .D(N1001), .SIN(dat_7_1[20]), .SMC(test_se), .C(
        net10451), .Q(dat_7_1[21]) );
  SDFFQX1 mem_reg_3__4_ ( .D(N1000), .SIN(dat_7_1[19]), .SMC(test_se), .C(
        net10451), .Q(dat_7_1[20]) );
  SDFFQX1 mem_reg_2__4_ ( .D(N1009), .SIN(dat_7_1[11]), .SMC(test_se), .C(
        net10446), .Q(dat_7_1[12]) );
  SDFFQX1 mem_reg_2__2_ ( .D(N1007), .SIN(dat_7_1[9]), .SMC(test_se), .C(
        net10446), .Q(dat_7_1[10]) );
  SDFFQX1 mem_reg_3__7_ ( .D(N1003), .SIN(dat_7_1[22]), .SMC(test_se), .C(
        net10451), .Q(dat_7_1[23]) );
  SDFFQX1 mem_reg_2__1_ ( .D(N1006), .SIN(dat_7_1[8]), .SMC(test_se), .C(
        net10446), .Q(dat_7_1[9]) );
  SDFFQX1 mem_reg_2__0_ ( .D(N1005), .SIN(dat_7_1[7]), .SMC(test_se), .C(
        net10446), .Q(dat_7_1[8]) );
  SDFFQX1 mem_reg_0__7_ ( .D(N1030), .SIN(rdat0[6]), .SMC(test_se), .C(
        net10435), .Q(rdat0[7]) );
  SDFFQX1 pshptr_reg_4_ ( .D(N1058), .SIN(ptr[3]), .SMC(test_se), .C(net10606), 
        .Q(ptr[4]) );
  SDFFQX1 mem_reg_0__4_ ( .D(N1027), .SIN(rdat0[3]), .SMC(test_se), .C(
        net10435), .Q(rdat0[4]) );
  SDFFQX1 mem_reg_0__1_ ( .D(N1024), .SIN(rdat0[0]), .SMC(test_se), .C(
        net10435), .Q(rdat0[1]) );
  SDFFQX1 mem_reg_0__5_ ( .D(N1028), .SIN(rdat0[4]), .SMC(test_se), .C(
        net10435), .Q(rdat0[5]) );
  SDFFQX1 pshptr_reg_2_ ( .D(N1056), .SIN(ptr[1]), .SMC(test_se), .C(net10606), 
        .Q(ptr[2]) );
  SDFFQX1 pshptr_reg_3_ ( .D(N1057), .SIN(ptr[2]), .SMC(test_se), .C(net10606), 
        .Q(ptr[3]) );
  SDFFQX1 mem_reg_0__3_ ( .D(N1026), .SIN(rdat0[2]), .SMC(test_se), .C(
        net10435), .Q(rdat0[3]) );
  SDFFQX1 mem_reg_0__2_ ( .D(N1025), .SIN(rdat0[1]), .SMC(test_se), .C(
        net10435), .Q(rdat0[2]) );
  SDFFQX1 mem_reg_0__0_ ( .D(N1023), .SIN(locked), .SMC(test_se), .C(net10435), 
        .Q(rdat0[0]) );
  SDFFQX1 mem_reg_0__6_ ( .D(N1029), .SIN(rdat0[5]), .SMC(test_se), .C(
        net10435), .Q(rdat0[6]) );
  SDFFQX1 pshptr_reg_1_ ( .D(N1055), .SIN(ptr[0]), .SMC(test_se), .C(net10606), 
        .Q(ptr[1]) );
  SDFFQX1 pshptr_reg_0_ ( .D(N1054), .SIN(mem_33__7_), .SMC(test_se), .C(
        net10606), .Q(ptr[0]) );
  SDFFQX1 pshptr_reg_5_ ( .D(N1059), .SIN(ptr[4]), .SMC(test_se), .C(net10606), 
        .Q(ptr[5]) );
  INVX1 U3 ( .A(ptr[0]), .Y(n514) );
  INVX1 U4 ( .A(ptr[4]), .Y(n512) );
  INVX1 U5 ( .A(ptr[5]), .Y(n428) );
  INVX1 U6 ( .A(n501), .Y(n1) );
  INVX1 U7 ( .A(n535), .Y(n2) );
  AND3XL U8 ( .A(ptr[0]), .B(ptr[4]), .C(n511), .Y(half) );
  NAND43X1 U9 ( .B(ptr[3]), .C(ptr[2]), .D(ptr[1]), .A(n428), .Y(n513) );
  OR4X1 U10 ( .A(ptx_pop), .B(n508), .C(prx_psh), .D(n3), .Y(n516) );
  AOI21X1 U11 ( .B(i_lockena), .C(n60), .A(locked), .Y(n3) );
  INVX1 U12 ( .A(n299), .Y(n286) );
  INVX1 U13 ( .A(n299), .Y(n298) );
  INVX1 U14 ( .A(r_psh), .Y(n575) );
  INVX1 U15 ( .A(n299), .Y(n275) );
  INVX1 U16 ( .A(n24), .Y(n23) );
  INVX1 U17 ( .A(n24), .Y(n22) );
  INVX1 U18 ( .A(n32), .Y(n31) );
  INVX1 U19 ( .A(n32), .Y(n30) );
  INVX1 U20 ( .A(n40), .Y(n39) );
  INVX1 U21 ( .A(n40), .Y(n38) );
  INVX1 U22 ( .A(n48), .Y(n47) );
  INVX1 U23 ( .A(n48), .Y(n46) );
  INVX1 U24 ( .A(n64), .Y(n299) );
  INVX1 U25 ( .A(n464), .Y(n508) );
  NOR21XL U26 ( .B(n250), .A(n14), .Y(n252) );
  NOR21XL U27 ( .B(n264), .A(n15), .Y(n266) );
  NOR21XL U28 ( .B(n287), .A(n15), .Y(n289) );
  NOR21XL U29 ( .B(n237), .A(n15), .Y(n239) );
  NAND2X1 U30 ( .A(n575), .B(n574), .Y(n60) );
  NOR21XL U31 ( .B(n138), .A(n14), .Y(n140) );
  NOR21XL U32 ( .B(n192), .A(n15), .Y(n194) );
  NOR21XL U33 ( .B(n300), .A(n14), .Y(n302) );
  NOR21XL U34 ( .B(n312), .A(n15), .Y(n314) );
  NOR21XL U35 ( .B(n381), .A(n14), .Y(n383) );
  NOR21XL U36 ( .B(n429), .A(n13), .Y(n431) );
  NOR21XL U37 ( .B(n80), .A(n15), .Y(n84) );
  NOR21XL U38 ( .B(n114), .A(n13), .Y(n116) );
  NOR21XL U39 ( .B(n127), .A(n13), .Y(n129) );
  NOR21XL U40 ( .B(n468), .A(n13), .Y(n470) );
  NOR21XL U41 ( .B(n153), .A(n13), .Y(n155) );
  NOR21XL U42 ( .B(n276), .A(n14), .Y(n278) );
  NOR21XL U43 ( .B(n324), .A(n15), .Y(n326) );
  NOR21XL U44 ( .B(n358), .A(n14), .Y(n360) );
  NOR21XL U45 ( .B(n166), .A(n15), .Y(n168) );
  NOR21XL U46 ( .B(n205), .A(n14), .Y(n207) );
  NOR21XL U47 ( .B(n216), .A(n16), .Y(n218) );
  NOR21XL U48 ( .B(n227), .A(n15), .Y(n229) );
  NAND21X1 U49 ( .B(n462), .A(n568), .Y(n460) );
  NOR2X1 U50 ( .A(n110), .B(n16), .Y(n102) );
  INVX1 U51 ( .A(n76), .Y(n555) );
  INVX1 U52 ( .A(n32), .Y(n29) );
  INVX1 U53 ( .A(n90), .Y(n32) );
  INVX1 U54 ( .A(n40), .Y(n37) );
  INVX1 U55 ( .A(n87), .Y(n40) );
  INVX1 U56 ( .A(n48), .Y(n45) );
  INVX1 U57 ( .A(n83), .Y(n48) );
  INVX1 U58 ( .A(n24), .Y(n21) );
  INVX1 U59 ( .A(n93), .Y(n24) );
  INVX1 U60 ( .A(n56), .Y(n54) );
  INVX1 U61 ( .A(n137), .Y(n99) );
  INVX1 U62 ( .A(n203), .Y(n190) );
  INVX1 U63 ( .A(n56), .Y(n55) );
  INVX1 U64 ( .A(n137), .Y(n126) );
  INVX1 U65 ( .A(n203), .Y(n191) );
  NAND2X1 U66 ( .A(fifowdat[3]), .B(n16), .Y(n64) );
  NAND2X1 U67 ( .A(n561), .B(n572), .Y(n391) );
  INVX1 U68 ( .A(n110), .Y(n569) );
  OAI21X1 U69 ( .B(n549), .C(n573), .A(n297), .Y(N833) );
  OAI21X1 U70 ( .B(n547), .C(n573), .A(n148), .Y(N941) );
  OAI21X1 U71 ( .B(n548), .C(n18), .A(n274), .Y(N851) );
  NAND2X1 U72 ( .A(n462), .B(n464), .Y(N1053) );
  INVX1 U73 ( .A(fifowdat[3]), .Y(n311) );
  INVX1 U74 ( .A(fifowdat[3]), .Y(n356) );
  INVX1 U75 ( .A(fifowdat[3]), .Y(n357) );
  NOR21XL U76 ( .B(srstz), .A(r_fiforst), .Y(n464) );
  NOR21XL U77 ( .B(n260), .A(n9), .Y(n250) );
  NOR21XL U78 ( .B(n274), .A(n11), .Y(n264) );
  NOR21XL U79 ( .B(n297), .A(n10), .Y(n287) );
  AOI211X1 U80 ( .C(n564), .D(n559), .A(n247), .B(n565), .Y(n237) );
  NAND2X1 U81 ( .A(n559), .B(n571), .Y(n260) );
  NAND2X1 U82 ( .A(n559), .B(n567), .Y(n274) );
  NAND2X1 U83 ( .A(n559), .B(n572), .Y(n297) );
  NOR21XL U84 ( .B(n478), .A(n13), .Y(n480) );
  NOR21XL U85 ( .B(n180), .A(n15), .Y(n182) );
  NOR21XL U86 ( .B(n334), .A(n13), .Y(n336) );
  NOR21XL U87 ( .B(n345), .A(n14), .Y(n347) );
  NOR21XL U88 ( .B(n370), .A(n13), .Y(n372) );
  NOR21XL U89 ( .B(n417), .A(n14), .Y(n419) );
  NOR21XL U90 ( .B(n5), .A(n13), .Y(n66) );
  NOR21XL U91 ( .B(n394), .A(n13), .Y(n396) );
  NOR21XL U92 ( .B(n407), .A(n14), .Y(n409) );
  NOR21XL U93 ( .B(n439), .A(n440), .Y(n429) );
  NOR21XL U94 ( .B(n310), .A(n549), .Y(n300) );
  NOR21XL U95 ( .B(n148), .A(n8), .Y(n138) );
  NOR21XL U96 ( .B(n202), .A(n7), .Y(n192) );
  NOR21XL U97 ( .B(n322), .A(n559), .Y(n312) );
  NOR21XL U98 ( .B(n391), .A(n392), .Y(n381) );
  NAND21X1 U99 ( .B(n100), .A(n503), .Y(n76) );
  NAND21X1 U100 ( .B(n462), .A(n463), .Y(n461) );
  OAI21X1 U101 ( .B(n562), .C(n100), .A(n111), .Y(n110) );
  XNOR2XL U102 ( .A(n4), .B(n568), .Y(n462) );
  INVX1 U103 ( .A(n19), .Y(n15) );
  INVX1 U104 ( .A(n19), .Y(n14) );
  INVX1 U105 ( .A(n19), .Y(n13) );
  AOI21X1 U106 ( .B(n555), .C(n572), .A(n98), .Y(n80) );
  AOI21X1 U107 ( .B(n557), .C(n571), .A(n547), .Y(n153) );
  AOI21X1 U108 ( .B(n553), .C(n559), .A(n548), .Y(n276) );
  AOI21X1 U109 ( .B(n555), .C(n571), .A(n546), .Y(n468) );
  AOI21X1 U110 ( .B(n557), .C(n563), .A(n556), .Y(n127) );
  AOI21X1 U111 ( .B(n124), .C(n556), .A(n555), .Y(n114) );
  AOI21X1 U112 ( .B(n563), .C(n559), .A(n565), .Y(n227) );
  AOI21X1 U113 ( .B(n563), .C(n561), .A(n558), .Y(n324) );
  AOI21X1 U114 ( .B(n567), .C(n561), .A(n368), .Y(n358) );
  AOI211X1 U115 ( .C(n124), .D(n565), .A(n557), .B(n556), .Y(n216) );
  AND2X1 U116 ( .A(n176), .B(n177), .Y(n166) );
  AND2X1 U117 ( .A(n6), .B(n215), .Y(n205) );
  INVX1 U118 ( .A(n19), .Y(n16) );
  INVX1 U119 ( .A(n344), .Y(n561) );
  INVX1 U120 ( .A(n100), .Y(n556) );
  INVX1 U121 ( .A(n137), .Y(n78) );
  INVX1 U122 ( .A(n203), .Y(n179) );
  INVX1 U123 ( .A(n56), .Y(n53) );
  INVX1 U124 ( .A(n74), .Y(n56) );
  INVX1 U125 ( .A(n543), .Y(n547) );
  INVX1 U126 ( .A(n463), .Y(n568) );
  INVX1 U127 ( .A(n467), .Y(n445) );
  INVX1 U128 ( .A(n493), .Y(n446) );
  INVX1 U129 ( .A(n71), .Y(n137) );
  INVX1 U130 ( .A(n68), .Y(n203) );
  NAND2X1 U131 ( .A(fifowdat[4]), .B(n16), .Y(n93) );
  NAND2X1 U132 ( .A(fifowdat[5]), .B(n16), .Y(n90) );
  NAND2X1 U133 ( .A(fifowdat[6]), .B(n16), .Y(n87) );
  NAND2X1 U134 ( .A(fifowdat[7]), .B(n16), .Y(n83) );
  NAND2X1 U135 ( .A(n557), .B(n567), .Y(n176) );
  NAND2X1 U136 ( .A(n564), .B(n557), .Y(n148) );
  NAND2X1 U137 ( .A(n557), .B(n572), .Y(n202) );
  NAND21X1 U138 ( .B(n17), .A(n100), .Y(n79) );
  NAND21X1 U139 ( .B(n558), .A(n20), .Y(n323) );
  OAI21BBX1 U140 ( .A(n524), .B(n561), .C(n498), .Y(N743) );
  OAI21BBX1 U141 ( .A(n322), .B(n20), .C(n310), .Y(N824) );
  INVX1 U142 ( .A(n534), .Y(n558) );
  INVX1 U143 ( .A(n533), .Y(n549) );
  INVX1 U144 ( .A(n112), .Y(n572) );
  INVX1 U145 ( .A(n77), .Y(n567) );
  INVX1 U146 ( .A(n19), .Y(n17) );
  INVX1 U147 ( .A(n20), .Y(n18) );
  INVX1 U148 ( .A(n536), .Y(n548) );
  INVX1 U149 ( .A(n124), .Y(n524) );
  OAI21X1 U150 ( .B(n11), .C(n573), .A(n260), .Y(N860) );
  OAI21X1 U151 ( .B(n76), .C(n124), .A(n79), .Y(N959) );
  OAI21BBX1 U152 ( .A(n20), .B(n6), .C(n202), .Y(N905) );
  NAND3X1 U153 ( .A(n111), .B(n79), .C(n125), .Y(N968) );
  INVX1 U154 ( .A(r_pop), .Y(n574) );
  NAND21X1 U155 ( .B(n124), .A(n20), .Y(n125) );
  INVX1 U156 ( .A(fifowdat[4]), .Y(n25) );
  INVX1 U157 ( .A(fifowdat[4]), .Y(n26) );
  INVX1 U158 ( .A(fifowdat[4]), .Y(n27) );
  INVX1 U159 ( .A(fifowdat[6]), .Y(n41) );
  INVX1 U160 ( .A(fifowdat[6]), .Y(n42) );
  INVX1 U161 ( .A(fifowdat[7]), .Y(n49) );
  INVX1 U162 ( .A(fifowdat[7]), .Y(n50) );
  INVX1 U163 ( .A(fifowdat[6]), .Y(n43) );
  INVX1 U164 ( .A(fifowdat[7]), .Y(n51) );
  INVX1 U165 ( .A(n63), .Y(fifowdat[3]) );
  INVX1 U166 ( .A(fifowdat[5]), .Y(n33) );
  INVX1 U167 ( .A(fifowdat[5]), .Y(n34) );
  INVX1 U168 ( .A(fifowdat[5]), .Y(n35) );
  INVX1 U169 ( .A(n248), .Y(n559) );
  AOI21BBXL U170 ( .B(n554), .C(n575), .A(prx_psh), .Y(n4) );
  INVX1 U171 ( .A(n4), .Y(fifopsh) );
  NAND21X1 U172 ( .B(n1), .A(n565), .Y(n100) );
  NAND21X1 U173 ( .B(n523), .A(n566), .Y(n344) );
  OR2X1 U174 ( .A(n447), .B(n461), .Y(n467) );
  NAND2X1 U175 ( .A(n495), .B(n525), .Y(n440) );
  AO21X1 U176 ( .B(n545), .C(n542), .A(n541), .Y(n543) );
  OAI21BBX1 U177 ( .A(n525), .B(n523), .C(n440), .Y(n417) );
  NAND21X1 U178 ( .B(n523), .A(n525), .Y(n496) );
  NAND21X1 U179 ( .B(n248), .A(n560), .Y(n310) );
  OR2X1 U180 ( .A(n427), .B(n460), .Y(n493) );
  AOI21X1 U181 ( .B(n555), .C(n553), .A(n520), .Y(n5) );
  AOI21X1 U182 ( .B(n565), .C(n113), .A(n556), .Y(n6) );
  OAI21AX1 U183 ( .B(n554), .C(n574), .A(ptx_pop), .Y(n463) );
  AOI21X1 U184 ( .B(n555), .C(n567), .A(n488), .Y(n478) );
  AOI21X1 U185 ( .B(n553), .C(n557), .A(n165), .Y(n180) );
  AOI21X1 U186 ( .B(n571), .C(n561), .A(n355), .Y(n345) );
  AOI211X1 U187 ( .C(n564), .D(n561), .A(n558), .B(n550), .Y(n334) );
  AOI211X1 U188 ( .C(n553), .D(n561), .A(n551), .B(n558), .Y(n370) );
  AND2X1 U189 ( .A(n12), .B(n404), .Y(n394) );
  AO21X1 U190 ( .B(n540), .C(n545), .A(n541), .Y(n177) );
  MUX2X1 U191 ( .D0(n451), .D1(n450), .S(n537), .Y(N1058) );
  OAI22X1 U192 ( .A(n465), .B(n461), .C(n449), .D(n460), .Y(n450) );
  AO21X1 U193 ( .B(n446), .C(n545), .A(n445), .Y(n451) );
  AND2X1 U194 ( .A(n448), .B(n545), .Y(n449) );
  NAND21X1 U195 ( .B(n344), .A(n560), .Y(n404) );
  NAND21X1 U196 ( .B(n150), .A(n560), .Y(n215) );
  OR2X1 U197 ( .A(n262), .B(n496), .Y(n439) );
  INVX1 U198 ( .A(n150), .Y(n557) );
  INVX1 U199 ( .A(n502), .Y(n565) );
  INVX1 U200 ( .A(n523), .Y(n503) );
  AOI21X1 U201 ( .B(n545), .C(n552), .A(n6), .Y(n7) );
  AOI21X1 U202 ( .B(n545), .C(n544), .A(n543), .Y(n8) );
  INVX1 U203 ( .A(n526), .Y(n407) );
  OAI211X1 U204 ( .C(n525), .D(n524), .A(n344), .B(n534), .Y(n526) );
  INVX1 U205 ( .A(n165), .Y(n541) );
  INVX1 U206 ( .A(n505), .Y(n546) );
  NAND21X1 U207 ( .B(n542), .A(n520), .Y(n505) );
  INVX1 U208 ( .A(n573), .Y(n19) );
  NAND2X1 U209 ( .A(fifowdat[0]), .B(n16), .Y(n74) );
  NAND2X1 U210 ( .A(fifowdat[1]), .B(n16), .Y(n71) );
  NAND2X1 U211 ( .A(fifowdat[2]), .B(n16), .Y(n68) );
  NAND2X1 U212 ( .A(n560), .B(n555), .Y(n111) );
  NAND21X1 U213 ( .B(n113), .A(n544), .Y(n124) );
  NAND21X1 U214 ( .B(n525), .A(n500), .Y(n534) );
  NAND21X1 U215 ( .B(n535), .A(n540), .Y(n77) );
  AO21X1 U216 ( .B(n537), .C(n535), .A(n534), .Y(n536) );
  AO21X1 U217 ( .B(n537), .C(n562), .A(n534), .Y(n533) );
  NAND21X1 U218 ( .B(n544), .A(n546), .Y(n522) );
  NAND21X1 U219 ( .B(n17), .A(n525), .Y(n498) );
  AOI21X1 U220 ( .B(n537), .C(n542), .A(n536), .Y(n9) );
  NAND21X1 U221 ( .B(n542), .A(n552), .Y(n112) );
  INVX1 U222 ( .A(n538), .Y(n247) );
  NAND21X1 U223 ( .B(n545), .A(n550), .Y(n538) );
  NAND21X1 U224 ( .B(n17), .A(n502), .Y(n226) );
  AO21X1 U225 ( .B(n551), .C(n529), .A(n558), .Y(n368) );
  AO21X1 U226 ( .B(n537), .C(n524), .A(n534), .Y(n322) );
  AOI21X1 U227 ( .B(n552), .C(n566), .A(n12), .Y(n392) );
  INVX1 U228 ( .A(n506), .Y(n507) );
  OAI211X1 U229 ( .C(n76), .D(n262), .A(n20), .B(n522), .Y(n506) );
  INVX1 U230 ( .A(n529), .Y(n540) );
  INVX1 U231 ( .A(n178), .Y(n571) );
  INVX1 U232 ( .A(n570), .Y(n553) );
  INVX1 U233 ( .A(n151), .Y(n563) );
  INVX1 U234 ( .A(n262), .Y(n564) );
  AOI21X1 U235 ( .B(n537), .C(n552), .A(n533), .Y(n10) );
  AOI21X1 U236 ( .B(n537), .C(n540), .A(n536), .Y(n11) );
  INVX1 U237 ( .A(n500), .Y(n566) );
  OAI32X1 U238 ( .A(n544), .B(empty), .C(n461), .D(n452), .E(n460), .Y(N1054)
         );
  XOR2X1 U239 ( .A(n544), .B(full), .Y(n452) );
  INVX1 U240 ( .A(n113), .Y(n562) );
  OAI221X1 U241 ( .A(n76), .B(n112), .C(n17), .D(n113), .E(n79), .Y(N977) );
  INVX1 U242 ( .A(n447), .Y(n465) );
  OAI22X1 U243 ( .A(n17), .B(n520), .C(n76), .D(n77), .Y(N995) );
  OAI22X1 U244 ( .A(n488), .B(n18), .C(n76), .D(n178), .Y(N1004) );
  OAI22X1 U245 ( .A(n546), .B(n18), .C(n76), .D(n262), .Y(N1013) );
  OAI22X1 U246 ( .A(n496), .B(n495), .C(n440), .D(n18), .Y(N734) );
  OAI22X1 U247 ( .A(n570), .B(n344), .C(n392), .D(n18), .Y(N770) );
  OAI22X1 U248 ( .A(n178), .B(n344), .C(n368), .D(n18), .Y(N788) );
  OAI22X1 U249 ( .A(n262), .B(n344), .C(n355), .D(n18), .Y(N797) );
  OAI22X1 U250 ( .A(n570), .B(n248), .C(n10), .D(n18), .Y(N842) );
  OAI22X1 U251 ( .A(n262), .B(n248), .C(n9), .D(n17), .Y(N869) );
  OAI22X1 U252 ( .A(n570), .B(n150), .C(n7), .D(n17), .Y(N914) );
  OAI22X1 U253 ( .A(n150), .B(n151), .C(n8), .D(n17), .Y(N950) );
  OAI22X1 U254 ( .A(n570), .B(n76), .C(n98), .D(n17), .Y(N986) );
  OAI22AX1 U255 ( .D(n522), .C(n18), .A(n76), .B(n151), .Y(N1022) );
  OAI22X1 U256 ( .A(n77), .B(n344), .C(n551), .D(n323), .Y(N779) );
  OAI22X1 U257 ( .A(n151), .B(n344), .C(n550), .D(n323), .Y(N806) );
  OAI22X1 U258 ( .A(n151), .B(n248), .C(n247), .D(n226), .Y(N878) );
  NOR3XL U259 ( .A(n552), .B(n562), .C(n100), .Y(n98) );
  OAI21X1 U260 ( .B(n124), .C(n248), .A(n323), .Y(N815) );
  OAI21X1 U261 ( .B(n124), .C(n150), .A(n226), .Y(N887) );
  OAI21X1 U262 ( .B(n17), .C(n165), .A(n176), .Y(N923) );
  INVX1 U263 ( .A(n406), .Y(n457) );
  NAND21X1 U264 ( .B(full), .A(n540), .Y(n406) );
  INVX1 U265 ( .A(n573), .Y(n20) );
  INVX1 U266 ( .A(n427), .Y(n448) );
  OAI211X1 U267 ( .C(n125), .D(n500), .A(n404), .B(n498), .Y(N752) );
  OAI21BBX1 U268 ( .A(n20), .B(n12), .C(n391), .Y(N761) );
  INVX1 U269 ( .A(n456), .Y(n441) );
  ENOX1 U270 ( .A(n150), .B(n178), .C(n177), .D(n20), .Y(N932) );
  INVX1 U271 ( .A(n91), .Y(fifowdat[4]) );
  INVX1 U272 ( .A(n85), .Y(fifowdat[6]) );
  INVX1 U273 ( .A(n81), .Y(fifowdat[7]) );
  MUX2IX1 U274 ( .D0(r_wdat[3]), .D1(prx_wdat[3]), .S(prx_psh), .Y(n63) );
  INVX1 U275 ( .A(n88), .Y(fifowdat[5]) );
  INVX1 U276 ( .A(fifowdat[0]), .Y(n57) );
  INVX1 U277 ( .A(fifowdat[0]), .Y(n59) );
  INVX1 U278 ( .A(fifowdat[1]), .Y(n149) );
  INVX1 U279 ( .A(fifowdat[1]), .Y(n152) );
  INVX1 U280 ( .A(fifowdat[2]), .Y(n204) );
  INVX1 U281 ( .A(fifowdat[2]), .Y(n249) );
  INVX1 U282 ( .A(fifowdat[0]), .Y(n61) );
  INVX1 U283 ( .A(fifowdat[1]), .Y(n163) );
  INVX1 U284 ( .A(fifowdat[2]), .Y(n261) );
  INVX1 U285 ( .A(n515), .Y(one) );
  NAND32X1 U286 ( .B(n514), .C(n513), .A(n512), .Y(n515) );
  NOR3XL U287 ( .A(n577), .B(n554), .C(n58), .Y(txreq) );
  INVX1 U288 ( .A(n519), .Y(n554) );
  NAND32X1 U289 ( .B(n523), .C(n499), .A(n501), .Y(n248) );
  NAND21X1 U290 ( .B(n4), .A(n494), .Y(n523) );
  NAND32X1 U291 ( .B(n535), .C(n542), .A(n521), .Y(n151) );
  NAND21X1 U292 ( .B(n537), .A(n531), .Y(n502) );
  NAND32X1 U293 ( .B(n502), .C(n501), .A(n503), .Y(n150) );
  AO21X1 U294 ( .B(n565), .C(n539), .A(n556), .Y(n165) );
  NAND32X1 U295 ( .B(n151), .C(n545), .A(n499), .Y(n495) );
  NOR21XL U296 ( .B(n519), .A(n518), .Y(ffack[0]) );
  NOR21XL U297 ( .B(n58), .A(n517), .Y(n518) );
  AND2XL U298 ( .A(one), .B(r_pop), .Y(n517) );
  NAND21X1 U299 ( .B(n568), .A(n510), .Y(n573) );
  INVX1 U300 ( .A(n530), .Y(n542) );
  INVX1 U301 ( .A(n539), .Y(n535) );
  INVX1 U302 ( .A(n501), .Y(n545) );
  INVX1 U303 ( .A(n499), .Y(n537) );
  NAND21X1 U304 ( .B(n444), .A(n467), .Y(N1057) );
  MUX2X1 U305 ( .D0(n446), .D1(n443), .S(n545), .Y(n444) );
  OAI22X1 U306 ( .A(n448), .B(n460), .C(n442), .D(n461), .Y(n443) );
  AND2X1 U307 ( .A(n441), .B(n539), .Y(n442) );
  INVX1 U308 ( .A(n504), .Y(n520) );
  NAND21X1 U309 ( .B(n100), .A(n539), .Y(n504) );
  OAI221X1 U310 ( .A(n500), .B(n493), .C(n502), .D(n467), .E(n466), .Y(N1059)
         );
  GEN2XL U311 ( .D(n465), .E(n499), .C(n461), .B(n460), .A(n531), .Y(n466) );
  AO2222XL U312 ( .A(r_pop), .B(empty), .C(r_psh), .D(full), .E(n577), .F(n576), .G(n554), .H(n60), .Y(ffack[1]) );
  NAND21X1 U313 ( .B(n501), .A(n537), .Y(n500) );
  NAND21X1 U314 ( .B(n2), .A(n542), .Y(n113) );
  NAND32X1 U315 ( .B(n535), .C(n521), .A(n530), .Y(n262) );
  NAND32X1 U316 ( .B(n542), .C(n539), .A(n521), .Y(n570) );
  NAND32X1 U317 ( .B(n542), .C(empty), .A(n521), .Y(n456) );
  NAND21X1 U318 ( .B(n521), .A(n542), .Y(n529) );
  NAND32X1 U319 ( .B(n535), .C(n530), .A(n521), .Y(n178) );
  NAND21X1 U320 ( .B(n539), .A(n457), .Y(n427) );
  INVX1 U321 ( .A(n497), .Y(n560) );
  NAND21X1 U322 ( .B(n113), .A(n521), .Y(n497) );
  NAND32X1 U323 ( .B(n545), .C(n456), .A(n539), .Y(n447) );
  INVX1 U324 ( .A(n527), .Y(n552) );
  NAND21X1 U325 ( .B(n539), .A(n544), .Y(n527) );
  INVX1 U326 ( .A(n521), .Y(n544) );
  INVX1 U327 ( .A(n531), .Y(n525) );
  AO21X1 U328 ( .B(n551), .C(n530), .A(n558), .Y(n355) );
  INVX1 U329 ( .A(n532), .Y(n550) );
  NAND21X1 U330 ( .B(n151), .A(n531), .Y(n532) );
  AND2X1 U331 ( .A(n369), .B(n556), .Y(n488) );
  AND2X1 U332 ( .A(n529), .B(n539), .Y(n369) );
  AOI21X1 U333 ( .B(n113), .C(n531), .A(n558), .Y(n12) );
  INVX1 U334 ( .A(n528), .Y(n551) );
  NAND21X1 U335 ( .B(n535), .A(n531), .Y(n528) );
  OAI22X1 U336 ( .A(n459), .B(n461), .C(n458), .D(n460), .Y(N1056) );
  XOR2X1 U337 ( .A(n456), .B(n535), .Y(n459) );
  OA22X1 U338 ( .A(n457), .B(n539), .C(n77), .D(full), .Y(n458) );
  OAI22X1 U339 ( .A(n455), .B(n461), .C(n454), .D(n460), .Y(N1055) );
  AND2X1 U340 ( .A(n456), .B(n529), .Y(n455) );
  XOR2X1 U341 ( .A(n530), .B(n453), .Y(n454) );
  AND2X1 U342 ( .A(n544), .B(n494), .Y(n453) );
  OAI31XL U343 ( .A(n494), .B(n4), .C(n18), .D(n439), .Y(N733) );
  OAI211X1 U344 ( .C(n125), .D(n501), .A(n215), .B(n226), .Y(N896) );
  INVX1 U345 ( .A(n58), .Y(n576) );
  INVX1 U346 ( .A(n516), .Y(ps_locked) );
  AND2X1 U347 ( .A(n510), .B(n509), .Y(obsd) );
  INVX1 U348 ( .A(srstz), .Y(n509) );
  MUX2IX1 U349 ( .D0(r_wdat[4]), .D1(prx_wdat[4]), .S(prx_psh), .Y(n91) );
  MUX2IX1 U350 ( .D0(r_wdat[6]), .D1(prx_wdat[6]), .S(prx_psh), .Y(n85) );
  MUX2IX1 U351 ( .D0(r_wdat[7]), .D1(prx_wdat[7]), .S(prx_psh), .Y(n81) );
  MUX2IX1 U352 ( .D0(r_wdat[5]), .D1(prx_wdat[5]), .S(prx_psh), .Y(n88) );
  INVX1 U353 ( .A(n494), .Y(full) );
  INVX1 U354 ( .A(n510), .Y(empty) );
  INVX1 U355 ( .A(n73), .Y(fifowdat[0]) );
  INVX1 U356 ( .A(n70), .Y(fifowdat[1]) );
  INVX1 U357 ( .A(n67), .Y(fifowdat[2]) );
  INVX1 U358 ( .A(n513), .Y(n511) );
  NAND21X1 U359 ( .B(r_unlock), .A(n516), .Y(n519) );
  OAI211X1 U360 ( .C(n237), .D(n59), .A(n246), .B(n54), .Y(N879) );
  NAND2X1 U361 ( .A(mem_17__0_), .B(n239), .Y(n246) );
  OAI211X1 U362 ( .C(n250), .D(n59), .A(n259), .B(n54), .Y(N870) );
  NAND2X1 U363 ( .A(mem_18__0_), .B(n252), .Y(n259) );
  OAI211X1 U364 ( .C(n264), .D(n59), .A(n273), .B(n54), .Y(N861) );
  NAND2X1 U365 ( .A(mem_19__0_), .B(n266), .Y(n273) );
  OAI211X1 U366 ( .C(n287), .D(n59), .A(n296), .B(n54), .Y(N843) );
  NAND2X1 U367 ( .A(mem_21__0_), .B(n289), .Y(n296) );
  OAI211X1 U368 ( .C(n237), .D(n152), .A(n245), .B(n99), .Y(N880) );
  NAND2X1 U369 ( .A(mem_17__1_), .B(n239), .Y(n245) );
  OAI211X1 U370 ( .C(n250), .D(n152), .A(n258), .B(n99), .Y(N871) );
  NAND2X1 U371 ( .A(mem_18__1_), .B(n252), .Y(n258) );
  OAI211X1 U372 ( .C(n264), .D(n152), .A(n272), .B(n99), .Y(N862) );
  NAND2X1 U373 ( .A(mem_19__1_), .B(n266), .Y(n272) );
  OAI211X1 U374 ( .C(n287), .D(n152), .A(n295), .B(n126), .Y(N844) );
  NAND2X1 U375 ( .A(mem_21__1_), .B(n289), .Y(n295) );
  OAI211X1 U376 ( .C(n237), .D(n249), .A(n244), .B(n190), .Y(N881) );
  NAND2X1 U377 ( .A(mem_17__2_), .B(n239), .Y(n244) );
  OAI211X1 U378 ( .C(n250), .D(n249), .A(n257), .B(n190), .Y(N872) );
  NAND2X1 U379 ( .A(mem_18__2_), .B(n252), .Y(n257) );
  OAI211X1 U380 ( .C(n264), .D(n249), .A(n271), .B(n190), .Y(N863) );
  NAND2X1 U381 ( .A(mem_19__2_), .B(n266), .Y(n271) );
  OAI211X1 U382 ( .C(n287), .D(n249), .A(n294), .B(n191), .Y(N845) );
  NAND2X1 U383 ( .A(mem_21__2_), .B(n289), .Y(n294) );
  OAI211X1 U384 ( .C(n237), .D(n356), .A(n243), .B(n286), .Y(N882) );
  NAND2X1 U385 ( .A(mem_17__3_), .B(n239), .Y(n243) );
  OAI211X1 U386 ( .C(n250), .D(n356), .A(n256), .B(n286), .Y(N873) );
  NAND2X1 U387 ( .A(mem_18__3_), .B(n252), .Y(n256) );
  OAI211X1 U388 ( .C(n264), .D(n356), .A(n270), .B(n286), .Y(N864) );
  NAND2X1 U389 ( .A(mem_19__3_), .B(n266), .Y(n270) );
  OAI211X1 U390 ( .C(n287), .D(n356), .A(n293), .B(n298), .Y(N846) );
  NAND2X1 U391 ( .A(mem_21__3_), .B(n289), .Y(n293) );
  OAI211X1 U392 ( .C(n237), .D(n26), .A(n242), .B(n22), .Y(N883) );
  NAND2X1 U393 ( .A(mem_17__4_), .B(n239), .Y(n242) );
  OAI211X1 U394 ( .C(n250), .D(n26), .A(n255), .B(n22), .Y(N874) );
  NAND2X1 U395 ( .A(mem_18__4_), .B(n252), .Y(n255) );
  OAI211X1 U396 ( .C(n264), .D(n26), .A(n269), .B(n22), .Y(N865) );
  NAND2X1 U397 ( .A(mem_19__4_), .B(n266), .Y(n269) );
  OAI211X1 U398 ( .C(n287), .D(n26), .A(n292), .B(n22), .Y(N847) );
  NAND2X1 U399 ( .A(mem_21__4_), .B(n289), .Y(n292) );
  OAI211X1 U400 ( .C(n237), .D(n34), .A(n241), .B(n30), .Y(N884) );
  NAND2X1 U401 ( .A(mem_17__5_), .B(n239), .Y(n241) );
  OAI211X1 U402 ( .C(n250), .D(n34), .A(n254), .B(n30), .Y(N875) );
  NAND2X1 U403 ( .A(mem_18__5_), .B(n252), .Y(n254) );
  OAI211X1 U404 ( .C(n264), .D(n34), .A(n268), .B(n30), .Y(N866) );
  NAND2X1 U405 ( .A(mem_19__5_), .B(n266), .Y(n268) );
  OAI211X1 U406 ( .C(n287), .D(n34), .A(n291), .B(n30), .Y(N848) );
  NAND2X1 U407 ( .A(mem_21__5_), .B(n289), .Y(n291) );
  OAI211X1 U408 ( .C(n237), .D(n42), .A(n240), .B(n38), .Y(N885) );
  NAND2X1 U409 ( .A(mem_17__6_), .B(n239), .Y(n240) );
  OAI211X1 U410 ( .C(n250), .D(n42), .A(n253), .B(n38), .Y(N876) );
  NAND2X1 U411 ( .A(mem_18__6_), .B(n252), .Y(n253) );
  OAI211X1 U412 ( .C(n264), .D(n42), .A(n267), .B(n38), .Y(N867) );
  NAND2X1 U413 ( .A(mem_19__6_), .B(n266), .Y(n267) );
  OAI211X1 U414 ( .C(n287), .D(n42), .A(n290), .B(n38), .Y(N849) );
  NAND2X1 U415 ( .A(mem_21__6_), .B(n289), .Y(n290) );
  OAI211X1 U416 ( .C(n237), .D(n50), .A(n238), .B(n46), .Y(N886) );
  NAND2X1 U417 ( .A(mem_17__7_), .B(n239), .Y(n238) );
  OAI211X1 U418 ( .C(n250), .D(n50), .A(n251), .B(n46), .Y(N877) );
  NAND2X1 U419 ( .A(mem_18__7_), .B(n252), .Y(n251) );
  OAI211X1 U420 ( .C(n264), .D(n50), .A(n265), .B(n46), .Y(N868) );
  NAND2X1 U421 ( .A(mem_19__7_), .B(n266), .Y(n265) );
  OAI211X1 U422 ( .C(n287), .D(n50), .A(n288), .B(n46), .Y(N850) );
  NAND2X1 U423 ( .A(mem_21__7_), .B(n289), .Y(n288) );
  NAND21XL U424 ( .B(n508), .A(ptr[2]), .Y(n539) );
  NAND21XL U425 ( .B(n508), .A(ptr[5]), .Y(n531) );
  NAND21XL U426 ( .B(n508), .A(ptr[1]), .Y(n530) );
  NAND21XL U427 ( .B(n508), .A(ptr[3]), .Y(n501) );
  NAND21XL U428 ( .B(n508), .A(ptr[4]), .Y(n499) );
  OAI211X1 U429 ( .C(n468), .D(n25), .A(n21), .B(n473), .Y(N1018) );
  NAND2X1 U430 ( .A(dat_7_1[12]), .B(n470), .Y(n473) );
  OAI211X1 U431 ( .C(n468), .D(n33), .A(n29), .B(n472), .Y(N1019) );
  NAND2X1 U432 ( .A(dat_7_1[13]), .B(n470), .Y(n472) );
  OAI211X1 U433 ( .C(n468), .D(n41), .A(n37), .B(n471), .Y(N1020) );
  NAND2X1 U434 ( .A(dat_7_1[14]), .B(n470), .Y(n471) );
  OAI211X1 U435 ( .C(n468), .D(n49), .A(n45), .B(n469), .Y(N1021) );
  NAND2X1 U436 ( .A(dat_7_1[15]), .B(n470), .Y(n469) );
  OAI211X1 U437 ( .C(n5), .D(n57), .A(n53), .B(n75), .Y(N996) );
  NAND2X1 U438 ( .A(dat_7_1[24]), .B(n66), .Y(n75) );
  OAI211X1 U439 ( .C(n5), .D(n149), .A(n78), .B(n72), .Y(N997) );
  NAND2X1 U440 ( .A(dat_7_1[25]), .B(n66), .Y(n72) );
  OAI211X1 U441 ( .C(n5), .D(n204), .A(n179), .B(n69), .Y(N998) );
  NAND2X1 U442 ( .A(dat_7_1[26]), .B(n66), .Y(n69) );
  OAI211X1 U443 ( .C(n5), .D(n311), .A(n275), .B(n65), .Y(N999) );
  NAND2X1 U444 ( .A(dat_7_1[27]), .B(n66), .Y(n65) );
  OAI211X1 U445 ( .C(n80), .D(n57), .A(n97), .B(n53), .Y(N987) );
  NAND2X1 U446 ( .A(dat_7_1[32]), .B(n84), .Y(n97) );
  OAI211X1 U447 ( .C(n569), .D(n57), .A(n109), .B(n53), .Y(N978) );
  NAND2X1 U448 ( .A(dat_7_1[40]), .B(n102), .Y(n109) );
  OAI211X1 U449 ( .C(n80), .D(n149), .A(n96), .B(n78), .Y(N988) );
  NAND2X1 U450 ( .A(dat_7_1[33]), .B(n84), .Y(n96) );
  OAI211X1 U451 ( .C(n569), .D(n149), .A(n108), .B(n78), .Y(N979) );
  NAND2X1 U452 ( .A(dat_7_1[41]), .B(n102), .Y(n108) );
  OAI211X1 U453 ( .C(n80), .D(n204), .A(n95), .B(n179), .Y(N989) );
  NAND2X1 U454 ( .A(dat_7_1[34]), .B(n84), .Y(n95) );
  OAI211X1 U455 ( .C(n569), .D(n204), .A(n107), .B(n179), .Y(N980) );
  NAND2X1 U456 ( .A(dat_7_1[42]), .B(n102), .Y(n107) );
  OAI211X1 U457 ( .C(n80), .D(n311), .A(n94), .B(n275), .Y(N990) );
  NAND2X1 U458 ( .A(dat_7_1[35]), .B(n84), .Y(n94) );
  OAI211X1 U459 ( .C(n569), .D(n311), .A(n106), .B(n275), .Y(N981) );
  NAND2X1 U460 ( .A(dat_7_1[43]), .B(n102), .Y(n106) );
  OAI211X1 U461 ( .C(n80), .D(n25), .A(n92), .B(n93), .Y(N991) );
  NAND2X1 U462 ( .A(dat_7_1[36]), .B(n84), .Y(n92) );
  OAI211X1 U463 ( .C(n569), .D(n25), .A(n105), .B(n93), .Y(N982) );
  NAND2X1 U464 ( .A(dat_7_1[44]), .B(n102), .Y(n105) );
  OAI211X1 U465 ( .C(n80), .D(n33), .A(n89), .B(n90), .Y(N992) );
  NAND2X1 U466 ( .A(dat_7_1[37]), .B(n84), .Y(n89) );
  OAI211X1 U467 ( .C(n569), .D(n33), .A(n104), .B(n90), .Y(N983) );
  NAND2X1 U468 ( .A(dat_7_1[45]), .B(n102), .Y(n104) );
  OAI211X1 U469 ( .C(n80), .D(n41), .A(n86), .B(n87), .Y(N993) );
  NAND2X1 U470 ( .A(dat_7_1[38]), .B(n84), .Y(n86) );
  OAI211X1 U471 ( .C(n569), .D(n41), .A(n103), .B(n87), .Y(N984) );
  NAND2X1 U472 ( .A(dat_7_1[46]), .B(n102), .Y(n103) );
  OAI211X1 U473 ( .C(n80), .D(n49), .A(n82), .B(n83), .Y(N994) );
  NAND2X1 U474 ( .A(dat_7_1[39]), .B(n84), .Y(n82) );
  OAI211X1 U475 ( .C(n569), .D(n49), .A(n101), .B(n83), .Y(N985) );
  NAND2X1 U476 ( .A(dat_7_1[47]), .B(n102), .Y(n101) );
  OAI211X1 U477 ( .C(n114), .D(n57), .A(n123), .B(n53), .Y(N969) );
  NAND2X1 U478 ( .A(dat_7_1[48]), .B(n116), .Y(n123) );
  OAI211X1 U479 ( .C(n127), .D(n57), .A(n136), .B(n53), .Y(N960) );
  NAND2X1 U480 ( .A(mem_8__0_), .B(n129), .Y(n136) );
  OAI211X1 U481 ( .C(n114), .D(n149), .A(n122), .B(n78), .Y(N970) );
  NAND2X1 U482 ( .A(dat_7_1[49]), .B(n116), .Y(n122) );
  OAI211X1 U483 ( .C(n127), .D(n149), .A(n135), .B(n78), .Y(N961) );
  NAND2X1 U484 ( .A(mem_8__1_), .B(n129), .Y(n135) );
  OAI211X1 U485 ( .C(n114), .D(n311), .A(n120), .B(n275), .Y(N972) );
  NAND2X1 U486 ( .A(dat_7_1[51]), .B(n116), .Y(n120) );
  OAI211X1 U487 ( .C(n114), .D(n33), .A(n118), .B(n31), .Y(N974) );
  NAND2X1 U488 ( .A(dat_7_1[53]), .B(n116), .Y(n118) );
  OAI211X1 U489 ( .C(n114), .D(n41), .A(n117), .B(n39), .Y(N975) );
  NAND2X1 U490 ( .A(dat_7_1[54]), .B(n116), .Y(n117) );
  OAI211X1 U491 ( .C(n127), .D(n41), .A(n130), .B(n39), .Y(N966) );
  NAND2X1 U492 ( .A(mem_8__6_), .B(n129), .Y(n130) );
  OAI211X1 U493 ( .C(n114), .D(n49), .A(n115), .B(n47), .Y(N976) );
  NAND2X1 U494 ( .A(dat_7_1[55]), .B(n116), .Y(n115) );
  OAI211X1 U495 ( .C(n114), .D(n204), .A(n121), .B(n179), .Y(N971) );
  NAND2X1 U496 ( .A(dat_7_1[50]), .B(n116), .Y(n121) );
  OAI211X1 U497 ( .C(n127), .D(n204), .A(n134), .B(n179), .Y(N962) );
  NAND2X1 U498 ( .A(mem_8__2_), .B(n129), .Y(n134) );
  OAI211X1 U499 ( .C(n127), .D(n311), .A(n133), .B(n275), .Y(N963) );
  NAND2X1 U500 ( .A(mem_8__3_), .B(n129), .Y(n133) );
  OAI211X1 U501 ( .C(n114), .D(n25), .A(n119), .B(n23), .Y(N973) );
  NAND2X1 U502 ( .A(dat_7_1[52]), .B(n116), .Y(n119) );
  OAI211X1 U503 ( .C(n127), .D(n25), .A(n132), .B(n23), .Y(N964) );
  NAND2X1 U504 ( .A(mem_8__4_), .B(n129), .Y(n132) );
  OAI211X1 U505 ( .C(n127), .D(n33), .A(n131), .B(n31), .Y(N965) );
  NAND2X1 U506 ( .A(mem_8__5_), .B(n129), .Y(n131) );
  OAI211X1 U507 ( .C(n127), .D(n49), .A(n128), .B(n47), .Y(N967) );
  NAND2X1 U508 ( .A(mem_8__7_), .B(n129), .Y(n128) );
  OAI211X1 U509 ( .C(n468), .D(n149), .A(n78), .B(n476), .Y(N1015) );
  NAND2X1 U510 ( .A(dat_7_1[9]), .B(n470), .Y(n476) );
  OAI211X1 U511 ( .C(n468), .D(n204), .A(n179), .B(n475), .Y(N1016) );
  NAND2X1 U512 ( .A(dat_7_1[10]), .B(n470), .Y(n475) );
  OAI211X1 U513 ( .C(n468), .D(n311), .A(n275), .B(n474), .Y(N1017) );
  NAND2X1 U514 ( .A(dat_7_1[11]), .B(n470), .Y(n474) );
  OAI211X1 U515 ( .C(n468), .D(n57), .A(n53), .B(n477), .Y(N1014) );
  NAND2X1 U516 ( .A(dat_7_1[8]), .B(n470), .Y(n477) );
  OAI211X1 U517 ( .C(n138), .D(n57), .A(n147), .B(n53), .Y(N951) );
  NAND2X1 U518 ( .A(mem_9__0_), .B(n140), .Y(n147) );
  OAI211X1 U519 ( .C(n153), .D(n57), .A(n162), .B(n53), .Y(N942) );
  NAND2X1 U520 ( .A(mem_10__0_), .B(n155), .Y(n162) );
  OAI211X1 U521 ( .C(n166), .D(n57), .A(n175), .B(n53), .Y(N933) );
  NAND2X1 U522 ( .A(mem_11__0_), .B(n168), .Y(n175) );
  OAI211X1 U523 ( .C(n180), .D(n57), .A(n189), .B(n54), .Y(N924) );
  NAND2X1 U524 ( .A(mem_12__0_), .B(n182), .Y(n189) );
  OAI211X1 U525 ( .C(n192), .D(n59), .A(n201), .B(n54), .Y(N915) );
  NAND2X1 U526 ( .A(mem_13__0_), .B(n194), .Y(n201) );
  OAI211X1 U527 ( .C(n205), .D(n59), .A(n214), .B(n54), .Y(N906) );
  NAND2X1 U528 ( .A(mem_14__0_), .B(n207), .Y(n214) );
  OAI211X1 U529 ( .C(n216), .D(n59), .A(n225), .B(n54), .Y(N897) );
  NAND2X1 U530 ( .A(mem_15__0_), .B(n218), .Y(n225) );
  OAI211X1 U531 ( .C(n227), .D(n59), .A(n236), .B(n54), .Y(N888) );
  NAND2X1 U532 ( .A(mem_16__0_), .B(n229), .Y(n236) );
  OAI211X1 U533 ( .C(n276), .D(n59), .A(n285), .B(n54), .Y(N852) );
  NAND2X1 U534 ( .A(mem_20__0_), .B(n278), .Y(n285) );
  OAI211X1 U535 ( .C(n300), .D(n59), .A(n309), .B(n55), .Y(N834) );
  NAND2X1 U536 ( .A(mem_22__0_), .B(n302), .Y(n309) );
  OAI211X1 U537 ( .C(n312), .D(n61), .A(n321), .B(n55), .Y(N825) );
  NAND2X1 U538 ( .A(mem_23__0_), .B(n314), .Y(n321) );
  OAI211X1 U539 ( .C(n324), .D(n61), .A(n333), .B(n55), .Y(N816) );
  NAND2X1 U540 ( .A(mem_24__0_), .B(n326), .Y(n333) );
  OAI211X1 U541 ( .C(n334), .D(n61), .A(n343), .B(n55), .Y(N807) );
  NAND2X1 U542 ( .A(mem_25__0_), .B(n336), .Y(n343) );
  OAI211X1 U543 ( .C(n345), .D(n61), .A(n354), .B(n55), .Y(N798) );
  NAND2X1 U544 ( .A(mem_26__0_), .B(n347), .Y(n354) );
  OAI211X1 U545 ( .C(n358), .D(n61), .A(n367), .B(n55), .Y(N789) );
  NAND2X1 U546 ( .A(mem_27__0_), .B(n360), .Y(n367) );
  OAI211X1 U547 ( .C(n370), .D(n61), .A(n379), .B(n55), .Y(N780) );
  NAND2X1 U548 ( .A(mem_28__0_), .B(n372), .Y(n379) );
  OAI211X1 U549 ( .C(n138), .D(n149), .A(n146), .B(n99), .Y(N952) );
  NAND2X1 U550 ( .A(mem_9__1_), .B(n140), .Y(n146) );
  OAI211X1 U551 ( .C(n153), .D(n149), .A(n161), .B(n78), .Y(N943) );
  NAND2X1 U552 ( .A(mem_10__1_), .B(n155), .Y(n161) );
  OAI211X1 U553 ( .C(n166), .D(n149), .A(n174), .B(n78), .Y(N934) );
  NAND2X1 U554 ( .A(mem_11__1_), .B(n168), .Y(n174) );
  OAI211X1 U555 ( .C(n180), .D(n149), .A(n188), .B(n99), .Y(N925) );
  NAND2X1 U556 ( .A(mem_12__1_), .B(n182), .Y(n188) );
  OAI211X1 U557 ( .C(n192), .D(n152), .A(n200), .B(n99), .Y(N916) );
  NAND2X1 U558 ( .A(mem_13__1_), .B(n194), .Y(n200) );
  OAI211X1 U559 ( .C(n205), .D(n152), .A(n213), .B(n99), .Y(N907) );
  NAND2X1 U560 ( .A(mem_14__1_), .B(n207), .Y(n213) );
  OAI211X1 U561 ( .C(n216), .D(n152), .A(n224), .B(n99), .Y(N898) );
  NAND2X1 U562 ( .A(mem_15__1_), .B(n218), .Y(n224) );
  OAI211X1 U563 ( .C(n227), .D(n152), .A(n235), .B(n99), .Y(N889) );
  NAND2X1 U564 ( .A(mem_16__1_), .B(n229), .Y(n235) );
  OAI211X1 U565 ( .C(n276), .D(n152), .A(n284), .B(n99), .Y(N853) );
  NAND2X1 U566 ( .A(mem_20__1_), .B(n278), .Y(n284) );
  OAI211X1 U567 ( .C(n300), .D(n152), .A(n308), .B(n126), .Y(N835) );
  NAND2X1 U568 ( .A(mem_22__1_), .B(n302), .Y(n308) );
  OAI211X1 U569 ( .C(n312), .D(n163), .A(n320), .B(n126), .Y(N826) );
  NAND2X1 U570 ( .A(mem_23__1_), .B(n314), .Y(n320) );
  OAI211X1 U571 ( .C(n324), .D(n163), .A(n332), .B(n126), .Y(N817) );
  NAND2X1 U572 ( .A(mem_24__1_), .B(n326), .Y(n332) );
  OAI211X1 U573 ( .C(n334), .D(n163), .A(n342), .B(n126), .Y(N808) );
  NAND2X1 U574 ( .A(mem_25__1_), .B(n336), .Y(n342) );
  OAI211X1 U575 ( .C(n345), .D(n163), .A(n353), .B(n126), .Y(N799) );
  NAND2X1 U576 ( .A(mem_26__1_), .B(n347), .Y(n353) );
  OAI211X1 U577 ( .C(n358), .D(n163), .A(n366), .B(n126), .Y(N790) );
  NAND2X1 U578 ( .A(mem_27__1_), .B(n360), .Y(n366) );
  OAI211X1 U579 ( .C(n370), .D(n163), .A(n378), .B(n126), .Y(N781) );
  NAND2X1 U580 ( .A(mem_28__1_), .B(n372), .Y(n378) );
  OAI211X1 U581 ( .C(n138), .D(n204), .A(n145), .B(n190), .Y(N953) );
  NAND2X1 U582 ( .A(mem_9__2_), .B(n140), .Y(n145) );
  OAI211X1 U583 ( .C(n153), .D(n204), .A(n160), .B(n179), .Y(N944) );
  NAND2X1 U584 ( .A(mem_10__2_), .B(n155), .Y(n160) );
  OAI211X1 U585 ( .C(n166), .D(n204), .A(n173), .B(n179), .Y(N935) );
  NAND2X1 U586 ( .A(mem_11__2_), .B(n168), .Y(n173) );
  OAI211X1 U587 ( .C(n180), .D(n204), .A(n187), .B(n190), .Y(N926) );
  NAND2X1 U588 ( .A(mem_12__2_), .B(n182), .Y(n187) );
  OAI211X1 U589 ( .C(n192), .D(n249), .A(n199), .B(n190), .Y(N917) );
  NAND2X1 U590 ( .A(mem_13__2_), .B(n194), .Y(n199) );
  OAI211X1 U591 ( .C(n205), .D(n249), .A(n212), .B(n190), .Y(N908) );
  NAND2X1 U592 ( .A(mem_14__2_), .B(n207), .Y(n212) );
  OAI211X1 U593 ( .C(n216), .D(n249), .A(n223), .B(n190), .Y(N899) );
  NAND2X1 U594 ( .A(mem_15__2_), .B(n218), .Y(n223) );
  OAI211X1 U595 ( .C(n227), .D(n249), .A(n234), .B(n190), .Y(N890) );
  NAND2X1 U596 ( .A(mem_16__2_), .B(n229), .Y(n234) );
  OAI211X1 U597 ( .C(n276), .D(n249), .A(n283), .B(n190), .Y(N854) );
  NAND2X1 U598 ( .A(mem_20__2_), .B(n278), .Y(n283) );
  OAI211X1 U599 ( .C(n300), .D(n249), .A(n307), .B(n191), .Y(N836) );
  NAND2X1 U600 ( .A(mem_22__2_), .B(n302), .Y(n307) );
  OAI211X1 U601 ( .C(n312), .D(n261), .A(n319), .B(n191), .Y(N827) );
  NAND2X1 U602 ( .A(mem_23__2_), .B(n314), .Y(n319) );
  OAI211X1 U603 ( .C(n324), .D(n261), .A(n331), .B(n191), .Y(N818) );
  NAND2X1 U604 ( .A(mem_24__2_), .B(n326), .Y(n331) );
  OAI211X1 U605 ( .C(n334), .D(n261), .A(n341), .B(n191), .Y(N809) );
  NAND2X1 U606 ( .A(mem_25__2_), .B(n336), .Y(n341) );
  OAI211X1 U607 ( .C(n345), .D(n261), .A(n352), .B(n191), .Y(N800) );
  NAND2X1 U608 ( .A(mem_26__2_), .B(n347), .Y(n352) );
  OAI211X1 U609 ( .C(n358), .D(n261), .A(n365), .B(n191), .Y(N791) );
  NAND2X1 U610 ( .A(mem_27__2_), .B(n360), .Y(n365) );
  OAI211X1 U611 ( .C(n370), .D(n261), .A(n377), .B(n191), .Y(N782) );
  NAND2X1 U612 ( .A(mem_28__2_), .B(n372), .Y(n377) );
  OAI211X1 U613 ( .C(n138), .D(n311), .A(n144), .B(n286), .Y(N954) );
  NAND2X1 U614 ( .A(mem_9__3_), .B(n140), .Y(n144) );
  OAI211X1 U615 ( .C(n153), .D(n311), .A(n159), .B(n275), .Y(N945) );
  NAND2X1 U616 ( .A(mem_10__3_), .B(n155), .Y(n159) );
  OAI211X1 U617 ( .C(n166), .D(n311), .A(n172), .B(n275), .Y(N936) );
  NAND2X1 U618 ( .A(mem_11__3_), .B(n168), .Y(n172) );
  OAI211X1 U619 ( .C(n180), .D(n311), .A(n186), .B(n286), .Y(N927) );
  NAND2X1 U620 ( .A(mem_12__3_), .B(n182), .Y(n186) );
  OAI211X1 U621 ( .C(n192), .D(n356), .A(n198), .B(n286), .Y(N918) );
  NAND2X1 U622 ( .A(mem_13__3_), .B(n194), .Y(n198) );
  OAI211X1 U623 ( .C(n205), .D(n356), .A(n211), .B(n286), .Y(N909) );
  NAND2X1 U624 ( .A(mem_14__3_), .B(n207), .Y(n211) );
  OAI211X1 U625 ( .C(n216), .D(n356), .A(n222), .B(n286), .Y(N900) );
  NAND2X1 U626 ( .A(mem_15__3_), .B(n218), .Y(n222) );
  OAI211X1 U627 ( .C(n227), .D(n356), .A(n233), .B(n286), .Y(N891) );
  NAND2X1 U628 ( .A(mem_16__3_), .B(n229), .Y(n233) );
  OAI211X1 U629 ( .C(n276), .D(n356), .A(n282), .B(n286), .Y(N855) );
  NAND2X1 U630 ( .A(mem_20__3_), .B(n278), .Y(n282) );
  OAI211X1 U631 ( .C(n300), .D(n356), .A(n306), .B(n298), .Y(N837) );
  NAND2X1 U632 ( .A(mem_22__3_), .B(n302), .Y(n306) );
  OAI211X1 U633 ( .C(n312), .D(n357), .A(n318), .B(n298), .Y(N828) );
  NAND2X1 U634 ( .A(mem_23__3_), .B(n314), .Y(n318) );
  OAI211X1 U635 ( .C(n324), .D(n357), .A(n330), .B(n298), .Y(N819) );
  NAND2X1 U636 ( .A(mem_24__3_), .B(n326), .Y(n330) );
  OAI211X1 U637 ( .C(n334), .D(n357), .A(n340), .B(n298), .Y(N810) );
  NAND2X1 U638 ( .A(mem_25__3_), .B(n336), .Y(n340) );
  OAI211X1 U639 ( .C(n345), .D(n357), .A(n351), .B(n298), .Y(N801) );
  NAND2X1 U640 ( .A(mem_26__3_), .B(n347), .Y(n351) );
  OAI211X1 U641 ( .C(n358), .D(n357), .A(n364), .B(n298), .Y(N792) );
  NAND2X1 U642 ( .A(mem_27__3_), .B(n360), .Y(n364) );
  OAI211X1 U643 ( .C(n370), .D(n357), .A(n376), .B(n298), .Y(N783) );
  NAND2X1 U644 ( .A(mem_28__3_), .B(n372), .Y(n376) );
  OAI211X1 U645 ( .C(n138), .D(n25), .A(n143), .B(n23), .Y(N955) );
  NAND2X1 U646 ( .A(mem_9__4_), .B(n140), .Y(n143) );
  OAI211X1 U647 ( .C(n153), .D(n25), .A(n158), .B(n23), .Y(N946) );
  NAND2X1 U648 ( .A(mem_10__4_), .B(n155), .Y(n158) );
  OAI211X1 U649 ( .C(n166), .D(n25), .A(n171), .B(n23), .Y(N937) );
  NAND2X1 U650 ( .A(mem_11__4_), .B(n168), .Y(n171) );
  OAI211X1 U651 ( .C(n180), .D(n25), .A(n185), .B(n23), .Y(N928) );
  NAND2X1 U652 ( .A(mem_12__4_), .B(n182), .Y(n185) );
  OAI211X1 U653 ( .C(n192), .D(n25), .A(n197), .B(n23), .Y(N919) );
  NAND2X1 U654 ( .A(mem_13__4_), .B(n194), .Y(n197) );
  OAI211X1 U655 ( .C(n205), .D(n26), .A(n210), .B(n23), .Y(N910) );
  NAND2X1 U656 ( .A(mem_14__4_), .B(n207), .Y(n210) );
  OAI211X1 U657 ( .C(n216), .D(n26), .A(n221), .B(n23), .Y(N901) );
  NAND2X1 U658 ( .A(mem_15__4_), .B(n218), .Y(n221) );
  OAI211X1 U659 ( .C(n227), .D(n26), .A(n232), .B(n23), .Y(N892) );
  NAND2X1 U660 ( .A(mem_16__4_), .B(n229), .Y(n232) );
  OAI211X1 U661 ( .C(n276), .D(n26), .A(n281), .B(n22), .Y(N856) );
  NAND2X1 U662 ( .A(mem_20__4_), .B(n278), .Y(n281) );
  OAI211X1 U663 ( .C(n300), .D(n26), .A(n305), .B(n22), .Y(N838) );
  NAND2X1 U664 ( .A(mem_22__4_), .B(n302), .Y(n305) );
  OAI211X1 U665 ( .C(n312), .D(n26), .A(n317), .B(n22), .Y(N829) );
  NAND2X1 U666 ( .A(mem_23__4_), .B(n314), .Y(n317) );
  OAI211X1 U667 ( .C(n324), .D(n27), .A(n329), .B(n22), .Y(N820) );
  NAND2X1 U668 ( .A(mem_24__4_), .B(n326), .Y(n329) );
  OAI211X1 U669 ( .C(n334), .D(n27), .A(n339), .B(n22), .Y(N811) );
  NAND2X1 U670 ( .A(mem_25__4_), .B(n336), .Y(n339) );
  OAI211X1 U671 ( .C(n345), .D(n27), .A(n350), .B(n22), .Y(N802) );
  NAND2X1 U672 ( .A(mem_26__4_), .B(n347), .Y(n350) );
  OAI211X1 U673 ( .C(n358), .D(n27), .A(n363), .B(n21), .Y(N793) );
  NAND2X1 U674 ( .A(mem_27__4_), .B(n360), .Y(n363) );
  OAI211X1 U675 ( .C(n370), .D(n27), .A(n375), .B(n21), .Y(N784) );
  NAND2X1 U676 ( .A(mem_28__4_), .B(n372), .Y(n375) );
  OAI211X1 U677 ( .C(n138), .D(n33), .A(n142), .B(n31), .Y(N956) );
  NAND2X1 U678 ( .A(mem_9__5_), .B(n140), .Y(n142) );
  OAI211X1 U679 ( .C(n153), .D(n33), .A(n157), .B(n31), .Y(N947) );
  NAND2X1 U680 ( .A(mem_10__5_), .B(n155), .Y(n157) );
  OAI211X1 U681 ( .C(n166), .D(n33), .A(n170), .B(n31), .Y(N938) );
  NAND2X1 U682 ( .A(mem_11__5_), .B(n168), .Y(n170) );
  OAI211X1 U683 ( .C(n180), .D(n33), .A(n184), .B(n31), .Y(N929) );
  NAND2X1 U684 ( .A(mem_12__5_), .B(n182), .Y(n184) );
  OAI211X1 U685 ( .C(n192), .D(n33), .A(n196), .B(n31), .Y(N920) );
  NAND2X1 U686 ( .A(mem_13__5_), .B(n194), .Y(n196) );
  OAI211X1 U687 ( .C(n205), .D(n34), .A(n209), .B(n31), .Y(N911) );
  NAND2X1 U688 ( .A(mem_14__5_), .B(n207), .Y(n209) );
  OAI211X1 U689 ( .C(n216), .D(n34), .A(n220), .B(n31), .Y(N902) );
  NAND2X1 U690 ( .A(mem_15__5_), .B(n218), .Y(n220) );
  OAI211X1 U691 ( .C(n227), .D(n34), .A(n231), .B(n31), .Y(N893) );
  NAND2X1 U692 ( .A(mem_16__5_), .B(n229), .Y(n231) );
  OAI211X1 U693 ( .C(n276), .D(n34), .A(n280), .B(n30), .Y(N857) );
  NAND2X1 U694 ( .A(mem_20__5_), .B(n278), .Y(n280) );
  OAI211X1 U695 ( .C(n300), .D(n34), .A(n304), .B(n30), .Y(N839) );
  NAND2X1 U696 ( .A(mem_22__5_), .B(n302), .Y(n304) );
  OAI211X1 U697 ( .C(n312), .D(n34), .A(n316), .B(n30), .Y(N830) );
  NAND2X1 U698 ( .A(mem_23__5_), .B(n314), .Y(n316) );
  OAI211X1 U699 ( .C(n324), .D(n35), .A(n328), .B(n30), .Y(N821) );
  NAND2X1 U700 ( .A(mem_24__5_), .B(n326), .Y(n328) );
  OAI211X1 U701 ( .C(n334), .D(n35), .A(n338), .B(n30), .Y(N812) );
  NAND2X1 U702 ( .A(mem_25__5_), .B(n336), .Y(n338) );
  OAI211X1 U703 ( .C(n345), .D(n35), .A(n349), .B(n30), .Y(N803) );
  NAND2X1 U704 ( .A(mem_26__5_), .B(n347), .Y(n349) );
  OAI211X1 U705 ( .C(n358), .D(n35), .A(n362), .B(n29), .Y(N794) );
  NAND2X1 U706 ( .A(mem_27__5_), .B(n360), .Y(n362) );
  OAI211X1 U707 ( .C(n370), .D(n35), .A(n374), .B(n29), .Y(N785) );
  NAND2X1 U708 ( .A(mem_28__5_), .B(n372), .Y(n374) );
  OAI211X1 U709 ( .C(n138), .D(n41), .A(n141), .B(n39), .Y(N957) );
  NAND2X1 U710 ( .A(mem_9__6_), .B(n140), .Y(n141) );
  OAI211X1 U711 ( .C(n153), .D(n41), .A(n156), .B(n39), .Y(N948) );
  NAND2X1 U712 ( .A(mem_10__6_), .B(n155), .Y(n156) );
  OAI211X1 U713 ( .C(n166), .D(n41), .A(n169), .B(n39), .Y(N939) );
  NAND2X1 U714 ( .A(mem_11__6_), .B(n168), .Y(n169) );
  OAI211X1 U715 ( .C(n180), .D(n41), .A(n183), .B(n39), .Y(N930) );
  NAND2X1 U716 ( .A(mem_12__6_), .B(n182), .Y(n183) );
  OAI211X1 U717 ( .C(n192), .D(n41), .A(n195), .B(n39), .Y(N921) );
  NAND2X1 U718 ( .A(mem_13__6_), .B(n194), .Y(n195) );
  OAI211X1 U719 ( .C(n205), .D(n42), .A(n208), .B(n39), .Y(N912) );
  NAND2X1 U720 ( .A(mem_14__6_), .B(n207), .Y(n208) );
  OAI211X1 U721 ( .C(n216), .D(n42), .A(n219), .B(n39), .Y(N903) );
  NAND2X1 U722 ( .A(mem_15__6_), .B(n218), .Y(n219) );
  OAI211X1 U723 ( .C(n227), .D(n42), .A(n230), .B(n39), .Y(N894) );
  NAND2X1 U724 ( .A(mem_16__6_), .B(n229), .Y(n230) );
  OAI211X1 U725 ( .C(n276), .D(n42), .A(n279), .B(n38), .Y(N858) );
  NAND2X1 U726 ( .A(mem_20__6_), .B(n278), .Y(n279) );
  OAI211X1 U727 ( .C(n300), .D(n42), .A(n303), .B(n38), .Y(N840) );
  NAND2X1 U728 ( .A(mem_22__6_), .B(n302), .Y(n303) );
  OAI211X1 U729 ( .C(n312), .D(n42), .A(n315), .B(n38), .Y(N831) );
  NAND2X1 U730 ( .A(mem_23__6_), .B(n314), .Y(n315) );
  OAI211X1 U731 ( .C(n324), .D(n43), .A(n327), .B(n38), .Y(N822) );
  NAND2X1 U732 ( .A(mem_24__6_), .B(n326), .Y(n327) );
  OAI211X1 U733 ( .C(n334), .D(n43), .A(n337), .B(n38), .Y(N813) );
  NAND2X1 U734 ( .A(mem_25__6_), .B(n336), .Y(n337) );
  OAI211X1 U735 ( .C(n345), .D(n43), .A(n348), .B(n38), .Y(N804) );
  NAND2X1 U736 ( .A(mem_26__6_), .B(n347), .Y(n348) );
  OAI211X1 U737 ( .C(n358), .D(n43), .A(n361), .B(n37), .Y(N795) );
  NAND2X1 U738 ( .A(mem_27__6_), .B(n360), .Y(n361) );
  OAI211X1 U739 ( .C(n370), .D(n43), .A(n373), .B(n37), .Y(N786) );
  NAND2X1 U740 ( .A(mem_28__6_), .B(n372), .Y(n373) );
  OAI211X1 U741 ( .C(n138), .D(n49), .A(n139), .B(n47), .Y(N958) );
  NAND2X1 U742 ( .A(mem_9__7_), .B(n140), .Y(n139) );
  OAI211X1 U743 ( .C(n153), .D(n49), .A(n154), .B(n47), .Y(N949) );
  NAND2X1 U744 ( .A(mem_10__7_), .B(n155), .Y(n154) );
  OAI211X1 U745 ( .C(n166), .D(n49), .A(n167), .B(n47), .Y(N940) );
  NAND2X1 U746 ( .A(mem_11__7_), .B(n168), .Y(n167) );
  OAI211X1 U747 ( .C(n180), .D(n49), .A(n181), .B(n47), .Y(N931) );
  NAND2X1 U748 ( .A(mem_12__7_), .B(n182), .Y(n181) );
  OAI211X1 U749 ( .C(n192), .D(n49), .A(n193), .B(n47), .Y(N922) );
  NAND2X1 U750 ( .A(mem_13__7_), .B(n194), .Y(n193) );
  OAI211X1 U751 ( .C(n205), .D(n50), .A(n206), .B(n47), .Y(N913) );
  NAND2X1 U752 ( .A(mem_14__7_), .B(n207), .Y(n206) );
  OAI211X1 U753 ( .C(n216), .D(n50), .A(n217), .B(n47), .Y(N904) );
  NAND2X1 U754 ( .A(mem_15__7_), .B(n218), .Y(n217) );
  OAI211X1 U755 ( .C(n227), .D(n50), .A(n228), .B(n47), .Y(N895) );
  NAND2X1 U756 ( .A(mem_16__7_), .B(n229), .Y(n228) );
  OAI211X1 U757 ( .C(n276), .D(n50), .A(n277), .B(n46), .Y(N859) );
  NAND2X1 U758 ( .A(mem_20__7_), .B(n278), .Y(n277) );
  OAI211X1 U759 ( .C(n300), .D(n50), .A(n301), .B(n46), .Y(N841) );
  NAND2X1 U760 ( .A(mem_22__7_), .B(n302), .Y(n301) );
  OAI211X1 U761 ( .C(n312), .D(n50), .A(n313), .B(n46), .Y(N832) );
  NAND2X1 U762 ( .A(mem_23__7_), .B(n314), .Y(n313) );
  OAI211X1 U763 ( .C(n324), .D(n51), .A(n325), .B(n46), .Y(N823) );
  NAND2X1 U764 ( .A(mem_24__7_), .B(n326), .Y(n325) );
  OAI211X1 U765 ( .C(n334), .D(n51), .A(n335), .B(n46), .Y(N814) );
  NAND2X1 U766 ( .A(mem_25__7_), .B(n336), .Y(n335) );
  OAI211X1 U767 ( .C(n345), .D(n51), .A(n346), .B(n46), .Y(N805) );
  NAND2X1 U768 ( .A(mem_26__7_), .B(n347), .Y(n346) );
  OAI211X1 U769 ( .C(n358), .D(n51), .A(n359), .B(n45), .Y(N796) );
  NAND2X1 U770 ( .A(mem_27__7_), .B(n360), .Y(n359) );
  OAI211X1 U771 ( .C(n370), .D(n51), .A(n371), .B(n45), .Y(N787) );
  NAND2X1 U772 ( .A(mem_28__7_), .B(n372), .Y(n371) );
  OAI211X1 U773 ( .C(n381), .D(n61), .A(n390), .B(n55), .Y(N771) );
  NAND2X1 U774 ( .A(mem_29__0_), .B(n383), .Y(n390) );
  OAI211X1 U775 ( .C(n394), .D(n61), .A(n403), .B(n55), .Y(N762) );
  NAND2X1 U776 ( .A(mem_30__0_), .B(n396), .Y(n403) );
  OAI211X1 U777 ( .C(n407), .D(n61), .A(n416), .B(n55), .Y(N753) );
  NAND2X1 U778 ( .A(mem_31__0_), .B(n409), .Y(n416) );
  OAI211X1 U779 ( .C(n417), .D(n61), .A(n426), .B(n74), .Y(N744) );
  NAND2X1 U780 ( .A(mem_32__0_), .B(n419), .Y(n426) );
  OAI211X1 U781 ( .C(n381), .D(n163), .A(n389), .B(n126), .Y(N772) );
  NAND2X1 U782 ( .A(mem_29__1_), .B(n383), .Y(n389) );
  OAI211X1 U783 ( .C(n394), .D(n163), .A(n402), .B(n126), .Y(N763) );
  NAND2X1 U784 ( .A(mem_30__1_), .B(n396), .Y(n402) );
  OAI211X1 U785 ( .C(n407), .D(n163), .A(n415), .B(n71), .Y(N754) );
  NAND2X1 U786 ( .A(mem_31__1_), .B(n409), .Y(n415) );
  OAI211X1 U787 ( .C(n417), .D(n163), .A(n425), .B(n71), .Y(N745) );
  NAND2X1 U788 ( .A(mem_32__1_), .B(n419), .Y(n425) );
  OAI211X1 U789 ( .C(n381), .D(n261), .A(n388), .B(n191), .Y(N773) );
  NAND2X1 U790 ( .A(mem_29__2_), .B(n383), .Y(n388) );
  OAI211X1 U791 ( .C(n394), .D(n261), .A(n401), .B(n191), .Y(N764) );
  NAND2X1 U792 ( .A(mem_30__2_), .B(n396), .Y(n401) );
  OAI211X1 U793 ( .C(n407), .D(n261), .A(n414), .B(n68), .Y(N755) );
  NAND2X1 U794 ( .A(mem_31__2_), .B(n409), .Y(n414) );
  OAI211X1 U795 ( .C(n417), .D(n261), .A(n424), .B(n68), .Y(N746) );
  NAND2X1 U796 ( .A(mem_32__2_), .B(n419), .Y(n424) );
  OAI211X1 U797 ( .C(n381), .D(n357), .A(n387), .B(n298), .Y(N774) );
  NAND2X1 U798 ( .A(mem_29__3_), .B(n383), .Y(n387) );
  OAI211X1 U799 ( .C(n394), .D(n357), .A(n400), .B(n298), .Y(N765) );
  NAND2X1 U800 ( .A(mem_30__3_), .B(n396), .Y(n400) );
  OAI211X1 U801 ( .C(n407), .D(n357), .A(n413), .B(n64), .Y(N756) );
  NAND2X1 U802 ( .A(mem_31__3_), .B(n409), .Y(n413) );
  OAI211X1 U803 ( .C(n417), .D(n357), .A(n423), .B(n64), .Y(N747) );
  NAND2X1 U804 ( .A(mem_32__3_), .B(n419), .Y(n423) );
  OAI211X1 U805 ( .C(n381), .D(n27), .A(n386), .B(n21), .Y(N775) );
  NAND2X1 U806 ( .A(mem_29__4_), .B(n383), .Y(n386) );
  OAI211X1 U807 ( .C(n394), .D(n27), .A(n399), .B(n21), .Y(N766) );
  NAND2X1 U808 ( .A(mem_30__4_), .B(n396), .Y(n399) );
  OAI211X1 U809 ( .C(n407), .D(n27), .A(n412), .B(n21), .Y(N757) );
  NAND2X1 U810 ( .A(mem_31__4_), .B(n409), .Y(n412) );
  OAI211X1 U811 ( .C(n417), .D(n27), .A(n422), .B(n21), .Y(N748) );
  NAND2X1 U812 ( .A(mem_32__4_), .B(n419), .Y(n422) );
  OAI211X1 U813 ( .C(n429), .D(n27), .A(n434), .B(n21), .Y(N739) );
  NAND2X1 U814 ( .A(mem_33__4_), .B(n431), .Y(n434) );
  OAI211X1 U815 ( .C(n381), .D(n35), .A(n385), .B(n29), .Y(N776) );
  NAND2X1 U816 ( .A(mem_29__5_), .B(n383), .Y(n385) );
  OAI211X1 U817 ( .C(n394), .D(n35), .A(n398), .B(n29), .Y(N767) );
  NAND2X1 U818 ( .A(mem_30__5_), .B(n396), .Y(n398) );
  OAI211X1 U819 ( .C(n407), .D(n35), .A(n411), .B(n29), .Y(N758) );
  NAND2X1 U820 ( .A(mem_31__5_), .B(n409), .Y(n411) );
  OAI211X1 U821 ( .C(n417), .D(n35), .A(n421), .B(n29), .Y(N749) );
  NAND2X1 U822 ( .A(mem_32__5_), .B(n419), .Y(n421) );
  OAI211X1 U823 ( .C(n429), .D(n35), .A(n433), .B(n29), .Y(N740) );
  NAND2X1 U824 ( .A(mem_33__5_), .B(n431), .Y(n433) );
  OAI211X1 U825 ( .C(n381), .D(n43), .A(n384), .B(n37), .Y(N777) );
  NAND2X1 U826 ( .A(mem_29__6_), .B(n383), .Y(n384) );
  OAI211X1 U827 ( .C(n394), .D(n43), .A(n397), .B(n37), .Y(N768) );
  NAND2X1 U828 ( .A(mem_30__6_), .B(n396), .Y(n397) );
  OAI211X1 U829 ( .C(n407), .D(n43), .A(n410), .B(n37), .Y(N759) );
  NAND2X1 U830 ( .A(mem_31__6_), .B(n409), .Y(n410) );
  OAI211X1 U831 ( .C(n417), .D(n43), .A(n420), .B(n37), .Y(N750) );
  NAND2X1 U832 ( .A(mem_32__6_), .B(n419), .Y(n420) );
  OAI211X1 U833 ( .C(n429), .D(n43), .A(n432), .B(n37), .Y(N741) );
  NAND2X1 U834 ( .A(mem_33__6_), .B(n431), .Y(n432) );
  OAI211X1 U835 ( .C(n381), .D(n51), .A(n382), .B(n45), .Y(N778) );
  NAND2X1 U836 ( .A(mem_29__7_), .B(n383), .Y(n382) );
  OAI211X1 U837 ( .C(n394), .D(n51), .A(n395), .B(n45), .Y(N769) );
  NAND2X1 U838 ( .A(mem_30__7_), .B(n396), .Y(n395) );
  OAI211X1 U839 ( .C(n407), .D(n51), .A(n408), .B(n45), .Y(N760) );
  NAND2X1 U840 ( .A(mem_31__7_), .B(n409), .Y(n408) );
  OAI211X1 U841 ( .C(n417), .D(n51), .A(n418), .B(n45), .Y(N751) );
  NAND2X1 U842 ( .A(mem_32__7_), .B(n419), .Y(n418) );
  OAI211X1 U843 ( .C(n429), .D(n51), .A(n430), .B(n45), .Y(N742) );
  NAND2X1 U844 ( .A(mem_33__7_), .B(n431), .Y(n430) );
  OAI211X1 U845 ( .C(n478), .D(n73), .A(n487), .B(n53), .Y(N1005) );
  NAND2X1 U846 ( .A(dat_7_1[16]), .B(n480), .Y(n487) );
  OAI211X1 U847 ( .C(n478), .D(n67), .A(n179), .B(n485), .Y(N1007) );
  NAND2X1 U848 ( .A(dat_7_1[18]), .B(n480), .Y(n485) );
  OAI211X1 U849 ( .C(n478), .D(n91), .A(n483), .B(n21), .Y(N1009) );
  NAND2X1 U850 ( .A(dat_7_1[20]), .B(n480), .Y(n483) );
  OAI211X1 U851 ( .C(n5), .D(n91), .A(n492), .B(n21), .Y(N1000) );
  NAND2X1 U852 ( .A(dat_7_1[28]), .B(n66), .Y(n492) );
  OAI211X1 U853 ( .C(n5), .D(n88), .A(n29), .B(n491), .Y(N1001) );
  NAND2X1 U854 ( .A(dat_7_1[29]), .B(n66), .Y(n491) );
  OAI211X1 U855 ( .C(n478), .D(n70), .A(n78), .B(n486), .Y(N1006) );
  NAND2X1 U856 ( .A(dat_7_1[17]), .B(n480), .Y(n486) );
  OAI211X1 U857 ( .C(n478), .D(n63), .A(n275), .B(n484), .Y(N1008) );
  NAND2X1 U858 ( .A(dat_7_1[19]), .B(n480), .Y(n484) );
  OAI211X1 U859 ( .C(n5), .D(n85), .A(n37), .B(n490), .Y(N1002) );
  NAND2X1 U860 ( .A(dat_7_1[30]), .B(n66), .Y(n490) );
  OAI211X1 U861 ( .C(n5), .D(n81), .A(n45), .B(n489), .Y(N1003) );
  NAND2X1 U862 ( .A(dat_7_1[31]), .B(n66), .Y(n489) );
  OAI211X1 U863 ( .C(n478), .D(n88), .A(n482), .B(n29), .Y(N1010) );
  NAND2X1 U864 ( .A(dat_7_1[21]), .B(n480), .Y(n482) );
  OAI211X1 U865 ( .C(n478), .D(n81), .A(n479), .B(n45), .Y(N1012) );
  NAND2X1 U866 ( .A(dat_7_1[23]), .B(n480), .Y(n479) );
  OAI211X1 U867 ( .C(n478), .D(n85), .A(n481), .B(n37), .Y(N1011) );
  NAND2X1 U868 ( .A(dat_7_1[22]), .B(n480), .Y(n481) );
  OAI211X1 U869 ( .C(n429), .D(n73), .A(n438), .B(n74), .Y(N735) );
  NAND2X1 U870 ( .A(mem_33__0_), .B(n431), .Y(n438) );
  OAI211X1 U871 ( .C(n429), .D(n70), .A(n437), .B(n78), .Y(N736) );
  NAND2X1 U872 ( .A(mem_33__1_), .B(n431), .Y(n437) );
  OAI211X1 U873 ( .C(n429), .D(n67), .A(n436), .B(n179), .Y(N737) );
  NAND2X1 U874 ( .A(mem_33__2_), .B(n431), .Y(n436) );
  OAI211X1 U875 ( .C(n429), .D(n63), .A(n435), .B(n275), .Y(N738) );
  NAND2X1 U876 ( .A(mem_33__3_), .B(n431), .Y(n435) );
  NAND21XL U877 ( .B(n508), .A(ptr[0]), .Y(n521) );
  MUX2X1 U878 ( .D0(fifowdat[2]), .D1(dat_7_1[2]), .S(n507), .Y(N1025) );
  MUX2X1 U879 ( .D0(fifowdat[3]), .D1(dat_7_1[3]), .S(n507), .Y(N1026) );
  MUX2X1 U880 ( .D0(fifowdat[5]), .D1(dat_7_1[5]), .S(n507), .Y(N1028) );
  MUX2X1 U881 ( .D0(fifowdat[6]), .D1(dat_7_1[6]), .S(n507), .Y(N1029) );
  MUX2X1 U882 ( .D0(fifowdat[7]), .D1(dat_7_1[7]), .S(n507), .Y(N1030) );
  MUX2X1 U883 ( .D0(fifowdat[0]), .D1(dat_7_1[0]), .S(n507), .Y(N1023) );
  MUX2X1 U884 ( .D0(fifowdat[1]), .D1(dat_7_1[1]), .S(n507), .Y(N1024) );
  MUX2X1 U885 ( .D0(fifowdat[4]), .D1(dat_7_1[4]), .S(n507), .Y(N1027) );
  NAND2X1 U886 ( .A(r_psh), .B(r_last), .Y(n58) );
  MUX2IX1 U887 ( .D0(r_wdat[0]), .D1(prx_wdat[0]), .S(prx_psh), .Y(n73) );
  MUX2IX1 U888 ( .D0(r_wdat[1]), .D1(prx_wdat[1]), .S(prx_psh), .Y(n70) );
  MUX2IX1 U889 ( .D0(r_wdat[2]), .D1(prx_wdat[2]), .S(prx_psh), .Y(n67) );
  NAND21X1 U890 ( .B(n428), .A(n405), .Y(n494) );
  NAND42XL U891 ( .C(ptr[1]), .D(ptr[2]), .A(n512), .B(n393), .Y(n405) );
  INVXL U892 ( .A(ptr[3]), .Y(n393) );
  NAND32XL U893 ( .B(ptr[4]), .C(n513), .A(n514), .Y(n510) );
  INVX1 U894 ( .A(i_ccidle), .Y(n577) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phycrc_a0 ( crc32_3_0, rx_good, i_shfidat, i_start, i_shfi4, i_shfo4, 
        clk, test_si, test_so, test_se );
  output [3:0] crc32_3_0;
  input [3:0] i_shfidat;
  input i_start, i_shfi4, i_shfo4, clk, test_si, test_se;
  output rx_good, test_so;
  wire   crc32_r_30_, crc32_r_29_, crc32_r_28_, crc32_r_27_, crc32_r_26_,
         crc32_r_25_, crc32_r_24_, crc32_r_23_, crc32_r_22_, crc32_r_21_,
         crc32_r_20_, crc32_r_19_, crc32_r_18_, crc32_r_17_, crc32_r_16_,
         crc32_r_15_, crc32_r_14_, crc32_r_13_, crc32_r_12_, crc32_r_11_,
         crc32_r_10_, crc32_r_9_, crc32_r_8_, crc32_r_7_, crc32_r_6_,
         crc32_r_5_, crc32_r_4_, crc32_r_3_, crc32_r_2_, crc32_r_1_,
         crc32_r_0_, N188, N189, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, net10623, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n58, n121, n122, n123, n124, n125, n126, n127;

  SNPS_CLOCK_GATE_HIGH_phycrc_a0 clk_gate_crc32_r_reg ( .CLK(clk), .EN(N188), 
        .ENCLK(net10623), .TE(test_se) );
  SDFFQX1 crc32_r_reg_26_ ( .D(N215), .SIN(crc32_r_25_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_26_) );
  SDFFQX1 crc32_r_reg_16_ ( .D(N205), .SIN(crc32_r_15_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_16_) );
  SDFFQX1 crc32_r_reg_27_ ( .D(N216), .SIN(crc32_r_26_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_27_) );
  SDFFQX1 crc32_r_reg_5_ ( .D(N194), .SIN(crc32_r_4_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_5_) );
  SDFFQX1 crc32_r_reg_0_ ( .D(N189), .SIN(test_si), .SMC(test_se), .C(net10623), .Q(crc32_r_0_) );
  SDFFQX1 crc32_r_reg_4_ ( .D(N193), .SIN(crc32_r_3_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_4_) );
  SDFFQX1 crc32_r_reg_14_ ( .D(N203), .SIN(crc32_r_13_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_14_) );
  SDFFQX1 crc32_r_reg_25_ ( .D(N214), .SIN(crc32_r_24_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_25_) );
  SDFFQX1 crc32_r_reg_3_ ( .D(N192), .SIN(crc32_r_2_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_3_) );
  SDFFQX1 crc32_r_reg_24_ ( .D(N213), .SIN(crc32_r_23_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_24_) );
  SDFFQX1 crc32_r_reg_21_ ( .D(N210), .SIN(crc32_r_20_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_21_) );
  SDFFQX1 crc32_r_reg_17_ ( .D(N206), .SIN(crc32_r_16_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_17_) );
  SDFFQX1 crc32_r_reg_8_ ( .D(N197), .SIN(crc32_r_7_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_8_) );
  SDFFQX1 crc32_r_reg_1_ ( .D(N190), .SIN(crc32_r_0_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_1_) );
  SDFFQX1 crc32_r_reg_10_ ( .D(N199), .SIN(crc32_r_9_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_10_) );
  SDFFQX1 crc32_r_reg_6_ ( .D(N195), .SIN(crc32_r_5_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_6_) );
  SDFFQX1 crc32_r_reg_11_ ( .D(N200), .SIN(crc32_r_10_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_11_) );
  SDFFQX1 crc32_r_reg_15_ ( .D(N204), .SIN(crc32_r_14_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_15_) );
  SDFFQX1 crc32_r_reg_12_ ( .D(N201), .SIN(crc32_r_11_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_12_) );
  SDFFQX1 crc32_r_reg_18_ ( .D(N207), .SIN(crc32_r_17_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_18_) );
  SDFFQX1 crc32_r_reg_20_ ( .D(N209), .SIN(crc32_r_19_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_20_) );
  SDFFQX1 crc32_r_reg_9_ ( .D(N198), .SIN(crc32_r_8_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_9_) );
  SDFFQX1 crc32_r_reg_7_ ( .D(N196), .SIN(crc32_r_6_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_7_) );
  SDFFQX1 crc32_r_reg_22_ ( .D(N211), .SIN(crc32_r_21_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_22_) );
  SDFFQX1 crc32_r_reg_2_ ( .D(N191), .SIN(crc32_r_1_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_2_) );
  SDFFQX1 crc32_r_reg_13_ ( .D(N202), .SIN(crc32_r_12_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_13_) );
  SDFFQX1 crc32_r_reg_23_ ( .D(N212), .SIN(crc32_r_22_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_23_) );
  SDFFQX1 crc32_r_reg_28_ ( .D(N217), .SIN(crc32_r_27_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_28_) );
  SDFFQX1 crc32_r_reg_29_ ( .D(N218), .SIN(crc32_r_28_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_29_) );
  SDFFQX1 crc32_r_reg_19_ ( .D(N208), .SIN(crc32_r_18_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_19_) );
  SDFFQX1 crc32_r_reg_31_ ( .D(N220), .SIN(crc32_r_30_), .SMC(test_se), .C(
        net10623), .Q(test_so) );
  SDFFQX1 crc32_r_reg_30_ ( .D(N219), .SIN(crc32_r_29_), .SMC(test_se), .C(
        net10623), .Q(crc32_r_30_) );
  INVX1 U3 ( .A(n18), .Y(n1) );
  XNOR2XL U4 ( .A(i_shfidat[2]), .B(n119), .Y(n56) );
  INVX1 U5 ( .A(n17), .Y(n2) );
  XNOR2XL U6 ( .A(i_shfidat[3]), .B(n120), .Y(n71) );
  INVX1 U7 ( .A(n19), .Y(n3) );
  XNOR2XL U8 ( .A(i_shfidat[1]), .B(n117), .Y(n51) );
  INVX1 U9 ( .A(n15), .Y(n4) );
  XNOR2XL U10 ( .A(i_shfidat[0]), .B(n114), .Y(n62) );
  INVX1 U11 ( .A(n62), .Y(n5) );
  INVX1 U12 ( .A(n62), .Y(n6) );
  AND2X1 U13 ( .A(i_shfo4), .B(n12), .Y(n60) );
  INVX1 U14 ( .A(n60), .Y(n7) );
  INVX1 U15 ( .A(n60), .Y(n8) );
  INVX1 U16 ( .A(n78), .Y(n9) );
  INVX1 U17 ( .A(n78), .Y(n10) );
  INVX1 U18 ( .A(n78), .Y(n16) );
  INVX1 U19 ( .A(n11), .Y(n12) );
  NAND2X1 U20 ( .A(n12), .B(n7), .Y(N188) );
  INVX1 U21 ( .A(n11), .Y(n14) );
  INVX1 U22 ( .A(n11), .Y(n13) );
  NAND21X1 U23 ( .B(n81), .A(n80), .Y(n63) );
  NAND2X1 U24 ( .A(i_start), .B(n19), .Y(n49) );
  NAND21X1 U25 ( .B(n12), .A(n81), .Y(n46) );
  OAI21X1 U26 ( .B(n14), .C(n115), .A(n9), .Y(N191) );
  XNOR2XL U27 ( .A(n17), .B(n116), .Y(n115) );
  XNOR2XL U28 ( .A(n18), .B(n19), .Y(n116) );
  OAI21X1 U29 ( .B(n14), .C(n118), .A(n10), .Y(N190) );
  XNOR2XL U30 ( .A(n17), .B(n18), .Y(n118) );
  INVX1 U31 ( .A(i_start), .Y(n15) );
  AOI21X1 U32 ( .B(n18), .C(n4), .A(n78), .Y(n55) );
  AOI21X1 U33 ( .B(n17), .C(n4), .A(n78), .Y(n74) );
  NOR2X1 U34 ( .A(i_shfi4), .B(n12), .Y(n78) );
  AND2X1 U35 ( .A(n80), .B(n16), .Y(n48) );
  NOR2X1 U36 ( .A(n12), .B(n4), .Y(n52) );
  OR2X1 U37 ( .A(i_start), .B(i_shfi4), .Y(n11) );
  OAI21X1 U38 ( .B(n14), .C(n17), .A(n16), .Y(N189) );
  INVX1 U39 ( .A(n51), .Y(n19) );
  AOI21AX1 U40 ( .B(n15), .C(n51), .A(n49), .Y(n68) );
  NOR2X1 U41 ( .A(n5), .B(i_start), .Y(n81) );
  INVX1 U42 ( .A(n56), .Y(n18) );
  NAND2X1 U43 ( .A(i_start), .B(n5), .Y(n80) );
  OAI21X1 U44 ( .B(n14), .C(n112), .A(n9), .Y(N192) );
  XNOR2XL U45 ( .A(n18), .B(n113), .Y(n112) );
  XNOR2XL U46 ( .A(n19), .B(n6), .Y(n113) );
  INVX1 U47 ( .A(n71), .Y(n17) );
  OAI21BX1 U48 ( .C(n7), .B(n6), .A(N188), .Y(n47) );
  OAI21X1 U49 ( .B(n14), .C(n3), .A(n7), .Y(n53) );
  OAI21X1 U50 ( .B(n14), .C(n56), .A(n7), .Y(n57) );
  OAI21X1 U51 ( .B(n14), .C(n71), .A(n7), .Y(n75) );
  NOR4XL U52 ( .A(n22), .B(n27), .C(n20), .D(n30), .Y(n41) );
  NOR4XL U53 ( .A(n31), .B(n21), .C(n32), .D(n26), .Y(n40) );
  NOR4XL U54 ( .A(n23), .B(n25), .C(n29), .D(n24), .Y(n38) );
  NOR2X1 U55 ( .A(crc32_r_30_), .B(i_start), .Y(n117) );
  NOR2X1 U56 ( .A(test_so), .B(i_start), .Y(n114) );
  OAI221X1 U57 ( .A(n13), .B(n106), .C(n26), .D(n7), .E(n9), .Y(N194) );
  XNOR2XL U58 ( .A(n107), .B(n71), .Y(n106) );
  XNOR2XL U59 ( .A(n56), .B(n108), .Y(n107) );
  OAI22X1 U60 ( .A(n26), .B(n6), .C(crc32_r_1_), .D(n63), .Y(n108) );
  OAI221X1 U61 ( .A(n13), .B(n98), .C(n23), .D(n7), .E(n10), .Y(N197) );
  XNOR2XL U62 ( .A(n99), .B(n71), .Y(n98) );
  XNOR2XL U63 ( .A(n56), .B(n100), .Y(n99) );
  OAI22X1 U64 ( .A(n23), .B(n6), .C(crc32_r_4_), .D(n63), .Y(n100) );
  OAI221X1 U65 ( .A(n13), .B(n90), .C(n8), .D(n122), .E(n16), .Y(N200) );
  XNOR2XL U66 ( .A(n91), .B(n71), .Y(n90) );
  XNOR2XL U67 ( .A(n56), .B(n92), .Y(n91) );
  OAI22X1 U68 ( .A(n6), .B(n122), .C(crc32_r_7_), .D(n63), .Y(n92) );
  OAI221X1 U69 ( .A(n12), .B(n84), .C(n8), .D(n35), .E(n9), .Y(N202) );
  XNOR2XL U70 ( .A(n85), .B(n56), .Y(n84) );
  XNOR2XL U71 ( .A(n51), .B(n86), .Y(n85) );
  OAI22X1 U72 ( .A(n6), .B(n35), .C(crc32_r_9_), .D(n63), .Y(n86) );
  OAI221X1 U73 ( .A(n13), .B(n101), .C(n28), .D(n7), .E(n10), .Y(N196) );
  XNOR2XL U74 ( .A(n102), .B(n71), .Y(n101) );
  XNOR2XL U75 ( .A(n51), .B(n103), .Y(n102) );
  OAI22X1 U76 ( .A(n28), .B(n5), .C(crc32_r_3_), .D(n63), .Y(n103) );
  OAI221X1 U77 ( .A(n13), .B(n93), .C(n29), .D(n7), .E(n16), .Y(N199) );
  XNOR2XL U78 ( .A(n94), .B(n71), .Y(n93) );
  XNOR2XL U79 ( .A(n51), .B(n95), .Y(n94) );
  OAI22X1 U80 ( .A(n29), .B(n5), .C(crc32_r_6_), .D(n63), .Y(n95) );
  OAI221X1 U81 ( .A(n13), .B(n109), .C(n22), .D(n7), .E(n9), .Y(N193) );
  XNOR2XL U82 ( .A(n110), .B(n71), .Y(n109) );
  XNOR2XL U83 ( .A(n51), .B(n111), .Y(n110) );
  OAI22X1 U84 ( .A(n22), .B(n6), .C(crc32_r_0_), .D(n63), .Y(n111) );
  OAI221X1 U85 ( .A(n13), .B(n87), .C(n24), .D(n8), .E(n10), .Y(N201) );
  XNOR2XL U86 ( .A(n88), .B(n71), .Y(n87) );
  XNOR2XL U87 ( .A(n89), .B(n18), .Y(n88) );
  AOI22X1 U88 ( .A(n68), .B(n24), .C(n51), .D(crc32_r_8_), .Y(n89) );
  NOR2X1 U89 ( .A(crc32_r_29_), .B(i_start), .Y(n119) );
  OAI221X1 U90 ( .A(n12), .B(n64), .C(n8), .D(n58), .E(n16), .Y(N214) );
  XNOR2XL U91 ( .A(n19), .B(n65), .Y(n64) );
  OAI22X1 U92 ( .A(n6), .B(n58), .C(crc32_r_21_), .D(n63), .Y(n65) );
  INVX1 U93 ( .A(crc32_r_21_), .Y(n58) );
  OAI221X1 U94 ( .A(n13), .B(n59), .C(n123), .D(n8), .E(n9), .Y(N215) );
  XNOR2XL U95 ( .A(n17), .B(n61), .Y(n59) );
  OAI22X1 U96 ( .A(n6), .B(n123), .C(crc32_r_22_), .D(n63), .Y(n61) );
  INVX1 U97 ( .A(crc32_r_22_), .Y(n123) );
  OAI221X1 U98 ( .A(n12), .B(n82), .C(n27), .D(n8), .E(n10), .Y(N203) );
  XNOR2XL U99 ( .A(n19), .B(n83), .Y(n82) );
  OAI22X1 U100 ( .A(n27), .B(n6), .C(crc32_r_10_), .D(n63), .Y(n83) );
  OAI221X1 U101 ( .A(n13), .B(n96), .C(n25), .D(n8), .E(n16), .Y(N198) );
  XNOR2XL U102 ( .A(n97), .B(n56), .Y(n96) );
  AOI22X1 U103 ( .A(n68), .B(n25), .C(n51), .D(crc32_r_5_), .Y(n97) );
  OAI221X1 U104 ( .A(n12), .B(n66), .C(n8), .D(n121), .E(n9), .Y(N213) );
  XNOR2XL U105 ( .A(n67), .B(n56), .Y(n66) );
  AOI22X1 U106 ( .A(n68), .B(n121), .C(crc32_r_20_), .D(n51), .Y(n67) );
  INVX1 U107 ( .A(crc32_r_20_), .Y(n121) );
  OAI221X1 U108 ( .A(n13), .B(n104), .C(n8), .D(n125), .E(n10), .Y(N195) );
  XNOR2XL U109 ( .A(n105), .B(n56), .Y(n104) );
  AOI22X1 U110 ( .A(n68), .B(n125), .C(crc32_r_2_), .D(n51), .Y(n105) );
  INVX1 U111 ( .A(crc32_r_2_), .Y(n125) );
  NAND2X1 U112 ( .A(n73), .B(n74), .Y(N211) );
  AOI32X1 U113 ( .A(n52), .B(n32), .C(n2), .D(crc32_r_18_), .E(n75), .Y(n73)
         );
  NAND2X1 U114 ( .A(n77), .B(n55), .Y(N206) );
  AOI32X1 U115 ( .A(n52), .B(n124), .C(n1), .D(crc32_r_13_), .E(n57), .Y(n77)
         );
  INVX1 U116 ( .A(crc32_r_13_), .Y(n124) );
  NAND2X1 U117 ( .A(n54), .B(n55), .Y(N216) );
  AOI32X1 U118 ( .A(n52), .B(n126), .C(n1), .D(crc32_r_23_), .E(n57), .Y(n54)
         );
  INVX1 U119 ( .A(crc32_r_23_), .Y(n126) );
  NAND2X1 U120 ( .A(n79), .B(n74), .Y(N205) );
  AOI32X1 U121 ( .A(n52), .B(n30), .C(n2), .D(crc32_r_12_), .E(n75), .Y(n79)
         );
  OAI221X1 U122 ( .A(crc32_r_15_), .B(n46), .C(n21), .D(n47), .E(n48), .Y(N208) );
  OAI221X1 U123 ( .A(crc32_r_25_), .B(n46), .C(n33), .D(n47), .E(n48), .Y(N218) );
  INVX1 U124 ( .A(crc32_r_25_), .Y(n33) );
  OAI221X1 U125 ( .A(crc32_r_11_), .B(n46), .C(n20), .D(n47), .E(n48), .Y(N204) );
  OAI221X1 U126 ( .A(n12), .B(n69), .C(n8), .D(n127), .E(n16), .Y(N212) );
  INVX1 U127 ( .A(crc32_r_19_), .Y(n127) );
  XNOR2XL U128 ( .A(n70), .B(n71), .Y(n69) );
  XNOR2XL U129 ( .A(n72), .B(n56), .Y(n70) );
  NOR2X1 U130 ( .A(crc32_r_19_), .B(i_start), .Y(n72) );
  NOR2X1 U131 ( .A(crc32_r_28_), .B(i_start), .Y(n120) );
  NAND3X1 U132 ( .A(n49), .B(n10), .C(n50), .Y(N217) );
  AOI32X1 U133 ( .A(n3), .B(n34), .C(n52), .D(crc32_r_24_), .E(n53), .Y(n50)
         );
  INVX1 U134 ( .A(crc32_r_24_), .Y(n34) );
  NAND3X1 U135 ( .A(n49), .B(n16), .C(n76), .Y(N207) );
  AOI32X1 U136 ( .A(n3), .B(n31), .C(n52), .D(crc32_r_14_), .E(n53), .Y(n76)
         );
  OAI21BBX1 U137 ( .A(N188), .B(crc32_r_26_), .C(n15), .Y(N219) );
  OAI21BBX1 U138 ( .A(N188), .B(crc32_r_27_), .C(n15), .Y(N220) );
  OAI21BBX1 U139 ( .A(N188), .B(crc32_r_16_), .C(n15), .Y(N209) );
  OAI21BBX1 U140 ( .A(N188), .B(crc32_r_17_), .C(n15), .Y(N210) );
  NOR2X1 U141 ( .A(n36), .B(n37), .Y(rx_good) );
  NAND4X1 U142 ( .A(n38), .B(n39), .C(n40), .D(n41), .Y(n37) );
  NAND4X1 U143 ( .A(n42), .B(n43), .C(n44), .D(n45), .Y(n36) );
  AND4X1 U144 ( .A(crc32_r_24_), .B(crc32_r_25_), .C(crc32_r_26_), .D(
        crc32_r_3_), .Y(n39) );
  NOR4XL U145 ( .A(crc32_r_9_), .B(crc32_r_7_), .C(crc32_r_2_), .D(crc32_r_29_), .Y(n45) );
  NOR4XL U146 ( .A(crc32_r_28_), .B(crc32_r_27_), .C(crc32_r_23_), .D(
        crc32_r_22_), .Y(n44) );
  NOR4XL U147 ( .A(crc32_r_21_), .B(crc32_r_20_), .C(crc32_r_19_), .D(
        crc32_r_17_), .Y(n43) );
  NOR4XL U148 ( .A(crc32_r_16_), .B(crc32_r_13_), .C(crc32_3_0[1]), .D(
        crc32_3_0[0]), .Y(n42) );
  INVX1 U149 ( .A(crc32_r_30_), .Y(crc32_3_0[1]) );
  INVX1 U150 ( .A(test_so), .Y(crc32_3_0[0]) );
  INVX1 U151 ( .A(crc32_r_6_), .Y(n29) );
  INVX1 U152 ( .A(crc32_r_1_), .Y(n26) );
  INVX1 U153 ( .A(crc32_r_10_), .Y(n27) );
  INVX1 U154 ( .A(crc32_r_8_), .Y(n24) );
  INVX1 U155 ( .A(crc32_r_18_), .Y(n32) );
  INVX1 U156 ( .A(crc32_r_12_), .Y(n30) );
  INVX1 U157 ( .A(crc32_r_11_), .Y(n20) );
  INVX1 U158 ( .A(crc32_r_15_), .Y(n21) );
  INVX1 U159 ( .A(crc32_r_28_), .Y(crc32_3_0[3]) );
  INVX1 U160 ( .A(crc32_r_29_), .Y(crc32_3_0[2]) );
  INVX1 U161 ( .A(crc32_r_4_), .Y(n23) );
  INVX1 U162 ( .A(crc32_r_0_), .Y(n22) );
  INVX1 U163 ( .A(crc32_r_5_), .Y(n25) );
  INVX1 U164 ( .A(crc32_r_14_), .Y(n31) );
  INVX1 U165 ( .A(crc32_r_7_), .Y(n122) );
  INVX1 U166 ( .A(crc32_r_9_), .Y(n35) );
  INVX1 U167 ( .A(crc32_r_3_), .Y(n28) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phycrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phytx_a0 ( r_txnumk, r_txendk, r_txshrt, r_txauto, prx_cccnt, ptx_txact, 
        ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, i_rdat, i_txreq, i_one, 
        ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4, ptx_crcsidat, ptx_fsm, 
        pcc_crc30, clk, srstz, test_si, test_se );
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [1:0] prx_cccnt;
  input [7:0] i_rdat;
  output [3:0] ptx_crcsidat;
  output [2:0] ptx_fsm;
  input [3:0] pcc_crc30;
  input r_txendk, r_txshrt, i_txreq, i_one, clk, srstz, test_si, test_se;
  output ptx_txact, ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, ptx_crcstart,
         ptx_crcshfi4, ptx_crcshfo4;
  wire   hinib, N251, N254, N255, N268, N270, N271, N272, N273, N297, N298,
         N299, net10645, net10651, n237, n238, n120, n126, n134, n135, n137,
         n154, n156, n157, n171, n190, n191, n1, n2, n3, n4, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n121, n122, n123, n124, n125, n127, n128, n129, n130,
         n131, n132, n133, n136, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n155, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314;
  wire   [4:0] bytcnt;
  wire   [3:0] bitcnt;

  SNPS_CLOCK_GATE_HIGH_phytx_a0_0 clk_gate_bitcnt_reg ( .CLK(clk), .EN(N251), 
        .ENCLK(net10645), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phytx_a0_1 clk_gate_bytcnt_reg ( .CLK(clk), .EN(N268), 
        .ENCLK(net10651), .TE(test_se) );
  SDFFQX1 ptx_cc_reg ( .D(n238), .SIN(n25), .SMC(test_se), .C(clk), .Q(ptx_cc)
         );
  SDFFQX1 bitcnt_reg_1_ ( .D(n307), .SIN(bitcnt[0]), .SMC(test_se), .C(
        net10645), .Q(bitcnt[1]) );
  SDFFQX1 bitcnt_reg_0_ ( .D(n304), .SIN(test_si), .SMC(test_se), .C(net10645), 
        .Q(bitcnt[0]) );
  SDFFQX1 bytcnt_reg_4_ ( .D(N273), .SIN(bytcnt[3]), .SMC(test_se), .C(
        net10651), .Q(bytcnt[4]) );
  SDFFQX1 bitcnt_reg_3_ ( .D(N255), .SIN(bitcnt[2]), .SMC(test_se), .C(
        net10645), .Q(bitcnt[3]) );
  SDFFQX1 bytcnt_reg_1_ ( .D(N270), .SIN(bytcnt[0]), .SMC(test_se), .C(
        net10651), .Q(bytcnt[1]) );
  SDFFQX1 bytcnt_reg_3_ ( .D(N272), .SIN(bytcnt[2]), .SMC(test_se), .C(
        net10651), .Q(bytcnt[3]) );
  SDFFQX1 cs_txph_reg_0_ ( .D(N297), .SIN(bytcnt[4]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[0]) );
  SDFFQX1 hinib_reg ( .D(n237), .SIN(ptx_fsm[2]), .SMC(test_se), .C(net10645), 
        .Q(hinib) );
  SDFFQX1 bitcnt_reg_2_ ( .D(N254), .SIN(bitcnt[1]), .SMC(test_se), .C(
        net10645), .Q(bitcnt[2]) );
  SDFFQX1 cs_txph_reg_1_ ( .D(N298), .SIN(ptx_fsm[0]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[1]) );
  SDFFQX1 bytcnt_reg_0_ ( .D(n305), .SIN(bitcnt[3]), .SMC(test_se), .C(
        net10651), .Q(bytcnt[0]) );
  SDFFQX1 bytcnt_reg_2_ ( .D(N271), .SIN(bytcnt[1]), .SMC(test_se), .C(
        net10651), .Q(bytcnt[2]) );
  SDFFQX1 cs_txph_reg_2_ ( .D(N299), .SIN(ptx_fsm[1]), .SMC(test_se), .C(clk), 
        .Q(ptx_fsm[2]) );
  INVX2 U3 ( .A(n283), .Y(n48) );
  INVXL U4 ( .A(n280), .Y(n55) );
  INVXL U5 ( .A(n296), .Y(n26) );
  AND2XL U6 ( .A(r_txnumk[3]), .B(n147), .Y(n51) );
  NAND21XL U7 ( .B(r_txnumk[3]), .A(bytcnt[3]), .Y(n280) );
  NAND21XL U8 ( .B(bytcnt[0]), .A(r_txnumk[0]), .Y(n45) );
  NOR21X1 U9 ( .B(r_txnumk[1]), .A(bytcnt[1]), .Y(n46) );
  MUX2IX4 U10 ( .D0(i_rdat[0]), .D1(i_rdat[4]), .S(hinib), .Y(n174) );
  MUX2IX4 U11 ( .D0(i_rdat[2]), .D1(i_rdat[6]), .S(hinib), .Y(n169) );
  INVX2 U12 ( .A(n4), .Y(n19) );
  INVX2 U13 ( .A(n23), .Y(n103) );
  NAND42X2 U14 ( .C(n71), .D(n70), .A(n69), .B(n68), .Y(n82) );
  NAND21X4 U15 ( .B(n207), .A(n63), .Y(n204) );
  NOR41X2 U16 ( .D(n32), .A(n103), .B(n302), .C(n33), .Y(n31) );
  NAND31X1 U17 ( .C(n67), .A(n260), .B(n296), .Y(n68) );
  INVX1 U18 ( .A(r_txendk), .Y(n11) );
  NOR21X1 U19 ( .B(r_txnumk[4]), .A(n44), .Y(n57) );
  NOR21XL U20 ( .B(bytcnt[4]), .A(n43), .Y(n44) );
  AND4X1 U21 ( .A(r_txnumk[2]), .B(r_txnumk[3]), .C(r_txnumk[0]), .D(
        r_txnumk[1]), .Y(n43) );
  NAND32X1 U22 ( .B(n55), .C(n54), .A(n53), .Y(n56) );
  INVX2 U23 ( .A(i_rdat[5]), .Y(n102) );
  NAND2X1 U24 ( .A(n100), .B(n1), .Y(n2) );
  INVX1 U25 ( .A(n104), .Y(n32) );
  INVX1 U26 ( .A(ptx_fsm[0]), .Y(n122) );
  INVX1 U27 ( .A(n132), .Y(n207) );
  NAND21X1 U28 ( .B(ptx_fsm[1]), .A(n122), .Y(n228) );
  INVX1 U29 ( .A(bytcnt[3]), .Y(n147) );
  NAND21X1 U30 ( .B(n39), .A(prx_cccnt[0]), .Y(n266) );
  INVXL U31 ( .A(i_rdat[0]), .Y(n20) );
  NAND2X1 U32 ( .A(n2), .B(n3), .Y(n4) );
  NAND2X1 U33 ( .A(n189), .B(n179), .Y(n3) );
  NAND21X2 U34 ( .B(ptx_crcsidat[1]), .A(n61), .Y(n67) );
  MUX2IX2 U35 ( .D0(n60), .D1(ptx_crcsidat[2]), .S(n19), .Y(n61) );
  INVX2 U36 ( .A(i_rdat[1]), .Y(n97) );
  INVX1 U37 ( .A(i_rdat[4]), .Y(n98) );
  INVXL U38 ( .A(n179), .Y(n1) );
  INVX2 U39 ( .A(i_rdat[3]), .Y(n189) );
  NOR2X1 U40 ( .A(ptx_fsm[2]), .B(n228), .Y(n39) );
  INVX1 U41 ( .A(n39), .Y(ptx_txact) );
  INVXL U42 ( .A(i_rdat[6]), .Y(n101) );
  INVXL U43 ( .A(i_rdat[2]), .Y(n96) );
  INVX1 U44 ( .A(n288), .Y(n296) );
  INVX1 U45 ( .A(bitcnt[2]), .Y(n24) );
  INVXL U46 ( .A(n19), .Y(n205) );
  INVX1 U47 ( .A(n205), .Y(ptx_crcsidat[3]) );
  INVX1 U48 ( .A(ptx_crcsidat[0]), .Y(n6) );
  INVXL U49 ( .A(n169), .Y(ptx_crcsidat[2]) );
  INVX1 U50 ( .A(n10), .Y(n7) );
  NAND2X1 U51 ( .A(n204), .B(n16), .Y(n14) );
  NAND3X2 U52 ( .A(n22), .B(n21), .C(n56), .Y(n58) );
  NOR21X1 U53 ( .B(n288), .A(n64), .Y(n70) );
  INVX1 U54 ( .A(n204), .Y(n13) );
  OA33X1 U55 ( .A(n66), .B(n65), .C(n64), .D(n288), .E(r_txauto[6]), .F(
        bitcnt[0]), .Y(n69) );
  BUFX1 U56 ( .A(n302), .Y(n8) );
  NOR41XL U57 ( .D(n32), .A(n7), .B(n8), .C(n33), .Y(n9) );
  INVXL U58 ( .A(n103), .Y(n10) );
  INVX2 U59 ( .A(n57), .Y(n21) );
  NAND21X2 U60 ( .B(n11), .A(i_one), .Y(n22) );
  NAND21X2 U61 ( .B(n288), .A(n62), .Y(n63) );
  NAND21X2 U62 ( .B(n290), .A(n58), .Y(n288) );
  BUFXL U63 ( .A(n204), .Y(n12) );
  NAND2X1 U64 ( .A(n13), .B(bitcnt[1]), .Y(n15) );
  NAND2X2 U65 ( .A(n14), .B(n15), .Y(n302) );
  INVX1 U66 ( .A(bitcnt[1]), .Y(n16) );
  NAND21X1 U67 ( .B(n8), .A(n301), .Y(n303) );
  BUFXL U68 ( .A(n20), .Y(n17) );
  INVXL U69 ( .A(n17), .Y(n18) );
  NAND21X2 U70 ( .B(n169), .A(n174), .Y(n60) );
  INVX2 U71 ( .A(i_rdat[7]), .Y(n100) );
  NAND2X2 U72 ( .A(n67), .B(r_txauto[6]), .Y(n62) );
  NAND6XL U73 ( .A(n99), .B(n98), .C(n97), .D(n96), .E(n189), .F(i_one), .Y(
        n104) );
  XOR2X1 U74 ( .A(n204), .B(n24), .Y(n23) );
  INVX1 U75 ( .A(n179), .Y(n25) );
  NAND21XL U76 ( .B(n264), .A(ptx_txact), .Y(n265) );
  INVXL U77 ( .A(ptx_fsm[2]), .Y(n109) );
  INVXL U78 ( .A(n287), .Y(n54) );
  NAND21X1 U79 ( .B(r_txnumk[2]), .A(bytcnt[2]), .Y(n282) );
  AO44X1 U80 ( .A(n23), .B(n299), .C(n298), .D(n300), .E(n297), .F(n296), .G(
        n295), .H(n294), .Y(n301) );
  INVXL U81 ( .A(bytcnt[1]), .Y(n142) );
  NAND21XL U82 ( .B(n296), .A(n236), .Y(n247) );
  INVX2 U83 ( .A(n199), .Y(n233) );
  NAND21XL U84 ( .B(n9), .A(n105), .Y(n106) );
  NAND4XL U85 ( .A(n102), .B(n101), .C(n100), .D(n17), .Y(n33) );
  NAND2XL U86 ( .A(n34), .B(r_txauto[6]), .Y(n295) );
  INVX1 U87 ( .A(n73), .Y(n294) );
  OAI211XL U88 ( .C(n140), .D(n146), .A(n306), .B(n139), .Y(n171) );
  OAI211XL U89 ( .C(n116), .D(n167), .A(n115), .B(n114), .Y(n291) );
  AOI211XL U90 ( .C(n148), .D(n147), .A(n171), .B(n150), .Y(N272) );
  NAND32XL U91 ( .B(n260), .C(n16), .A(n275), .Y(n79) );
  AOI31XL U92 ( .A(n233), .B(n91), .C(n142), .D(ptx_goidle), .Y(n92) );
  MUX2X1 U93 ( .D0(n262), .D1(n263), .S(n27), .Y(n264) );
  XNOR2XL U94 ( .A(n24), .B(n261), .Y(n27) );
  NAND31XL U95 ( .C(n6), .A(r_txauto[6]), .B(n168), .Y(n206) );
  AO21XL U96 ( .B(n259), .C(n260), .A(n165), .Y(n208) );
  NAND21XL U97 ( .B(n228), .A(n284), .Y(n105) );
  MUX2AXL U98 ( .D0(n28), .D1(n254), .S(n253), .Y(n256) );
  OAI21X1 U99 ( .B(n252), .C(n251), .A(n250), .Y(n28) );
  OA21XL U100 ( .B(n120), .C(n234), .A(n233), .Y(n235) );
  NAND21XL U101 ( .B(r_txauto[6]), .A(n168), .Y(n192) );
  NAND32XL U102 ( .B(n167), .C(n109), .A(n122), .Y(n131) );
  AO21XL U103 ( .B(n260), .C(n16), .A(n259), .Y(n261) );
  OR2XL U104 ( .A(n147), .B(n148), .Y(n146) );
  NAND21X1 U105 ( .B(r_txnumk[1]), .A(bytcnt[1]), .Y(n283) );
  NAND32X1 U106 ( .B(n52), .C(n51), .A(n50), .Y(n53) );
  NAND32X1 U107 ( .B(ptx_fsm[0]), .C(n167), .A(n109), .Y(n290) );
  INVX1 U108 ( .A(n72), .Y(n83) );
  INVX1 U109 ( .A(n74), .Y(n300) );
  OAI21BBX1 U110 ( .A(n179), .B(n16), .C(n29), .Y(n250) );
  MUX2IX1 U111 ( .D0(n158), .D1(n165), .S(n155), .Y(n29) );
  INVX1 U112 ( .A(n247), .Y(n223) );
  INVX1 U113 ( .A(n42), .Y(n41) );
  INVX1 U114 ( .A(n266), .Y(n298) );
  INVX1 U115 ( .A(n77), .Y(n275) );
  NAND21X1 U116 ( .B(n266), .A(n274), .Y(n77) );
  NAND21X1 U117 ( .B(n275), .A(n274), .Y(N251) );
  INVX1 U118 ( .A(n133), .Y(n277) );
  INVX1 U119 ( .A(n173), .Y(n193) );
  AND2X1 U120 ( .A(n217), .B(n247), .Y(n184) );
  AND2X1 U121 ( .A(n241), .B(n193), .Y(n185) );
  INVX1 U122 ( .A(n217), .Y(n220) );
  INVX1 U123 ( .A(n107), .Y(n138) );
  INVX1 U124 ( .A(n190), .Y(n310) );
  INVX1 U125 ( .A(srstz), .Y(n42) );
  INVX1 U126 ( .A(n171), .Y(n149) );
  INVX1 U127 ( .A(n76), .Y(n274) );
  NAND32X1 U128 ( .B(i_txreq), .C(n107), .A(n105), .Y(n76) );
  INVX1 U129 ( .A(i_txreq), .Y(n267) );
  AND2X1 U130 ( .A(n41), .B(n291), .Y(N298) );
  AND2X1 U131 ( .A(n278), .B(n279), .Y(ptx_crcshfo4) );
  INVX1 U132 ( .A(n276), .Y(n284) );
  NAND32XL U133 ( .B(n266), .C(n81), .A(n10), .Y(n133) );
  NAND21X1 U134 ( .B(n170), .A(n216), .Y(n173) );
  NAND21X1 U135 ( .B(n173), .A(n248), .Y(n217) );
  OAI31XL U136 ( .A(n75), .B(n26), .C(n276), .D(n133), .Y(n107) );
  INVX1 U137 ( .A(n295), .Y(n75) );
  INVX1 U138 ( .A(n159), .Y(n168) );
  INVX1 U139 ( .A(n206), .Y(n255) );
  NAND21X1 U140 ( .B(n277), .A(n276), .Y(n279) );
  INVX1 U141 ( .A(n170), .Y(n236) );
  AND2X1 U142 ( .A(n218), .B(n245), .Y(n219) );
  INVX1 U143 ( .A(n172), .Y(n245) );
  NAND21X1 U144 ( .B(n248), .A(n193), .Y(n172) );
  INVX1 U145 ( .A(n209), .Y(n225) );
  NAND21X1 U146 ( .B(n254), .A(n253), .Y(n209) );
  INVX1 U147 ( .A(n183), .Y(n241) );
  INVX1 U148 ( .A(n208), .Y(n253) );
  INVX1 U149 ( .A(n192), .Y(n258) );
  INVX1 U150 ( .A(n157), .Y(n309) );
  AND2X1 U151 ( .A(n41), .B(n289), .Y(N299) );
  INVX1 U152 ( .A(n106), .Y(n121) );
  INVX1 U153 ( .A(n134), .Y(n311) );
  INVX1 U154 ( .A(n188), .Y(n249) );
  NAND21X1 U155 ( .B(n215), .A(n218), .Y(n188) );
  INVX1 U156 ( .A(n81), .Y(n85) );
  MUX2AXL U157 ( .D0(n126), .D1(n30), .S(n194), .Y(n161) );
  NAND2X1 U158 ( .A(n309), .B(n135), .Y(n30) );
  INVX1 U159 ( .A(n131), .Y(n278) );
  NAND4X1 U160 ( .A(n135), .B(n126), .C(n134), .D(n191), .Y(n190) );
  NOR3XL U161 ( .A(n137), .B(n120), .C(n157), .Y(n191) );
  AND2X1 U162 ( .A(n311), .B(n314), .Y(n162) );
  INVX1 U163 ( .A(n126), .Y(n313) );
  INVX1 U164 ( .A(n135), .Y(n178) );
  INVX1 U165 ( .A(n146), .Y(n150) );
  INVX1 U166 ( .A(n289), .Y(n292) );
  INVX2 U167 ( .A(n82), .Y(n297) );
  INVX1 U168 ( .A(n166), .Y(ptx_crcsidat[1]) );
  INVX1 U169 ( .A(n282), .Y(n49) );
  NAND4XL U170 ( .A(n102), .B(n98), .C(n101), .D(n100), .Y(n34) );
  NAND32X1 U171 ( .B(n122), .C(n167), .A(n109), .Y(n199) );
  NAND21XL U172 ( .B(n266), .A(n83), .Y(n73) );
  INVX1 U173 ( .A(n290), .Y(n299) );
  OAI22X1 U174 ( .A(n138), .B(n290), .C(n136), .D(n133), .Y(n139) );
  AND3XL U175 ( .A(n199), .B(n132), .C(n131), .Y(n136) );
  AND2X1 U176 ( .A(n121), .B(n119), .Y(n124) );
  OAI211XL U177 ( .C(r_txauto[3]), .D(n190), .A(i_txreq), .B(n39), .Y(n119) );
  INVX1 U178 ( .A(n271), .Y(n293) );
  OA22XL U179 ( .A(n9), .B(n199), .C(n118), .D(n113), .Y(n114) );
  AOI221XL U180 ( .A(n278), .B(n117), .C(n299), .D(n118), .E(n111), .Y(n116)
         );
  AOI32XL U181 ( .A(n308), .B(i_txreq), .C(n39), .D(n207), .E(n112), .Y(n115)
         );
  AOI211X1 U182 ( .C(n281), .D(n142), .A(n171), .B(n141), .Y(N270) );
  INVX1 U183 ( .A(n143), .Y(n141) );
  INVX1 U184 ( .A(n151), .Y(n305) );
  NAND2X1 U185 ( .A(n306), .B(n171), .Y(N268) );
  AO21X1 U186 ( .B(n275), .C(n16), .A(n304), .Y(n272) );
  INVX1 U187 ( .A(n79), .Y(n273) );
  OA21XL U188 ( .B(r_txnumk[0]), .C(n281), .A(n280), .Y(n286) );
  AND2X1 U189 ( .A(n41), .B(n271), .Y(N297) );
  AND3XL U190 ( .A(n299), .B(n26), .C(n279), .Y(ptx_crcshfi4) );
  NAND21X1 U191 ( .B(n142), .A(n91), .Y(n117) );
  AND4XL U192 ( .A(n284), .B(n299), .C(n283), .D(n282), .Y(n285) );
  INVX1 U193 ( .A(n93), .Y(n111) );
  NAND43X1 U194 ( .B(n207), .C(n299), .D(n278), .A(n92), .Y(n93) );
  AOI21BXL U195 ( .C(n112), .B(n207), .A(n111), .Y(n35) );
  OAI211X1 U196 ( .C(n110), .D(n109), .A(n121), .B(n118), .Y(n289) );
  AND2X1 U197 ( .A(n35), .B(n131), .Y(n110) );
  GEN2XL U198 ( .D(n231), .E(n230), .C(n229), .B(n228), .A(n227), .Y(n263) );
  AND4X1 U199 ( .A(n232), .B(n206), .C(n226), .D(n208), .Y(n231) );
  AND4X1 U200 ( .A(n226), .B(n250), .C(n225), .D(n224), .Y(n227) );
  MUX2BXL U201 ( .D0(n213), .D1(n212), .S(n232), .Y(n229) );
  AOI211X1 U202 ( .C(n258), .D(n257), .A(n256), .B(n255), .Y(n262) );
  NAND32X1 U203 ( .B(n108), .C(n290), .A(n107), .Y(n118) );
  INVXL U204 ( .A(i_one), .Y(n108) );
  AO21X1 U205 ( .B(i_rdat[4]), .C(n258), .A(n242), .Y(n252) );
  OAI31XL U206 ( .A(n249), .B(n248), .C(n247), .D(n246), .Y(n251) );
  AOI221XL U207 ( .A(n215), .B(n223), .C(i_rdat[2]), .D(n258), .E(n177), .Y(
        n230) );
  MUX2X1 U208 ( .D0(n176), .D1(n175), .S(n218), .Y(n177) );
  AND2XL U209 ( .A(n245), .B(n26), .Y(n176) );
  OAI22XL U210 ( .A(n244), .B(n173), .C(n26), .D(n217), .Y(n175) );
  AOI31XL U211 ( .A(n245), .B(n296), .C(n244), .D(n243), .Y(n246) );
  AOI211XL U212 ( .C(n18), .D(n258), .A(n187), .B(n186), .Y(n213) );
  OAI211XL U213 ( .C(n182), .D(n199), .A(n181), .B(n208), .Y(n187) );
  MUX2BXL U214 ( .D0(n185), .D1(n184), .S(n218), .Y(n186) );
  AOI221XL U215 ( .A(n194), .B(n120), .C(n179), .D(n178), .E(n313), .Y(n182)
         );
  MUX2IX1 U216 ( .D0(n36), .D1(n37), .S(n253), .Y(n257) );
  NAND2XL U217 ( .A(i_rdat[6]), .B(n232), .Y(n36) );
  MUX2IX1 U218 ( .D0(i_rdat[5]), .D1(i_rdat[7]), .S(n232), .Y(n37) );
  AOI221XL U219 ( .A(n223), .B(n222), .C(i_rdat[1]), .D(n258), .E(n221), .Y(
        n224) );
  OAI22X1 U220 ( .A(n216), .B(n248), .C(n215), .D(n214), .Y(n222) );
  MUX2X1 U221 ( .D0(n220), .D1(n219), .S(n241), .Y(n221) );
  AND2X1 U222 ( .A(n218), .B(n216), .Y(n214) );
  OR2XL U223 ( .A(n260), .B(n12), .Y(n152) );
  INVX1 U224 ( .A(n243), .Y(n181) );
  NAND32X1 U225 ( .B(n211), .C(n210), .A(n225), .Y(n212) );
  GEN2XL U226 ( .D(n249), .E(n203), .C(n26), .B(n202), .A(n201), .Y(n210) );
  OAI22X1 U227 ( .A(n192), .B(n189), .C(n249), .D(n217), .Y(n211) );
  OAI22XL U228 ( .A(n200), .B(n199), .C(n247), .D(n203), .Y(n201) );
  INVX1 U229 ( .A(n250), .Y(n232) );
  AND2X1 U230 ( .A(n193), .B(n244), .Y(n202) );
  GEN2XL U231 ( .D(n241), .E(n240), .C(n239), .B(n236), .A(n235), .Y(n242) );
  NAND3X1 U232 ( .A(r_txauto[1]), .B(n314), .C(r_txauto[2]), .Y(n126) );
  INVX1 U233 ( .A(r_txauto[0]), .Y(n314) );
  NAND2X1 U234 ( .A(r_txauto[1]), .B(n312), .Y(n134) );
  NAND31XL U235 ( .C(n207), .A(n38), .B(n206), .Y(n254) );
  NAND3XL U236 ( .A(r_txauto[6]), .B(n205), .C(n12), .Y(n38) );
  NOR3XL U237 ( .A(r_txauto[0]), .B(r_txauto[1]), .C(n312), .Y(n157) );
  NAND3X1 U238 ( .A(r_txauto[2]), .B(r_txauto[1]), .C(r_txauto[0]), .Y(n135)
         );
  INVX1 U239 ( .A(r_txauto[2]), .Y(n312) );
  INVX1 U240 ( .A(n239), .Y(n216) );
  INVX1 U241 ( .A(n203), .Y(n248) );
  INVX1 U242 ( .A(n244), .Y(n215) );
  NOR3XL U243 ( .A(n312), .B(r_txauto[1]), .C(n314), .Y(n137) );
  AOI211X1 U244 ( .C(n120), .D(n198), .A(n197), .B(n234), .Y(n200) );
  INVX1 U245 ( .A(n240), .Y(n218) );
  NOR3XL U246 ( .A(r_txauto[1]), .B(r_txauto[2]), .C(n314), .Y(n120) );
  INVX1 U247 ( .A(n198), .Y(n194) );
  INVX1 U248 ( .A(r_txauto[4]), .Y(n113) );
  INVX1 U249 ( .A(r_txauto[3]), .Y(n308) );
  AND4X1 U250 ( .A(n293), .B(n292), .C(n291), .D(n290), .Y(ptx_pspyld) );
  NOR2XL U251 ( .A(bitcnt[0]), .B(n132), .Y(n71) );
  MUX2X2 U252 ( .D0(n97), .D1(n102), .S(hinib), .Y(n166) );
  NAND21X1 U253 ( .B(r_txnumk[4]), .A(bytcnt[4]), .Y(n287) );
  NOR21XL U254 ( .B(r_txnumk[2]), .A(bytcnt[2]), .Y(n52) );
  NAND32X1 U255 ( .B(n49), .C(n48), .A(n47), .Y(n50) );
  NAND21X1 U256 ( .B(n46), .A(n45), .Y(n47) );
  INVX1 U257 ( .A(r_txauto[6]), .Y(n65) );
  INVXL U258 ( .A(n67), .Y(n66) );
  AND4XL U259 ( .A(n95), .B(n233), .C(r_txendk), .D(n298), .Y(n99) );
  AND4XL U260 ( .A(bitcnt[3]), .B(n147), .C(bytcnt[0]), .D(n94), .Y(n95) );
  AND4X1 U261 ( .A(n140), .B(n144), .C(bitcnt[0]), .D(n142), .Y(n94) );
  INVXL U262 ( .A(ptx_fsm[1]), .Y(n167) );
  NAND32XL U263 ( .B(ptx_fsm[1]), .C(n122), .A(n109), .Y(n132) );
  NAND21XL U264 ( .B(n207), .A(bitcnt[0]), .Y(n64) );
  INVXL U265 ( .A(bytcnt[2]), .Y(n144) );
  INVXL U266 ( .A(bytcnt[4]), .Y(n140) );
  NAND21XL U267 ( .B(bitcnt[3]), .A(bitcnt[2]), .Y(n72) );
  INVXL U268 ( .A(bitcnt[0]), .Y(n260) );
  NAND21XL U269 ( .B(n260), .A(bitcnt[3]), .Y(n74) );
  NOR21XL U270 ( .B(n267), .A(n130), .Y(n306) );
  NAND31X1 U271 ( .C(n129), .A(n128), .B(n127), .Y(n130) );
  NOR21XL U272 ( .B(n289), .A(ptx_fsm[2]), .Y(n129) );
  XNOR2XL U273 ( .A(ptx_fsm[1]), .B(n291), .Y(n128) );
  NAND21XL U274 ( .B(bytcnt[0]), .A(n149), .Y(n151) );
  OAI211X1 U275 ( .C(r_txauto[5]), .D(n125), .A(n124), .B(n123), .Y(n271) );
  OA22X1 U276 ( .A(r_txauto[4]), .B(n118), .C(n131), .D(n117), .Y(n125) );
  OA22XL U277 ( .A(n35), .B(n122), .C(n310), .D(n132), .Y(n123) );
  XOR2XL U278 ( .A(ptx_fsm[0]), .B(n293), .Y(n127) );
  OAI22XL U279 ( .A(n171), .B(n145), .C(n144), .D(n151), .Y(N271) );
  MUX2XL U280 ( .D0(n143), .D1(bytcnt[1]), .S(bytcnt[2]), .Y(n145) );
  OA21XL U281 ( .B(bytcnt[4]), .C(n150), .A(n149), .Y(N273) );
  GEN2XL U282 ( .D(n275), .E(n24), .C(n272), .B(bitcnt[3]), .A(n80), .Y(N255)
         );
  AND2XL U283 ( .A(n273), .B(n83), .Y(n80) );
  MUX2XL U284 ( .D0(n273), .D1(n272), .S(bitcnt[2]), .Y(N254) );
  MUX2AXL U285 ( .D0(n40), .D1(n304), .S(bitcnt[1]), .Y(n307) );
  NAND2XL U286 ( .A(n275), .B(bitcnt[0]), .Y(n40) );
  INVX1 U287 ( .A(n78), .Y(n304) );
  NAND21XL U288 ( .B(bitcnt[0]), .A(n275), .Y(n78) );
  INVXL U289 ( .A(n174), .Y(ptx_crcsidat[0]) );
  MUX2XL U290 ( .D0(n87), .D1(n25), .S(n86), .Y(n237) );
  AOI211XL U291 ( .C(n10), .D(n85), .A(i_txreq), .B(n84), .Y(n86) );
  AND3X1 U292 ( .A(n138), .B(n284), .C(n267), .Y(n87) );
  AND4XL U293 ( .A(n83), .B(n155), .C(n297), .D(n228), .Y(n84) );
  MUX2X1 U294 ( .D0(n270), .D1(ptx_cc), .S(n269), .Y(n238) );
  NAND21X1 U295 ( .B(n42), .A(ptx_cc), .Y(n270) );
  AND3X1 U296 ( .A(n41), .B(n268), .C(n267), .Y(n269) );
  MUX2XL U297 ( .D0(n266), .D1(n265), .S(prx_cccnt[1]), .Y(n268) );
  OAI21BBX1 U298 ( .A(r_txshrt), .B(n277), .C(n117), .Y(n112) );
  INVX1 U299 ( .A(n88), .Y(n91) );
  NAND5XL U300 ( .A(bytcnt[0]), .B(n277), .C(n144), .D(n140), .E(n147), .Y(n88) );
  GEN2XL U301 ( .D(n137), .E(n25), .C(n197), .B(n233), .A(n255), .Y(n243) );
  AND2XL U302 ( .A(n25), .B(n152), .Y(n158) );
  INVX1 U303 ( .A(n153), .Y(n165) );
  NAND21XL U304 ( .B(n152), .A(n25), .Y(n153) );
  MUX2XL U305 ( .D0(n19), .D1(pcc_crc30[3]), .S(n278), .Y(n239) );
  MUX2BXL U306 ( .D0(n166), .D1(pcc_crc30[1]), .S(n278), .Y(n244) );
  MUX2BXL U307 ( .D0(n169), .D1(pcc_crc30[2]), .S(n278), .Y(n203) );
  MUX2BXL U308 ( .D0(n6), .D1(pcc_crc30[0]), .S(n278), .Y(n240) );
  OAI221XL U309 ( .A(n154), .B(n25), .C(n156), .D(bytcnt[0]), .E(n196), .Y(
        n234) );
  AOI21X1 U310 ( .B(n311), .C(r_txauto[0]), .A(n157), .Y(n154) );
  AOI21X1 U311 ( .B(n314), .C(n311), .A(n137), .Y(n156) );
  MUX2X1 U312 ( .D0(n195), .D1(n126), .S(n194), .Y(n196) );
  NAND21XL U313 ( .B(n135), .A(n25), .Y(n195) );
  INVX1 U314 ( .A(n180), .Y(n197) );
  OAI211XL U315 ( .C(bytcnt[0]), .D(n25), .A(n198), .B(n157), .Y(n180) );
  INVX1 U316 ( .A(n90), .Y(ptx_goidle) );
  NAND5XL U317 ( .A(ptx_fsm[2]), .B(ptx_fsm[0]), .C(n298), .D(n167), .E(n89), 
        .Y(n90) );
  INVX1 U318 ( .A(ptx_cc), .Y(n89) );
  OAI21X1 U319 ( .B(n164), .C(n163), .A(n233), .Y(n226) );
  MUX2XL U320 ( .D0(n178), .D1(n160), .S(n25), .Y(n164) );
  GEN2XL U321 ( .D(n137), .E(n179), .C(n162), .B(bytcnt[0]), .A(n161), .Y(n163) );
  AND2X1 U322 ( .A(r_txauto[0]), .B(n311), .Y(n160) );
  NAND21XL U323 ( .B(n281), .A(hinib), .Y(n198) );
  INVXL U324 ( .A(bytcnt[0]), .Y(n281) );
  INVXL U325 ( .A(hinib), .Y(n179) );
  NAND21XL U326 ( .B(n142), .A(bytcnt[0]), .Y(n143) );
  NAND21XL U327 ( .B(n143), .A(bytcnt[2]), .Y(n148) );
  INVXL U328 ( .A(n8), .Y(n155) );
  NAND21XL U329 ( .B(n8), .A(n300), .Y(n81) );
  NAND32XL U330 ( .B(n8), .C(n82), .A(n294), .Y(n276) );
  NAND21XL U331 ( .B(n12), .A(n25), .Y(n259) );
  NAND32XL U332 ( .B(n167), .C(n12), .A(n199), .Y(n170) );
  NAND21XL U333 ( .B(n207), .A(n12), .Y(n159) );
  AND4XL U334 ( .A(n26), .B(n287), .C(n286), .D(n285), .Y(ptx_crcstart) );
  NAND21XL U335 ( .B(n26), .A(n215), .Y(n183) );
  NAND21X1 U336 ( .B(n31), .A(n303), .Y(ptx_fifopop) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyidd_a0 ( i_trans, i_goidle, o_ccidle, o_goidle, o_gobusy, clk, srstz, 
        test_si, test_so, test_se );
  input i_trans, i_goidle, clk, srstz, test_si, test_se;
  output o_ccidle, o_goidle, o_gobusy, test_so;
  wire   ttranwin_6_, ttranwin_5_, ttranwin_4_, ttranwin_3_, ttranwin_2_,
         ttranwin_1_, ttranwin_0_, N11, N12, N13, N14, N15, N16, N17, N18, N46,
         N47, N48, N49, N50, N51, N52, N53, N55, N56, N57, N58, N59, N60, N61,
         N62, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, net10668, net10674, net10679, n55, n56,
         n57, n17, n18, n19, n20, n21, n22, n23, n24, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n25, n26, n27, n28;
  wire   [1:0] ntrancnt;
  wire   [7:0] trans0;
  wire   [7:0] ttranwin_minus;
  wire   [7:0] trans1;

  SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 clk_gate_trans1_reg ( .CLK(clk), .EN(N90), 
        .ENCLK(net10668), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 clk_gate_trans0_reg ( .CLK(clk), .EN(N91), 
        .ENCLK(net10674), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 clk_gate_ttranwin_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net10679), .TE(test_se) );
  phyidd_a0_DW01_sub_0 sub_47 ( .A(trans1), .B(trans0), .CI(1'b0), .DIFF({N53, 
        N52, N51, N50, N49, N48, N47, N46}), .CO() );
  phyidd_a0_DW01_sub_1 sub_24 ( .A({n24, n23, n22, n21, n20, n19, n18, n17}), 
        .B(trans0), .CI(1'b0), .DIFF(ttranwin_minus), .CO() );
  phyidd_a0_DW01_inc_0 add_23 ( .A({test_so, ttranwin_6_, ttranwin_5_, 
        ttranwin_4_, ttranwin_3_, ttranwin_2_, ttranwin_1_, ttranwin_0_}), 
        .SUM({N18, N17, N16, N15, N14, N13, N12, N11}) );
  SDFFQX1 trans1_reg_7_ ( .D(N80), .SIN(trans1[6]), .SMC(test_se), .C(net10668), .Q(trans1[7]) );
  SDFFQX1 trans0_reg_7_ ( .D(N62), .SIN(trans0[6]), .SMC(test_se), .C(net10674), .Q(trans0[7]) );
  SDFFQX1 trans1_reg_6_ ( .D(N79), .SIN(trans1[5]), .SMC(test_se), .C(net10668), .Q(trans1[6]) );
  SDFFQX1 trans1_reg_5_ ( .D(N78), .SIN(trans1[4]), .SMC(test_se), .C(net10668), .Q(trans1[5]) );
  SDFFQX1 trans0_reg_6_ ( .D(N61), .SIN(trans0[5]), .SMC(test_se), .C(net10674), .Q(trans0[6]) );
  SDFFQX1 trans1_reg_4_ ( .D(N77), .SIN(trans1[3]), .SMC(test_se), .C(net10668), .Q(trans1[4]) );
  SDFFQX1 ntrancnt_reg_1_ ( .D(n56), .SIN(ntrancnt[0]), .SMC(test_se), .C(clk), 
        .Q(ntrancnt[1]) );
  SDFFQX1 ntrancnt_reg_0_ ( .D(n57), .SIN(o_ccidle), .SMC(test_se), .C(clk), 
        .Q(ntrancnt[0]) );
  SDFFQX1 trans0_reg_5_ ( .D(N60), .SIN(trans0[4]), .SMC(test_se), .C(net10674), .Q(trans0[5]) );
  SDFFQX1 trans0_reg_4_ ( .D(N59), .SIN(trans0[3]), .SMC(test_se), .C(net10674), .Q(trans0[4]) );
  SDFFQX1 trans1_reg_3_ ( .D(N76), .SIN(trans1[2]), .SMC(test_se), .C(net10668), .Q(trans1[3]) );
  SDFFQX1 trans1_reg_2_ ( .D(N75), .SIN(trans1[1]), .SMC(test_se), .C(net10668), .Q(trans1[2]) );
  SDFFQX1 trans0_reg_3_ ( .D(N58), .SIN(trans0[2]), .SMC(test_se), .C(net10674), .Q(trans0[3]) );
  SDFFQX1 trans1_reg_1_ ( .D(N74), .SIN(trans1[0]), .SMC(test_se), .C(net10668), .Q(trans1[1]) );
  SDFFQX1 trans1_reg_0_ ( .D(N73), .SIN(trans0[7]), .SMC(test_se), .C(net10668), .Q(trans1[0]) );
  SDFFQX1 trans0_reg_2_ ( .D(N57), .SIN(trans0[1]), .SMC(test_se), .C(net10674), .Q(trans0[2]) );
  SDFFQX1 trans0_reg_1_ ( .D(N56), .SIN(trans0[0]), .SMC(test_se), .C(net10674), .Q(trans0[1]) );
  SDFFQX1 ttranwin_reg_7_ ( .D(N89), .SIN(ttranwin_6_), .SMC(test_se), .C(
        net10679), .Q(test_so) );
  SDFFQX1 ttranwin_reg_6_ ( .D(N88), .SIN(ttranwin_5_), .SMC(test_se), .C(
        net10679), .Q(ttranwin_6_) );
  SDFFQX1 trans0_reg_0_ ( .D(N55), .SIN(ntrancnt[1]), .SMC(test_se), .C(
        net10674), .Q(trans0[0]) );
  SDFFQX1 ttranwin_reg_5_ ( .D(N87), .SIN(ttranwin_4_), .SMC(test_se), .C(
        net10679), .Q(ttranwin_5_) );
  SDFFQX1 ttranwin_reg_4_ ( .D(N86), .SIN(ttranwin_3_), .SMC(test_se), .C(
        net10679), .Q(ttranwin_4_) );
  SDFFQX1 ttranwin_reg_1_ ( .D(N83), .SIN(ttranwin_0_), .SMC(test_se), .C(
        net10679), .Q(ttranwin_1_) );
  SDFFQX1 ttranwin_reg_2_ ( .D(N84), .SIN(ttranwin_1_), .SMC(test_se), .C(
        net10679), .Q(ttranwin_2_) );
  SDFFQX1 ttranwin_reg_3_ ( .D(N85), .SIN(ttranwin_2_), .SMC(test_se), .C(
        net10679), .Q(ttranwin_3_) );
  SDFFQX1 ttranwin_reg_0_ ( .D(N82), .SIN(trans1[7]), .SMC(test_se), .C(
        net10679), .Q(ttranwin_0_) );
  SDFFQX1 ccidle_reg ( .D(n55), .SIN(test_si), .SMC(test_se), .C(clk), .Q(
        o_ccidle) );
  BUFX3 U5 ( .A(n48), .Y(n1) );
  NAND2X1 U6 ( .A(ntrancnt[1]), .B(n16), .Y(n2) );
  INVX1 U7 ( .A(n12), .Y(n5) );
  OAI22X1 U8 ( .A(n48), .B(n10), .C(n49), .D(n31), .Y(N87) );
  OAI22X1 U9 ( .A(n48), .B(n9), .C(n30), .D(n49), .Y(N88) );
  INVX1 U10 ( .A(n43), .Y(o_goidle) );
  OAI22X1 U11 ( .A(n48), .B(n11), .C(n49), .D(n32), .Y(N86) );
  OAI22X1 U12 ( .A(n48), .B(n14), .C(n49), .D(n33), .Y(N85) );
  OAI22X1 U13 ( .A(n48), .B(n15), .C(n49), .D(n34), .Y(N84) );
  OAI22X1 U14 ( .A(n48), .B(n25), .C(n49), .D(n35), .Y(N83) );
  NOR2X1 U15 ( .A(n38), .B(n7), .Y(n37) );
  INVX1 U16 ( .A(n40), .Y(n12) );
  NAND2X1 U17 ( .A(N12), .B(n44), .Y(n35) );
  OAI22X1 U18 ( .A(n12), .B(n8), .C(n29), .D(n45), .Y(N80) );
  OAI22X1 U19 ( .A(n48), .B(n8), .C(n29), .D(n49), .Y(N89) );
  INVX1 U20 ( .A(n36), .Y(n17) );
  INVX1 U21 ( .A(ttranwin_minus[5]), .Y(n10) );
  INVX1 U22 ( .A(ttranwin_minus[6]), .Y(n9) );
  NAND2X1 U23 ( .A(N13), .B(n44), .Y(n34) );
  NAND2X1 U24 ( .A(N14), .B(n44), .Y(n33) );
  OAI22X1 U25 ( .A(n12), .B(n10), .C(n45), .D(n31), .Y(N78) );
  OAI22X1 U26 ( .A(n12), .B(n9), .C(n30), .D(n2), .Y(N79) );
  AOI21X1 U27 ( .B(n27), .C(n28), .A(i_goidle), .Y(n43) );
  NOR3XL U28 ( .A(n7), .B(n45), .C(n28), .Y(o_gobusy) );
  INVX1 U29 ( .A(ttranwin_minus[4]), .Y(n11) );
  NOR2X1 U30 ( .A(N17), .B(n27), .Y(n30) );
  NAND2X1 U31 ( .A(N16), .B(n44), .Y(n31) );
  NAND2X1 U32 ( .A(N15), .B(n44), .Y(n32) );
  INVX1 U33 ( .A(i_trans), .Y(n7) );
  OAI22X1 U34 ( .A(n12), .B(n11), .C(n2), .D(n32), .Y(N77) );
  ENOX1 U35 ( .A(n30), .B(n46), .C(N52), .D(n40), .Y(N61) );
  NAND31X1 U36 ( .C(n47), .A(i_trans), .B(n5), .Y(n48) );
  OA33X1 U37 ( .A(n47), .B(i_trans), .C(n27), .D(n47), .E(n41), .F(n7), .Y(n49) );
  INVX1 U38 ( .A(ttranwin_minus[2]), .Y(n15) );
  INVX1 U39 ( .A(ttranwin_minus[3]), .Y(n14) );
  NAND31X1 U40 ( .C(o_gobusy), .A(n6), .B(n43), .Y(n38) );
  OA21X1 U41 ( .B(n44), .C(i_trans), .A(srstz), .Y(n6) );
  OAI22AX1 U42 ( .D(n37), .C(n41), .A(n38), .B(n13), .Y(n56) );
  OAI22X1 U43 ( .A(n48), .B(n26), .C(n49), .D(n36), .Y(N82) );
  OAI22X1 U44 ( .A(n12), .B(n15), .C(n45), .D(n34), .Y(N75) );
  OAI22X1 U45 ( .A(n12), .B(n14), .C(n2), .D(n33), .Y(N76) );
  OAI31XL U46 ( .A(n16), .B(n37), .C(n38), .D(n39), .Y(n57) );
  OAI21X1 U47 ( .B(n40), .C(n16), .A(n37), .Y(n39) );
  ENOX1 U48 ( .A(n46), .B(n31), .C(N51), .D(n40), .Y(N60) );
  INVX1 U49 ( .A(n44), .Y(n27) );
  OAI211X1 U50 ( .C(n41), .D(n7), .A(n1), .B(n50), .Y(N81) );
  AOI21X1 U51 ( .B(n44), .C(n7), .A(n47), .Y(n50) );
  INVX1 U52 ( .A(ttranwin_minus[1]), .Y(n25) );
  OAI22X1 U53 ( .A(n12), .B(n26), .C(n45), .D(n36), .Y(N73) );
  OAI22X1 U54 ( .A(n12), .B(n25), .C(n2), .D(n35), .Y(N74) );
  OAI31XL U55 ( .A(n46), .B(n7), .C(n47), .D(n48), .Y(N91) );
  OAI31XL U56 ( .A(n47), .B(n45), .C(n7), .D(n1), .Y(N90) );
  ENOX1 U57 ( .A(n46), .B(n33), .C(N49), .D(n40), .Y(N58) );
  ENOX1 U58 ( .A(n46), .B(n32), .C(N50), .D(n40), .Y(N59) );
  OAI211X1 U59 ( .C(o_gobusy), .D(n28), .A(n43), .B(srstz), .Y(n55) );
  ENOX1 U60 ( .A(n46), .B(n35), .C(N47), .D(n40), .Y(N56) );
  ENOX1 U61 ( .A(n46), .B(n34), .C(N48), .D(n40), .Y(N57) );
  NOR2X1 U62 ( .A(n16), .B(n13), .Y(n40) );
  AND2X1 U63 ( .A(n46), .B(n2), .Y(n41) );
  INVX1 U64 ( .A(n34), .Y(n19) );
  INVX1 U65 ( .A(n33), .Y(n20) );
  INVX1 U66 ( .A(n32), .Y(n21) );
  INVX1 U67 ( .A(n31), .Y(n22) );
  INVX1 U68 ( .A(n35), .Y(n18) );
  INVX1 U69 ( .A(n30), .Y(n23) );
  NAND2X1 U70 ( .A(N11), .B(n44), .Y(n36) );
  INVX1 U71 ( .A(ttranwin_minus[7]), .Y(n8) );
  INVX1 U72 ( .A(n29), .Y(n24) );
  NAND4X1 U73 ( .A(test_so), .B(ttranwin_6_), .C(n51), .D(n52), .Y(n44) );
  NOR2X1 U74 ( .A(ttranwin_1_), .B(ttranwin_0_), .Y(n51) );
  NOR4XL U75 ( .A(ttranwin_5_), .B(ttranwin_4_), .C(ttranwin_3_), .D(
        ttranwin_2_), .Y(n52) );
  ENOX1 U76 ( .A(n29), .B(n46), .C(N53), .D(n40), .Y(N62) );
  OAI31XL U77 ( .A(n28), .B(ntrancnt[0]), .C(n7), .D(srstz), .Y(n47) );
  INVX1 U78 ( .A(o_ccidle), .Y(n28) );
  NOR2X1 U79 ( .A(N18), .B(n27), .Y(n29) );
  NAND2X1 U80 ( .A(ntrancnt[1]), .B(n16), .Y(n45) );
  INVX1 U81 ( .A(ttranwin_minus[0]), .Y(n26) );
  INVX1 U82 ( .A(ntrancnt[0]), .Y(n16) );
  ENOX1 U83 ( .A(n46), .B(n36), .C(N46), .D(n40), .Y(N55) );
  NAND2X1 U84 ( .A(ntrancnt[0]), .B(n13), .Y(n46) );
  INVX1 U85 ( .A(ntrancnt[1]), .Y(n13) );
endmodule


module phyidd_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module phyidd_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n17), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n10), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(A[0]), .Y(n18) );
  INVX1 U2 ( .A(B[2]), .Y(n14) );
  INVX1 U3 ( .A(B[3]), .Y(n15) );
  INVX1 U4 ( .A(B[4]), .Y(n13) );
  INVX1 U5 ( .A(B[5]), .Y(n11) );
  INVX1 U6 ( .A(B[1]), .Y(n17) );
  NAND21X1 U7 ( .B(n16), .A(n18), .Y(carry[1]) );
  INVX1 U8 ( .A(B[6]), .Y(n12) );
  INVX1 U9 ( .A(B[7]), .Y(n10) );
  INVX1 U10 ( .A(B[0]), .Y(n16) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module phyidd_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n18), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n10), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(B[2]), .Y(n14) );
  INVX1 U2 ( .A(B[3]), .Y(n15) );
  INVX1 U3 ( .A(B[4]), .Y(n13) );
  INVX1 U4 ( .A(B[5]), .Y(n11) );
  INVX1 U5 ( .A(B[1]), .Y(n18) );
  NAND21X1 U6 ( .B(n17), .A(n16), .Y(carry[1]) );
  INVX1 U7 ( .A(A[0]), .Y(n16) );
  INVX1 U8 ( .A(B[6]), .Y(n12) );
  INVX1 U9 ( .A(B[7]), .Y(n10) );
  INVX1 U10 ( .A(B[0]), .Y(n17) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_a0 ( i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, 
        r_rxdb_opt, r_ords_ena, r_pshords, r_rgdcrc, prx_cccnt, prx_rst, 
        prx_setsta, prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, 
        prx_fifopsh, prx_fifowdat, pff_txreq, pid_gobusy, pid_goidle, 
        pid_ccidle, pcc_rxgood, prx_crcstart, prx_crcshfi4, prx_crcsidat, 
        prx_rxcode, prx_adpn, prx_rcvdords, prx_eoprcvd, prx_fsm, clk, srstz, 
        test_si, test_so, test_se );
  input [1:0] r_rxdb_opt;
  input [6:0] r_ords_ena;
  output [1:0] prx_cccnt;
  output [1:0] prx_rst;
  output [6:0] prx_setsta;
  output [7:0] prx_fifowdat;
  output [3:0] prx_crcsidat;
  output [4:0] prx_rxcode;
  output [5:0] prx_adpn;
  output [2:0] prx_rcvdords;
  output [3:0] prx_fsm;
  input i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_pshords,
         r_rgdcrc, pff_txreq, pid_gobusy, pid_goidle, pid_ccidle, pcc_rxgood,
         clk, srstz, test_si, test_se;
  output prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, prx_fifopsh,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd, test_so;
  wire   N31, N32, db_gohi, db_golo, k0_det, cctrans, shrtrans, N70, N71, N72,
         N73, N74, N75, N76, N96, N153, N154, N155, N156, N157, N236, N239,
         N246, N247, N248, N249, N250, N275, N276, N277, N278, N279, net10696,
         net10702, net10707, net10712, net10717, net10722, net10727, n214,
         n314, n313, n282, n283, n284, n289, n75, n119, n120, n122, n131, n139,
         n142, n143, n147, n148, n152, n153, n154, n155, n156, n157, n162,
         n163, n175, n176, n178, n179, n181, n182, n183, n185, n186, n220,
         n221, n1, n2, n5, n7, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n121, n123, n124, n125, n126, n127, n128, n129, n130, n132, n133,
         n134, n135, n136, n137, n138, n140, n141, n144, n145, n146, n149,
         n150, n151, n158, n159, n160, n161, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n177, n180, n184, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n215, n216, n217, n218, n219, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n285, n286, n287, n288, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312;
  wire   [5:0] cccnt;
  wire   [2:0] ps_dat5b;
  wire   [2:0] bcnt;
  wire   [7:3] ordsbuf;

  phyrx_db u0_phyrx_db ( .clk(clk), .srstz(n35), .x_cc(i_cc), .ptx_txact(
        ptx_txact), .r_rxdb_opt(r_rxdb_opt), .gohi(db_gohi), .golo(db_golo), 
        .gotrans(prx_trans), .test_si(n289), .test_so(test_so), .test_se(
        test_se) );
  phyrx_adp u0_phyrx_adp ( .clk(clk), .srstz(n36), .gohi(db_gohi), .golo(
        db_golo), .gobusy(pid_gobusy), .goidle(pid_goidle), .i_ccidle(
        pid_ccidle), .k0_det(k0_det), .r_adprx_en(r_adprx_en), .r_adp2nd(
        r_adp2nd), .adp_val(prx_adpn), .d_cc(prx_d_cc), .cctrans(cctrans), 
        .test_si(shrtrans), .test_so(n289), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 clk_gate_cccnt_reg ( .CLK(clk), .EN(N70), 
        .ENCLK(net10696), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 clk_gate_cs_dat5b_reg ( .CLK(clk), .EN(N153), 
        .ENCLK(net10702), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 clk_gate_bcnt_reg ( .CLK(clk), .EN(N236), 
        .ENCLK(net10707), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 clk_gate_cs_dat4b_reg ( .CLK(clk), .EN(n220), 
        .ENCLK(net10712), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 clk_gate_ordsbuf_reg ( .CLK(clk), .EN(n221), 
        .ENCLK(net10717), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 clk_gate_ordsbuf_reg_0 ( .CLK(clk), .EN(N250), .ENCLK(net10722), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 clk_gate_cs_bmni_reg ( .CLK(clk), .EN(N275), 
        .ENCLK(net10727), .TE(test_se) );
  SDFFQX1 ordsbuf_reg_4_ ( .D(prx_crcsidat[0]), .SIN(ordsbuf[3]), .SMC(test_se), .C(net10717), .Q(ordsbuf[4]) );
  SDFFQX1 ordsbuf_reg_5_ ( .D(prx_fifowdat[5]), .SIN(ordsbuf[4]), .SMC(test_se), .C(net10717), .Q(ordsbuf[5]) );
  SDFFQX1 ordsbuf_reg_3_ ( .D(N249), .SIN(prx_rcvdords[2]), .SMC(test_se), .C(
        net10722), .Q(ordsbuf[3]) );
  SDFFQX1 ordsbuf_reg_7_ ( .D(prx_fifowdat[7]), .SIN(ordsbuf[6]), .SMC(test_se), .C(net10717), .Q(ordsbuf[7]) );
  SDFFQX1 ordsbuf_reg_6_ ( .D(prx_crcsidat[2]), .SIN(ordsbuf[5]), .SMC(test_se), .C(net10717), .Q(ordsbuf[6]) );
  SDFFQX1 cs_dat4b_reg_2_ ( .D(prx_fifowdat[6]), .SIN(prx_fifowdat[1]), .SMC(
        test_se), .C(net10712), .Q(n313) );
  SDFFQX1 cs_dat4b_reg_1_ ( .D(prx_fifowdat[5]), .SIN(prx_fifowdat[0]), .SMC(
        test_se), .C(net10712), .Q(prx_fifowdat[1]) );
  SDFFQX1 cs_dat4b_reg_0_ ( .D(prx_crcsidat[0]), .SIN(prx_fsm[3]), .SMC(
        test_se), .C(net10712), .Q(prx_fifowdat[0]) );
  SDFFQX1 cs_dat4b_reg_3_ ( .D(prx_crcsidat[3]), .SIN(prx_fifowdat[2]), .SMC(
        test_se), .C(net10712), .Q(prx_rxcode[3]) );
  SDFFQX1 cs_dat4b_reg_4_ ( .D(N96), .SIN(prx_rxcode[3]), .SMC(test_se), .C(
        net10712), .Q(prx_rxcode[4]) );
  SDFFQX1 cs_dat5b_reg_0_ ( .D(N154), .SIN(prx_rxcode[4]), .SMC(test_se), .C(
        net10702), .Q(ps_dat5b[0]) );
  SDFFQX1 cs_dat5b_reg_2_ ( .D(N156), .SIN(ps_dat5b[1]), .SMC(test_se), .C(
        net10702), .Q(ps_dat5b[2]) );
  SDFFQX1 cs_dat5b_reg_1_ ( .D(N155), .SIN(ps_dat5b[0]), .SMC(test_se), .C(
        net10702), .Q(ps_dat5b[1]) );
  SDFFQX1 cs_dat5b_reg_3_ ( .D(N157), .SIN(ps_dat5b[2]), .SMC(test_se), .C(
        net10702), .Q(prx_bmc) );
  SDFFQX1 bcnt_reg_2_ ( .D(N239), .SIN(bcnt[1]), .SMC(test_se), .C(net10707), 
        .Q(bcnt[2]) );
  SDFFQX1 cs_bmni_reg_0_ ( .D(N276), .SIN(cccnt[5]), .SMC(test_se), .C(
        net10727), .Q(prx_fsm[0]) );
  SDFFQX1 cccnt_reg_3_ ( .D(N74), .SIN(cccnt[2]), .SMC(test_se), .C(net10696), 
        .Q(cccnt[3]) );
  SDFFQX1 cccnt_reg_2_ ( .D(N73), .SIN(cccnt[1]), .SMC(test_se), .C(net10696), 
        .Q(cccnt[2]) );
  SDFFQX1 ordsbuf_reg_1_ ( .D(N247), .SIN(prx_rcvdords[0]), .SMC(test_se), .C(
        net10722), .Q(prx_rcvdords[1]) );
  MUX2X1 U297 ( .D0(r_ords_ena[1]), .D1(r_ords_ena[2]), .S(N31), .Y(n283) );
  NOR21XL U292 ( .B(r_ords_ena[0]), .A(n299), .Y(n284) );
  MUX4X1 U291 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[4]), .D2(r_ords_ena[5]), 
        .D3(r_ords_ena[6]), .S0(N31), .S1(N32), .Y(n282) );
  SDFFQX1 ordsbuf_reg_2_ ( .D(N248), .SIN(prx_rcvdords[1]), .SMC(test_se), .C(
        net10722), .Q(prx_rcvdords[2]) );
  SDFFQX1 cs_bmni_reg_3_ ( .D(N279), .SIN(prx_fsm[2]), .SMC(test_se), .C(
        net10727), .Q(n314) );
  SDFFQX1 cccnt_reg_1_ ( .D(N72), .SIN(cccnt[0]), .SMC(test_se), .C(net10696), 
        .Q(cccnt[1]) );
  SDFFQX1 cs_bmni_reg_2_ ( .D(N278), .SIN(prx_fsm[1]), .SMC(test_se), .C(
        net10727), .Q(prx_fsm[2]) );
  SDFFQX1 bcnt_reg_1_ ( .D(n307), .SIN(bcnt[0]), .SMC(test_se), .C(net10707), 
        .Q(bcnt[1]) );
  SDFFQX1 shrtrans_reg ( .D(n214), .SIN(ordsbuf[7]), .SMC(test_se), .C(clk), 
        .Q(shrtrans) );
  SDFFQX1 cccnt_reg_4_ ( .D(N75), .SIN(cccnt[3]), .SMC(test_se), .C(net10696), 
        .Q(cccnt[4]) );
  SDFFQX1 bcnt_reg_0_ ( .D(n295), .SIN(test_si), .SMC(test_se), .C(net10707), 
        .Q(bcnt[0]) );
  SDFFQX1 cccnt_reg_0_ ( .D(N71), .SIN(bcnt[2]), .SMC(test_se), .C(net10696), 
        .Q(cccnt[0]) );
  SDFFQX1 cccnt_reg_5_ ( .D(N76), .SIN(cccnt[4]), .SMC(test_se), .C(net10696), 
        .Q(cccnt[5]) );
  SDFFQX1 cs_bmni_reg_1_ ( .D(N277), .SIN(prx_fsm[0]), .SMC(test_se), .C(
        net10727), .Q(prx_fsm[1]) );
  SDFFQX1 ordsbuf_reg_0_ ( .D(N246), .SIN(prx_bmc), .SMC(test_se), .C(net10722), .Q(prx_rcvdords[0]) );
  INVX2 U3 ( .A(cctrans), .Y(n51) );
  INVX1 U4 ( .A(n252), .Y(n22) );
  NOR2X1 U5 ( .A(cccnt[4]), .B(cccnt[3]), .Y(n23) );
  MUX2X1 U6 ( .D0(n227), .D1(n226), .S(prx_rcvdords[1]), .Y(n228) );
  INVX1 U7 ( .A(n207), .Y(n246) );
  INVX1 U8 ( .A(n104), .Y(n105) );
  INVX1 U9 ( .A(prx_fsm[0]), .Y(n109) );
  NAND21X1 U10 ( .B(n190), .A(cccnt[0]), .Y(n271) );
  INVX1 U11 ( .A(cccnt[2]), .Y(n48) );
  INVX1 U12 ( .A(cccnt[5]), .Y(n40) );
  INVX1 U13 ( .A(prx_fsm[1]), .Y(n249) );
  NAND21X1 U14 ( .B(bcnt[1]), .A(n41), .Y(n244) );
  INVX1 U15 ( .A(bcnt[0]), .Y(n41) );
  INVX1 U16 ( .A(cccnt[1]), .Y(n190) );
  NAND21X1 U17 ( .B(n314), .A(n105), .Y(n207) );
  INVX1 U18 ( .A(n271), .Y(n193) );
  NAND21X1 U19 ( .B(n48), .A(n193), .Y(n196) );
  INVX1 U20 ( .A(shrtrans), .Y(n242) );
  AOI222XL U21 ( .A(prx_bmc), .B(n70), .C(ps_dat5b[0]), .D(n69), .E(n68), .F(
        ps_dat5b[1]), .Y(n1) );
  OR2X1 U22 ( .A(n155), .B(n122), .Y(n2) );
  INVX1 U23 ( .A(cccnt[3]), .Y(n195) );
  INVXL U24 ( .A(n1), .Y(prx_crcsidat[2]) );
  INVXL U25 ( .A(n1), .Y(prx_fifowdat[6]) );
  INVXL U26 ( .A(n313), .Y(n5) );
  INVXL U27 ( .A(n5), .Y(prx_fifowdat[2]) );
  INVXL U28 ( .A(n314), .Y(n7) );
  INVXL U29 ( .A(n7), .Y(prx_fsm[3]) );
  INVXL U30 ( .A(prx_fifowdat[4]), .Y(n9) );
  INVXL U31 ( .A(n9), .Y(prx_crcsidat[0]) );
  INVX1 U32 ( .A(n15), .Y(n11) );
  AND3X1 U33 ( .A(bcnt[2]), .B(n254), .C(n13), .Y(n12) );
  AND2X2 U34 ( .A(n255), .B(n12), .Y(prx_fifopsh) );
  INVX1 U35 ( .A(n244), .Y(n254) );
  NAND2X1 U36 ( .A(n253), .B(n22), .Y(n13) );
  OR2XL U37 ( .A(n15), .B(n17), .Y(n14) );
  INVX1 U38 ( .A(n50), .Y(n17) );
  BUFXL U39 ( .A(n51), .Y(n15) );
  NOR2X2 U40 ( .A(n51), .B(n17), .Y(n16) );
  INVX1 U41 ( .A(n72), .Y(n18) );
  AND2X1 U42 ( .A(prx_bmc), .B(ps_dat5b[2]), .Y(n78) );
  INVXL U43 ( .A(ptx_txact), .Y(n310) );
  BUFX3 U44 ( .A(n313), .Y(prx_rxcode[2]) );
  BUFX3 U45 ( .A(prx_fifowdat[1]), .Y(prx_rxcode[1]) );
  BUFX3 U46 ( .A(prx_fifowdat[0]), .Y(prx_rxcode[0]) );
  INVX1 U47 ( .A(n106), .Y(n108) );
  NAND43XL U48 ( .B(n240), .C(n110), .D(n169), .A(n245), .Y(n111) );
  INVXL U49 ( .A(n245), .Y(n215) );
  OAI211XL U50 ( .C(n48), .D(n191), .A(n42), .B(n23), .Y(n241) );
  INVXL U51 ( .A(n45), .Y(n42) );
  OAI32XL U52 ( .A(n244), .B(n74), .C(n187), .D(n74), .E(n205), .Y(n220) );
  AND2XL U53 ( .A(n191), .B(n190), .Y(n192) );
  AO21XL U54 ( .B(n200), .C(n191), .A(n37), .Y(N71) );
  NAND21XL U55 ( .B(n249), .A(n166), .Y(n161) );
  NAND32XL U56 ( .B(n7), .C(n249), .A(n251), .Y(n206) );
  NAND21XL U57 ( .B(cccnt[5]), .A(n49), .Y(n50) );
  NAND31XL U58 ( .C(n48), .A(cccnt[3]), .B(cccnt[4]), .Y(n49) );
  INVXL U59 ( .A(prx_fsm[2]), .Y(n251) );
  INVX1 U60 ( .A(n116), .Y(n285) );
  INVX1 U61 ( .A(n37), .Y(n36) );
  INVX1 U62 ( .A(n37), .Y(n35) );
  INVX1 U63 ( .A(n157), .Y(n302) );
  INVX1 U64 ( .A(n238), .Y(n239) );
  NAND21X1 U65 ( .B(n157), .A(n293), .Y(n116) );
  INVX1 U66 ( .A(N32), .Y(n308) );
  INVX1 U67 ( .A(n236), .Y(n266) );
  INVX1 U68 ( .A(n160), .Y(n170) );
  NAND2X1 U69 ( .A(n233), .B(n35), .Y(n165) );
  NAND21X1 U70 ( .B(n218), .A(n217), .Y(N236) );
  NAND21X1 U71 ( .B(n219), .A(n20), .Y(N153) );
  INVX1 U72 ( .A(n76), .Y(n219) );
  NAND21X1 U73 ( .B(n74), .A(n20), .Y(n76) );
  AND2X1 U74 ( .A(n219), .B(n77), .Y(N157) );
  OR2X1 U75 ( .A(pid_goidle), .B(n165), .Y(n209) );
  NAND21X1 U76 ( .B(n221), .A(n236), .Y(N250) );
  INVX1 U77 ( .A(n216), .Y(n221) );
  NAND21X1 U78 ( .B(n237), .A(n215), .Y(n216) );
  INVX1 U79 ( .A(srstz), .Y(n37) );
  INVX1 U80 ( .A(n270), .Y(prx_cccnt[0]) );
  NAND21X1 U81 ( .B(n248), .A(n247), .Y(n253) );
  NAND21X1 U82 ( .B(n246), .A(n245), .Y(n247) );
  INVX1 U83 ( .A(r_pshords), .Y(n248) );
  INVX1 U84 ( .A(n259), .Y(n77) );
  INVX1 U85 ( .A(n241), .Y(n43) );
  INVX1 U86 ( .A(n222), .Y(n200) );
  OR2X1 U87 ( .A(n9), .B(n224), .Y(n157) );
  NAND32X1 U88 ( .B(n96), .C(n97), .A(n152), .Y(n149) );
  INVX1 U89 ( .A(n139), .Y(n96) );
  AOI21X1 U90 ( .B(n153), .C(n154), .A(n2), .Y(n152) );
  AOI31X1 U91 ( .A(n292), .B(n297), .C(n302), .D(n291), .Y(n153) );
  NAND2X1 U92 ( .A(n235), .B(n266), .Y(n238) );
  NAND21X1 U93 ( .B(n237), .A(n21), .Y(n233) );
  OR2X1 U94 ( .A(n117), .B(n19), .Y(n278) );
  AOI21X1 U95 ( .B(n294), .C(n302), .A(n293), .Y(n19) );
  NAND32X1 U96 ( .B(n223), .C(n37), .A(n222), .Y(N70) );
  INVX1 U97 ( .A(n220), .Y(n237) );
  NAND21X1 U98 ( .B(n117), .A(n285), .Y(n279) );
  INVX1 U99 ( .A(n88), .Y(n304) );
  AO21X1 U100 ( .B(n120), .C(n280), .A(n122), .Y(n146) );
  AO21X1 U101 ( .B(n263), .C(n220), .A(prx_setsta[6]), .Y(prx_fiforst) );
  INVX1 U102 ( .A(n179), .Y(n309) );
  NAND21X1 U103 ( .B(n224), .A(n303), .Y(n179) );
  AO21X1 U104 ( .B(n124), .C(n2), .A(n102), .Y(N32) );
  NAND21X1 U105 ( .B(n99), .A(n98), .Y(n102) );
  INVX1 U106 ( .A(n97), .Y(n98) );
  INVX1 U107 ( .A(n149), .Y(n99) );
  NOR2X1 U108 ( .A(n299), .B(n75), .Y(prx_rst[0]) );
  NOR2X1 U109 ( .A(N31), .B(n75), .Y(prx_rst[1]) );
  INVX1 U110 ( .A(N31), .Y(n299) );
  NAND21X1 U111 ( .B(n308), .A(n103), .Y(n75) );
  NAND21X1 U112 ( .B(n237), .A(n246), .Y(n236) );
  INVX1 U113 ( .A(n261), .Y(n74) );
  INVX1 U114 ( .A(n103), .Y(n125) );
  AOI21X1 U115 ( .B(n164), .C(n161), .A(n212), .Y(N278) );
  AO21X1 U116 ( .B(n264), .C(n235), .A(n160), .Y(n164) );
  NAND2X1 U117 ( .A(n75), .B(n246), .Y(n160) );
  INVX1 U118 ( .A(n117), .Y(n303) );
  INVX1 U119 ( .A(n273), .Y(n293) );
  INVX1 U120 ( .A(n172), .Y(n217) );
  NAND21X1 U121 ( .B(n220), .A(n35), .Y(n172) );
  INVX1 U122 ( .A(n188), .Y(n218) );
  INVX1 U123 ( .A(n95), .Y(n86) );
  INVX1 U124 ( .A(n280), .Y(n281) );
  NAND43X1 U125 ( .B(pid_goidle), .C(n21), .D(n237), .A(n36), .Y(n212) );
  NOR2X1 U126 ( .A(n165), .B(pid_gobusy), .Y(n20) );
  INVX1 U127 ( .A(n90), .Y(n275) );
  INVX1 U128 ( .A(n311), .Y(n183) );
  INVX1 U129 ( .A(n290), .Y(n291) );
  INVX1 U130 ( .A(n288), .Y(n292) );
  INVX1 U131 ( .A(n143), .Y(n305) );
  AO21X1 U132 ( .B(n294), .C(n305), .A(n293), .Y(n148) );
  INVX1 U133 ( .A(n129), .Y(n240) );
  INVX1 U134 ( .A(n111), .Y(n208) );
  INVX1 U135 ( .A(n161), .Y(n110) );
  INVX1 U136 ( .A(n197), .Y(n199) );
  AND2X1 U137 ( .A(n215), .B(prx_fifowdat[3]), .Y(N249) );
  NAND32X1 U138 ( .B(n196), .C(n40), .A(n23), .Y(n270) );
  NAND32X1 U139 ( .B(n109), .C(n249), .A(n108), .Y(n245) );
  NAND32X1 U140 ( .B(n249), .C(n251), .A(n109), .Y(n104) );
  NAND32XL U141 ( .B(n15), .C(n242), .A(n202), .Y(n259) );
  INVX1 U142 ( .A(n55), .Y(n66) );
  NAND21X1 U143 ( .B(n65), .A(n77), .Y(n55) );
  NAND21X1 U144 ( .B(n59), .A(n66), .Y(n58) );
  NAND32X1 U145 ( .B(n65), .C(n63), .A(n259), .Y(n71) );
  INVX1 U146 ( .A(n114), .Y(prx_fifowdat[3]) );
  NAND21X1 U147 ( .B(pff_txreq), .A(n38), .Y(n223) );
  OAI31XL U148 ( .A(n197), .B(n272), .C(n40), .D(n39), .Y(n222) );
  INVX1 U149 ( .A(n223), .Y(n39) );
  AO21X1 U150 ( .B(n240), .C(n220), .A(n239), .Y(prx_crcstart) );
  NAND21X1 U151 ( .B(prx_crcsidat[2]), .A(n304), .Y(n224) );
  AND3X1 U152 ( .A(prx_eoprcvd), .B(pcc_rxgood), .C(n267), .Y(prx_setsta[3])
         );
  OAI221X1 U153 ( .A(n143), .B(n123), .C(n296), .D(n279), .E(n150), .Y(n122)
         );
  OA21X1 U154 ( .B(n296), .C(n278), .A(n116), .Y(n123) );
  INVX1 U155 ( .A(n234), .Y(prx_eoprcvd) );
  NAND32X1 U156 ( .B(n233), .C(n7), .A(n269), .Y(n234) );
  OAI31XL U157 ( .A(n198), .B(n199), .C(n222), .D(n36), .Y(N74) );
  AND2XL U158 ( .A(n196), .B(n195), .Y(n198) );
  OAI31XL U159 ( .A(n192), .B(n193), .C(n222), .D(n36), .Y(N72) );
  NAND43X1 U160 ( .B(n159), .C(n158), .D(n151), .A(n150), .Y(n235) );
  INVX1 U161 ( .A(n137), .Y(n159) );
  INVX1 U162 ( .A(n138), .Y(n158) );
  OAI211X1 U163 ( .C(n290), .D(n149), .A(n146), .B(n277), .Y(n151) );
  NAND2X1 U164 ( .A(prx_fifowdat[7]), .B(prx_fifowdat[5]), .Y(n88) );
  GEN2XL U165 ( .D(n306), .E(n301), .C(n300), .B(n296), .A(n175), .Y(n155) );
  AO21X1 U166 ( .B(n285), .C(n306), .A(n281), .Y(n175) );
  INVX1 U167 ( .A(n279), .Y(n300) );
  INVX1 U168 ( .A(n278), .Y(n301) );
  NOR2X1 U169 ( .A(n162), .B(n163), .Y(n139) );
  OAI21X1 U170 ( .B(n181), .C(n296), .A(n182), .Y(n163) );
  AOI31X1 U171 ( .A(n304), .B(n1), .C(n183), .D(n119), .Y(n182) );
  AOI32X1 U172 ( .A(n185), .B(n9), .C(n309), .D(n303), .E(n183), .Y(n181) );
  INVX1 U173 ( .A(n277), .Y(n119) );
  INVX1 U174 ( .A(n256), .Y(prx_setsta[6]) );
  NAND32X1 U175 ( .B(n267), .C(n268), .A(prx_eoprcvd), .Y(n256) );
  OAI211X1 U176 ( .C(n297), .D(n302), .A(n156), .B(n305), .Y(n154) );
  OAI31XL U177 ( .A(n287), .B(n157), .C(n286), .D(n288), .Y(n156) );
  NOR41XL U178 ( .D(N96), .A(n1), .B(prx_crcsidat[0]), .C(prx_fifowdat[5]), 
        .Y(n21) );
  OAI211X1 U179 ( .C(n142), .D(n122), .A(n124), .B(n149), .Y(N31) );
  AOI21BX1 U180 ( .C(n162), .B(n163), .A(n155), .Y(n142) );
  OAI211X1 U181 ( .C(n95), .D(n288), .A(n94), .B(n137), .Y(n97) );
  NAND32X1 U182 ( .B(prx_crcsidat[0]), .C(n89), .A(n304), .Y(n94) );
  GEN2XL U183 ( .D(n286), .E(n140), .C(n288), .B(n87), .A(n1), .Y(n89) );
  NAND21X1 U184 ( .B(n287), .A(n86), .Y(n87) );
  OAI31XL U185 ( .A(n21), .B(n237), .C(n7), .D(n238), .Y(prx_crcshfi4) );
  AND2X1 U186 ( .A(n266), .B(n265), .Y(prx_setsta[2]) );
  AND2X1 U187 ( .A(n264), .B(n266), .Y(prx_setsta[1]) );
  INVX1 U188 ( .A(n265), .Y(n264) );
  OAI31XL U189 ( .A(n139), .B(n2), .C(n101), .D(n100), .Y(n103) );
  INVX1 U190 ( .A(n102), .Y(n100) );
  NAND21X1 U191 ( .B(n265), .A(n170), .Y(n126) );
  OAI22X1 U192 ( .A(n209), .B(n211), .C(n171), .D(n212), .Y(N276) );
  AOI211X1 U193 ( .C(n170), .D(n265), .A(n169), .B(n168), .Y(n171) );
  INVX1 U194 ( .A(n206), .Y(n168) );
  INVX1 U195 ( .A(n101), .Y(n124) );
  AOI31X1 U196 ( .A(n206), .B(n129), .C(n128), .D(n212), .Y(N279) );
  OA21X1 U197 ( .B(n263), .C(n127), .A(n126), .Y(n128) );
  AND2X1 U198 ( .A(prx_eoprcvd), .B(n268), .Y(prx_setsta[4]) );
  OAI22XL U199 ( .A(n125), .B(n207), .C(n5), .D(n245), .Y(N248) );
  OAI22XL U200 ( .A(n296), .B(n245), .C(n308), .D(n207), .Y(N247) );
  OAI22XL U201 ( .A(n144), .B(n245), .C(n299), .D(n207), .Y(N246) );
  NAND32X1 U202 ( .B(n114), .C(n144), .A(n5), .Y(n117) );
  NAND21X1 U203 ( .B(r_ordrs4), .A(n80), .Y(n273) );
  INVX1 U204 ( .A(n115), .Y(n80) );
  NAND21X1 U205 ( .B(n286), .A(n93), .Y(n95) );
  OR3XL U206 ( .A(n143), .B(n229), .C(n141), .Y(n280) );
  OAI211X1 U207 ( .C(n177), .D(n174), .A(n261), .B(n173), .Y(n188) );
  INVX1 U208 ( .A(n258), .Y(n177) );
  AND2X1 U209 ( .A(n217), .B(n257), .Y(n173) );
  NAND32X1 U210 ( .B(n176), .C(n141), .A(n229), .Y(n150) );
  NAND21X1 U211 ( .B(n312), .A(n115), .Y(n294) );
  INVX1 U212 ( .A(n205), .Y(k0_det) );
  INVX1 U213 ( .A(n184), .Y(n295) );
  NAND21X1 U214 ( .B(n91), .A(n312), .Y(n288) );
  NAND21X1 U215 ( .B(n273), .A(n274), .Y(n311) );
  NAND32X1 U216 ( .B(n140), .C(n141), .A(n229), .Y(n290) );
  NAND32X1 U217 ( .B(n296), .C(n114), .A(n144), .Y(n90) );
  NAND32X1 U218 ( .B(n176), .C(n145), .A(n144), .Y(n277) );
  AO21X1 U219 ( .B(n274), .C(n294), .A(n293), .Y(n185) );
  NAND32X1 U220 ( .B(n144), .C(n145), .A(n274), .Y(n120) );
  NAND5XL U221 ( .A(n232), .B(prx_fifowdat[3]), .C(n134), .D(n133), .E(n132), 
        .Y(n145) );
  NAND2X1 U222 ( .A(n178), .B(n298), .Y(n143) );
  INVX1 U223 ( .A(n140), .Y(n93) );
  INVX1 U224 ( .A(n127), .Y(n169) );
  INVX1 U225 ( .A(n174), .Y(n263) );
  INVX1 U226 ( .A(n85), .Y(n287) );
  NAND21X1 U227 ( .B(n312), .A(n91), .Y(n85) );
  OAI211X1 U228 ( .C(n213), .D(n212), .A(n211), .B(n210), .Y(N275) );
  AND3XL U229 ( .A(n208), .B(n207), .C(n206), .Y(n213) );
  INVX1 U230 ( .A(n209), .Y(n210) );
  INVX1 U231 ( .A(n286), .Y(n297) );
  INVX1 U232 ( .A(n176), .Y(n306) );
  INVX1 U233 ( .A(pcc_rxgood), .Y(n268) );
  NAND43X1 U234 ( .B(n143), .C(n90), .D(n115), .A(n133), .Y(n138) );
  NAND21XL U235 ( .B(n7), .A(n105), .Y(n129) );
  NAND32X1 U236 ( .B(n167), .C(n257), .A(n310), .Y(n211) );
  INVX1 U237 ( .A(pid_gobusy), .Y(n167) );
  OR2XL U238 ( .A(n195), .B(n196), .Y(n197) );
  AND4X1 U239 ( .A(n263), .B(n262), .C(n261), .D(n260), .Y(prx_setsta[0]) );
  INVX1 U240 ( .A(n257), .Y(prx_idle) );
  NOR32XL U241 ( .B(n251), .C(prx_fsm[3]), .A(n250), .Y(n252) );
  XOR2XL U242 ( .A(n249), .B(prx_fsm[0]), .Y(n250) );
  AO21XL U243 ( .B(cccnt[1]), .C(cccnt[2]), .A(cccnt[5]), .Y(n45) );
  NAND21X1 U244 ( .B(prx_fsm[2]), .A(n7), .Y(n106) );
  INVXL U245 ( .A(cccnt[0]), .Y(n191) );
  NAND32X1 U246 ( .B(ps_dat5b[2]), .C(n259), .A(n53), .Y(n57) );
  GEN2XL U247 ( .D(ps_dat5b[2]), .E(n63), .C(n262), .B(n58), .A(n61), .Y(n56)
         );
  MUX2X1 U248 ( .D0(n52), .D1(ps_dat5b[1]), .S(ps_dat5b[0]), .Y(n53) );
  NAND21X1 U249 ( .B(n77), .A(prx_bmc), .Y(n262) );
  INVX1 U250 ( .A(n47), .Y(n202) );
  GEN2XL U251 ( .D(cccnt[2]), .E(n46), .C(n45), .B(n44), .A(n43), .Y(n47) );
  NAND21XL U252 ( .B(cccnt[0]), .A(shrtrans), .Y(n46) );
  AO21XL U253 ( .B(cccnt[4]), .C(cccnt[3]), .A(cccnt[5]), .Y(n44) );
  INVX1 U254 ( .A(ps_dat5b[1]), .Y(n63) );
  AND2X1 U255 ( .A(n18), .B(n63), .Y(n52) );
  INVX1 U256 ( .A(prx_bmc), .Y(n72) );
  INVX1 U257 ( .A(n54), .Y(n59) );
  NAND21X1 U258 ( .B(n72), .A(ps_dat5b[1]), .Y(n54) );
  INVX1 U259 ( .A(ps_dat5b[2]), .Y(n65) );
  INVX1 U260 ( .A(ps_dat5b[0]), .Y(n61) );
  MUX2IXL U261 ( .D0(prx_rxcode[4]), .D1(prx_rxcode[3]), .S(n314), .Y(n114) );
  MUX2XL U262 ( .D0(N96), .D1(prx_crcsidat[3]), .S(n314), .Y(prx_fifowdat[7])
         );
  AO21X1 U263 ( .B(n25), .C(n63), .A(n62), .Y(N96) );
  GEN2XL U264 ( .D(n63), .E(n61), .C(n72), .B(n259), .A(n60), .Y(n62) );
  AND3X1 U265 ( .A(ps_dat5b[0]), .B(n66), .C(n59), .Y(n60) );
  INVX1 U266 ( .A(n71), .Y(n69) );
  INVX1 U267 ( .A(n262), .Y(n68) );
  AO21X1 U268 ( .B(n25), .C(ps_dat5b[0]), .A(n67), .Y(n70) );
  OR2X1 U269 ( .A(n73), .B(n24), .Y(prx_fifowdat[5]) );
  AOI21X1 U270 ( .B(ps_dat5b[0]), .C(n72), .A(n71), .Y(n24) );
  MUX2X1 U271 ( .D0(n66), .D1(n65), .S(ps_dat5b[1]), .Y(n67) );
  OAI31XL U272 ( .A(ps_dat5b[1]), .B(n259), .C(n61), .D(n58), .Y(n73) );
  XNOR2XL U273 ( .A(n259), .B(ps_dat5b[2]), .Y(n25) );
  AO21X1 U274 ( .B(n201), .C(n200), .A(n37), .Y(N75) );
  XOR2XL U275 ( .A(cccnt[4]), .B(n199), .Y(n201) );
  AO21X1 U276 ( .B(n194), .C(n200), .A(n37), .Y(N73) );
  XOR2XL U277 ( .A(cccnt[2]), .B(n193), .Y(n194) );
  NOR2X1 U278 ( .A(n259), .B(n27), .Y(prx_crcsidat[3]) );
  XNOR2XL U279 ( .A(ps_dat5b[1]), .B(n78), .Y(n27) );
  OAI211X1 U280 ( .C(prx_crcsidat[0]), .D(n64), .A(n263), .B(N96), .Y(n205) );
  AND2X1 U281 ( .A(prx_bmc), .B(n73), .Y(n64) );
  GEN2XL U282 ( .D(n199), .E(cccnt[4]), .C(cccnt[5]), .B(n200), .A(n37), .Y(
        N76) );
  OAI211X1 U283 ( .C(n157), .D(n311), .A(n186), .B(n120), .Y(n162) );
  OAI211X1 U284 ( .C(n302), .D(n183), .A(n185), .B(n276), .Y(n186) );
  AND2X1 U285 ( .A(n275), .B(prx_fifowdat[2]), .Y(n276) );
  MUX2AXL U286 ( .D0(n282), .D1(n131), .S(n125), .Y(n265) );
  AOI22X1 U287 ( .A(n284), .B(n308), .C(n283), .D(N32), .Y(n131) );
  NAND32X1 U288 ( .B(n83), .C(n147), .A(n138), .Y(n101) );
  AND3X1 U289 ( .A(n293), .B(n305), .C(n81), .Y(n83) );
  AND4X1 U290 ( .A(n296), .B(n9), .C(n148), .D(n309), .Y(n147) );
  OAI32X1 U293 ( .A(n88), .B(prx_crcsidat[0]), .C(prx_fifowdat[6]), .D(
        prx_fifowdat[1]), .E(n117), .Y(n81) );
  AND2X1 U294 ( .A(n113), .B(n112), .Y(N277) );
  INVX1 U295 ( .A(n212), .Y(n113) );
  OAI211XL U296 ( .C(prx_fsm[0]), .D(n206), .A(n126), .B(n208), .Y(n112) );
  INVX1 U298 ( .A(r_rgdcrc), .Y(n267) );
  OR2XL U299 ( .A(prx_rcvdords[2]), .B(n84), .Y(n115) );
  NAND43X1 U300 ( .B(prx_fifowdat[1]), .C(n114), .D(n144), .A(prx_fifowdat[2]), 
        .Y(n286) );
  NAND21XL U301 ( .B(bcnt[0]), .A(n218), .Y(n184) );
  NAND32X1 U302 ( .B(n79), .C(n132), .A(n229), .Y(n84) );
  INVX1 U303 ( .A(ordsbuf[3]), .Y(n79) );
  MUX3XL U304 ( .D0(r_ords_ena[0]), .D1(r_ords_ena[2]), .D2(n230), .S0(
        prx_rcvdords[1]), .S1(prx_rcvdords[2]), .Y(n231) );
  AND2X1 U305 ( .A(r_ords_ena[4]), .B(n229), .Y(n230) );
  MUX2IXL U306 ( .D0(n28), .D1(n29), .S(prx_rcvdords[0]), .Y(n269) );
  AOI21X1 U307 ( .B(r_ords_ena[5]), .C(n232), .A(n228), .Y(n28) );
  AOI21X1 U308 ( .B(r_ords_ena[6]), .C(n232), .A(n231), .Y(n29) );
  NAND5XL U309 ( .A(n303), .B(n121), .C(n225), .D(n134), .E(prx_rcvdords[0]), 
        .Y(n141) );
  OAI22X1 U310 ( .A(n189), .B(n188), .C(n187), .D(n184), .Y(N239) );
  MUX2BXL U311 ( .D0(n187), .D1(n180), .S(bcnt[1]), .Y(n189) );
  AND2XL U312 ( .A(bcnt[0]), .B(n187), .Y(n180) );
  MUX2AXL U313 ( .D0(n30), .D1(n295), .S(bcnt[1]), .Y(n307) );
  NAND2XL U314 ( .A(bcnt[0]), .B(n218), .Y(n30) );
  INVXL U315 ( .A(prx_rcvdords[0]), .Y(n132) );
  NOR32XL U316 ( .B(ordsbuf[4]), .C(ordsbuf[7]), .A(ordsbuf[6]), .Y(n178) );
  NAND21XL U317 ( .B(n84), .A(prx_rcvdords[2]), .Y(n91) );
  NAND21XL U318 ( .B(prx_fsm[3]), .A(n169), .Y(n174) );
  NAND32XL U319 ( .B(prx_fsm[2]), .C(n109), .A(n249), .Y(n127) );
  INVX1 U320 ( .A(n118), .Y(n134) );
  NAND21X1 U321 ( .B(n296), .A(ordsbuf[3]), .Y(n118) );
  NAND5XL U322 ( .A(n93), .B(n313), .C(n275), .D(n92), .E(n121), .Y(n137) );
  INVX1 U323 ( .A(n91), .Y(n92) );
  INVXL U324 ( .A(prx_rcvdords[1]), .Y(n229) );
  INVX1 U325 ( .A(prx_fifowdat[0]), .Y(n144) );
  INVX1 U326 ( .A(n136), .Y(n274) );
  NAND43X1 U327 ( .B(ordsbuf[4]), .C(n135), .D(n298), .A(ordsbuf[6]), .Y(n136)
         );
  INVX1 U328 ( .A(ordsbuf[7]), .Y(n135) );
  INVX1 U329 ( .A(r_ordrs4), .Y(n312) );
  NAND2X1 U330 ( .A(n178), .B(ordsbuf[5]), .Y(n176) );
  INVX1 U331 ( .A(prx_fifowdat[1]), .Y(n296) );
  INVXL U332 ( .A(prx_rcvdords[2]), .Y(n225) );
  INVX1 U333 ( .A(n82), .Y(n133) );
  NAND21X1 U334 ( .B(r_exist1st), .A(n5), .Y(n82) );
  INVX1 U335 ( .A(n130), .Y(n232) );
  NAND21XL U336 ( .B(n225), .A(prx_rcvdords[1]), .Y(n130) );
  AND2X1 U337 ( .A(n219), .B(prx_bmc), .Y(N156) );
  AND2X1 U338 ( .A(n219), .B(ps_dat5b[1]), .Y(N154) );
  AND2X1 U339 ( .A(n219), .B(ps_dat5b[2]), .Y(N155) );
  AND2X1 U340 ( .A(r_ords_ena[1]), .B(n225), .Y(n226) );
  INVX1 U341 ( .A(ordsbuf[5]), .Y(n298) );
  NAND41X1 U342 ( .D(ordsbuf[5]), .A(ordsbuf[4]), .B(ordsbuf[6]), .C(
        ordsbuf[7]), .Y(n140) );
  AND2XL U343 ( .A(r_ords_ena[3]), .B(prx_rcvdords[2]), .Y(n227) );
  INVXL U344 ( .A(bcnt[2]), .Y(n187) );
  INVX1 U345 ( .A(r_exist1st), .Y(n121) );
  AND2X1 U346 ( .A(n36), .B(n204), .Y(n214) );
  AND2XL U347 ( .A(n202), .B(n242), .Y(n203) );
  AND3XL U348 ( .A(pid_goidle), .B(n314), .C(n269), .Y(prx_setsta[5]) );
  NAND21XL U349 ( .B(prx_fsm[1]), .A(n166), .Y(n257) );
  NOR5XL U350 ( .A(cccnt[2]), .B(cccnt[3]), .C(cccnt[5]), .D(n272), .E(n271), 
        .Y(prx_cccnt[1]) );
  INVX1 U351 ( .A(n107), .Y(n166) );
  NAND21XL U352 ( .B(prx_fsm[0]), .A(n108), .Y(n107) );
  INVXL U353 ( .A(cccnt[4]), .Y(n272) );
  NAND21XL U354 ( .B(bcnt[1]), .A(n187), .Y(n258) );
  OA21X1 U355 ( .B(prx_bmc), .C(n259), .A(n258), .Y(n260) );
  BUFX3 U356 ( .A(prx_fifowdat[5]), .Y(prx_crcsidat[1]) );
  OAI211X1 U357 ( .C(prx_bmc), .D(n71), .A(n57), .B(n56), .Y(prx_fifowdat[4])
         );
  NAND21XL U358 ( .B(n77), .A(n14), .Y(n261) );
  NAND21X1 U359 ( .B(n16), .A(n243), .Y(n255) );
  MUX2XL U360 ( .D0(shrtrans), .D1(n203), .S(n11), .Y(n204) );
  MUX2IXL U361 ( .D0(n11), .D1(prx_cccnt[0]), .S(ptx_txact), .Y(n38) );
  NAND31XL U362 ( .C(n242), .A(n241), .B(cctrans), .Y(n243) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_adp ( clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, 
        r_adprx_en, r_adp2nd, adp_val, d_cc, cctrans, test_si, test_so, 
        test_se );
  output [5:0] adp_val;
  input clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, r_adprx_en,
         r_adp2nd, test_si, test_se;
  output d_cc, cctrans, test_so;
  wire   dcnt_n_2_, dcnt_n_1_, dcnt_n_0_, N49, N50, N51, N52, N53, N55, N97,
         N98, N99, N100, N101, N102, N103, N104, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N169, N170, N171, N172, N173, net10744, net10750, net10755, net10760,
         n115, n39, n41, n62, n64, n65, n66, n67, n68, n69, n70, n75, n91, n92,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n40, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n63, n71, n72, n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n150, n151, n152, n153, n154, n155, n156, n157,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7;
  wire   [7:0] dcnt_h;
  wire   [5:0] adp_v0;
  wire   [5:0] dcnt_e;

  SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 clk_gate_adp_n_reg ( .CLK(clk), .EN(N49), 
        .ENCLK(net10744), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 clk_gate_dcnt_e_reg ( .CLK(clk), .EN(N130), 
        .ENCLK(net10750), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 clk_gate_dcnt_h_reg ( .CLK(clk), .EN(N137), 
        .ENCLK(net10755), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 clk_gate_dcnt_n_reg ( .CLK(clk), .EN(N169), 
        .ENCLK(net10760), .TE(test_se) );
  phyrx_adp_DW01_inc_0 add_385 ( .A(dcnt_h), .SUM({N104, N103, N102, N101, 
        N100, N99, N98, N97}) );
  phyrx_adp_DW_div_tc_6 div_338 ( .a({n8, dcnt_h}), .b({1'b0, 1'b1, 1'b1, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, adp_v0}), .remainder({SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7}), .divide_by_0() );
  SDFFQX1 adp_n_reg_5_ ( .D(N55), .SIN(adp_val[4]), .SMC(test_se), .C(net10744), .Q(adp_val[5]) );
  SDFFQX1 dcnt_h_reg_6_ ( .D(N144), .SIN(dcnt_h[5]), .SMC(test_se), .C(
        net10755), .Q(dcnt_h[6]) );
  SDFFQX1 dcnt_h_reg_3_ ( .D(N141), .SIN(dcnt_h[2]), .SMC(test_se), .C(
        net10755), .Q(dcnt_h[3]) );
  SDFFQX1 dcnt_h_reg_4_ ( .D(N142), .SIN(dcnt_h[3]), .SMC(test_se), .C(
        net10755), .Q(dcnt_h[4]) );
  SDFFQX1 dcnt_h_reg_5_ ( .D(N143), .SIN(dcnt_h[4]), .SMC(test_se), .C(
        net10755), .Q(dcnt_h[5]) );
  SDFFQX1 dcnt_h_reg_1_ ( .D(N139), .SIN(dcnt_h[0]), .SMC(test_se), .C(
        net10755), .Q(dcnt_h[1]) );
  SDFFQX1 dcnt_h_reg_2_ ( .D(N140), .SIN(dcnt_h[1]), .SMC(test_se), .C(
        net10755), .Q(dcnt_h[2]) );
  SDFFQX1 dcnt_h_reg_0_ ( .D(N138), .SIN(dcnt_e[5]), .SMC(test_se), .C(
        net10755), .Q(dcnt_h[0]) );
  SDFFQX1 dcnt_h_reg_7_ ( .D(N145), .SIN(dcnt_h[6]), .SMC(test_se), .C(
        net10755), .Q(dcnt_h[7]) );
  SDFFQX1 adp_n_reg_4_ ( .D(n150), .SIN(adp_val[3]), .SMC(test_se), .C(
        net10744), .Q(adp_val[4]) );
  SDFFQX1 dcnt_n_reg_1_ ( .D(N171), .SIN(dcnt_n_0_), .SMC(test_se), .C(
        net10760), .Q(dcnt_n_1_) );
  SDFFQX1 dcnt_e_reg_4_ ( .D(N135), .SIN(dcnt_e[3]), .SMC(test_se), .C(
        net10750), .Q(dcnt_e[4]) );
  SDFFQX1 dcnt_e_reg_5_ ( .D(N136), .SIN(dcnt_e[4]), .SMC(test_se), .C(
        net10750), .Q(dcnt_e[5]) );
  SDFFQX1 dcnt_e_reg_2_ ( .D(N133), .SIN(dcnt_e[1]), .SMC(test_se), .C(
        net10750), .Q(dcnt_e[2]) );
  SDFFQX1 dcnt_e_reg_3_ ( .D(N134), .SIN(dcnt_e[2]), .SMC(test_se), .C(
        net10750), .Q(dcnt_e[3]) );
  SDFFQX1 adp_n_reg_2_ ( .D(N52), .SIN(adp_val[1]), .SMC(test_se), .C(net10744), .Q(adp_val[2]) );
  SDFFQX1 dcnt_n_reg_2_ ( .D(N172), .SIN(dcnt_n_1_), .SMC(test_se), .C(
        net10760), .Q(dcnt_n_2_) );
  SDFFQX1 dcnt_e_reg_1_ ( .D(N132), .SIN(dcnt_e[0]), .SMC(test_se), .C(
        net10750), .Q(dcnt_e[1]) );
  SDFFQX1 dcnt_n_reg_3_ ( .D(N173), .SIN(dcnt_n_2_), .SMC(test_se), .C(
        net10760), .Q(test_so) );
  SDFFQX1 adp_n_reg_0_ ( .D(N50), .SIN(test_si), .SMC(test_se), .C(net10744), 
        .Q(adp_val[0]) );
  SDFFQX1 cs_d_cc_reg ( .D(n115), .SIN(adp_val[5]), .SMC(test_se), .C(clk), 
        .Q(d_cc) );
  SDFFQX1 adp_n_reg_3_ ( .D(N53), .SIN(adp_val[2]), .SMC(test_se), .C(net10744), .Q(adp_val[3]) );
  SDFFQX1 dcnt_e_reg_0_ ( .D(N131), .SIN(d_cc), .SMC(test_se), .C(net10750), 
        .Q(dcnt_e[0]) );
  SDFFQX1 adp_n_reg_1_ ( .D(N51), .SIN(adp_val[0]), .SMC(test_se), .C(net10744), .Q(adp_val[1]) );
  SDFFQX1 dcnt_n_reg_0_ ( .D(N170), .SIN(n8), .SMC(test_se), .C(net10760), .Q(
        dcnt_n_0_) );
  NAND31X2 U5 ( .C(n148), .A(n147), .B(n146), .Y(cctrans) );
  INVXL U6 ( .A(n144), .Y(n6) );
  XOR2X1 U7 ( .A(n27), .B(dcnt_n_1_), .Y(n28) );
  INVX1 U8 ( .A(adp_val[1]), .Y(n27) );
  NOR2X1 U9 ( .A(dcnt_e[4]), .B(n22), .Y(n16) );
  INVX1 U10 ( .A(n136), .Y(n148) );
  INVX1 U11 ( .A(dcnt_e[3]), .Y(n140) );
  INVX1 U12 ( .A(dcnt_e[4]), .Y(n139) );
  INVX1 U13 ( .A(d_cc), .Y(n81) );
  NAND4X1 U14 ( .A(n17), .B(n18), .C(n3), .D(n28), .Y(n121) );
  XNOR2XL U15 ( .A(dcnt_n_2_), .B(adp_val[2]), .Y(n17) );
  XNOR2XL U16 ( .A(test_so), .B(adp_val[3]), .Y(n18) );
  NAND42X1 U17 ( .C(adp_val[0]), .D(adp_val[2]), .A(n27), .B(n23), .Y(n24) );
  NAND2X1 U18 ( .A(n137), .B(n24), .Y(n125) );
  XNOR2XL U19 ( .A(dcnt_n_0_), .B(adp_val[0]), .Y(n3) );
  BUFXL U20 ( .A(gohi), .Y(n4) );
  NAND31X4 U21 ( .C(n145), .A(n144), .B(d_cc), .Y(n146) );
  OAI31X1 U22 ( .A(n141), .B(n140), .C(n139), .D(n138), .Y(n144) );
  BUFXL U23 ( .A(golo), .Y(n5) );
  NAND32X2 U24 ( .B(d_cc), .C(n6), .A(n143), .Y(n147) );
  INVX1 U25 ( .A(dcnt_h[7]), .Y(n7) );
  INVX1 U26 ( .A(n7), .Y(n8) );
  INVXL U27 ( .A(n137), .Y(n138) );
  INVXL U28 ( .A(adp_val[3]), .Y(n23) );
  NAND21XL U29 ( .B(n20), .A(n106), .Y(n120) );
  AND2X2 U30 ( .A(gohi), .B(n142), .Y(n143) );
  NAND32X2 U31 ( .B(n121), .C(n125), .A(n118), .Y(n136) );
  AO21XL U32 ( .B(n103), .C(n131), .A(n102), .Y(N131) );
  AOI21XL U33 ( .B(n33), .C(n74), .A(n52), .Y(n14) );
  OAI211XL U34 ( .C(n131), .D(n130), .A(n129), .B(n128), .Y(N137) );
  AND2XL U35 ( .A(n121), .B(srstz), .Y(n122) );
  NAND32X1 U36 ( .B(dcnt_e[2]), .C(dcnt_e[1]), .A(n140), .Y(n73) );
  INVX1 U37 ( .A(n22), .Y(n78) );
  NAND21XL U38 ( .B(dcnt_e[0]), .A(n56), .Y(n22) );
  XOR2X1 U39 ( .A(n139), .B(dcnt_e[5]), .Y(n71) );
  NAND31XL U40 ( .C(n120), .A(n121), .B(n108), .Y(n123) );
  INVX1 U41 ( .A(srstz), .Y(n20) );
  NAND21X1 U42 ( .B(n101), .A(n151), .Y(n93) );
  OR2X1 U43 ( .A(n94), .B(n93), .Y(n98) );
  INVX1 U44 ( .A(n75), .Y(n80) );
  NAND21X1 U45 ( .B(n99), .A(n98), .Y(n39) );
  MUX2X1 U46 ( .D0(n97), .D1(n96), .S(n95), .Y(n99) );
  AND2X1 U47 ( .A(n94), .B(n93), .Y(n97) );
  INVX1 U48 ( .A(n92), .Y(n95) );
  INVX1 U49 ( .A(n42), .Y(n36) );
  INVX1 U50 ( .A(n104), .Y(n151) );
  INVX1 U51 ( .A(n41), .Y(n101) );
  INVX1 U52 ( .A(n96), .Y(n94) );
  OAI31XL U53 ( .A(n92), .B(n151), .C(n41), .D(n39), .Y(n91) );
  INVX1 U54 ( .A(n37), .Y(n38) );
  NAND21X1 U55 ( .B(n151), .A(n92), .Y(n100) );
  INVX1 U56 ( .A(n102), .Y(n51) );
  INVX1 U57 ( .A(k0_det), .Y(n132) );
  NOR3XL U58 ( .A(goidle), .B(gobusy), .C(n20), .Y(n75) );
  NAND21X1 U59 ( .B(n16), .A(n71), .Y(n137) );
  INVX1 U60 ( .A(n125), .Y(n106) );
  INVX1 U61 ( .A(n73), .Y(n56) );
  NAND21X1 U62 ( .B(adp_v0[5]), .A(adp_v0[4]), .Y(n42) );
  AO21X1 U63 ( .B(adp_v0[4]), .C(n42), .A(n38), .Y(n92) );
  AO21X1 U64 ( .B(n42), .C(n34), .A(n38), .Y(n41) );
  INVX1 U65 ( .A(adp_v0[1]), .Y(n34) );
  NAND32X1 U66 ( .B(n36), .C(adp_v0[0]), .A(n37), .Y(n104) );
  AO21X1 U67 ( .B(n42), .C(n40), .A(n38), .Y(n96) );
  INVX1 U68 ( .A(adp_v0[2]), .Y(n40) );
  OAI21BBX1 U69 ( .A(n9), .B(adp_v0[4]), .C(adp_v0[5]), .Y(n37) );
  OR3XL U70 ( .A(adp_v0[1]), .B(adp_v0[3]), .C(adp_v0[2]), .Y(n9) );
  XOR2X1 U71 ( .A(n10), .B(n11), .Y(n90) );
  AOI21X1 U72 ( .B(adp_v0[3]), .C(n37), .A(n36), .Y(n10) );
  NAND2X1 U73 ( .A(n98), .B(n92), .Y(n11) );
  NOR21XL U74 ( .B(n135), .A(n39), .Y(N52) );
  MUX2IX1 U75 ( .D0(n12), .D1(n13), .S(n101), .Y(N51) );
  NAND2X1 U76 ( .A(n150), .B(n104), .Y(n12) );
  NAND2X1 U77 ( .A(n135), .B(n100), .Y(n13) );
  AND2X1 U78 ( .A(n135), .B(n90), .Y(N53) );
  INVX1 U79 ( .A(n89), .Y(n150) );
  NAND21X1 U80 ( .B(n95), .A(n135), .Y(n89) );
  AND2X1 U81 ( .A(n135), .B(n104), .Y(N50) );
  AO21X1 U82 ( .B(n103), .C(n32), .A(n80), .Y(n102) );
  AO21X1 U83 ( .B(n63), .C(n61), .A(k0_det), .Y(n126) );
  INVX1 U84 ( .A(n72), .Y(n61) );
  INVX1 U85 ( .A(n52), .Y(n103) );
  INVX1 U86 ( .A(n79), .Y(n88) );
  NAND32X1 U87 ( .B(n80), .C(n129), .A(n81), .Y(n79) );
  OR2X1 U88 ( .A(n102), .B(n14), .Y(N132) );
  NOR3XL U89 ( .A(n81), .B(n80), .C(n129), .Y(n15) );
  OAI31XL U90 ( .A(n53), .B(n58), .C(n52), .D(n51), .Y(N136) );
  AND2X1 U91 ( .A(n127), .B(n75), .Y(n128) );
  INVX1 U92 ( .A(n126), .Y(n127) );
  NAND32X1 U93 ( .B(n73), .C(n72), .A(n71), .Y(n130) );
  NAND21X1 U94 ( .B(n135), .A(srstz), .Y(N49) );
  AND2X1 U95 ( .A(n135), .B(n58), .Y(N55) );
  OAI211X1 U96 ( .C(n125), .D(n124), .A(n123), .B(n122), .Y(N169) );
  AND3X1 U97 ( .A(n113), .B(n112), .C(n111), .Y(N171) );
  INVX1 U98 ( .A(n123), .Y(n113) );
  AOI211X1 U99 ( .C(n111), .D(n114), .A(n109), .B(n123), .Y(N172) );
  INVX1 U100 ( .A(n44), .Y(n63) );
  INVX1 U101 ( .A(n68), .Y(n155) );
  INVX1 U102 ( .A(n66), .Y(n154) );
  INVX1 U103 ( .A(n70), .Y(n152) );
  INVX1 U104 ( .A(n64), .Y(n153) );
  INVX1 U105 ( .A(n112), .Y(n119) );
  INVX1 U106 ( .A(n50), .Y(n48) );
  INVX1 U107 ( .A(n47), .Y(n35) );
  OAI21BX1 U108 ( .C(adp_val[4]), .B(n125), .A(golo), .Y(n145) );
  NAND21XL U109 ( .B(adp_val[4]), .A(n106), .Y(n142) );
  XOR2X1 U110 ( .A(n81), .B(adp_val[4]), .Y(n118) );
  NAND21XL U111 ( .B(n74), .A(dcnt_e[2]), .Y(n141) );
  NAND21XL U112 ( .B(n131), .A(dcnt_e[1]), .Y(n74) );
  INVXL U113 ( .A(dcnt_e[0]), .Y(n131) );
  GEN2XL U114 ( .D(dcnt_e[3]), .E(n47), .C(n48), .B(n103), .A(n46), .Y(N134)
         );
  OAI31XL U115 ( .A(n45), .B(n133), .C(n44), .D(n51), .Y(n46) );
  AOI211X1 U116 ( .C(n43), .D(n41), .A(n91), .B(n90), .Y(n45) );
  INVX1 U117 ( .A(n100), .Y(n43) );
  NAND43X1 U118 ( .B(dcnt_e[3]), .C(n126), .D(n78), .A(n77), .Y(n129) );
  NOR32XL U119 ( .B(n130), .C(n141), .A(n76), .Y(n77) );
  AND2XL U120 ( .A(dcnt_e[5]), .B(n139), .Y(n76) );
  NAND43X1 U121 ( .B(n63), .C(n133), .D(n134), .A(n31), .Y(n52) );
  NAND32XL U122 ( .B(r_adp2nd), .C(n73), .A(n30), .Y(n31) );
  GEN2XL U123 ( .D(n153), .E(dcnt_h[6]), .C(n62), .B(n88), .A(n82), .Y(N144)
         );
  AND2X1 U124 ( .A(N103), .B(n15), .Y(n82) );
  GEN2XL U125 ( .D(dcnt_h[1]), .E(dcnt_h[0]), .C(n85), .B(n88), .A(n84), .Y(
        N139) );
  INVX1 U126 ( .A(n156), .Y(n85) );
  AND2X1 U127 ( .A(N98), .B(n15), .Y(n84) );
  GEN2XL U128 ( .D(dcnt_h[2]), .E(n156), .C(n70), .B(n88), .A(n86), .Y(N140)
         );
  AND2X1 U129 ( .A(N99), .B(n15), .Y(n86) );
  AO22AXL U130 ( .A(N102), .B(n15), .C(n88), .D(n65), .Y(N143) );
  AOI21X1 U131 ( .B(dcnt_h[5]), .C(n154), .A(n64), .Y(n65) );
  AO22AXL U132 ( .A(N101), .B(n15), .C(n88), .D(n67), .Y(N142) );
  AOI21X1 U133 ( .B(dcnt_h[4]), .C(n155), .A(n66), .Y(n67) );
  AO22AXL U134 ( .A(N100), .B(n15), .C(n88), .D(n69), .Y(N141) );
  AOI21X1 U135 ( .B(dcnt_h[3]), .C(n152), .A(n68), .Y(n69) );
  AO22X1 U136 ( .A(N97), .B(n15), .C(n88), .D(n83), .Y(N138) );
  AO22X1 U137 ( .A(N104), .B(n15), .C(n88), .D(n87), .Y(N145) );
  XOR2X1 U138 ( .A(dcnt_h[7]), .B(n62), .Y(n87) );
  OAI211X1 U139 ( .C(n132), .D(n32), .A(n59), .B(n157), .Y(n133) );
  GEN2XL U140 ( .D(dcnt_e[4]), .E(n50), .C(n53), .B(n103), .A(n102), .Y(N135)
         );
  GEN2XL U141 ( .D(dcnt_e[2]), .E(n33), .C(n35), .B(n103), .A(n102), .Y(N133)
         );
  OAI221X1 U142 ( .A(n134), .B(n133), .C(n32), .D(n132), .E(n75), .Y(N130) );
  NAND2XL U143 ( .A(n19), .B(n136), .Y(n59) );
  MUX2IXL U144 ( .D0(n26), .D1(n25), .S(d_cc), .Y(n19) );
  NAND21X1 U145 ( .B(n60), .A(n157), .Y(n72) );
  INVX1 U146 ( .A(i_ccidle), .Y(n157) );
  INVX1 U147 ( .A(n59), .Y(n60) );
  INVX1 U148 ( .A(n57), .Y(n135) );
  NAND5XL U149 ( .A(dcnt_e[0]), .B(srstz), .C(n56), .D(n71), .E(n55), .Y(n57)
         );
  MUX2XL U150 ( .D0(n4), .D1(n5), .S(d_cc), .Y(n55) );
  NAND5XL U151 ( .A(n119), .B(n118), .C(n117), .D(n116), .E(n114), .Y(n124) );
  MUX2XL U152 ( .D0(n4), .D1(n5), .S(adp_val[4]), .Y(n116) );
  OAI22XL U153 ( .A(n120), .B(n124), .C(dcnt_n_0_), .D(n123), .Y(N170) );
  AND2X1 U154 ( .A(n54), .B(srstz), .Y(n115) );
  XOR2XL U155 ( .A(n59), .B(d_cc), .Y(n54) );
  NAND31XL U156 ( .C(dcnt_n_2_), .A(n117), .B(n119), .Y(n108) );
  AND2X1 U157 ( .A(n110), .B(n113), .Y(N173) );
  XOR2XL U158 ( .A(test_so), .B(n109), .Y(n110) );
  NAND21X1 U159 ( .B(dcnt_h[1]), .A(n83), .Y(n156) );
  NAND32XL U160 ( .B(dcnt_e[5]), .C(n73), .A(n30), .Y(n44) );
  NOR2X1 U161 ( .A(n152), .B(dcnt_h[3]), .Y(n68) );
  NOR2X1 U162 ( .A(n155), .B(dcnt_h[4]), .Y(n66) );
  NOR2X1 U163 ( .A(n154), .B(dcnt_h[5]), .Y(n64) );
  NOR2X1 U164 ( .A(n156), .B(dcnt_h[2]), .Y(n70) );
  INVX1 U165 ( .A(n21), .Y(n30) );
  NAND21XL U166 ( .B(n139), .A(dcnt_e[0]), .Y(n21) );
  INVX1 U167 ( .A(dcnt_h[0]), .Y(n83) );
  INVX1 U168 ( .A(r_adprx_en), .Y(n32) );
  INVX1 U169 ( .A(n29), .Y(n134) );
  NAND21XL U170 ( .B(dcnt_e[5]), .A(n16), .Y(n29) );
  NOR2X1 U171 ( .A(n153), .B(dcnt_h[6]), .Y(n62) );
  NAND21XL U172 ( .B(dcnt_e[1]), .A(n131), .Y(n33) );
  NAND21XL U173 ( .B(dcnt_n_1_), .A(n107), .Y(n112) );
  NAND21XL U174 ( .B(dcnt_e[3]), .A(n35), .Y(n50) );
  NAND21XL U175 ( .B(n107), .A(dcnt_n_1_), .Y(n111) );
  OR2XL U176 ( .A(dcnt_e[2]), .B(n33), .Y(n47) );
  INVX1 U177 ( .A(n105), .Y(n109) );
  NAND21XL U178 ( .B(n111), .A(dcnt_n_2_), .Y(n105) );
  INVXL U179 ( .A(dcnt_n_0_), .Y(n107) );
  INVX1 U180 ( .A(n49), .Y(n53) );
  NAND21XL U181 ( .B(dcnt_e[4]), .A(n48), .Y(n49) );
  INVXL U182 ( .A(test_so), .Y(n117) );
  INVXL U183 ( .A(dcnt_n_2_), .Y(n114) );
  INVXL U184 ( .A(dcnt_e[5]), .Y(n58) );
  INVXL U185 ( .A(n145), .Y(n25) );
  AND2XL U186 ( .A(n4), .B(n142), .Y(n26) );
endmodule


module phyrx_adp_DW_div_tc_6 ( a, b, quotient, remainder, divide_by_0 );
  input [8:0] a;
  input [3:0] b;
  output [8:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   u_div_SumTmp_1__0_, u_div_SumTmp_1__2_, u_div_SumTmp_2__0_,
         u_div_SumTmp_3__0_, u_div_SumTmp_4__0_, u_div_SumTmp_5__0_,
         u_div_CryTmp_0__2_, u_div_CryTmp_0__3_, u_div_CryTmp_0__4_,
         u_div_CryTmp_1__4_, u_div_CryTmp_2__4_, u_div_CryTmp_3__4_,
         u_div_CryTmp_4__4_, u_div_CryTmp_5__4_, u_div_PartRem_1__2_,
         u_div_PartRem_1__3_, u_div_PartRem_2__3_, u_div_PartRem_3__3_,
         u_div_PartRem_4__3_, u_div_PartRem_5__3_, u_div_PartRem_7__0_,
         u_div_PartRem_7__1_, n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12,
         n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32;
  wire   [5:1] u_div_QIncCry;
  wire   [5:0] u_div_QInv;
  wire   [6:1] u_div_AIncCry;
  wire   [6:0] u_div_AInv;

  HAD1X1 u_div_u_ha_AInc_6 ( .A(u_div_AInv[6]), .B(u_div_AIncCry[6]), .CO(
        u_div_PartRem_7__1_), .SO(u_div_PartRem_7__0_) );
  HAD1X1 u_div_u_ha_AInc_5 ( .A(u_div_AInv[5]), .B(u_div_AIncCry[5]), .CO(
        u_div_AIncCry[6]), .SO(u_div_SumTmp_5__0_) );
  HAD1X1 u_div_u_ha_AInc_4 ( .A(u_div_AInv[4]), .B(u_div_AIncCry[4]), .CO(
        u_div_AIncCry[5]), .SO(u_div_SumTmp_4__0_) );
  HAD1X1 u_div_u_ha_AInc_3 ( .A(u_div_AInv[3]), .B(u_div_AIncCry[3]), .CO(
        u_div_AIncCry[4]), .SO(u_div_SumTmp_3__0_) );
  HAD1X1 u_div_u_ha_AInc_2 ( .A(u_div_AInv[2]), .B(u_div_AIncCry[2]), .CO(
        u_div_AIncCry[3]), .SO(u_div_SumTmp_2__0_) );
  HAD1X1 u_div_u_ha_AInc_1 ( .A(u_div_AInv[1]), .B(u_div_AIncCry[1]), .CO(
        u_div_AIncCry[2]), .SO(u_div_SumTmp_1__0_) );
  HAD1X1 u_div_u_ha_QInc_4 ( .A(u_div_QInv[4]), .B(u_div_QIncCry[4]), .CO(
        u_div_QIncCry[5]), .SO(quotient[4]) );
  HAD1X1 u_div_u_ha_QInc_3 ( .A(u_div_QInv[3]), .B(u_div_QIncCry[3]), .CO(
        u_div_QIncCry[4]), .SO(quotient[3]) );
  HAD1X1 u_div_u_ha_QInc_2 ( .A(u_div_QInv[2]), .B(u_div_QIncCry[2]), .CO(
        u_div_QIncCry[3]), .SO(quotient[2]) );
  HAD1X1 u_div_u_ha_QInc_1 ( .A(u_div_QInv[1]), .B(u_div_QIncCry[1]), .CO(
        u_div_QIncCry[2]), .SO(quotient[1]) );
  HAD1X1 u_div_u_ha_QInc_0 ( .A(u_div_QInv[0]), .B(a[7]), .CO(u_div_QIncCry[1]), .SO(quotient[0]) );
  AND2X1 u_div_u_ha_AInc_0 ( .A(u_div_AInv[0]), .B(a[8]), .Y(u_div_AIncCry[1])
         );
  XOR2X1 u_div_u_ha_QInc_5 ( .A(u_div_QInv[5]), .B(u_div_QIncCry[5]), .Y(
        quotient[5]) );
  XOR2X1 U1 ( .A(n26), .B(n25), .Y(u_div_SumTmp_1__2_) );
  INVX1 U2 ( .A(n18), .Y(n28) );
  INVX1 U3 ( .A(n19), .Y(n27) );
  INVX1 U4 ( .A(n20), .Y(n25) );
  NAND21X1 U5 ( .B(u_div_PartRem_3__3_), .A(n2), .Y(u_div_CryTmp_2__4_) );
  MUX2IX1 U6 ( .D0(n18), .D1(n6), .S(u_div_CryTmp_3__4_), .Y(
        u_div_PartRem_3__3_) );
  NAND2X1 U7 ( .A(n27), .B(n12), .Y(n2) );
  XNOR2XL U8 ( .A(n11), .B(n28), .Y(n6) );
  MUX2AXL U9 ( .D0(n10), .D1(n10), .S(u_div_CryTmp_4__4_), .Y(n18) );
  MUX2AXL U10 ( .D0(n11), .D1(n11), .S(u_div_CryTmp_3__4_), .Y(n19) );
  NAND21X1 U11 ( .B(u_div_PartRem_4__3_), .A(n1), .Y(u_div_CryTmp_3__4_) );
  MUX2IX1 U12 ( .D0(n17), .D1(n5), .S(u_div_CryTmp_4__4_), .Y(
        u_div_PartRem_4__3_) );
  NAND2X1 U13 ( .A(n28), .B(n11), .Y(n1) );
  XNOR2XL U14 ( .A(n10), .B(n31), .Y(n5) );
  MUX2AXL U15 ( .D0(n12), .D1(n12), .S(u_div_CryTmp_2__4_), .Y(n20) );
  MUX2AXL U16 ( .D0(n21), .D1(n21), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__2_) );
  INVX1 U17 ( .A(n21), .Y(n26) );
  INVX1 U18 ( .A(u_div_CryTmp_0__3_), .Y(n23) );
  NOR21XL U19 ( .B(u_div_CryTmp_0__2_), .A(n24), .Y(u_div_CryTmp_0__3_) );
  MUX2IX1 U20 ( .D0(n32), .D1(n32), .S(u_div_CryTmp_1__4_), .Y(
        u_div_CryTmp_0__2_) );
  INVX1 U21 ( .A(u_div_PartRem_1__2_), .Y(n24) );
  INVX1 U22 ( .A(n17), .Y(n31) );
  NAND21X1 U23 ( .B(u_div_PartRem_2__3_), .A(n4), .Y(u_div_CryTmp_1__4_) );
  MUX2IX1 U24 ( .D0(n19), .D1(n7), .S(u_div_CryTmp_2__4_), .Y(
        u_div_PartRem_2__3_) );
  NAND2X1 U25 ( .A(n25), .B(n26), .Y(n4) );
  XNOR2XL U26 ( .A(n12), .B(n27), .Y(n7) );
  MUX2IX1 U27 ( .D0(u_div_SumTmp_2__0_), .D1(u_div_SumTmp_2__0_), .S(
        u_div_CryTmp_2__4_), .Y(n21) );
  MUX2AXL U28 ( .D0(u_div_PartRem_7__0_), .D1(u_div_PartRem_7__0_), .S(
        u_div_CryTmp_5__4_), .Y(n17) );
  AND2X1 U29 ( .A(u_div_PartRem_7__1_), .B(u_div_PartRem_7__0_), .Y(
        u_div_CryTmp_5__4_) );
  NAND21X1 U30 ( .B(u_div_PartRem_5__3_), .A(n3), .Y(u_div_CryTmp_4__4_) );
  MUX2IX1 U31 ( .D0(n29), .D1(n8), .S(u_div_CryTmp_5__4_), .Y(
        u_div_PartRem_5__3_) );
  NAND2X1 U32 ( .A(n31), .B(n10), .Y(n3) );
  INVX1 U33 ( .A(u_div_PartRem_7__1_), .Y(n29) );
  MUX2X1 U34 ( .D0(u_div_SumTmp_5__0_), .D1(u_div_SumTmp_5__0_), .S(
        u_div_CryTmp_5__4_), .Y(n10) );
  MUX2X1 U35 ( .D0(u_div_SumTmp_4__0_), .D1(u_div_SumTmp_4__0_), .S(
        u_div_CryTmp_4__4_), .Y(n11) );
  MUX2X1 U36 ( .D0(u_div_SumTmp_3__0_), .D1(u_div_SumTmp_3__0_), .S(
        u_div_CryTmp_3__4_), .Y(n12) );
  XNOR2XL U37 ( .A(u_div_PartRem_7__0_), .B(u_div_PartRem_7__1_), .Y(n8) );
  INVX1 U38 ( .A(u_div_SumTmp_1__0_), .Y(n32) );
  XOR2X1 U39 ( .A(a[7]), .B(u_div_CryTmp_4__4_), .Y(u_div_QInv[4]) );
  XOR2X1 U40 ( .A(a[8]), .B(a[6]), .Y(u_div_AInv[6]) );
  XNOR2XL U41 ( .A(a[7]), .B(n30), .Y(u_div_QInv[5]) );
  INVX1 U42 ( .A(u_div_CryTmp_5__4_), .Y(n30) );
  XOR2X1 U43 ( .A(a[7]), .B(u_div_CryTmp_0__4_), .Y(u_div_QInv[0]) );
  NAND21X1 U44 ( .B(u_div_PartRem_1__3_), .A(n23), .Y(u_div_CryTmp_0__4_) );
  MUX2AXL U45 ( .D0(n20), .D1(u_div_SumTmp_1__2_), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__3_) );
  XOR2X1 U46 ( .A(a[8]), .B(a[1]), .Y(u_div_AInv[1]) );
  XOR2X1 U47 ( .A(a[8]), .B(a[0]), .Y(u_div_AInv[0]) );
  XOR2X1 U48 ( .A(a[8]), .B(a[2]), .Y(u_div_AInv[2]) );
  XOR2X1 U49 ( .A(a[8]), .B(a[3]), .Y(u_div_AInv[3]) );
  XOR2X1 U50 ( .A(a[8]), .B(a[4]), .Y(u_div_AInv[4]) );
  XOR2X1 U51 ( .A(a[8]), .B(a[5]), .Y(u_div_AInv[5]) );
  XOR2X1 U52 ( .A(a[7]), .B(u_div_CryTmp_1__4_), .Y(u_div_QInv[1]) );
  XOR2X1 U53 ( .A(a[7]), .B(u_div_CryTmp_2__4_), .Y(u_div_QInv[2]) );
  XOR2X1 U54 ( .A(a[7]), .B(u_div_CryTmp_3__4_), .Y(u_div_QInv[3]) );
endmodule


module phyrx_adp_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_db ( clk, srstz, x_cc, ptx_txact, r_rxdb_opt, gohi, golo, gotrans, 
        test_si, test_so, test_se );
  input [1:0] r_rxdb_opt;
  input clk, srstz, x_cc, ptx_txact, test_si, test_se;
  output gohi, golo, gotrans, test_so;
  wire   cc_buf_6_, cc_buf_5_, cc_buf_4_, cc_buf_3_, cc_buf_1_, N11, N12, N13,
         N14, N15, N16, N17, N18, net168382, net81680, net81685, net81687,
         net81696, net81697, net81701, net81703, net81721, net81723, net81724,
         net81725, net92135, net92162, net92165, net95574, net98443, net99302,
         net99737, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52;

  SDFFQX1 cc_buf_reg_3_ ( .D(N14), .SIN(net98443), .SMC(test_se), .C(clk), .Q(
        cc_buf_3_) );
  SDFFQX1 cc_buf_reg_5_ ( .D(N16), .SIN(cc_buf_4_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_5_) );
  SDFFQX1 cc_buf_reg_4_ ( .D(N15), .SIN(cc_buf_3_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_4_) );
  SDFFQXX2 cc_buf_reg_0_ ( .D(N11), .SIN(test_si), .SMC(test_se), .C(clk), .Q(
        net168382), .XQ(net81721) );
  SDFFQX4 cc_buf_reg_2_ ( .D(N13), .SIN(n6), .SMC(test_se), .C(clk), .Q(
        net98443) );
  SDFFQX2 cc_buf_reg_7_ ( .D(N18), .SIN(cc_buf_6_), .SMC(test_se), .C(clk), 
        .Q(test_so) );
  SDFFQX2 cc_buf_reg_1_ ( .D(N12), .SIN(n28), .SMC(test_se), .C(clk), .Q(
        cc_buf_1_) );
  SDFFQX1 cc_buf_reg_6_ ( .D(N17), .SIN(cc_buf_5_), .SMC(test_se), .C(clk), 
        .Q(cc_buf_6_) );
  OAI21BX1 U3 ( .C(n39), .B(cc_buf_5_), .A(n38), .Y(n43) );
  NAND2XL U4 ( .A(n48), .B(r_rxdb_opt[1]), .Y(n32) );
  NAND21X1 U5 ( .B(net81701), .A(n44), .Y(n52) );
  INVXL U6 ( .A(cc_buf_6_), .Y(n19) );
  INVXL U7 ( .A(cc_buf_1_), .Y(n1) );
  INVX1 U8 ( .A(net81680), .Y(net99737) );
  INVX1 U9 ( .A(r_rxdb_opt[0]), .Y(n29) );
  AND2XL U10 ( .A(net92135), .B(cc_buf_6_), .Y(n12) );
  NAND21X2 U11 ( .B(n15), .A(n16), .Y(net99302) );
  INVX1 U12 ( .A(cc_buf_4_), .Y(n39) );
  INVX1 U13 ( .A(net81697), .Y(n17) );
  NAND2X1 U14 ( .A(n36), .B(n37), .Y(n41) );
  NAND2X1 U15 ( .A(n6), .B(net98443), .Y(n37) );
  INVX1 U16 ( .A(n26), .Y(net95574) );
  XOR3X1 U17 ( .A(net98443), .B(n28), .C(n5), .Y(n25) );
  INVX1 U18 ( .A(cc_buf_3_), .Y(net81685) );
  AND2X1 U19 ( .A(cc_buf_6_), .B(test_so), .Y(n21) );
  AND2X2 U20 ( .A(n18), .B(n19), .Y(n20) );
  AND3X1 U21 ( .A(net81687), .B(net99302), .C(n35), .Y(n34) );
  NAND2X1 U22 ( .A(n32), .B(n33), .Y(n31) );
  OR2X1 U23 ( .A(r_rxdb_opt[1]), .B(net92162), .Y(n33) );
  INVX2 U24 ( .A(cc_buf_1_), .Y(n26) );
  OR2X1 U25 ( .A(net95574), .B(net98443), .Y(n36) );
  INVX3 U26 ( .A(n22), .Y(n7) );
  NAND2X1 U27 ( .A(n10), .B(n9), .Y(net81696) );
  NAND2X2 U28 ( .A(net81723), .B(net98443), .Y(n16) );
  INVX1 U29 ( .A(net81724), .Y(n15) );
  INVXL U30 ( .A(n11), .Y(n30) );
  XOR2X1 U31 ( .A(n2), .B(n1), .Y(n24) );
  XNOR2X1 U32 ( .A(net98443), .B(net168382), .Y(n2) );
  INVX3 U33 ( .A(test_so), .Y(n18) );
  XOR2X2 U34 ( .A(cc_buf_6_), .B(net92165), .Y(n3) );
  XOR2X1 U35 ( .A(n3), .B(n41), .Y(n46) );
  NAND31XL U36 ( .C(net81685), .A(net98443), .B(n15), .Y(net81680) );
  NAND31XL U37 ( .C(net98443), .A(net81685), .B(n14), .Y(net81725) );
  NAND2XL U38 ( .A(n46), .B(n45), .Y(n4) );
  INVXL U39 ( .A(n26), .Y(n5) );
  INVX1 U40 ( .A(n26), .Y(n6) );
  XNOR2X1 U41 ( .A(net99302), .B(n7), .Y(n27) );
  XOR3X1 U42 ( .A(n11), .B(net81696), .C(net81697), .Y(n49) );
  OAI21BX1 U43 ( .C(n43), .B(cc_buf_3_), .A(n42), .Y(n45) );
  NAND2X1 U44 ( .A(n8), .B(n22), .Y(n9) );
  NAND2X1 U45 ( .A(n7), .B(net99302), .Y(n10) );
  INVX3 U46 ( .A(net99302), .Y(n8) );
  NOR2X2 U47 ( .A(n46), .B(n45), .Y(n11) );
  NAND21XL U48 ( .B(n18), .A(n25), .Y(n13) );
  NAND21X1 U49 ( .B(n12), .A(n13), .Y(net81687) );
  NAND21X2 U50 ( .B(n21), .A(n23), .Y(n22) );
  AND2XL U51 ( .A(net81724), .B(net81723), .Y(gotrans) );
  NAND21X1 U52 ( .B(n20), .A(n24), .Y(n23) );
  INVXL U53 ( .A(net81723), .Y(n14) );
  NOR21X1 U54 ( .B(n17), .A(n27), .Y(net81701) );
  NAND21X1 U55 ( .B(n17), .A(n27), .Y(net81703) );
  BUFXL U56 ( .A(net168382), .Y(n28) );
  XNOR2X1 U57 ( .A(net168382), .B(n18), .Y(net92165) );
  MUX2IX1 U58 ( .D0(n50), .D1(net99737), .S(n29), .Y(n51) );
  AND4X2 U59 ( .A(n49), .B(r_rxdb_opt[1]), .C(n30), .D(n4), .Y(n47) );
  NAND21X1 U60 ( .B(n34), .A(n51), .Y(gohi) );
  AND2XL U61 ( .A(n49), .B(n48), .Y(n50) );
  NOR2X2 U62 ( .A(n47), .B(n31), .Y(golo) );
  INVXL U63 ( .A(n52), .Y(n35) );
  NAND21X1 U64 ( .B(n5), .A(net81721), .Y(net81723) );
  NAND21X1 U65 ( .B(net81721), .A(n5), .Y(net81724) );
  XNOR2XL U66 ( .A(n41), .B(net92165), .Y(net92135) );
  NAND21X1 U67 ( .B(n11), .A(net81703), .Y(n44) );
  INVX1 U68 ( .A(net81725), .Y(net92162) );
  NAND21X1 U69 ( .B(n43), .A(cc_buf_3_), .Y(n42) );
  AND2X1 U70 ( .A(x_cc), .B(srstz), .Y(N11) );
  OAI21BBX1 U71 ( .A(net99302), .B(net81687), .C(n52), .Y(n48) );
  NAND21X1 U72 ( .B(n40), .A(n42), .Y(net81697) );
  INVX1 U73 ( .A(n38), .Y(n40) );
  NAND21X1 U74 ( .B(n39), .A(cc_buf_5_), .Y(n38) );
  AND2XL U75 ( .A(srstz), .B(net98443), .Y(N14) );
  AND2XL U76 ( .A(srstz), .B(cc_buf_5_), .Y(N17) );
  AND2XL U77 ( .A(srstz), .B(cc_buf_3_), .Y(N15) );
  AND2XL U78 ( .A(srstz), .B(cc_buf_6_), .Y(N18) );
  AND2XL U79 ( .A(srstz), .B(cc_buf_4_), .Y(N16) );
  AND2XL U80 ( .A(srstz), .B(n28), .Y(N12) );
  NOR32XL U81 ( .B(srstz), .C(n5), .A(ptx_txact), .Y(N13) );
endmodule


module i2cslv_a0 ( i_sda, i_scl, o_sda, i_deva, i_inc, i_fwnak, i_fwack, o_we, 
        o_re, o_r_early, o_idle, o_dec, o_busev, o_ofs, o_lt_ofs, o_wdat, 
        o_lt_buf, o_dbgpo, i_rdat, i_rd_mem, i_clk, i_rstz, i_prefetch, 
        test_si, test_se );
  input [7:1] i_deva;
  output [3:0] o_busev;
  output [7:0] o_ofs;
  output [7:0] o_lt_ofs;
  output [7:0] o_wdat;
  output [7:0] o_lt_buf;
  output [7:0] o_dbgpo;
  input [7:0] i_rdat;
  input i_sda, i_scl, i_inc, i_fwnak, i_fwack, i_rd_mem, i_clk, i_rstz,
         i_prefetch, test_si, test_se;
  output o_sda, o_we, o_re, o_r_early, o_idle, o_dec;
  wire   i2c_scl, sdafall, cs_rwb, N74, N75, N76, N77, N78, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, ps_rwbuf_0_, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, net10777, net10783, net10788, net10793,
         net10798, n118, n119, n120, n121, n16, n17, n18, n19, n20, n62, n85,
         n86, n87, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179;
  wire   [1:0] cs_sta;

  INVX1 U63 ( .A(n20), .Y(n17) );
  INVX1 U64 ( .A(n20), .Y(n18) );
  INVX1 U65 ( .A(n20), .Y(n19) );
  INVX1 U67 ( .A(n20), .Y(n16) );
  INVX1 U68 ( .A(i_rstz), .Y(n20) );
  i2cdbnc_a0_1 db_scl ( .i_clk(i_clk), .i_rstz(n16), .i_i2c(i_scl), .r_opt({
        1'b1, 1'b0}), .o_i2c(i2c_scl), .rise(o_dbgpo[6]), .fall(o_dbgpo[7]), 
        .test_si(cs_sta[1]), .test_se(test_se) );
  i2cdbnc_a0_0 db_sda ( .i_clk(i_clk), .i_rstz(n16), .i_i2c(i_sda), .r_opt({
        1'b0, 1'b0}), .o_i2c(ps_rwbuf_0_), .rise(o_dbgpo[5]), .fall(sdafall), 
        .test_si(i2c_scl), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 clk_gate_cs_bit_reg ( .CLK(i_clk), .EN(N74), 
        .ENCLK(net10777), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 clk_gate_adcnt_reg ( .CLK(i_clk), .EN(N114), 
        .ENCLK(net10783), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 clk_gate_rwbuf_reg ( .CLK(i_clk), .EN(N144), 
        .ENCLK(net10788), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 clk_gate_lt_buf_reg ( .CLK(i_clk), .EN(N179), .ENCLK(net10793), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 clk_gate_lt_ofs_reg ( .CLK(i_clk), .EN(
        o_busev[2]), .ENCLK(net10798), .TE(test_se) );
  SDFFQX1 lt_ofs_reg_7_ ( .D(o_wdat[7]), .SIN(o_lt_ofs[6]), .SMC(test_se), .C(
        net10798), .Q(o_lt_ofs[7]) );
  SDFFQX1 lt_buf_reg_7_ ( .D(N187), .SIN(o_lt_buf[6]), .SMC(test_se), .C(
        net10793), .Q(o_lt_buf[7]) );
  SDFFQX1 lt_ofs_reg_6_ ( .D(o_wdat[6]), .SIN(o_lt_ofs[5]), .SMC(test_se), .C(
        net10798), .Q(o_lt_ofs[6]) );
  SDFFQX1 lt_buf_reg_6_ ( .D(N186), .SIN(o_lt_buf[5]), .SMC(test_se), .C(
        net10793), .Q(o_lt_buf[6]) );
  SDFFQX1 lt_ofs_reg_5_ ( .D(o_wdat[5]), .SIN(o_lt_ofs[4]), .SMC(test_se), .C(
        net10798), .Q(o_lt_ofs[5]) );
  SDFFQX1 lt_buf_reg_5_ ( .D(N185), .SIN(o_lt_buf[4]), .SMC(test_se), .C(
        net10793), .Q(o_lt_buf[5]) );
  SDFFQX1 lt_ofs_reg_4_ ( .D(o_wdat[4]), .SIN(o_lt_ofs[3]), .SMC(test_se), .C(
        net10798), .Q(o_lt_ofs[4]) );
  SDFFQX1 lt_buf_reg_4_ ( .D(N184), .SIN(o_lt_buf[3]), .SMC(test_se), .C(
        net10793), .Q(o_lt_buf[4]) );
  SDFFQX1 lt_ofs_reg_3_ ( .D(o_wdat[3]), .SIN(o_lt_ofs[2]), .SMC(test_se), .C(
        net10798), .Q(o_lt_ofs[3]) );
  SDFFQX1 lt_buf_reg_3_ ( .D(N183), .SIN(o_lt_buf[2]), .SMC(test_se), .C(
        net10793), .Q(o_lt_buf[3]) );
  SDFFSQX1 sdat_reg ( .D(n118), .SIN(o_wdat[7]), .SMC(test_se), .C(i_clk), 
        .XS(n17), .Q(o_sda) );
  SDFFQX1 lt_ofs_reg_2_ ( .D(o_wdat[2]), .SIN(o_lt_ofs[1]), .SMC(test_se), .C(
        net10798), .Q(o_lt_ofs[2]) );
  SDFFQX1 lt_buf_reg_2_ ( .D(N182), .SIN(o_lt_buf[1]), .SMC(test_se), .C(
        net10793), .Q(o_lt_buf[2]) );
  SDFFQX1 lt_ofs_reg_0_ ( .D(o_wdat[0]), .SIN(o_lt_buf[7]), .SMC(test_se), .C(
        net10798), .Q(o_lt_ofs[0]) );
  SDFFQX1 lt_buf_reg_0_ ( .D(N180), .SIN(ps_rwbuf_0_), .SMC(test_se), .C(
        net10793), .Q(o_lt_buf[0]) );
  SDFFQX1 lt_ofs_reg_1_ ( .D(o_wdat[1]), .SIN(o_lt_ofs[0]), .SMC(test_se), .C(
        net10798), .Q(o_lt_ofs[1]) );
  SDFFQX1 lt_buf_reg_1_ ( .D(N181), .SIN(o_lt_buf[0]), .SMC(test_se), .C(
        net10793), .Q(o_lt_buf[1]) );
  SDFFRQX1 adcnt_reg_5_ ( .D(N111), .SIN(o_ofs[4]), .SMC(test_se), .C(net10783), .XR(n18), .Q(o_ofs[5]) );
  SDFFRQX1 adcnt_reg_1_ ( .D(N107), .SIN(o_ofs[0]), .SMC(test_se), .C(net10783), .XR(n18), .Q(o_ofs[1]) );
  SDFFRQX1 adcnt_reg_0_ ( .D(N106), .SIN(test_si), .SMC(test_se), .C(net10783), 
        .XR(n18), .Q(o_ofs[0]) );
  SDFFRQX1 adcnt_reg_2_ ( .D(N108), .SIN(o_ofs[1]), .SMC(test_se), .C(net10783), .XR(n18), .Q(o_ofs[2]) );
  SDFFRQX1 adcnt_reg_6_ ( .D(N112), .SIN(o_ofs[5]), .SMC(test_se), .C(net10783), .XR(n19), .Q(o_ofs[6]) );
  SDFFRQX1 adcnt_reg_3_ ( .D(N109), .SIN(o_ofs[2]), .SMC(test_se), .C(net10783), .XR(n18), .Q(o_ofs[3]) );
  SDFFRQX1 adcnt_reg_4_ ( .D(N110), .SIN(o_ofs[3]), .SMC(test_se), .C(net10783), .XR(n18), .Q(o_ofs[4]) );
  SDFFRQX1 cs_rwb_reg ( .D(n119), .SIN(o_dbgpo[3]), .SMC(test_se), .C(i_clk), 
        .XR(n18), .Q(cs_rwb) );
  SDFFSQX1 rwbuf_reg_6_ ( .D(N142), .SIN(o_wdat[5]), .SMC(test_se), .C(
        net10788), .XS(n17), .Q(o_wdat[6]) );
  SDFFSQX1 rwbuf_reg_3_ ( .D(N139), .SIN(o_wdat[2]), .SMC(test_se), .C(
        net10788), .XS(n17), .Q(o_wdat[3]) );
  SDFFSQX1 rwbuf_reg_4_ ( .D(N140), .SIN(o_wdat[3]), .SMC(test_se), .C(
        net10788), .XS(n17), .Q(o_wdat[4]) );
  SDFFSQX1 rwbuf_reg_7_ ( .D(N143), .SIN(o_wdat[6]), .SMC(test_se), .C(
        net10788), .XS(n16), .Q(o_wdat[7]) );
  SDFFSQX1 rwbuf_reg_1_ ( .D(N137), .SIN(o_wdat[0]), .SMC(test_se), .C(
        net10788), .XS(n18), .Q(o_wdat[1]) );
  SDFFSQX1 cs_bit_reg_3_ ( .D(N78), .SIN(o_dbgpo[2]), .SMC(test_se), .C(
        net10777), .XS(n17), .Q(o_dbgpo[3]) );
  SDFFSQX1 cs_bit_reg_2_ ( .D(N77), .SIN(o_dbgpo[1]), .SMC(test_se), .C(
        net10777), .XS(n17), .Q(o_dbgpo[2]) );
  SDFFSQX1 rwbuf_reg_0_ ( .D(N136), .SIN(o_lt_ofs[7]), .SMC(test_se), .C(
        net10788), .XS(n16), .Q(o_wdat[0]) );
  SDFFSQX1 rwbuf_reg_5_ ( .D(N141), .SIN(o_wdat[4]), .SMC(test_se), .C(
        net10788), .XS(n17), .Q(o_wdat[5]) );
  SDFFSQX1 rwbuf_reg_2_ ( .D(N138), .SIN(o_wdat[1]), .SMC(test_se), .C(
        net10788), .XS(n17), .Q(o_wdat[2]) );
  SDFFRQX1 cs_sta_reg_0_ ( .D(n120), .SIN(cs_rwb), .SMC(test_se), .C(i_clk), 
        .XR(n18), .Q(cs_sta[0]) );
  SDFFSQX1 cs_bit_reg_0_ ( .D(N75), .SIN(o_ofs[7]), .SMC(test_se), .C(net10777), .XS(n17), .Q(o_dbgpo[0]) );
  SDFFRQX1 adcnt_reg_7_ ( .D(N113), .SIN(o_ofs[6]), .SMC(test_se), .C(net10783), .XR(n18), .Q(o_ofs[7]) );
  SDFFRQX1 cs_sta_reg_1_ ( .D(n121), .SIN(cs_sta[0]), .SMC(test_se), .C(i_clk), 
        .XR(n19), .Q(cs_sta[1]) );
  SDFFSQX1 cs_bit_reg_1_ ( .D(N76), .SIN(o_dbgpo[0]), .SMC(test_se), .C(
        net10777), .XS(n17), .Q(o_dbgpo[1]) );
  MUX2X1 U3 ( .D0(n148), .D1(n147), .S(i_prefetch), .Y(o_r_early) );
  MUX2X1 U4 ( .D0(n150), .D1(n162), .S(i_prefetch), .Y(n152) );
  OR3XL U5 ( .A(o_dbgpo[1]), .B(n73), .C(n27), .Y(n165) );
  INVX1 U6 ( .A(o_dbgpo[7]), .Y(n178) );
  INVX1 U7 ( .A(o_dbgpo[3]), .Y(n135) );
  NAND21X1 U8 ( .B(o_dbgpo[3]), .A(n26), .Y(n164) );
  INVX1 U9 ( .A(n164), .Y(n149) );
  INVX1 U10 ( .A(n22), .Y(o_busev[1]) );
  INVX1 U11 ( .A(n69), .Y(n153) );
  INVX1 U12 ( .A(o_wdat[1]), .Y(n40) );
  INVX1 U13 ( .A(o_wdat[2]), .Y(n91) );
  INVX1 U14 ( .A(o_wdat[3]), .Y(n49) );
  INVX1 U15 ( .A(o_wdat[4]), .Y(n90) );
  INVX1 U16 ( .A(o_wdat[5]), .Y(n92) );
  INVX1 U17 ( .A(o_wdat[6]), .Y(n32) );
  INVX1 U18 ( .A(o_dbgpo[1]), .Y(n24) );
  NAND21X1 U19 ( .B(o_dbgpo[2]), .A(n135), .Y(n27) );
  INVX1 U20 ( .A(cs_rwb), .Y(n166) );
  INVX1 U21 ( .A(n129), .Y(o_we) );
  NAND5XL U22 ( .A(o_busev[1]), .B(n80), .C(n78), .D(n81), .E(n31), .Y(n34) );
  NAND32X1 U23 ( .B(cs_rwb), .C(n69), .A(n30), .Y(n129) );
  INVX1 U24 ( .A(n128), .Y(n30) );
  INVX1 U25 ( .A(cs_sta[0]), .Y(n122) );
  MUX2X1 U26 ( .D0(n149), .D1(n136), .S(cs_rwb), .Y(n137) );
  INVXL U27 ( .A(n35), .Y(n147) );
  INVX1 U28 ( .A(o_dbgpo[0]), .Y(n73) );
  XOR2X1 U29 ( .A(n49), .B(i_deva[4]), .Y(n81) );
  INVX1 U30 ( .A(o_wdat[7]), .Y(n93) );
  INVX1 U31 ( .A(ps_rwbuf_0_), .Y(n163) );
  NAND21XL U32 ( .B(n128), .A(n127), .Y(n138) );
  INVXL U33 ( .A(n142), .Y(o_dec) );
  INVXL U34 ( .A(n165), .Y(n162) );
  NAND31XL U35 ( .C(n166), .A(i_rd_mem), .B(n24), .Y(n28) );
  INVXL U36 ( .A(n77), .Y(n83) );
  XOR2X1 U37 ( .A(n32), .B(i_deva[7]), .Y(n80) );
  XOR2X1 U38 ( .A(n91), .B(i_deva[3]), .Y(n76) );
  XOR2X1 U39 ( .A(n33), .B(i_deva[1]), .Y(n75) );
  OR2XL U40 ( .A(o_dbgpo[2]), .B(n114), .Y(n14) );
  NAND21X1 U41 ( .B(cs_sta[1]), .A(n122), .Y(n102) );
  XOR2XL U42 ( .A(n93), .B(i_deva[7]), .Y(n94) );
  NAND43X1 U43 ( .B(n101), .C(n100), .D(n99), .A(n98), .Y(n144) );
  XOR2XL U44 ( .A(i_deva[6]), .B(o_wdat[6]), .Y(n100) );
  NAND31XL U45 ( .C(n135), .A(o_dbgpo[2]), .B(n12), .Y(n143) );
  NAND41XL U46 ( .D(cs_sta[0]), .A(cs_rwb), .B(n160), .C(n159), .Y(n161) );
  NAND31XL U47 ( .C(n53), .A(o_ofs[2]), .B(n52), .Y(n54) );
  INVXL U48 ( .A(o_ofs[1]), .Y(n43) );
  OAI21BBXL U49 ( .A(o_wdat[6]), .B(n127), .C(n1), .Y(N112) );
  MUX2IXL U50 ( .D0(n64), .D1(n65), .S(o_ofs[6]), .Y(n1) );
  INVXL U51 ( .A(o_ofs[0]), .Y(n44) );
  INVXL U52 ( .A(o_ofs[5]), .Y(n61) );
  OAI21BBXL U53 ( .A(o_wdat[4]), .B(n127), .C(n2), .Y(N110) );
  MUX2IX1 U54 ( .D0(n55), .D1(n56), .S(o_ofs[4]), .Y(n2) );
  OAI21BBXL U55 ( .A(o_wdat[2]), .B(n127), .C(n3), .Y(N108) );
  MUX2IXL U56 ( .D0(n46), .D1(n47), .S(o_ofs[2]), .Y(n3) );
  OAI21BBXL U57 ( .A(o_wdat[0]), .B(n127), .C(n4), .Y(N106) );
  MUX2IXL U58 ( .D0(n37), .D1(n38), .S(o_ofs[0]), .Y(n4) );
  INVX1 U59 ( .A(n138), .Y(o_busev[2]) );
  INVX1 U60 ( .A(n113), .Y(n21) );
  INVX1 U61 ( .A(n34), .Y(n130) );
  NAND21X1 U62 ( .B(n178), .A(n162), .Y(n128) );
  INVX1 U66 ( .A(n29), .Y(n133) );
  INVX1 U69 ( .A(n140), .Y(n106) );
  NAND21XL U70 ( .B(n178), .A(n141), .Y(n154) );
  NAND21X1 U71 ( .B(n149), .A(n13), .Y(n113) );
  AND2X1 U72 ( .A(n162), .B(n155), .Y(n156) );
  INVX1 U73 ( .A(n139), .Y(n13) );
  NAND21X1 U74 ( .B(n140), .A(n139), .Y(N74) );
  BUFX3 U75 ( .A(o_busev[3]), .Y(o_dbgpo[4]) );
  AND4X1 U76 ( .A(n75), .B(n79), .C(n77), .D(n76), .Y(n31) );
  AND3X1 U77 ( .A(n153), .B(n152), .C(n151), .Y(o_re) );
  INVX1 U78 ( .A(o_dbgpo[6]), .Y(n103) );
  INVX1 U79 ( .A(n102), .Y(n141) );
  NAND32X1 U80 ( .B(n165), .C(n103), .A(n141), .Y(n22) );
  AND3X1 U81 ( .A(n146), .B(o_dec), .C(n151), .Y(n148) );
  INVX1 U82 ( .A(n144), .Y(n146) );
  NAND21XL U83 ( .B(n164), .A(n141), .Y(n142) );
  INVX1 U84 ( .A(n14), .Y(n26) );
  NAND21X1 U85 ( .B(n163), .A(n130), .Y(n35) );
  INVX1 U86 ( .A(n145), .Y(n151) );
  NAND21X1 U87 ( .B(n166), .A(o_dbgpo[6]), .Y(n145) );
  AND2X1 U88 ( .A(n149), .B(n163), .Y(n150) );
  INVX1 U89 ( .A(n143), .Y(o_idle) );
  OAI31XL U90 ( .A(n28), .B(n171), .C(n27), .D(n176), .Y(n132) );
  NAND32XL U91 ( .B(n103), .C(n132), .A(n164), .Y(n29) );
  INVX1 U92 ( .A(i_rd_mem), .Y(n179) );
  NAND21X1 U93 ( .B(n175), .A(n174), .Y(n118) );
  NOR32XL U94 ( .B(n158), .C(n157), .A(n156), .Y(n175) );
  MUX2IXL U95 ( .D0(n173), .D1(n172), .S(o_dbgpo[7]), .Y(n174) );
  INVX1 U96 ( .A(n154), .Y(n158) );
  INVX1 U97 ( .A(i_rdat[7]), .Y(n177) );
  OAI22AX1 U98 ( .D(n132), .C(n177), .A(n32), .B(n29), .Y(N143) );
  INVX1 U99 ( .A(n85), .Y(n173) );
  EORX1 U100 ( .A(i_fwnak), .B(n86), .C(n87), .D(i_fwack), .Y(n85) );
  NAND2X1 U101 ( .A(i_fwack), .B(n87), .Y(n86) );
  OA21X1 U102 ( .B(n133), .C(n132), .A(n131), .Y(N144) );
  INVX1 U103 ( .A(n23), .Y(o_busev[0]) );
  INVX1 U104 ( .A(n62), .Y(o_busev[3]) );
  NAND21X1 U105 ( .B(o_busev[0]), .A(n62), .Y(n140) );
  NOR21XL U106 ( .B(n111), .A(n110), .Y(n125) );
  AND2X1 U107 ( .A(n154), .B(n106), .Y(n111) );
  NOR21XL U108 ( .B(n149), .A(n109), .Y(n110) );
  NOR21XL U109 ( .B(n108), .A(n107), .Y(n109) );
  AO21XL U110 ( .B(n153), .C(n54), .A(n141), .Y(n56) );
  AO21XL U111 ( .B(n153), .C(n63), .A(n141), .Y(n65) );
  NAND21XL U112 ( .B(i_prefetch), .A(n144), .Y(n155) );
  INVX1 U113 ( .A(n68), .Y(n127) );
  INVX1 U114 ( .A(n54), .Y(n60) );
  INVX1 U115 ( .A(n45), .Y(n52) );
  OR4XL U116 ( .A(o_dbgpo[7]), .B(n103), .C(n102), .D(n155), .Y(n108) );
  INVX1 U117 ( .A(n75), .Y(n88) );
  INVX1 U118 ( .A(n76), .Y(n84) );
  NAND32XL U119 ( .B(n178), .C(n171), .A(n143), .Y(n139) );
  AO21XL U120 ( .B(n153), .C(n36), .A(n141), .Y(n38) );
  INVX1 U121 ( .A(i_inc), .Y(n36) );
  AO21XL U122 ( .B(n153), .C(n45), .A(n141), .Y(n47) );
  AO21X1 U123 ( .B(n21), .C(n73), .A(n140), .Y(N75) );
  NAND21XL U124 ( .B(n130), .A(n129), .Y(N179) );
  OR2X1 U125 ( .A(n116), .B(n5), .Y(N76) );
  AOI21X1 U126 ( .B(n115), .C(n114), .A(n113), .Y(n5) );
  OAI22XL U127 ( .A(n166), .B(n165), .C(n164), .D(n163), .Y(n167) );
  INVX1 U128 ( .A(n131), .Y(n171) );
  OAI22XL U129 ( .A(n129), .B(n40), .C(n34), .D(n33), .Y(N181) );
  OAI22XL U130 ( .A(n129), .B(n91), .C(n34), .D(n40), .Y(N182) );
  OAI22XL U131 ( .A(n129), .B(n49), .C(n34), .D(n91), .Y(N183) );
  OAI22XL U132 ( .A(n129), .B(n90), .C(n34), .D(n49), .Y(N184) );
  OAI22XL U133 ( .A(n129), .B(n92), .C(n34), .D(n90), .Y(N185) );
  OAI22XL U134 ( .A(n129), .B(n32), .C(n34), .D(n92), .Y(N186) );
  OAI22XL U135 ( .A(n93), .B(n129), .C(n34), .D(n32), .Y(N187) );
  INVX1 U136 ( .A(n63), .Y(n66) );
  INVX1 U137 ( .A(n15), .Y(n116) );
  NAND21X1 U138 ( .B(n62), .A(n23), .Y(n15) );
  XOR2XL U139 ( .A(i_deva[3]), .B(o_wdat[3]), .Y(n101) );
  AND4X1 U140 ( .A(n97), .B(n96), .C(n95), .D(n94), .Y(n98) );
  NAND21X1 U141 ( .B(o_dbgpo[0]), .A(n24), .Y(n114) );
  XOR2X1 U142 ( .A(n92), .B(i_deva[6]), .Y(n77) );
  XOR2X1 U143 ( .A(n90), .B(i_deva[5]), .Y(n78) );
  XOR2X1 U144 ( .A(n40), .B(i_deva[2]), .Y(n79) );
  XOR2XL U145 ( .A(n92), .B(i_deva[5]), .Y(n95) );
  XOR2XL U146 ( .A(n91), .B(i_deva[2]), .Y(n96) );
  XOR2XL U147 ( .A(i_deva[1]), .B(o_wdat[1]), .Y(n99) );
  INVX1 U148 ( .A(o_wdat[0]), .Y(n33) );
  XOR2XL U149 ( .A(n90), .B(i_deva[4]), .Y(n97) );
  NAND21XL U150 ( .B(cs_sta[0]), .A(cs_sta[1]), .Y(n69) );
  INVX1 U151 ( .A(n115), .Y(n12) );
  NAND21XL U152 ( .B(n73), .A(o_dbgpo[1]), .Y(n115) );
  MUX2BXL U153 ( .D0(n177), .D1(o_sda), .S(n176), .Y(n87) );
  NAND6XL U154 ( .A(o_dbgpo[3]), .B(cs_rwb), .C(n26), .D(n131), .E(i_rd_mem), 
        .F(n25), .Y(n176) );
  AO22XL U155 ( .A(n133), .B(o_wdat[2]), .C(i_rdat[3]), .D(n132), .Y(N139) );
  AO22XL U156 ( .A(n133), .B(o_wdat[0]), .C(i_rdat[1]), .D(n132), .Y(N137) );
  AO22XL U157 ( .A(n133), .B(o_wdat[3]), .C(i_rdat[4]), .D(n132), .Y(N140) );
  AO22XL U158 ( .A(n133), .B(o_wdat[5]), .C(i_rdat[6]), .D(n132), .Y(N142) );
  AO22XL U159 ( .A(n133), .B(o_wdat[1]), .C(i_rdat[2]), .D(n132), .Y(N138) );
  AO22XL U160 ( .A(n133), .B(o_wdat[4]), .C(i_rdat[5]), .D(n132), .Y(N141) );
  NAND21XL U161 ( .B(i_rd_mem), .A(o_wdat[7]), .Y(n159) );
  NAND21X1 U162 ( .B(n179), .A(i_rdat[7]), .Y(n160) );
  NAND31X1 U163 ( .C(n171), .A(n170), .B(n169), .Y(n172) );
  NAND21X1 U164 ( .B(n168), .A(n167), .Y(n169) );
  NAND21XL U165 ( .B(n162), .A(n161), .Y(n170) );
  INVXL U166 ( .A(cs_sta[1]), .Y(n168) );
  OAI21BBX1 U167 ( .A(i_rdat[0]), .B(n132), .C(n6), .Y(N136) );
  NAND4XL U168 ( .A(o_dbgpo[6]), .B(ps_rwbuf_0_), .C(n164), .D(n166), .Y(n6)
         );
  NAND32XL U169 ( .B(n25), .C(o_dbgpo[7]), .A(sdafall), .Y(n23) );
  NAND3XL U170 ( .A(i2c_scl), .B(n178), .C(o_dbgpo[5]), .Y(n62) );
  AO21X1 U171 ( .B(n104), .C(n108), .A(n140), .Y(n117) );
  NAND5XL U172 ( .A(i_prefetch), .B(o_dbgpo[1]), .C(n135), .D(n134), .E(n89), 
        .Y(n104) );
  NAND43X1 U173 ( .B(n88), .C(n84), .D(n83), .A(n82), .Y(n89) );
  AND4XL U174 ( .A(n81), .B(n80), .C(n79), .D(n78), .Y(n82) );
  NAND21XL U175 ( .B(cs_sta[1]), .A(cs_sta[0]), .Y(n68) );
  NAND21XL U176 ( .B(n122), .A(cs_sta[1]), .Y(n131) );
  NAND32X1 U177 ( .B(n44), .C(n43), .A(i_inc), .Y(n45) );
  NAND31X1 U178 ( .C(n61), .A(o_ofs[4]), .B(n60), .Y(n63) );
  MUX2XL U179 ( .D0(n126), .D1(cs_sta[1]), .S(n125), .Y(n121) );
  NAND21X1 U180 ( .B(n124), .A(n123), .Y(n126) );
  AO21XL U181 ( .B(n157), .C(n122), .A(n140), .Y(n123) );
  INVX1 U182 ( .A(n117), .Y(n124) );
  AND2XL U183 ( .A(n60), .B(n153), .Y(n55) );
  AND2XL U184 ( .A(n66), .B(n153), .Y(n64) );
  MUX2XL U185 ( .D0(n112), .D1(cs_sta[0]), .S(n125), .Y(n120) );
  NAND21X1 U186 ( .B(n105), .A(n117), .Y(n112) );
  AND4XL U187 ( .A(n106), .B(n149), .C(n122), .D(n166), .Y(n105) );
  INVXL U188 ( .A(i2c_scl), .Y(n25) );
  INVX1 U189 ( .A(o_ofs[3]), .Y(n53) );
  NOR21XL U190 ( .B(o_dbgpo[7]), .A(cs_sta[1]), .Y(n107) );
  GEN2XL U191 ( .D(o_dbgpo[3]), .E(n14), .C(n149), .B(n13), .A(n140), .Y(N78)
         );
  GEN2XL U192 ( .D(o_dbgpo[2]), .E(n114), .C(n26), .B(n21), .A(n116), .Y(N77)
         );
  MUX2BXL U193 ( .D0(ps_rwbuf_0_), .D1(n7), .S(n8), .Y(n119) );
  NAND2XL U194 ( .A(cs_rwb), .B(n23), .Y(n7) );
  NAND2XL U195 ( .A(o_busev[1]), .B(n23), .Y(n8) );
  MUX2BXL U196 ( .D0(n162), .D1(n9), .S(i_prefetch), .Y(n136) );
  NAND3XL U197 ( .A(o_dbgpo[1]), .B(n135), .C(n134), .Y(n9) );
  NAND21XL U198 ( .B(n164), .A(cs_rwb), .Y(n157) );
  AO21XL U199 ( .B(o_wdat[0]), .C(o_we), .A(n147), .Y(N180) );
  AND2XL U200 ( .A(n52), .B(n153), .Y(n46) );
  AND2XL U201 ( .A(i_inc), .B(n153), .Y(n37) );
  NAND3X1 U202 ( .A(n154), .B(n10), .C(n138), .Y(N114) );
  NAND3XL U203 ( .A(n153), .B(o_dbgpo[7]), .C(n137), .Y(n10) );
  OAI222XL U204 ( .A(n72), .B(n71), .C(n70), .D(n69), .E(n93), .F(n68), .Y(
        N113) );
  MUX2BXL U205 ( .D0(n71), .D1(n67), .S(o_ofs[6]), .Y(n70) );
  INVX1 U206 ( .A(n65), .Y(n72) );
  AND2X1 U207 ( .A(n66), .B(n71), .Y(n67) );
  OAI222XL U208 ( .A(n42), .B(n43), .C(n41), .D(n69), .E(n68), .F(n40), .Y(
        N107) );
  MUX2BXL U209 ( .D0(n43), .D1(n39), .S(o_ofs[0]), .Y(n41) );
  INVX1 U210 ( .A(n38), .Y(n42) );
  AND2X1 U211 ( .A(i_inc), .B(n43), .Y(n39) );
  OAI222XL U212 ( .A(n59), .B(n61), .C(n58), .D(n69), .E(n68), .F(n92), .Y(
        N111) );
  MUX2BXL U213 ( .D0(n61), .D1(n57), .S(o_ofs[4]), .Y(n58) );
  INVX1 U214 ( .A(n56), .Y(n59) );
  AND2X1 U215 ( .A(n60), .B(n61), .Y(n57) );
  OAI222XL U216 ( .A(n51), .B(n53), .C(n50), .D(n69), .E(n68), .F(n49), .Y(
        N109) );
  MUX2BXL U217 ( .D0(n53), .D1(n48), .S(o_ofs[2]), .Y(n50) );
  INVX1 U218 ( .A(n47), .Y(n51) );
  AND2X1 U219 ( .A(n52), .B(n53), .Y(n48) );
  INVXL U220 ( .A(o_ofs[7]), .Y(n71) );
  INVX1 U221 ( .A(n74), .Y(n134) );
  NAND21XL U222 ( .B(o_dbgpo[2]), .A(n73), .Y(n74) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2cdbnc_a0_0 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall, test_si, 
        test_se );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c, test_si, test_se;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n9, n1, n2, n3, n4, n5;

  SDFFSQX1 d_i2c_reg_2_ ( .D(N19), .SIN(N19), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(d_i2c_2_) );
  SDFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .SIN(test_si), .SMC(test_se), .C(i_clk), 
        .XS(i_rstz), .Q(N18) );
  SDFFSQX1 d_i2c_reg_1_ ( .D(N18), .SIN(N18), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(N19) );
  SDFFSQXX1 r_i2c_reg ( .D(n9), .SIN(d_i2c_2_), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(o_i2c), .XQ() );
  NOR21XL U3 ( .B(o_i2c), .A(n5), .Y(fall) );
  NOR42XL U4 ( .C(N19), .D(N18), .A(o_i2c), .B(n4), .Y(rise) );
  NOR2X1 U5 ( .A(r_opt[0]), .B(d_i2c_2_), .Y(n4) );
  OAI211X1 U6 ( .C(r_opt[1]), .D(n3), .A(n2), .B(n1), .Y(n5) );
  INVX1 U7 ( .A(N18), .Y(n2) );
  INVX1 U8 ( .A(N19), .Y(n1) );
  INVX1 U9 ( .A(d_i2c_2_), .Y(n3) );
  AO21XL U10 ( .B(o_i2c), .C(n5), .A(rise), .Y(n9) );
endmodule


module i2cdbnc_a0_1 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall, test_si, 
        test_se );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c, test_si, test_se;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n6, n1, n2, n3;

  SDFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .SIN(test_si), .SMC(test_se), .C(i_clk), 
        .XS(i_rstz), .Q(N18) );
  SDFFSQX1 d_i2c_reg_1_ ( .D(N18), .SIN(N18), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(N19) );
  SDFFSQXX1 r_i2c_reg ( .D(n6), .SIN(d_i2c_2_), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(o_i2c), .XQ() );
  SDFFSQX1 d_i2c_reg_2_ ( .D(N19), .SIN(N19), .SMC(test_se), .C(i_clk), .XS(
        i_rstz), .Q(d_i2c_2_) );
  NOR42XL U3 ( .C(N19), .D(N18), .A(o_i2c), .B(n2), .Y(rise) );
  INVX1 U4 ( .A(n3), .Y(fall) );
  NOR2XL U5 ( .A(d_i2c_2_), .B(r_opt[0]), .Y(n2) );
  NAND42XL U6 ( .C(N18), .D(N19), .A(n1), .B(o_i2c), .Y(n3) );
  NAND21XL U7 ( .B(r_opt[1]), .A(d_i2c_2_), .Y(n1) );
  AO21XL U8 ( .B(o_i2c), .C(n3), .A(rise), .Y(n6) );
endmodule


module regbank_a0 ( srci, lg_pulse_len, dm_fault, cc1_di, cc2_di, di_rd_det, 
        i_tmrf, i_vcbyval, dnchk_en, r_pwrv_upd, aswkup, lg_dischg, gating_pwr, 
        ps_pwrdn, r_sleep, r_pwrdn, r_ocdrv_enz, r_osc_stop, r_osc_lo, 
        r_osc_gate, r_fw_pwrv, r_cvcwr, r_cvofs, r_otpi_gate, r_pwrctl, 
        r_pwr_i, r_cvctl, r_srcctl, r_dpdmctl, r_ccrx, r_cctrx, r_ccctl, 
        r_fcpwr, r_fcpre, fcp_r_dat, fcp_r_sta, fcp_r_msk, fcp_r_ctl, 
        fcp_r_crc, fcp_r_acc, fcp_r_tui, r_accctl, r_bclk_sel, r_dacwr, 
        r_dac_en, r_sar_en, r_adofs, r_isofs, x_daclsb, r_comp_opt, dac_r_ctl, 
        dac_r_comp, dac_r_cmpsta, dac_r_vs, REVID, atpg_en, sfr_r, sfr_w, 
        set_hold, bkpt_hold, cpurst, sfr_addr, sfr_wdat, sfr_rdat, ff_p0, 
        di_p0, ictlr_idle, ictlr_inc, r_inst_ofs, r_psrd, r_pswr, r_fortxdat, 
        r_fortxrdy, r_fortxen, r_ana_tm, r_gpio_tm, r_gpio_ie, r_gpio_oe, 
        r_gpio_pu, r_gpio_pd, r_gpio_s0, r_gpio_s1, r_gpio_s2, r_gpio_s3, 
        r_regtrm, i_pc, i_goidle, i_gobusy, i_i2c_idle, bus_idle, i2c_stretch, 
        i_i2c_rwbuf, i_i2c_ltbuf, i_i2c_ofs, o_intr, r_auto_gdcrc, r_exist1st, 
        r_ordrs4, r_fifopsh, r_fifopop, r_unlock, r_first, r_last, r_fiforst, 
        r_set_cpmsgid, r_txendk, r_txnumk, r_txshrt, r_auto_discard, 
        r_hold_mcu, r_txauto, r_rxords_ena, r_spec, r_dat_spec, r_dat_portrole, 
        r_dat_datarole, r_discard, r_pshords, r_pg0_sel, r_strtch, r_i2c_attr, 
        r_i2c_ninc, r_hwi2c_en, r_i2c_fwnak, r_i2c_fwack, r_i2c_deva, i2c_ev, 
        prl_c0set, prl_cany0, prl_discard, prl_GCTxDone, prl_cpmsgid, pff_ack, 
        prx_rst, pff_obsd, pff_full, pff_empty, ptx_ack, pff_ptr, prx_adpn, 
        pff_rdat, pff_rxpart, prx_rcvinf, ptx_fsm, prx_fsm, prl_fsm, 
        prx_setsta, clk_1p0m, clk_500, clk, xrstz, xclk, dbgpo, srstz, prstz, 
        test_si2, test_si1, test_so2, test_so1, test_se );
  input [5:0] srci;
  input [1:0] lg_pulse_len;
  output [11:0] r_fw_pwrv;
  output [1:0] r_cvcwr;
  input [15:0] r_cvofs;
  output [7:4] r_pwrctl;
  output [7:0] r_pwr_i;
  output [7:0] r_cvctl;
  output [7:0] r_srcctl;
  output [7:0] r_dpdmctl;
  output [7:0] r_ccrx;
  output [7:0] r_cctrx;
  output [7:0] r_ccctl;
  output [6:0] r_fcpwr;
  input [7:0] fcp_r_dat;
  input [7:0] fcp_r_sta;
  input [7:0] fcp_r_msk;
  input [7:0] fcp_r_ctl;
  input [7:0] fcp_r_crc;
  input [7:0] fcp_r_acc;
  input [7:0] fcp_r_tui;
  input [7:0] r_accctl;
  output [14:0] r_dacwr;
  input [7:0] r_dac_en;
  input [7:0] r_sar_en;
  input [7:0] r_adofs;
  input [7:0] r_isofs;
  input [5:0] x_daclsb;
  output [7:0] r_comp_opt;
  input [7:0] dac_r_ctl;
  input [7:0] dac_r_comp;
  input [7:0] dac_r_cmpsta;
  input [63:0] dac_r_vs;
  input [6:0] REVID;
  input [7:0] sfr_addr;
  input [7:0] sfr_wdat;
  output [7:0] sfr_rdat;
  input [7:0] ff_p0;
  input [7:0] di_p0;
  output [14:0] r_inst_ofs;
  output [3:0] r_ana_tm;
  output [1:0] r_gpio_ie;
  output [6:0] r_gpio_oe;
  output [6:0] r_gpio_pu;
  output [6:0] r_gpio_pd;
  output [2:0] r_gpio_s0;
  output [2:0] r_gpio_s1;
  output [2:0] r_gpio_s2;
  output [2:0] r_gpio_s3;
  output [55:0] r_regtrm;
  input [15:0] i_pc;
  input [7:0] i_i2c_rwbuf;
  input [7:0] i_i2c_ltbuf;
  input [7:0] i_i2c_ofs;
  output [4:0] o_intr;
  output [1:0] r_auto_gdcrc;
  output [4:0] r_txnumk;
  output [6:0] r_txauto;
  output [6:0] r_rxords_ena;
  output [1:0] r_spec;
  output [1:0] r_dat_spec;
  output [3:0] r_pg0_sel;
  output [7:1] r_i2c_deva;
  input [7:0] i2c_ev;
  input [2:0] prl_cpmsgid;
  input [1:0] pff_ack;
  input [1:0] prx_rst;
  input [5:0] pff_ptr;
  input [5:0] prx_adpn;
  input [7:0] pff_rdat;
  input [15:0] pff_rxpart;
  input [4:0] prx_rcvinf;
  input [2:0] ptx_fsm;
  input [3:0] prx_fsm;
  input [3:0] prl_fsm;
  input [6:0] prx_setsta;
  output [31:0] dbgpo;
  input dm_fault, cc1_di, cc2_di, di_rd_det, i_tmrf, i_vcbyval, dnchk_en,
         atpg_en, sfr_r, sfr_w, set_hold, bkpt_hold, cpurst, ictlr_idle,
         ictlr_inc, i_goidle, i_gobusy, i_i2c_idle, prl_c0set, prl_cany0,
         prl_discard, prl_GCTxDone, pff_obsd, pff_full, pff_empty, ptx_ack,
         clk_1p0m, clk_500, clk, xrstz, xclk, test_si2, test_si1, test_se;
  output r_pwrv_upd, aswkup, lg_dischg, gating_pwr, ps_pwrdn, r_sleep, r_pwrdn,
         r_ocdrv_enz, r_osc_stop, r_osc_lo, r_osc_gate, r_otpi_gate, r_fcpre,
         r_bclk_sel, r_psrd, r_pswr, r_fortxdat, r_fortxrdy, r_fortxen,
         r_gpio_tm, bus_idle, i2c_stretch, r_exist1st, r_ordrs4, r_fifopsh,
         r_fifopop, r_unlock, r_first, r_last, r_fiforst, r_set_cpmsgid,
         r_txendk, r_txshrt, r_auto_discard, r_hold_mcu, r_dat_portrole,
         r_dat_datarole, r_discard, r_pshords, r_strtch, r_i2c_attr,
         r_i2c_ninc, r_hwi2c_en, r_i2c_fwnak, r_i2c_fwack, srstz, prstz,
         test_so2, test_so1;
  wire   we_246, we_245, we_232, we_231, we_230, we_228, we_222, we_217,
         we_215, we_214, we_213, we_211, we_209, we_203, we_191, we_187,
         we_182, we_181, we_176, we_175, we_172, we_171, we_148, we_143,
         regF4_7_, regF4_3, regE3_0, regD4_6_, regD4_5_, regD4_4_, regD4_3_,
         regD4_2_, regD4_1_, regD4_0_, regD3_7_, regD3_3, reg25_0_, reg19_7_,
         reg12_1, reg11_7_, reg11_4, regAD_7, N26, N27, N28, N29, N30, N32,
         N33, N34, N35, N36, N37, N38, N39, upd01, phyrst, upd12, upd18, upd19,
         upd20, upd21, lt_reg26_0, i2c_mode_upd, i2c_mode_wdat, upd31, N84,
         as_p0_chg, dmf_wkup, p0_chg_clr, di_rd_det_clr, dm_fault_clr,
         pwrdn_rstz, osc_low_clr, osc_low_rstz, r_pos_gate, osc_gate_n_2_,
         osc_gate_n_1_, osc_gate_n_0_, m_ovp, m_ovp_sta, setAE_7, m_scp,
         m_scp_sta, s_ovp, s_ovp_sta, s_scp, s_scp_sta, lg_pulse_12m, N108,
         N109, N110, N111, N112, N113, net10815, net10821, n1218, n1219, n1220,
         n1221, n20, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n75, n83, n86, n99, n100, n102,
         n103, n104, n106, n109, n114, n116, n117, n118, n119, n121, n122,
         n123, n124, n126, n127, n128, n129, n133, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n173, n174, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n1, n2, n3, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n21, n22, n23, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n76, n77,
         n78, n79, n80, n81, n82, n84, n85, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n101, n105, n107, n108, n110, n111, n112,
         n113, n115, n120, n125, n130, n131, n132, n134, n135, n159, n160,
         n172, n175, n176, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462,
         SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464,
         SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466,
         SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468,
         SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470,
         SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472,
         SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474,
         SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476,
         SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478,
         SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480,
         SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482,
         SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484,
         SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486,
         SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488,
         SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490,
         SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492,
         SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494,
         SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496,
         SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498,
         SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500,
         SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502,
         SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504,
         SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506,
         SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508,
         SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510,
         SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512,
         SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514,
         SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516,
         SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518,
         SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520,
         SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522,
         SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524,
         SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526,
         SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528,
         SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530,
         SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532,
         SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534,
         SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536,
         SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538,
         SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540,
         SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542,
         SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544,
         SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546,
         SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548,
         SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550,
         SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552,
         SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554,
         SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556,
         SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558,
         SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560,
         SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562,
         SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564,
         SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566,
         SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568,
         SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570,
         SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572,
         SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574,
         SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576,
         SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578,
         SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580,
         SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582,
         SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584,
         SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586,
         SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588,
         SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590,
         SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592,
         SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594,
         SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596,
         SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598,
         SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600,
         SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602,
         SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604,
         SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606,
         SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608,
         SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610,
         SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612,
         SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614,
         SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616,
         SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618,
         SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620,
         SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622,
         SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624,
         SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626,
         SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628,
         SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630,
         SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632,
         SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634,
         SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636,
         SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638,
         SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640,
         SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642,
         SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644,
         SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646,
         SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648,
         SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650,
         SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652,
         SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654,
         SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656,
         SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658,
         SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660,
         SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662,
         SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664,
         SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666,
         SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668,
         SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670,
         SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672,
         SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674,
         SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676,
         SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678,
         SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680,
         SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682,
         SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684,
         SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686,
         SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688,
         SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690,
         SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692,
         SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694,
         SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696,
         SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698,
         SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700,
         SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702,
         SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704,
         SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706,
         SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708,
         SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710,
         SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712,
         SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714,
         SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716,
         SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718,
         SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720,
         SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722,
         SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724,
         SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726,
         SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728,
         SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730,
         SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732,
         SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734,
         SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736,
         SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738,
         SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740,
         SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742,
         SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744,
         SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746,
         SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748,
         SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750,
         SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752,
         SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754,
         SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756,
         SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758,
         SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760,
         SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762,
         SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764,
         SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766,
         SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768,
         SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770,
         SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772,
         SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774,
         SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776,
         SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778,
         SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780,
         SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782,
         SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784,
         SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786,
         SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788,
         SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790,
         SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792,
         SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794,
         SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796,
         SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798,
         SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800,
         SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802,
         SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804,
         SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806,
         SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808,
         SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810,
         SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812,
         SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814,
         SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816,
         SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818,
         SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820,
         SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822,
         SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824,
         SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826,
         SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828,
         SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830,
         SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832,
         SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834,
         SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836,
         SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838,
         SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840,
         SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842,
         SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844,
         SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846,
         SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848,
         SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850,
         SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852,
         SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854,
         SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856,
         SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858,
         SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860,
         SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862,
         SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864,
         SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866,
         SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868,
         SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870,
         SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872,
         SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874,
         SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876,
         SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878,
         SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880,
         SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882,
         SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884,
         SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886,
         SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888,
         SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890,
         SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892,
         SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894,
         SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896,
         SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898,
         SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900,
         SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902,
         SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904,
         SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906,
         SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908,
         SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910,
         SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912,
         SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914,
         SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916,
         SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918,
         SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920,
         SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922,
         SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924,
         SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926,
         SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928,
         SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930,
         SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932,
         SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934,
         SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936,
         SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938,
         SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940,
         SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942,
         SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944,
         SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946,
         SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948,
         SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950,
         SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952,
         SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954,
         SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956,
         SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958,
         SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960,
         SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962,
         SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964,
         SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966,
         SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968,
         SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970,
         SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972,
         SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974,
         SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976,
         SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978,
         SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980,
         SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982,
         SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984,
         SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986,
         SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988,
         SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990,
         SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992,
         SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994,
         SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996,
         SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998,
         SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000,
         SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002,
         SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004,
         SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006,
         SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008,
         SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010,
         SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012,
         SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014,
         SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016,
         SYNOPSYS_UNCONNECTED_1017;
  wire   [167:161] we;
  wire   [3:2] regE3;
  wire   [7:0] regDF;
  wire   [7:0] regDE;
  wire   [7:0] reg31;
  wire   [7:0] reg30;
  wire   [7:0] reg28;
  wire   [7:0] reg27;
  wire   [7:1] reg21;
  wire   [4:0] reg20;
  wire   [7:3] reg12;
  wire   [7:0] reg06;
  wire   [7:0] reg05;
  wire   [7:0] regAF;
  wire   [7:0] regAE;
  wire   [5:0] regAD;
  wire   [7:0] regAC;
  wire   [7:0] regAB;
  wire   [7:0] reg94;
  wire   [7:0] irqAE;
  wire   [7:0] irqDF;
  wire   [7:0] irq28;
  wire   [7:0] irq04;
  wire   [7:0] irq03;
  wire   [1:0] drstz;
  wire   [4:0] rstcnt;
  wire   [1:0] r_phyrst;
  wire   [7:0] wd01;
  wire   [7:0] clr03;
  wire   [7:0] set03;
  wire   [7:0] clr04;
  wire   [7:0] set04;
  wire   [7:0] wd12;
  wire   [14:0] inst_ofs_plus;
  wire   [7:0] wd18;
  wire   [7:0] wd19;
  wire   [7:0] wd20;
  wire   [7:0] wd21;
  wire   [7:0] clr28;
  wire   [2:0] oscdwn_shft;
  wire   [7:0] d_p0;
  wire   [7:0] setDF;
  wire   [7:0] clrDF;
  wire   [7:0] clrAE;
  wire   [5:0] setAE;
  wire   [4:0] lg_pulse_cnt;
  wire   [3:0] lt_regE4_3_0;
  wire   [4:2] add_180_carry;

  AND2X1 U0_MASK_0 ( .A(oscdwn_shft[2]), .B(as_p0_chg), .Y(p0_chg_clr) );
  AND2X1 U0_MASK_2 ( .A(regD4_6_), .B(di_rd_det), .Y(di_rd_det_clr) );
  AND2X1 U0_MASK_3 ( .A(test_so2), .B(dmf_wkup), .Y(dm_fault_clr) );
  AND2X1 U0_MASK_4 ( .A(regD4_5_), .B(aswkup), .Y(osc_low_clr) );
  HAD1X1 add_180_U1_1_1 ( .A(N29), .B(N30), .CO(add_180_carry[2]), .SO(N32) );
  HAD1X1 add_180_U1_1_2 ( .A(N28), .B(add_180_carry[2]), .CO(add_180_carry[3]), 
        .SO(N33) );
  HAD1X1 add_180_U1_1_3 ( .A(N27), .B(add_180_carry[3]), .CO(add_180_carry[4]), 
        .SO(N34) );
  glreg_a0_79 u0_reg00 ( .clk(clk), .arstz(n40), .we(we_176), .wdat({n254, 
        n248, n238, n232, n220, n213, n207, n159}), .rdat({r_txendk, r_txauto}), .test_si(n279), .test_se(test_se) );
  glreg_a0_78 u0_reg01 ( .clk(clk), .arstz(n48), .we(upd01), .wdat(wd01), 
        .rdat({r_last, r_first, r_unlock, r_txnumk}), .test_si(r_txendk), 
        .test_se(test_se) );
  glsta_a0_6 u0_reg03 ( .clk(clk), .arstz(n41), .rst0(phyrst), .set2({
        set03[7:4], n75, set03[2:0]}), .clr1(clr03), .rdat(dbgpo[7:0]), .irq(
        irq03), .test_si(r_last), .test_se(test_se) );
  glsta_a0_5 u0_reg04 ( .clk(clk), .arstz(n42), .rst0(n21), .set2(set04), 
        .clr1(clr04), .rdat(dbgpo[15:8]), .irq(irq04), .test_si(dbgpo[7]), 
        .test_se(test_se) );
  glreg_a0_77 u0_reg05 ( .clk(clk), .arstz(n51), .we(we_181), .wdat({n255, 
        n248, n238, n232, n220, n213, n207, n135}), .rdat(reg05), .test_si(
        dbgpo[15]), .test_se(test_se) );
  glreg_a0_76 u0_reg06 ( .clk(clk), .arstz(n52), .we(we_182), .wdat({n255, 
        n248, n241, n232, n220, n214, n207, n159}), .rdat(reg06), .test_si(
        reg05[7]), .test_se(test_se) );
  glreg_a0_75 u0_reg11 ( .clk(clk), .arstz(n53), .we(we_187), .wdat({n255, 
        n249, sfr_wdat[5], n232, n220, n213, n208, n159}), .rdat({reg11_7_, 
        r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0]}), .test_si(r_dpdmctl[7]), .test_se(test_se) );
  glreg_a0_74 u0_reg12 ( .clk(clk), .arstz(n54), .we(upd12), .wdat(wd12), 
        .rdat({reg12, r_txshrt, reg12_1, r_pshords}), .test_si(reg11_7_), 
        .test_se(test_se) );
  glreg_WIDTH5_2 u0_reg14 ( .clk(clk), .arstz(n84), .we(r_set_cpmsgid), .wdat(
        {n256, n249, n238, n232, n221}), .rdat({r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1]}), .test_si(reg12[7]), 
        .test_se(test_se) );
  glreg_a0_73 u0_reg15 ( .clk(clk), .arstz(n56), .we(we_191), .wdat({n255, 
        n250, n239, n233, n220, n214, n208, n159}), .rdat(dbgpo[31:24]), 
        .test_si(r_auto_gdcrc[0]), .test_se(test_se) );
  glreg_a0_72 u0_reg18 ( .clk(clk), .arstz(n57), .we(upd18), .wdat(wd18), 
        .rdat(r_inst_ofs[7:0]), .test_si(dbgpo[31]), .test_se(test_se) );
  glreg_a0_71 u0_reg19 ( .clk(clk), .arstz(n59), .we(upd19), .wdat(wd19), 
        .rdat({reg19_7_, r_inst_ofs[14:8]}), .test_si(r_inst_ofs[7]), 
        .test_se(test_se) );
  glreg_a0_70 u0_reg20 ( .clk(clk), .arstz(n67), .we(upd20), .wdat(wd20), 
        .rdat({r_dat_spec, r_dat_datarole, reg20}), .test_si(n16), .test_se(
        test_se) );
  glreg_a0_69 u0_reg21 ( .clk(clk), .arstz(n74), .we(upd21), .wdat(wd21), 
        .rdat({reg21, r_dat_portrole}), .test_si(r_dat_spec[1]), .test_se(
        test_se) );
  glreg_6_00000018 u0_reg25 ( .clk(clk), .arstz(n79), .we(n205), .wdat({n238, 
        n231, n219, n215, n208, n160}), .rdat({r_i2c_attr, r_pg0_sel, reg25_0_}), .test_si(reg21[7]), .test_se(test_se) );
  glreg_1_1_1 u0_reg26 ( .clk(clk), .arstz(n92), .we(n204), .wdat(n135), 
        .rdat(lt_reg26_0), .test_si(r_i2c_attr), .test_se(test_se) );
  glreg_1_1_0 u1_reg26 ( .clk(clk), .arstz(n92), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat(r_hwi2c_en), .test_si(n274), .test_se(test_se)
         );
  glreg_7_70 u2_reg26 ( .clk(clk), .arstz(n76), .we(n204), .wdat({n254, n248, 
        sfr_wdat[5], n232, n220, n214, n208}), .rdat(r_i2c_deva), .test_si(
        n271), .test_se(test_se) );
  glreg_a0_68 u0_reg27 ( .clk(clk), .arstz(n73), .we(we_203), .wdat({n255, 
        n249, n238, n232, n220, n214, n208, n159}), .rdat(reg27), .test_si(
        lt_reg26_0), .test_se(test_se) );
  glsta_a0_4 u0_reg28 ( .clk(clk), .arstz(n71), .rst0(1'b0), .set2(i2c_ev), 
        .clr1(clr28), .rdat(reg28), .irq(irq28), .test_si(reg27[7]), .test_se(
        test_se) );
  glreg_a0_67 u0_reg31 ( .clk(clk), .arstz(n72), .we(upd31), .wdat(i_pc[15:8]), 
        .rdat(reg31), .test_si(reg28[7]), .test_se(test_se) );
  glreg_8_00000001 u0_regD1 ( .clk(clk), .arstz(n39), .we(we_209), .wdat({n255, 
        n249, n238, n232, n220, n214, n208, n135}), .rdat({r_exist1st, 
        r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, r_gpio_oe[6], r_gpio_pu[6], 
        r_gpio_pd[6]}), .test_si(regAF[7]), .test_se(test_se) );
  glreg_8_00000011 u0_regD3 ( .clk(clk), .arstz(n37), .we(we_211), .wdat({n255, 
        n249, n238, n231, n220, n214, n208, n135}), .rdat({regD3_7_, 
        r_gpio_oe[5], r_gpio_pu[5], r_gpio_pd[5], regD3_3, r_gpio_oe[4], 
        r_gpio_pu[4], r_gpio_pd[4]}), .test_si(r_exist1st), .test_se(test_se)
         );
  glreg_WIDTH3 u4_regD4 ( .clk(clk), .arstz(n92), .we(n368), .wdat({n255, n249, 
        n238}), .rdat({test_so2, regD4_6_, regD4_5_}), .test_si(regD4_4_), 
        .test_se(test_se) );
  glreg_WIDTH2_2 u3_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n368), .wdat({
        n231, n219}), .rdat({regD4_4_, regD4_3_}), .test_si(regD4_2_), 
        .test_se(test_se) );
  glreg_WIDTH1_5 u2_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n368), .wdat(
        n213), .rdat(regD4_2_), .test_si(r_i2c_deva[7]), .test_se(test_se) );
  glreg_WIDTH1_4 u1_regD4 ( .clk(clk), .arstz(osc_low_rstz), .we(n368), .wdat(
        n207), .rdat(regD4_1_), .test_si(r_hwi2c_en), .test_se(test_se) );
  glreg_WIDTH1_3 u0_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n9), .wdat(n135), .rdat(regD4_0_), .test_si(regD3_7_), .test_se(test_se) );
  glreg_8_000000f0 u0_regD5 ( .clk(clk), .arstz(n33), .we(we_213), .wdat({n254, 
        n248, n241, n231, n221, n214, n208, n159}), .rdat({r_gpio_pu[3:0], 
        r_gpio_pd[3:0]}), .test_si(regD4_0_), .test_se(test_se) );
  glreg_8_00000098 u0_regD6 ( .clk(clk), .arstz(n34), .we(we_214), .wdat({n254, 
        n249, n238, n231, n219, n214, n208, n159}), .rdat({r_gpio_oe[1], 
        r_gpio_s1, r_gpio_oe[0], r_gpio_s0}), .test_si(r_gpio_pu[3]), 
        .test_se(test_se) );
  glreg_8_00000032 u0_regD7 ( .clk(clk), .arstz(n35), .we(we_215), .wdat({n255, 
        n249, n241, n231, n221, n214, n207, n159}), .rdat({r_gpio_oe[3], 
        r_gpio_s3, r_gpio_oe[2], r_gpio_s2}), .test_si(r_gpio_oe[1]), 
        .test_se(test_se) );
  glreg_a0_66 u0_regD9 ( .clk(clk), .arstz(n63), .we(we_217), .wdat({n255, 
        n249, n238, n232, n221, n214, n208, n159}), .rdat({r_ana_tm, 
        r_fortxdat, r_fortxrdy, r_fortxen, r_sleep}), .test_si(r_gpio_oe[3]), 
        .test_se(test_se) );
  glreg_a0_65 u0_regDE ( .clk(clk), .arstz(n70), .we(we_222), .wdat({n256, 
        n249, n239, n232, n221, n215, n209, n159}), .rdat(regDE), .test_si(
        r_ana_tm[3]), .test_se(test_se) );
  glsta_a0_3 u0_regDF ( .clk(clk), .arstz(n69), .rst0(1'b0), .set2(setDF), 
        .clr1(clrDF), .rdat(regDF), .irq(irqDF), .test_si(regDE[7]), .test_se(
        test_se) );
  glreg_a0_64 u0_reg8F ( .clk(clk), .arstz(n68), .we(we_143), .wdat({n256, 
        n250, n239, n233, n221, n215, n209, n160}), .rdat(r_dpdmctl), 
        .test_si(reg06[7]), .test_se(test_se) );
  glreg_WIDTH4 u0_reg94 ( .clk(clk), .arstz(n87), .we(we_148), .wdat({n250, 
        n239, n233, n221}), .rdat(reg94[6:3]), .test_si(reg31[7]), .test_se(
        test_se) );
  glreg_a0_63 u0_regA1 ( .clk(clk), .arstz(n66), .we(we[161]), .wdat({n256, 
        n250, n239, n233, n221, n215, n209, n160}), .rdat(r_regtrm[7:0]), 
        .test_si(reg94[6]), .test_se(test_se) );
  glreg_a0_62 u0_regA2 ( .clk(clk), .arstz(n65), .we(we[162]), .wdat({n256, 
        n250, n239, n233, n221, n215, n209, n160}), .rdat(r_regtrm[15:8]), 
        .test_si(r_regtrm[7]), .test_se(test_se) );
  glreg_a0_61 u0_regA3 ( .clk(clk), .arstz(n64), .we(we[163]), .wdat({n256, 
        n250, n239, n233, n222, n215, n209, n160}), .rdat(r_regtrm[23:16]), 
        .test_si(r_regtrm[15]), .test_se(test_se) );
  glreg_a0_60 u0_regA4 ( .clk(clk), .arstz(n58), .we(we[164]), .wdat({n256, 
        n250, n239, n233, n222, n215, n209, n160}), .rdat(r_regtrm[31:24]), 
        .test_si(r_regtrm[23]), .test_se(test_se) );
  glreg_a0_59 u0_regA5 ( .clk(clk), .arstz(n62), .we(we[165]), .wdat({n256, 
        n250, n239, n233, n222, n215, n209, n160}), .rdat(r_regtrm[39:32]), 
        .test_si(r_regtrm[31]), .test_se(test_se) );
  glreg_a0_58 u0_regA6 ( .clk(clk), .arstz(n61), .we(we[166]), .wdat({n256, 
        n250, n239, n233, n222, n215, n209, n160}), .rdat(r_regtrm[47:40]), 
        .test_si(r_regtrm[39]), .test_se(test_se) );
  glreg_a0_57 u0_regA7 ( .clk(clk), .arstz(n60), .we(we[167]), .wdat({n256, 
        n250, n240, n233, n222, n215, n209, n160}), .rdat(r_regtrm[55:48]), 
        .test_si(r_regtrm[47]), .test_se(test_se) );
  glreg_a0_56 u0_regAB ( .clk(clk), .arstz(n55), .we(we_171), .wdat({n257, 
        n251, n240, n234, n222, n216, n209, n160}), .rdat(regAB), .test_si(
        r_regtrm[55]), .test_se(test_se) );
  glreg_8_00000028 u0_regAC ( .clk(clk), .arstz(n36), .we(we_172), .wdat({n257, 
        n251, n241, n234, n219, n216, n210, n172}), .rdat(regAC), .test_si(
        regAB[7]), .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_2 u2_ovp_db ( .o_dbc(reg94[2]), .o_chg(), .i_org(
        srci[2]), .clk(clk_500), .rstz(n81), .test_si(n272), .test_so(n271), 
        .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_1 u1_ocp_db ( .o_dbc(reg94[1]), .o_chg(), .i_org(
        srci[1]), .clk(clk_500), .rstz(n80), .test_si(n276), .test_so(n275), 
        .test_se(test_se) );
  dbnc_WIDTH4_TIMEOUT14_0 u1_uvp_db ( .o_dbc(reg94[0]), .o_chg(), .i_org(
        srci[0]), .clk(clk_500), .rstz(n82), .test_si(n273), .test_so(n272), 
        .test_se(test_se) );
  dbnc_WIDTH5_TIMEOUT30 u1_ovp_db ( .o_dbc(m_ovp), .o_chg(m_ovp_sta), .i_org(
        srci[2]), .clk(clk_1p0m), .rstz(n78), .test_si(n275), .test_so(n274), 
        .test_se(test_se) );
  dbnc_WIDTH2_4 u0_otpi_db ( .o_dbc(regAD[3]), .o_chg(setAE[3]), .i_org(
        srci[5]), .clk(clk_1p0m), .rstz(n87), .test_si(n282), .test_so(n281), 
        .test_se(test_se) );
  dbnc_WIDTH2_3 u0_ocp_db ( .o_dbc(regAD[1]), .o_chg(setAE[1]), .i_org(srci[1]), .clk(clk_1p0m), .rstz(n88), .test_si(n283), .test_so(n282), .test_se(test_se) );
  dbnc_WIDTH2_2 u0_uvp_db ( .o_dbc(regAD[0]), .o_chg(setAE[0]), .i_org(srci[0]), .clk(clk_1p0m), .rstz(n91), .test_si(n278), .test_so(n277), .test_se(test_se) );
  dbnc_WIDTH2_1 u1_scp_db ( .o_dbc(m_scp), .o_chg(m_scp_sta), .i_org(srci[3]), 
        .clk(clk_1p0m), .rstz(n88), .test_si(r_fw_pwrv[3]), .test_so(n273), 
        .test_se(test_se) );
  dbnc_WIDTH2_0 u0_dmf_db ( .o_dbc(regAD_7), .o_chg(setAE_7), .i_org(dm_fault), 
        .clk(clk_1p0m), .rstz(n91), .test_si(n284), .test_so(n283), .test_se(
        test_se) );
  dbnc_WIDTH2_TIMEOUT2_14 u0_otps_db ( .o_dbc(reg94[7]), .o_chg(), .i_org(
        srci[5]), .clk(clk), .rstz(n85), .test_si(n281), .test_so(n280), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_13 u0_cc1_db ( .o_dbc(regF4_3), .o_chg(), .i_org(cc1_di), .clk(clk), .rstz(n89), .test_si(rstcnt[4]), .test_so(n285), .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_12 u0_cc2_db ( .o_dbc(regF4_7_), .o_chg(), .i_org(
        cc2_di), .clk(clk), .rstz(n85), .test_si(n285), .test_so(n284), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_11 u0_ovp_db ( .o_dbc(s_ovp), .o_chg(s_ovp_sta), 
        .i_org(srci[2]), .clk(clk), .rstz(n89), .test_si(n280), .test_so(n279), 
        .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_10 u0_scp_db ( .o_dbc(s_scp), .o_chg(s_scp_sta), 
        .i_org(srci[3]), .clk(clk), .rstz(n90), .test_si(r_cctrx[7]), 
        .test_so(n278), .test_se(test_se) );
  dbnc_WIDTH2_TIMEOUT2_9 u0_v5oc_db ( .o_dbc(regAD[5]), .o_chg(setAE[5]), 
        .i_org(srci[4]), .clk(clk), .rstz(n90), .test_si(n277), .test_so(n276), 
        .test_se(test_se) );
  glsta_a0_2 u0_regAE ( .clk(clk), .arstz(n50), .rst0(1'b0), .set2({setAE_7, 
        1'b0, setAE}), .clr1(clrAE), .rdat(regAE), .irq(irqAE), .test_si(
        regAC[7]), .test_se(test_se) );
  glreg_a0_55 u0_regAF ( .clk(clk), .arstz(n49), .we(we_175), .wdat({n257, 
        n251, n240, n234, n222, n216, n210, n172}), .rdat(regAF), .test_si(
        regAE[7]), .test_se(test_se) );
  glreg_WIDTH7_2 u0_regE3 ( .clk(clk), .arstz(n77), .we(n206), .wdat({n257, 
        n251, n240, n234, n222, n216, n172}), .rdat({r_srcctl[7:4], regE3, 
        regE3_0}), .test_si(regDF[7]), .test_se(test_se) );
  glreg_4_00000004 u1_regE4 ( .clk(clk), .arstz(n84), .we(r_pwrv_upd), .wdat(
        lt_regE4_3_0), .rdat(r_fw_pwrv[3:0]), .test_si(regD4_1_), .test_se(
        test_se) );
  glreg_8_00000004 u0_regE4 ( .clk(clk), .arstz(n38), .we(we_228), .wdat({n257, 
        n251, n240, n234, n222, n213, n210, n172}), .rdat({r_pwrctl, 
        lt_regE4_3_0}), .test_si(r_srcctl[7]), .test_se(test_se) );
  glreg_8_0000001f u0_regE5 ( .clk(clk), .arstz(n32), .we(r_pwrv_upd), .wdat({
        n257, n251, n240, n231, n219, n213, n207, n135}), .rdat(
        r_fw_pwrv[11:4]), .test_si(r_pwrctl[7]), .test_se(test_se) );
  glreg_a0_54 u0_regE6 ( .clk(clk), .arstz(n47), .we(we_230), .wdat({n257, 
        n251, n240, n234, n223, n216, n210, n172}), .rdat(r_ccrx), .test_si(
        r_fw_pwrv[11]), .test_se(test_se) );
  glreg_a0_53 u0_regE7 ( .clk(clk), .arstz(n46), .we(we_231), .wdat({n257, 
        n251, n240, n234, n223, n216, n210, n172}), .rdat(r_ccctl), .test_si(
        r_ccrx[7]), .test_se(test_se) );
  glreg_a0_52 u0_regE8 ( .clk(clk), .arstz(n45), .we(we_232), .wdat({n257, 
        n251, n240, n234, n222, n216, n210, n172}), .rdat(r_comp_opt), 
        .test_si(r_ccctl[7]), .test_se(test_se) );
  glreg_a0_51 u0_regF5 ( .clk(clk), .arstz(n44), .we(we_245), .wdat({n257, 
        n251, n240, n234, n220, n216, n210, n172}), .rdat(r_cvctl), .test_si(
        r_comp_opt[7]), .test_se(test_se) );
  glreg_a0_50 u0_regF6 ( .clk(clk), .arstz(n43), .we(we_246), .wdat({n254, 
        n248, n241, n231, n221, n213, n207, n135}), .rdat(r_cctrx), .test_si(
        r_cvctl[7]), .test_se(test_se) );
  SNPS_CLOCK_GATE_HIGH_regbank_a0_1 clk_gate_rstcnt_reg ( .CLK(clk), .EN(N26), 
        .ENCLK(net10815), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_regbank_a0_0 clk_gate_lg_pulse_cnt_reg ( .CLK(clk_1p0m), 
        .EN(N108), .ENCLK(net10821), .TE(test_se) );
  regbank_a0_DW01_add_0 add_526 ( .A(regAC), .B(regAB), .CI(1'b0), .SUM(
        r_pwr_i), .CO() );
  regbank_a0_DW01_inc_0 add_304 ( .A({1'b0, r_inst_ofs}), .SUM({
        SYNOPSYS_UNCONNECTED_1, inst_ofs_plus}) );
  regbank_a0_DW_rightsh_2 srl_133 ( .A({dac_r_vs, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, r_cctrx, r_cvctl, regF4_7_, x_daclsb[5:3], regF4_3, 
        x_daclsb[2:0], r_sar_en, r_dac_en, dac_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_comp_opt, r_ccctl, r_ccrx, r_fw_pwrv[11:4], r_pwrctl, r_fw_pwrv[3:0], 
        r_srcctl[7:4], regE3, r_srcctl[1], regE3_0, dac_r_cmpsta, dac_r_comp, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, regDF, regDE, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_ana_tm, r_fortxdat, 
        r_fortxrdy, r_fortxen, r_sleep, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, r_gpio_oe[3], r_gpio_s3, r_gpio_oe[2], r_gpio_s2, 
        r_gpio_oe[1], r_gpio_s1, r_gpio_oe[0], r_gpio_s0, r_gpio_pu[3:0], 
        r_gpio_pd[3:0], test_so2, regD4_6_, regD4_5_, regD4_4_, regD4_3_, 
        regD4_2_, regD4_1_, regD4_0_, regD3_7_, r_gpio_oe[5], r_gpio_pu[5], 
        r_gpio_pd[5], regD3_3, r_gpio_oe[4], r_gpio_pu[4], r_gpio_pd[4], 
        i_i2c_rwbuf, r_exist1st, r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, 
        r_gpio_oe[6], r_gpio_pu[6], r_gpio_pd[6], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, reg31, reg30, i_i2c_ltbuf, reg28, reg27, r_i2c_deva, 
        r_hwi2c_en, 1'b0, 1'b0, r_i2c_attr, r_pg0_sel, reg25_0_, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, prx_rcvinf[4], REVID, 
        prx_rcvinf[3], ptx_fsm, prx_fsm, reg21, r_dat_portrole, r_dat_spec, 
        r_dat_datarole, reg20, n16, r_inst_ofs, i_i2c_ofs, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, dbgpo[31:24], r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1], prl_cpmsgid, prl_cany0, 
        prx_rcvinf[2:0], prl_fsm, reg12, r_txshrt, reg12_1, r_pshords, 
        reg11_7_, r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0], 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, pff_empty, 
        pff_full, pff_ptr, reg06, reg05, dbgpo[15:0], pff_rdat, r_last, 
        r_first, r_unlock, r_txnumk, r_txendk, r_txauto, regAF, regAE, regAD_7, 
        1'b0, regAD, regAC, regAB, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_regtrm, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, fcp_r_crc, fcp_r_dat, fcp_r_msk, fcp_r_sta, 
        fcp_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, fcp_r_acc, r_accctl, fcp_r_tui, reg94, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, r_isofs, r_adofs, r_dpdmctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_cvofs, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .DATA_TC(1'b0), .SH({sfr_addr[6:0], 1'b0, 
        1'b0, 1'b0}), .B({SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, 
        SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, 
        SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, 
        SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, 
        SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, 
        SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, 
        SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, 
        SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, 
        SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, 
        SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, 
        SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, 
        SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, 
        SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, 
        SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, 
        SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, 
        SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, 
        SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, 
        SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, 
        SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, 
        SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, 
        SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, 
        SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, 
        SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, 
        SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, 
        SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, 
        SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, 
        SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, 
        SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, 
        SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, 
        SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, 
        SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, 
        SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, 
        SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, 
        SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, 
        SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, 
        SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, 
        SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, 
        SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, 
        SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, 
        SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, 
        SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, 
        SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, 
        SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, 
        SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, 
        SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, 
        SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, 
        SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, 
        SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, 
        SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, 
        SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, 
        SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, 
        SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, 
        SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, 
        SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, 
        SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, 
        SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, 
        SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, 
        SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, 
        SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, 
        SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, 
        SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, 
        SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, 
        SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, 
        SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, 
        SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, 
        SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, 
        SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, 
        SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, 
        SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, 
        SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, 
        SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, 
        SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, 
        SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, 
        SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, 
        SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, 
        SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, 
        SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, 
        SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, 
        SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, 
        SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, 
        SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, 
        SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, 
        SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, 
        SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, 
        SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, 
        SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, 
        SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, 
        SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, 
        SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, 
        SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, 
        SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, 
        SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, 
        SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, 
        SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, 
        SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, 
        SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, 
        SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, 
        SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, 
        SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, 
        SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, 
        SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, 
        SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, 
        SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, 
        SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, 
        SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, 
        SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, 
        SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, 
        SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, 
        SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, 
        SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, 
        SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, 
        SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, 
        SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, 
        SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, 
        SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, 
        SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, 
        SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, 
        SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, 
        SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, 
        SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, 
        SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, 
        SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, 
        SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, 
        SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, 
        SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, 
        SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, 
        SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, 
        SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, 
        SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, 
        SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, 
        SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, 
        SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, 
        SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, 
        SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, 
        SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, 
        SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, 
        SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, 
        SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, 
        SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, 
        SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, 
        SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, 
        SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, 
        SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, 
        SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, 
        SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, 
        SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, 
        SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, 
        SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, 
        SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, 
        SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, 
        SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, 
        SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, 
        SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, 
        SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, 
        SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, 
        SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, 
        SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, 
        SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, 
        SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, 
        SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, 
        SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, 
        SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, 
        SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, 
        SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, 
        SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, 
        SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, 
        SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, 
        SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, 
        SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, 
        SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, 
        SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, 
        SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, 
        SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, 
        SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, 
        SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, 
        SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, 
        SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, 
        SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, 
        SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, 
        SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, 
        SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, 
        SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, 
        SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, 
        SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, 
        SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, 
        SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, 
        SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, 
        SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, 
        SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, 
        SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, 
        SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, 
        SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, 
        SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, 
        SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, 
        SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, 
        SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, 
        SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, 
        SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, 
        SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, 
        SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, 
        SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, 
        SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, 
        SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, 
        SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, 
        SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, 
        SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, 
        SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, 
        SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, 
        SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, 
        SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, 
        SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, 
        SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, 
        SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, 
        SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, 
        SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, 
        SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, 
        SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, 
        SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, 
        SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, 
        SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, 
        SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, 
        SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, 
        SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, 
        SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, 
        SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, 
        SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, 
        SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, 
        SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, 
        SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, 
        SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, 
        SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, 
        SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, 
        SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, 
        SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, 
        SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, 
        SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, 
        SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, 
        SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, 
        SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, 
        SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, 
        SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, 
        SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, 
        SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, 
        SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, 
        SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, 
        SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, 
        SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, 
        SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, 
        SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, 
        SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, 
        SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, 
        SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, 
        SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, 
        SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, 
        SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, 
        SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, 
        SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, 
        SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, 
        SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, 
        SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, 
        SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, 
        SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, 
        SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, 
        SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, 
        SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, 
        SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, 
        SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, 
        SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, 
        SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, 
        SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, 
        SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, 
        SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, 
        SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, 
        SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, 
        SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, 
        SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, 
        SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, 
        SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, 
        SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, 
        SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017, sfr_rdat}) );
  SDFFRQX1 r_phyrst_reg_0_ ( .D(n1221), .SIN(oscdwn_shft[2]), .SMC(test_se), 
        .C(clk), .XR(n2), .Q(r_phyrst[0]) );
  SDFFRQX1 lg_pulse_cnt_reg_3_ ( .D(N112), .SIN(lg_pulse_cnt[2]), .SMC(test_se), .C(net10821), .XR(n92), .Q(lg_pulse_cnt[3]) );
  SDFFRQX1 lg_pulse_cnt_reg_4_ ( .D(N113), .SIN(lg_pulse_cnt[3]), .SMC(test_se), .C(net10821), .XR(n92), .Q(lg_pulse_cnt[4]) );
  SDFFRQX1 lg_pulse_cnt_reg_1_ ( .D(N110), .SIN(lg_pulse_cnt[0]), .SMC(test_se), .C(net10821), .XR(n92), .Q(lg_pulse_cnt[1]) );
  SDFFRQX1 lg_pulse_cnt_reg_2_ ( .D(N111), .SIN(lg_pulse_cnt[1]), .SMC(test_se), .C(net10821), .XR(n92), .Q(lg_pulse_cnt[2]) );
  SDFFRQX1 rstcnt_reg_0_ ( .D(N39), .SIN(r_phyrst[1]), .SMC(test_se), .C(
        net10815), .XR(n3), .Q(rstcnt[0]) );
  SDFFRQX1 lg_pulse_cnt_reg_0_ ( .D(N109), .SIN(lg_pulse_12m), .SMC(test_se), 
        .C(net10821), .XR(n93), .Q(lg_pulse_cnt[0]) );
  SDFFRQX1 d_p0_reg_7_ ( .D(ff_p0[7]), .SIN(d_p0[6]), .SMC(test_se), .C(clk), 
        .XR(n93), .Q(d_p0[7]) );
  SDFFRQX1 d_p0_reg_6_ ( .D(ff_p0[6]), .SIN(d_p0[5]), .SMC(test_se), .C(clk), 
        .XR(n93), .Q(d_p0[6]) );
  SDFFRQX1 d_p0_reg_5_ ( .D(ff_p0[5]), .SIN(d_p0[4]), .SMC(test_se), .C(clk), 
        .XR(n93), .Q(d_p0[5]) );
  SDFFRQX1 d_p0_reg_4_ ( .D(ff_p0[4]), .SIN(d_p0[3]), .SMC(test_se), .C(clk), 
        .XR(n93), .Q(d_p0[4]) );
  SDFFRQX1 d_p0_reg_3_ ( .D(ff_p0[3]), .SIN(d_p0[2]), .SMC(test_se), .C(clk), 
        .XR(n93), .Q(d_p0[3]) );
  SDFFRQX1 d_p0_reg_2_ ( .D(ff_p0[2]), .SIN(d_p0[1]), .SMC(test_se), .C(clk), 
        .XR(n93), .Q(d_p0[2]) );
  SDFFRQX1 d_p0_reg_1_ ( .D(ff_p0[1]), .SIN(d_p0[0]), .SMC(test_se), .C(clk), 
        .XR(n93), .Q(d_p0[1]) );
  SDFFRQX1 d_p0_reg_0_ ( .D(ff_p0[0]), .SIN(test_si2), .SMC(test_se), .C(clk), 
        .XR(n93), .Q(d_p0[0]) );
  SDFFRQX1 r_phyrst_reg_1_ ( .D(n1220), .SIN(r_phyrst[0]), .SMC(test_se), .C(
        clk), .XR(n2), .Q(r_phyrst[1]) );
  SDFFNRQX1 osc_gate_n_reg_3_ ( .D(osc_gate_n_2_), .SIN(osc_gate_n_2_), .SMC(
        test_se), .XC(xclk), .XR(n3), .Q(test_so1) );
  SDFFNRQX1 osc_gate_n_reg_0_ ( .D(r_pos_gate), .SIN(test_si1), .SMC(test_se), 
        .XC(xclk), .XR(n2), .Q(osc_gate_n_0_) );
  SDFFNRQX1 osc_gate_n_reg_1_ ( .D(osc_gate_n_0_), .SIN(osc_gate_n_0_), .SMC(
        test_se), .XC(xclk), .XR(n3), .Q(osc_gate_n_1_) );
  SDFFNRQX1 osc_gate_n_reg_2_ ( .D(osc_gate_n_1_), .SIN(osc_gate_n_1_), .SMC(
        test_se), .XC(xclk), .XR(n2), .Q(osc_gate_n_2_) );
  SDFFQX1 oscdwn_shft_reg_1_ ( .D(oscdwn_shft[0]), .SIN(oscdwn_shft[0]), .SMC(
        test_se), .C(clk), .Q(oscdwn_shft[1]) );
  SDFFRQX1 drstz_reg_1_ ( .D(drstz[0]), .SIN(drstz[0]), .SMC(test_se), .C(clk), 
        .XR(n3), .Q(drstz[1]) );
  SDFFRQX1 rstcnt_reg_1_ ( .D(N38), .SIN(rstcnt[0]), .SMC(test_se), .C(
        net10815), .XR(n2), .Q(rstcnt[1]) );
  SDFFRQX1 rstcnt_reg_2_ ( .D(N37), .SIN(rstcnt[1]), .SMC(test_se), .C(
        net10815), .XR(n3), .Q(rstcnt[2]) );
  SDFFRQX1 rstcnt_reg_4_ ( .D(N35), .SIN(rstcnt[3]), .SMC(test_se), .C(
        net10815), .XR(n2), .Q(rstcnt[4]) );
  SDFFRQX1 rstcnt_reg_3_ ( .D(N36), .SIN(rstcnt[2]), .SMC(test_se), .C(
        net10815), .XR(n3), .Q(rstcnt[3]) );
  SDFFQX1 oscdwn_shft_reg_2_ ( .D(n367), .SIN(oscdwn_shft[1]), .SMC(test_se), 
        .C(clk), .Q(oscdwn_shft[2]) );
  SDFFRQX1 lg_pulse_reg ( .D(n1219), .SIN(lg_pulse_cnt[4]), .SMC(test_se), .C(
        clk_1p0m), .XR(n113), .Q(lg_dischg) );
  SDFFRQX1 lg_pulse_12m_reg ( .D(n1218), .SIN(drstz[1]), .SMC(test_se), .C(clk), .XR(n93), .Q(lg_pulse_12m) );
  INVX1 U354 ( .A(n20), .Y(srstz) );
  SDFFQX1 oscdwn_shft_reg_0_ ( .D(N84), .SIN(lg_dischg), .SMC(test_se), .C(clk), .Q(oscdwn_shft[0]) );
  SDFFRQX1 drstz_reg_0_ ( .D(1'b1), .SIN(d_p0[7]), .SMC(test_se), .C(clk), 
        .XR(n2), .Q(drstz[0]) );
  MUX2X1 U8 ( .D0(pff_rxpart[5]), .D1(n241), .S(n268), .Y(wd20[5]) );
  INVXL U9 ( .A(xrstz), .Y(n1) );
  INVXL U10 ( .A(n1), .Y(n2) );
  INVXL U11 ( .A(n1), .Y(n3) );
  INVXL U12 ( .A(n314), .Y(n9) );
  BUFXL U13 ( .A(sfr_addr[5]), .Y(n10) );
  BUFXL U14 ( .A(n10), .Y(n11) );
  BUFXL U15 ( .A(sfr_addr[6]), .Y(n12) );
  INVX1 U16 ( .A(n263), .Y(n13) );
  INVX1 U17 ( .A(n312), .Y(n14) );
  INVX1 U18 ( .A(reg19_7_), .Y(n15) );
  INVX1 U19 ( .A(n15), .Y(n16) );
  INVX1 U20 ( .A(n365), .Y(n17) );
  BUFX3 U21 ( .A(n369), .Y(n18) );
  BUFX3 U22 ( .A(n100), .Y(n19) );
  BUFX3 U23 ( .A(phyrst), .Y(n21) );
  BUFXL U24 ( .A(pff_ptr[4]), .Y(dbgpo[20]) );
  BUFXL U25 ( .A(pff_ptr[0]), .Y(dbgpo[16]) );
  BUFXL U26 ( .A(pff_ptr[1]), .Y(dbgpo[17]) );
  BUFXL U27 ( .A(pff_ptr[3]), .Y(dbgpo[19]) );
  BUFXL U28 ( .A(pff_ptr[2]), .Y(dbgpo[18]) );
  BUFXL U29 ( .A(pff_ptr[5]), .Y(dbgpo[21]) );
  INVXL U30 ( .A(n10), .Y(n132) );
  MUX2XL U31 ( .D0(i_pc[1]), .D1(prx_adpn[1]), .S(reg19_7_), .Y(reg30[1]) );
  INVX1 U32 ( .A(n225), .Y(n219) );
  INVX1 U33 ( .A(n245), .Y(n240) );
  INVX1 U34 ( .A(n245), .Y(n239) );
  INVX1 U35 ( .A(n244), .Y(n238) );
  INVX1 U36 ( .A(n224), .Y(n223) );
  INVX1 U37 ( .A(n243), .Y(n241) );
  INVX1 U38 ( .A(n228), .Y(n222) );
  INVX1 U39 ( .A(n227), .Y(n221) );
  INVX1 U40 ( .A(n226), .Y(n220) );
  BUFX3 U41 ( .A(n230), .Y(n225) );
  BUFX3 U42 ( .A(n247), .Y(n242) );
  NOR3XL U43 ( .A(n133), .B(n237), .C(n217), .Y(r_discard) );
  BUFX3 U44 ( .A(n230), .Y(n224) );
  INVX1 U45 ( .A(n259), .Y(n254) );
  INVX1 U46 ( .A(n253), .Y(n248) );
  INVX1 U47 ( .A(n237), .Y(n231) );
  INVX1 U48 ( .A(n237), .Y(n234) );
  INVX1 U49 ( .A(n212), .Y(n207) );
  INVX1 U50 ( .A(n237), .Y(n233) );
  INVX1 U51 ( .A(n237), .Y(n232) );
  BUFX3 U52 ( .A(n247), .Y(n243) );
  BUFX3 U53 ( .A(n243), .Y(n244) );
  INVX1 U54 ( .A(n237), .Y(n235) );
  INVX1 U55 ( .A(n176), .Y(n135) );
  INVX1 U56 ( .A(n218), .Y(n213) );
  INVX1 U57 ( .A(n253), .Y(n251) );
  INVX1 U58 ( .A(n259), .Y(n257) );
  INVX1 U59 ( .A(n253), .Y(n250) );
  INVX1 U60 ( .A(n259), .Y(n256) );
  INVX1 U61 ( .A(n253), .Y(n249) );
  INVX1 U62 ( .A(n259), .Y(n255) );
  INVX1 U63 ( .A(n176), .Y(n172) );
  INVX1 U64 ( .A(n218), .Y(n216) );
  INVX1 U65 ( .A(n212), .Y(n210) );
  BUFX3 U66 ( .A(n243), .Y(n245) );
  BUFX3 U67 ( .A(n226), .Y(n227) );
  BUFX3 U68 ( .A(n230), .Y(n226) );
  BUFX3 U69 ( .A(n226), .Y(n228) );
  BUFX3 U70 ( .A(n226), .Y(n229) );
  BUFX3 U71 ( .A(n243), .Y(n246) );
  INVX1 U72 ( .A(n212), .Y(n209) );
  INVX1 U73 ( .A(n218), .Y(n215) );
  INVX1 U74 ( .A(n176), .Y(n160) );
  INVX1 U75 ( .A(n212), .Y(n208) );
  INVX1 U76 ( .A(n217), .Y(n214) );
  INVX1 U77 ( .A(n176), .Y(n159) );
  INVX1 U78 ( .A(atpg_en), .Y(n260) );
  INVX1 U79 ( .A(sfr_wdat[3]), .Y(n230) );
  AND2X1 U80 ( .A(n335), .B(n351), .Y(r_dacwr[5]) );
  AND2X1 U81 ( .A(n335), .B(n338), .Y(r_dacwr[2]) );
  AND2X1 U82 ( .A(n335), .B(n346), .Y(r_dacwr[7]) );
  AND2X1 U83 ( .A(n335), .B(n349), .Y(r_dacwr[4]) );
  AND2X1 U84 ( .A(n335), .B(n345), .Y(r_dacwr[3]) );
  AND2X1 U85 ( .A(n335), .B(n340), .Y(r_dacwr[1]) );
  INVX1 U86 ( .A(n327), .Y(r_fifopsh) );
  INVX1 U87 ( .A(sfr_wdat[5]), .Y(n247) );
  INVX1 U88 ( .A(sfr_wdat[6]), .Y(n252) );
  NAND4X1 U89 ( .A(n254), .B(n175), .C(n248), .D(n163), .Y(n133) );
  NOR2X1 U90 ( .A(n225), .B(n128), .Y(n163) );
  INVX1 U91 ( .A(sfr_wdat[4]), .Y(n236) );
  INVX1 U92 ( .A(sfr_wdat[1]), .Y(n211) );
  INVX1 U93 ( .A(sfr_wdat[7]), .Y(n258) );
  INVX1 U94 ( .A(sfr_wdat[2]), .Y(n217) );
  INVX1 U95 ( .A(sfr_wdat[0]), .Y(n175) );
  INVX1 U96 ( .A(n330), .Y(n206) );
  NAND21X1 U97 ( .B(n117), .A(n131), .Y(n102) );
  AND2X1 U98 ( .A(n348), .B(n351), .Y(r_fcpwr[4]) );
  AND2X1 U99 ( .A(n205), .B(n254), .Y(r_i2c_fwack) );
  AND2X1 U100 ( .A(n320), .B(n241), .Y(clr28[5]) );
  AND2X1 U101 ( .A(n320), .B(n207), .Y(clr28[1]) );
  AND2X1 U102 ( .A(n325), .B(n241), .Y(clr04[5]) );
  AND2X1 U103 ( .A(n325), .B(n207), .Y(clr04[1]) );
  AND2X1 U104 ( .A(n320), .B(n231), .Y(clr28[4]) );
  AND2X1 U105 ( .A(n320), .B(n135), .Y(clr28[0]) );
  AND2X1 U106 ( .A(n325), .B(n231), .Y(clr04[4]) );
  AND2X1 U107 ( .A(n325), .B(n135), .Y(clr04[0]) );
  AND2X1 U108 ( .A(n320), .B(n248), .Y(clr28[6]) );
  AND2X1 U109 ( .A(n320), .B(n213), .Y(clr28[2]) );
  AND2X1 U110 ( .A(n325), .B(n248), .Y(clr04[6]) );
  AND2X1 U111 ( .A(n325), .B(n213), .Y(clr04[2]) );
  AND2X1 U112 ( .A(n320), .B(n254), .Y(clr28[7]) );
  AND2X1 U113 ( .A(n320), .B(n219), .Y(clr28[3]) );
  AND2X1 U114 ( .A(n325), .B(n254), .Y(clr04[7]) );
  AND2X1 U115 ( .A(n325), .B(n219), .Y(clr04[3]) );
  INVX1 U116 ( .A(n366), .Y(n364) );
  INVX1 U117 ( .A(n374), .Y(n204) );
  NOR2X1 U118 ( .A(n243), .B(n174), .Y(clrAE[5]) );
  NOR2X1 U119 ( .A(n211), .B(n174), .Y(clrAE[1]) );
  NOR2X1 U120 ( .A(n244), .B(n177), .Y(clr03[5]) );
  NOR2X1 U121 ( .A(n212), .B(n177), .Y(clr03[1]) );
  NOR2X1 U122 ( .A(n242), .B(n173), .Y(clrDF[5]) );
  NOR2X1 U123 ( .A(n211), .B(n173), .Y(clrDF[1]) );
  NOR2X1 U124 ( .A(n237), .B(n174), .Y(clrAE[4]) );
  NOR2X1 U125 ( .A(n176), .B(n174), .Y(clrAE[0]) );
  NOR2X1 U126 ( .A(n237), .B(n177), .Y(clr03[4]) );
  NOR2X1 U127 ( .A(n176), .B(n177), .Y(clr03[0]) );
  NOR2X1 U128 ( .A(n237), .B(n173), .Y(clrDF[4]) );
  NOR2X1 U129 ( .A(n175), .B(n173), .Y(clrDF[0]) );
  NOR2X1 U130 ( .A(n253), .B(n174), .Y(clrAE[6]) );
  NOR2X1 U131 ( .A(n218), .B(n174), .Y(clrAE[2]) );
  NOR2X1 U132 ( .A(n253), .B(n177), .Y(clr03[6]) );
  NOR2X1 U133 ( .A(n218), .B(n177), .Y(clr03[2]) );
  NOR2X1 U134 ( .A(n253), .B(n173), .Y(clrDF[6]) );
  NOR2X1 U135 ( .A(n217), .B(n173), .Y(clrDF[2]) );
  NOR2X1 U136 ( .A(n259), .B(n174), .Y(clrAE[7]) );
  NOR2X1 U137 ( .A(n227), .B(n174), .Y(clrAE[3]) );
  NOR2X1 U138 ( .A(n259), .B(n177), .Y(clr03[7]) );
  NOR2X1 U139 ( .A(n228), .B(n177), .Y(clr03[3]) );
  NOR2X1 U140 ( .A(n259), .B(n173), .Y(clrDF[7]) );
  NOR2X1 U141 ( .A(n226), .B(n173), .Y(clrDF[3]) );
  INVX1 U142 ( .A(n291), .Y(n362) );
  AO21X1 U143 ( .B(n338), .C(n360), .A(n125), .Y(upd18) );
  INVX1 U144 ( .A(sfr_wdat[7]), .Y(n259) );
  AND2X1 U145 ( .A(n322), .B(n346), .Y(we_191) );
  AND2X1 U146 ( .A(n302), .B(n346), .Y(we_175) );
  AND2X1 U147 ( .A(n302), .B(n349), .Y(we_172) );
  AND2X1 U148 ( .A(n348), .B(n340), .Y(r_dacwr[14]) );
  AND2X1 U149 ( .A(n348), .B(n349), .Y(we_148) );
  AND2X1 U150 ( .A(n351), .B(n356), .Y(we_181) );
  AND2X1 U151 ( .A(n315), .B(n346), .Y(we_215) );
  AND2X1 U152 ( .A(n315), .B(n351), .Y(we_213) );
  AND2X1 U153 ( .A(n315), .B(n345), .Y(we_211) );
  AND2X1 U154 ( .A(n315), .B(n340), .Y(we_209) );
  AND2X1 U155 ( .A(n340), .B(n311), .Y(we_217) );
  AND2X1 U156 ( .A(n345), .B(n302), .Y(we_171) );
  AND2X1 U157 ( .A(n345), .B(n322), .Y(we_187) );
  INVX1 U158 ( .A(sfr_wdat[6]), .Y(n253) );
  INVX1 U159 ( .A(sfr_wdat[4]), .Y(n237) );
  INVX1 U160 ( .A(sfr_wdat[1]), .Y(n212) );
  INVX1 U161 ( .A(n359), .Y(n302) );
  INVX1 U162 ( .A(sfr_wdat[0]), .Y(n176) );
  INVX1 U163 ( .A(sfr_wdat[2]), .Y(n218) );
  INVX1 U164 ( .A(n131), .Y(n125) );
  INVX1 U165 ( .A(n131), .Y(n130) );
  INVX1 U166 ( .A(n120), .Y(n92) );
  INVX1 U167 ( .A(n120), .Y(n93) );
  INVX1 U168 ( .A(n110), .Y(n84) );
  INVX1 U169 ( .A(n94), .Y(n91) );
  INVX1 U170 ( .A(n115), .Y(n50) );
  INVX1 U171 ( .A(n97), .Y(n69) );
  INVX1 U172 ( .A(n95), .Y(n71) );
  INVX1 U173 ( .A(n107), .Y(n42) );
  INVX1 U174 ( .A(n107), .Y(n41) );
  INVX1 U175 ( .A(n107), .Y(n43) );
  INVX1 U176 ( .A(n105), .Y(n44) );
  INVX1 U177 ( .A(n105), .Y(n45) );
  INVX1 U178 ( .A(n105), .Y(n46) );
  INVX1 U179 ( .A(n115), .Y(n47) );
  INVX1 U180 ( .A(n98), .Y(n49) );
  INVX1 U181 ( .A(n94), .Y(n90) );
  INVX1 U182 ( .A(n94), .Y(n89) );
  INVX1 U183 ( .A(n95), .Y(n85) );
  INVX1 U184 ( .A(n95), .Y(n88) );
  INVX1 U185 ( .A(n101), .Y(n55) );
  INVX1 U186 ( .A(n115), .Y(n60) );
  INVX1 U187 ( .A(n97), .Y(n61) );
  INVX1 U188 ( .A(n98), .Y(n62) );
  INVX1 U189 ( .A(n101), .Y(n58) );
  INVX1 U190 ( .A(n98), .Y(n64) );
  INVX1 U191 ( .A(n94), .Y(n65) );
  INVX1 U192 ( .A(n120), .Y(n66) );
  INVX1 U193 ( .A(n95), .Y(n87) );
  INVX1 U194 ( .A(n97), .Y(n68) );
  INVX1 U195 ( .A(n97), .Y(n70) );
  INVX1 U196 ( .A(n98), .Y(n63) );
  INVX1 U197 ( .A(n111), .Y(n72) );
  INVX1 U198 ( .A(n110), .Y(n73) );
  INVX1 U199 ( .A(n96), .Y(n74) );
  INVX1 U200 ( .A(n95), .Y(n67) );
  INVX1 U201 ( .A(n107), .Y(n59) );
  INVX1 U202 ( .A(n101), .Y(n57) );
  INVX1 U203 ( .A(n101), .Y(n56) );
  INVX1 U204 ( .A(n115), .Y(n54) );
  INVX1 U205 ( .A(n98), .Y(n53) );
  INVX1 U206 ( .A(n107), .Y(n52) );
  INVX1 U207 ( .A(n105), .Y(n51) );
  INVX1 U208 ( .A(n111), .Y(n48) );
  INVX1 U209 ( .A(n120), .Y(n76) );
  INVX1 U210 ( .A(n101), .Y(n77) );
  INVX1 U211 ( .A(n96), .Y(n78) );
  INVX1 U212 ( .A(n96), .Y(n79) );
  INVX1 U213 ( .A(n108), .Y(n82) );
  INVX1 U214 ( .A(n96), .Y(n80) );
  INVX1 U215 ( .A(n96), .Y(n81) );
  AND2X1 U216 ( .A(n336), .B(n340), .Y(r_dacwr[8]) );
  INVX1 U217 ( .A(n314), .Y(n368) );
  NAND21X1 U218 ( .B(n323), .A(n315), .Y(n314) );
  INVX1 U219 ( .A(n288), .Y(n340) );
  INVX1 U220 ( .A(n313), .Y(n315) );
  NAND32X1 U221 ( .B(n312), .C(n333), .A(n132), .Y(n313) );
  AND2X1 U222 ( .A(n335), .B(n13), .Y(r_dacwr[6]) );
  INVX1 U223 ( .A(n323), .Y(n349) );
  INVX1 U224 ( .A(n357), .Y(n345) );
  INVX1 U225 ( .A(n289), .Y(n338) );
  INVX1 U226 ( .A(n361), .Y(n351) );
  INVX1 U227 ( .A(n83), .Y(n346) );
  AND2X1 U228 ( .A(n335), .B(n339), .Y(r_dacwr[0]) );
  INVX1 U229 ( .A(n334), .Y(n335) );
  NAND21X1 U230 ( .B(n333), .A(n332), .Y(n334) );
  OAI31XL U231 ( .A(n127), .B(n128), .C(n129), .D(n376), .Y(r_fiforst) );
  NAND2X1 U232 ( .A(n175), .B(n217), .Y(n129) );
  NAND4X1 U233 ( .A(n224), .B(n236), .C(n252), .D(n258), .Y(n127) );
  NAND43X1 U234 ( .B(n83), .C(n355), .D(n241), .A(n211), .Y(n128) );
  NAND21X1 U235 ( .B(n355), .A(n338), .Y(n327) );
  AND2X1 U236 ( .A(n347), .B(n358), .Y(r_fcpwr[3]) );
  INVX1 U237 ( .A(prl_c0set), .Y(n376) );
  INVX1 U238 ( .A(n99), .Y(n303) );
  INVX1 U239 ( .A(n355), .Y(n356) );
  NAND21X1 U240 ( .B(n357), .A(n337), .Y(n330) );
  NAND21X1 U241 ( .B(n357), .A(n356), .Y(n177) );
  NAND21X1 U242 ( .B(n359), .A(n358), .Y(n174) );
  NAND21X1 U243 ( .B(n289), .A(n329), .Y(n374) );
  NAND21X1 U244 ( .B(n321), .A(n349), .Y(n366) );
  INVX1 U245 ( .A(n266), .Y(n297) );
  INVX1 U246 ( .A(n319), .Y(n320) );
  NAND21X1 U247 ( .B(n323), .A(n329), .Y(n319) );
  INVX1 U248 ( .A(n324), .Y(n325) );
  NAND21X1 U249 ( .B(n323), .A(n356), .Y(n324) );
  INVX1 U250 ( .A(n265), .Y(n205) );
  NAND21X1 U251 ( .B(n288), .A(n329), .Y(n265) );
  NAND21X1 U252 ( .B(n270), .A(n345), .Y(n117) );
  AND2X1 U253 ( .A(n338), .B(n337), .Y(r_dacwr[12]) );
  OR2X1 U254 ( .A(n86), .B(n83), .Y(n173) );
  AND2X1 U255 ( .A(n347), .B(n349), .Y(r_fcpwr[1]) );
  AND2X1 U256 ( .A(n347), .B(n346), .Y(r_fcpwr[5]) );
  NAND21X1 U257 ( .B(n361), .A(n360), .Y(n100) );
  NAND21XL U258 ( .B(n355), .A(n340), .Y(n291) );
  INVX1 U259 ( .A(n267), .Y(n268) );
  NAND21X1 U260 ( .B(n323), .A(n360), .Y(n267) );
  INVX1 U261 ( .A(n287), .Y(r_set_cpmsgid) );
  NAND21X1 U262 ( .B(n321), .A(n358), .Y(n287) );
  INVX1 U263 ( .A(n300), .Y(r_pwrv_upd) );
  NAND21X1 U264 ( .B(n361), .A(n337), .Y(n300) );
  AND2X1 U265 ( .A(n336), .B(n349), .Y(r_dacwr[11]) );
  AND3X1 U266 ( .A(n339), .B(n297), .C(n332), .Y(we_232) );
  AND3X1 U267 ( .A(n352), .B(n312), .C(n346), .Y(we_143) );
  AND2X1 U268 ( .A(n348), .B(n358), .Y(r_fcpwr[6]) );
  AND2X1 U269 ( .A(n336), .B(n358), .Y(we_246) );
  AND2X1 U270 ( .A(n337), .B(n358), .Y(we_230) );
  AND2X1 U271 ( .A(n305), .B(n358), .Y(we[166]) );
  AND2X1 U272 ( .A(n315), .B(n358), .Y(we_214) );
  AND2X1 U273 ( .A(n358), .B(n311), .Y(we_222) );
  AND2X1 U274 ( .A(n358), .B(n356), .Y(we_182) );
  AND2X1 U275 ( .A(n347), .B(n351), .Y(r_fcpwr[2]) );
  AND2X1 U276 ( .A(n347), .B(n345), .Y(r_fcpwr[0]) );
  AND2X1 U277 ( .A(n339), .B(n348), .Y(r_dacwr[13]) );
  AND2X1 U278 ( .A(n337), .B(n349), .Y(we_228) );
  AND2X1 U279 ( .A(n305), .B(n349), .Y(we[164]) );
  AND2X1 U280 ( .A(n339), .B(n356), .Y(we_176) );
  AND2X1 U281 ( .A(n305), .B(n346), .Y(we[167]) );
  AND2X1 U282 ( .A(n305), .B(n351), .Y(we[165]) );
  AND2X1 U283 ( .A(n305), .B(n345), .Y(we[163]) );
  AND2X1 U284 ( .A(n305), .B(n338), .Y(we[162]) );
  AND2XL U285 ( .A(n305), .B(n340), .Y(we[161]) );
  AND2X1 U286 ( .A(n336), .B(n345), .Y(r_dacwr[10]) );
  AND2X1 U287 ( .A(n336), .B(n338), .Y(r_dacwr[9]) );
  AND2X1 U288 ( .A(n336), .B(n351), .Y(we_245) );
  AND2X1 U289 ( .A(n329), .B(n345), .Y(we_203) );
  AND2X1 U290 ( .A(n337), .B(n346), .Y(we_231) );
  INVX1 U291 ( .A(n308), .Y(n348) );
  NAND21X1 U292 ( .B(n312), .A(n343), .Y(n308) );
  NAND21X1 U293 ( .B(n309), .A(n301), .Y(n359) );
  INVX1 U294 ( .A(n270), .Y(n360) );
  INVX1 U295 ( .A(n321), .Y(n322) );
  INVX1 U296 ( .A(n310), .Y(n352) );
  NAND32XL U297 ( .B(n309), .C(n11), .A(n134), .Y(n310) );
  INVX1 U298 ( .A(n86), .Y(n311) );
  INVX1 U299 ( .A(ictlr_inc), .Y(n131) );
  INVX1 U300 ( .A(n111), .Y(n32) );
  INVX1 U301 ( .A(n111), .Y(n33) );
  INVX1 U302 ( .A(n110), .Y(n35) );
  INVX1 U303 ( .A(n111), .Y(n34) );
  INVX1 U304 ( .A(n110), .Y(n36) );
  INVX1 U305 ( .A(n110), .Y(n37) );
  INVX1 U306 ( .A(n108), .Y(n38) );
  INVX1 U307 ( .A(n108), .Y(n39) );
  INVX1 U308 ( .A(n108), .Y(n40) );
  INVX1 U309 ( .A(n112), .Y(n107) );
  INVX1 U310 ( .A(n113), .Y(n105) );
  INVX1 U311 ( .A(n203), .Y(n94) );
  INVX1 U312 ( .A(n112), .Y(n95) );
  INVX1 U313 ( .A(n113), .Y(n97) );
  INVX1 U314 ( .A(n203), .Y(n98) );
  INVX1 U315 ( .A(n203), .Y(n96) );
  INVX1 U316 ( .A(n112), .Y(n101) );
  NAND32X1 U317 ( .B(n316), .C(n299), .A(n328), .Y(n323) );
  NAND32X1 U318 ( .B(n292), .C(n328), .A(n295), .Y(n288) );
  INVX1 U319 ( .A(n294), .Y(n336) );
  NAND32XL U320 ( .B(n132), .C(n333), .A(n350), .Y(n294) );
  INVX1 U321 ( .A(n350), .Y(n312) );
  INVX1 U322 ( .A(n295), .Y(n316) );
  NAND21X1 U323 ( .B(n292), .A(n298), .Y(n357) );
  NAND21X1 U324 ( .B(n299), .A(n298), .Y(n83) );
  NAND32X1 U325 ( .B(n299), .C(n328), .A(n295), .Y(n361) );
  NAND32X1 U326 ( .B(n292), .C(n295), .A(n328), .Y(n289) );
  INVX1 U327 ( .A(n263), .Y(n358) );
  NAND32X1 U328 ( .B(n299), .C(n295), .A(n328), .Y(n263) );
  INVX1 U329 ( .A(n293), .Y(n339) );
  NAND32X1 U330 ( .B(n316), .C(n292), .A(n328), .Y(n293) );
  INVX1 U331 ( .A(n269), .Y(n298) );
  NAND21X1 U332 ( .B(n328), .A(n316), .Y(n269) );
  INVX1 U333 ( .A(n296), .Y(n332) );
  NAND21XL U334 ( .B(n350), .A(n11), .Y(n296) );
  INVX1 U335 ( .A(n326), .Y(r_fifopop) );
  NAND21X1 U336 ( .B(n138), .A(n376), .Y(phyrst) );
  NAND32X1 U337 ( .B(n303), .C(n306), .A(n350), .Y(n355) );
  AND3X1 U338 ( .A(n342), .B(n341), .C(n348), .Y(r_fcpre) );
  OA21X1 U339 ( .B(prx_rst[0]), .C(prx_rst[1]), .A(set03[1]), .Y(set03[7]) );
  INVX1 U340 ( .A(n200), .Y(n373) );
  INVX1 U341 ( .A(n264), .Y(n329) );
  NAND32XL U342 ( .B(n350), .C(n11), .A(n297), .Y(n264) );
  INVX1 U343 ( .A(n306), .Y(n309) );
  NAND4X1 U344 ( .A(n117), .B(n118), .C(n119), .D(n131), .Y(upd19) );
  INVX1 U345 ( .A(n197), .Y(n372) );
  INVX1 U346 ( .A(n307), .Y(n343) );
  NAND32XL U347 ( .B(n11), .C(n306), .A(n134), .Y(n307) );
  MUX2X1 U348 ( .D0(pff_rxpart[1]), .D1(n210), .S(n268), .Y(wd20[1]) );
  INVX1 U349 ( .A(n344), .Y(n347) );
  NAND21X1 U350 ( .B(n350), .A(n343), .Y(n344) );
  ENOX1 U351 ( .A(n100), .B(n259), .C(pff_rxpart[15]), .D(n100), .Y(wd21[7])
         );
  INVX1 U352 ( .A(n328), .Y(n341) );
  AND3X1 U353 ( .A(n352), .B(n351), .C(n14), .Y(r_cvcwr[1]) );
  AND3X1 U355 ( .A(n352), .B(n349), .C(n14), .Y(r_cvcwr[0]) );
  INVX1 U356 ( .A(n261), .Y(n337) );
  NAND32XL U357 ( .B(n266), .C(n132), .A(n350), .Y(n261) );
  INVX1 U358 ( .A(n116), .Y(n75) );
  NAND32XL U359 ( .B(n266), .C(n11), .A(n350), .Y(n270) );
  NAND21X1 U360 ( .B(n306), .A(n301), .Y(n321) );
  NAND32X1 U361 ( .B(n350), .C(n333), .A(n132), .Y(n86) );
  INVX1 U362 ( .A(n286), .Y(n301) );
  NAND21X1 U363 ( .B(n350), .A(n99), .Y(n286) );
  INVX1 U364 ( .A(n304), .Y(n305) );
  NAND32X1 U365 ( .B(n312), .C(n303), .A(n306), .Y(n304) );
  XOR2X1 U366 ( .A(N34), .B(N35), .Y(N36) );
  XNOR2XL U367 ( .A(n393), .B(N32), .Y(N38) );
  XNOR2XL U368 ( .A(N34), .B(n393), .Y(N37) );
  INVX1 U369 ( .A(N33), .Y(n393) );
  INVX1 U370 ( .A(n94), .Y(n113) );
  INVX1 U371 ( .A(n112), .Y(n111) );
  INVX1 U372 ( .A(n112), .Y(n110) );
  INVX1 U373 ( .A(n112), .Y(n108) );
  BUFX3 U374 ( .A(pff_empty), .Y(dbgpo[23]) );
  BUFX3 U375 ( .A(pff_full), .Y(dbgpo[22]) );
  NAND2X1 U376 ( .A(n317), .B(sfr_w), .Y(n292) );
  NAND21XL U377 ( .B(n317), .A(sfr_w), .Y(n299) );
  NAND21XL U378 ( .B(n262), .A(sfr_addr[4]), .Y(n306) );
  NAND21XL U379 ( .B(n262), .A(sfr_addr[2]), .Y(n317) );
  NAND21XL U380 ( .B(n262), .A(sfr_addr[3]), .Y(n350) );
  NAND21XL U381 ( .B(n262), .A(sfr_addr[0]), .Y(n328) );
  NAND21XL U382 ( .B(n262), .A(sfr_addr[1]), .Y(n295) );
  NOR2X1 U383 ( .A(n395), .B(n370), .Y(r_osc_lo) );
  INVX1 U384 ( .A(n171), .Y(bus_idle) );
  AND2X1 U385 ( .A(pff_ack[0]), .B(n18), .Y(set04[4]) );
  AND2X1 U386 ( .A(pff_ack[1]), .B(n369), .Y(set04[5]) );
  NAND5XL U387 ( .A(sfr_r), .B(n316), .C(n356), .D(n317), .E(n328), .Y(n326)
         );
  NAND41X1 U388 ( .D(n133), .A(n218), .B(n162), .C(n237), .Y(n119) );
  INVX1 U389 ( .A(n318), .Y(n342) );
  NAND32X1 U390 ( .B(n317), .C(n375), .A(n316), .Y(n318) );
  INVX1 U391 ( .A(sfr_r), .Y(n375) );
  NAND2X1 U392 ( .A(n394), .B(n119), .Y(n138) );
  AND2X1 U393 ( .A(n205), .B(n248), .Y(r_i2c_fwnak) );
  AOI21X1 U394 ( .B(n377), .C(n378), .A(n166), .Y(n200) );
  OAI33XL U395 ( .A(n197), .B(n198), .C(n390), .D(n378), .E(n377), .F(n373), 
        .Y(N113) );
  AND2X1 U396 ( .A(prx_setsta[2]), .B(n369), .Y(set03[2]) );
  AND2X1 U397 ( .A(prx_setsta[1]), .B(n369), .Y(set03[1]) );
  NAND2X1 U398 ( .A(n104), .B(n364), .Y(n103) );
  NAND2X1 U399 ( .A(n166), .B(n165), .Y(n197) );
  OAI22X1 U400 ( .A(n258), .B(n102), .C(n131), .D(n15), .Y(wd19[7]) );
  NAND2X1 U401 ( .A(n166), .B(n197), .Y(N108) );
  MUX2IX1 U402 ( .D0(n290), .D1(n258), .S(n362), .Y(wd01[7]) );
  NAND21X1 U403 ( .B(n380), .A(n327), .Y(n290) );
  AND2X1 U404 ( .A(n109), .B(n22), .Y(wd01[6]) );
  MUX2IX1 U405 ( .D0(n363), .D1(n253), .S(n362), .Y(n22) );
  NAND43X1 U406 ( .B(set_hold), .C(cpurst), .D(n364), .A(n104), .Y(upd12) );
  AO21X1 U407 ( .B(n326), .C(n327), .A(n363), .Y(n109) );
  MUX2X1 U408 ( .D0(pff_rxpart[0]), .D1(n172), .S(n268), .Y(wd20[0]) );
  MUX2X1 U409 ( .D0(pff_rxpart[2]), .D1(n216), .S(n268), .Y(wd20[2]) );
  MUX2X1 U410 ( .D0(pff_rxpart[3]), .D1(n223), .S(n268), .Y(wd20[3]) );
  MUX2X1 U411 ( .D0(pff_rxpart[6]), .D1(sfr_wdat[6]), .S(n268), .Y(wd20[6]) );
  MUX2X1 U412 ( .D0(pff_rxpart[7]), .D1(sfr_wdat[7]), .S(n268), .Y(wd20[7]) );
  MUX2X1 U413 ( .D0(pff_rxpart[4]), .D1(n235), .S(n268), .Y(wd20[4]) );
  NAND21X1 U414 ( .B(n268), .A(n114), .Y(upd20) );
  OAI21X1 U415 ( .B(n191), .C(n171), .A(n118), .Y(N26) );
  AND2X1 U416 ( .A(n121), .B(n397), .Y(n191) );
  NAND4X1 U417 ( .A(n135), .B(n213), .C(n192), .D(n193), .Y(n118) );
  NOR4XL U418 ( .A(n254), .B(n219), .C(n252), .D(n236), .Y(n193) );
  NOR21XL U419 ( .B(n162), .A(n128), .Y(n192) );
  ENOX1 U420 ( .A(n19), .B(n236), .C(pff_rxpart[12]), .D(n100), .Y(wd21[4]) );
  ENOX1 U421 ( .A(n19), .B(n212), .C(pff_rxpart[9]), .D(n100), .Y(wd21[1]) );
  ENOX1 U422 ( .A(n19), .B(n218), .C(pff_rxpart[10]), .D(n100), .Y(wd21[2]) );
  ENOX1 U423 ( .A(n19), .B(n253), .C(pff_rxpart[14]), .D(n100), .Y(wd21[6]) );
  ENOX1 U424 ( .A(n19), .B(n245), .C(pff_rxpart[13]), .D(n100), .Y(wd21[5]) );
  ENOX1 U425 ( .A(n19), .B(n229), .C(pff_rxpart[11]), .D(n100), .Y(wd21[3]) );
  ENOX1 U426 ( .A(n212), .B(n102), .C(inst_ofs_plus[9]), .D(n130), .Y(wd19[1])
         );
  ENOX1 U427 ( .A(n218), .B(n102), .C(inst_ofs_plus[10]), .D(n130), .Y(wd19[2]) );
  ENOX1 U428 ( .A(n176), .B(n102), .C(inst_ofs_plus[8]), .D(n130), .Y(wd19[0])
         );
  ENOX1 U429 ( .A(n229), .B(n102), .C(inst_ofs_plus[11]), .D(ictlr_inc), .Y(
        wd19[3]) );
  ENOX1 U430 ( .A(n236), .B(n102), .C(inst_ofs_plus[12]), .D(ictlr_inc), .Y(
        wd19[4]) );
  ENOX1 U431 ( .A(n246), .B(n102), .C(inst_ofs_plus[13]), .D(ictlr_inc), .Y(
        wd19[5]) );
  AO22AXL U432 ( .A(r_pshords), .B(n103), .C(sfr_wdat[0]), .D(n103), .Y(
        wd12[0]) );
  OAI211X1 U433 ( .C(n380), .D(n327), .A(n109), .B(n291), .Y(upd01) );
  NAND2X1 U434 ( .A(n114), .B(n19), .Y(upd21) );
  AND2X1 U435 ( .A(pff_obsd), .B(n369), .Y(set04[3]) );
  AND2X1 U436 ( .A(prx_setsta[4]), .B(n18), .Y(set03[4]) );
  AND4X1 U437 ( .A(n329), .B(n342), .C(n328), .D(n15), .Y(upd31) );
  NAND2X1 U438 ( .A(prx_setsta[3]), .B(n369), .Y(n116) );
  ENOX1 U439 ( .A(n125), .B(n236), .C(inst_ofs_plus[4]), .D(n125), .Y(wd18[4])
         );
  ENOX1 U440 ( .A(n125), .B(n253), .C(inst_ofs_plus[6]), .D(n130), .Y(wd18[6])
         );
  ENOX1 U441 ( .A(n125), .B(n259), .C(inst_ofs_plus[7]), .D(n130), .Y(wd18[7])
         );
  ENOX1 U442 ( .A(n125), .B(n229), .C(inst_ofs_plus[3]), .D(n130), .Y(wd18[3])
         );
  ENOX1 U443 ( .A(n125), .B(n246), .C(inst_ofs_plus[5]), .D(n130), .Y(wd18[5])
         );
  ENOX1 U444 ( .A(n125), .B(n212), .C(inst_ofs_plus[1]), .D(n130), .Y(wd18[1])
         );
  ENOX1 U445 ( .A(n125), .B(n218), .C(inst_ofs_plus[2]), .D(n130), .Y(wd18[2])
         );
  AND2X1 U446 ( .A(i_gobusy), .B(n18), .Y(set04[2]) );
  XNOR2XL U447 ( .A(n397), .B(add_180_carry[4]), .Y(N35) );
  AND2X1 U448 ( .A(prl_GCTxDone), .B(n18), .Y(set04[6]) );
  XNOR2XL U449 ( .A(N30), .B(N32), .Y(N39) );
  NOR2X1 U450 ( .A(n18), .B(i_goidle), .Y(n164) );
  AND2X1 U451 ( .A(prl_discard), .B(n369), .Y(set04[7]) );
  NAND2X1 U452 ( .A(n198), .B(n390), .Y(n165) );
  INVX1 U453 ( .A(n201), .Y(n391) );
  INVX1 U454 ( .A(n202), .Y(n392) );
  NAND2X1 U455 ( .A(n126), .B(n370), .Y(N84) );
  XNOR2XL U456 ( .A(di_p0[5]), .B(n383), .Y(n187) );
  XNOR2XL U457 ( .A(di_p0[3]), .B(n385), .Y(n185) );
  XNOR2XL U458 ( .A(di_p0[7]), .B(n382), .Y(n189) );
  XNOR2XL U459 ( .A(di_p0[2]), .B(n387), .Y(n186) );
  XNOR2XL U460 ( .A(di_p0[4]), .B(n384), .Y(n188) );
  XNOR2XL U461 ( .A(di_p0[6]), .B(n381), .Y(n190) );
  NAND2X1 U462 ( .A(n260), .B(aswkup), .Y(pwrdn_rstz) );
  AND2X1 U463 ( .A(dnchk_en), .B(dm_fault), .Y(dmf_wkup) );
  INVX1 U464 ( .A(n120), .Y(n112) );
  INVX1 U465 ( .A(n203), .Y(n120) );
  INVX1 U466 ( .A(n203), .Y(n115) );
  MUX2XL U467 ( .D0(i_pc[2]), .D1(prx_adpn[2]), .S(n16), .Y(reg30[2]) );
  MUX2XL U468 ( .D0(i_pc[0]), .D1(prx_adpn[0]), .S(reg19_7_), .Y(reg30[0]) );
  MUX2X1 U469 ( .D0(s_ovp), .D1(m_ovp), .S(reg94[4]), .Y(regAD[2]) );
  AND3X1 U470 ( .A(n9), .B(n219), .C(n367), .Y(ps_pwrdn) );
  NAND32X1 U471 ( .B(bkpt_hold), .C(reg12[3]), .A(n126), .Y(r_hold_mcu) );
  NAND21X1 U472 ( .B(lg_dischg), .A(n331), .Y(r_srcctl[1]) );
  INVX1 U473 ( .A(lg_pulse_12m), .Y(n331) );
  NOR2X1 U474 ( .A(regD4_2_), .B(regD4_0_), .Y(n126) );
  AOI222XL U475 ( .A(reg28[7]), .B(reg27[7]), .C(reg28[4]), .D(reg27[4]), .E(
        reg28[6]), .F(reg27[6]), .Y(n169) );
  NAND3X1 U476 ( .A(n167), .B(n168), .C(n169), .Y(i2c_stretch) );
  AOI22X1 U477 ( .A(reg28[2]), .B(reg27[2]), .C(reg28[3]), .D(reg27[3]), .Y(
        n167) );
  AOI22X1 U478 ( .A(reg28[0]), .B(reg27[0]), .C(reg28[1]), .D(reg27[1]), .Y(
        n168) );
  MUX2XL U479 ( .D0(i_pc[3]), .D1(prx_adpn[3]), .S(n16), .Y(reg30[3]) );
  NOR21XL U480 ( .B(regD4_0_), .A(n395), .Y(r_osc_stop) );
  INVX1 U481 ( .A(oscdwn_shft[2]), .Y(n395) );
  INVX1 U482 ( .A(regD4_1_), .Y(n370) );
  INVX1 U483 ( .A(n354), .Y(n367) );
  OAI211X1 U484 ( .C(ictlr_idle), .D(n353), .A(oscdwn_shft[1]), .B(bus_idle), 
        .Y(n354) );
  AND2X1 U485 ( .A(regD4_1_), .B(n126), .Y(n353) );
  MUX2X1 U486 ( .D0(s_scp), .D1(m_scp), .S(reg94[5]), .Y(regAD[4]) );
  AOI21X1 U487 ( .B(n137), .C(drstz[1]), .A(atpg_en), .Y(n20) );
  OAI211X1 U488 ( .C(rstcnt[2]), .D(rstcnt[1]), .A(n396), .B(rstcnt[4]), .Y(
        n137) );
  INVX1 U489 ( .A(rstcnt[3]), .Y(n396) );
  NAND41X1 U490 ( .D(prl_cany0), .A(prx_rcvinf[4]), .B(i_i2c_idle), .C(n196), 
        .Y(n171) );
  MUX2X1 U491 ( .D0(i_pc[5]), .D1(prx_adpn[5]), .S(n16), .Y(reg30[5]) );
  MUX2XL U492 ( .D0(i_pc[4]), .D1(prx_adpn[4]), .S(n16), .Y(reg30[4]) );
  INVX1 U493 ( .A(regD3_7_), .Y(r_gpio_ie[1]) );
  AND2X1 U494 ( .A(i_pc[7]), .B(n15), .Y(reg30[7]) );
  NAND4X1 U495 ( .A(n151), .B(n152), .C(n153), .D(n154), .Y(o_intr[1]) );
  AOI22X1 U496 ( .A(reg06[6]), .B(irq04[6]), .C(reg06[7]), .D(irq04[7]), .Y(
        n151) );
  AOI22X1 U497 ( .A(reg06[0]), .B(irq04[0]), .C(reg06[1]), .D(irq04[1]), .Y(
        n154) );
  AOI22X1 U498 ( .A(reg06[4]), .B(irq04[4]), .C(reg06[5]), .D(irq04[5]), .Y(
        n152) );
  OR4X1 U499 ( .A(osc_gate_n_1_), .B(osc_gate_n_0_), .C(test_so1), .D(
        osc_gate_n_2_), .Y(r_osc_gate) );
  NOR21XL U500 ( .B(regD4_2_), .A(n395), .Y(r_pos_gate) );
  AND3X1 U501 ( .A(n16), .B(n346), .C(n329), .Y(r_pswr) );
  AND2X1 U502 ( .A(regE3[2]), .B(n122), .Y(r_srcctl[2]) );
  AND2X1 U503 ( .A(regE3[3]), .B(n122), .Y(r_srcctl[3]) );
  AND4X1 U504 ( .A(n16), .B(n342), .C(n329), .D(n341), .Y(r_psrd) );
  AOI22X1 U505 ( .A(regAF[5]), .B(regAE[5]), .C(regAD[5]), .D(i_vcbyval), .Y(
        n122) );
  OAI32X1 U506 ( .A(n389), .B(r_phyrst[1]), .C(n379), .D(r_phyrst[0]), .E(n161), .Y(n1221) );
  INVX1 U507 ( .A(n164), .Y(n379) );
  AOI21X1 U508 ( .B(reg11_7_), .C(set03[7]), .A(n138), .Y(n161) );
  NOR21XL U509 ( .B(regE3_0), .A(gating_pwr), .Y(r_srcctl[0]) );
  NOR21XL U510 ( .B(regD4_3_), .A(n395), .Y(r_pwrdn) );
  AOI21X1 U511 ( .B(n207), .C(n206), .A(lg_pulse_12m), .Y(n166) );
  AND2X1 U512 ( .A(reg94[7]), .B(reg94[6]), .Y(r_otpi_gate) );
  AO22X1 U513 ( .A(regAF[4]), .B(regAE[4]), .C(regAF[2]), .D(regAE[2]), .Y(
        gating_pwr) );
  GEN2XL U514 ( .D(lg_pulse_cnt[2]), .E(n392), .C(n201), .B(n372), .A(n200), 
        .Y(N111) );
  NOR21XL U515 ( .B(regD4_4_), .A(n395), .Y(r_ocdrv_enz) );
  NAND4X1 U516 ( .A(n155), .B(n156), .C(n157), .D(n158), .Y(o_intr[0]) );
  AOI22X1 U517 ( .A(reg05[4]), .B(irq03[4]), .C(reg05[5]), .D(irq03[5]), .Y(
        n156) );
  AOI22X1 U518 ( .A(reg05[2]), .B(irq03[2]), .C(reg05[3]), .D(irq03[3]), .Y(
        n157) );
  AOI22X1 U519 ( .A(reg05[0]), .B(irq03[0]), .C(reg05[1]), .D(irq03[1]), .Y(
        n158) );
  AOI22X1 U520 ( .A(reg05[6]), .B(irq03[6]), .C(reg05[7]), .D(irq03[7]), .Y(
        n155) );
  OAI22X1 U521 ( .A(n199), .B(n197), .C(n377), .D(n373), .Y(N112) );
  AOI21X1 U522 ( .B(lg_pulse_cnt[3]), .C(n391), .A(n198), .Y(n199) );
  GEN2XL U523 ( .D(lg_pulse_cnt[1]), .E(lg_pulse_cnt[0]), .C(n202), .B(n372), 
        .A(n371), .Y(N110) );
  INVX1 U524 ( .A(n166), .Y(n371) );
  ENOX1 U525 ( .A(n176), .B(n374), .C(n374), .D(lt_reg26_0), .Y(i2c_mode_wdat)
         );
  AOI21X1 U526 ( .B(n170), .C(n374), .A(n171), .Y(i2c_mode_upd) );
  XNOR2XL U527 ( .A(r_hwi2c_en), .B(lt_reg26_0), .Y(n170) );
  OAI21BBX1 U528 ( .A(n165), .B(lg_dischg), .C(n166), .Y(n1219) );
  OAI21X1 U529 ( .B(lg_pulse_cnt[0]), .C(n197), .A(n166), .Y(N109) );
  OAI21BX1 U530 ( .C(reg12[3]), .B(n104), .A(n106), .Y(wd12[3]) );
  AOI32X1 U531 ( .A(set_hold), .B(n104), .C(n366), .D(n219), .E(n365), .Y(n106) );
  INVX1 U532 ( .A(n103), .Y(n365) );
  MUX2XL U533 ( .D0(r_txnumk[2]), .D1(n216), .S(n362), .Y(wd01[2]) );
  MUX2XL U534 ( .D0(r_txnumk[0]), .D1(n172), .S(n362), .Y(wd01[0]) );
  MUX2XL U535 ( .D0(r_txnumk[1]), .D1(n210), .S(n362), .Y(wd01[1]) );
  MUX2XL U536 ( .D0(r_txnumk[3]), .D1(n223), .S(n362), .Y(wd01[3]) );
  MUX2XL U537 ( .D0(r_txnumk[4]), .D1(n235), .S(n362), .Y(wd01[4]) );
  MUX2X1 U538 ( .D0(r_unlock), .D1(n241), .S(n362), .Y(wd01[5]) );
  NAND2X1 U539 ( .A(n23), .B(n104), .Y(wd12[4]) );
  MUX2IX1 U540 ( .D0(reg12[4]), .D1(n234), .S(n364), .Y(n23) );
  OAI22X1 U541 ( .A(n212), .B(n330), .C(lg_dischg), .D(n331), .Y(n1218) );
  ENOX1 U542 ( .A(n19), .B(n176), .C(pff_rxpart[8]), .D(n100), .Y(wd21[0]) );
  ENOX1 U543 ( .A(n252), .B(n102), .C(inst_ofs_plus[14]), .D(ictlr_inc), .Y(
        wd19[6]) );
  ENOX1 U544 ( .A(n252), .B(n103), .C(reg12[6]), .D(n103), .Y(wd12[6]) );
  ENOX1 U545 ( .A(n259), .B(n103), .C(reg12[7]), .D(n103), .Y(wd12[7]) );
  ENOX1 U546 ( .A(n212), .B(n17), .C(reg12_1), .D(n103), .Y(wd12[1]) );
  ENOX1 U547 ( .A(n218), .B(n17), .C(r_txshrt), .D(n103), .Y(wd12[2]) );
  ENOX1 U548 ( .A(n246), .B(n17), .C(reg12[5]), .D(n103), .Y(wd12[5]) );
  AOI22X1 U549 ( .A(reg06[2]), .B(irq04[2]), .C(reg06[3]), .D(irq04[3]), .Y(
        n153) );
  NOR21XL U550 ( .B(prx_setsta[6]), .A(prl_cany0), .Y(set03[6]) );
  AND2X1 U551 ( .A(i_pc[6]), .B(n15), .Y(reg30[6]) );
  AOI21BBXL U552 ( .B(r_auto_gdcrc[1]), .C(n116), .A(set03[6]), .Y(n114) );
  AO21X1 U553 ( .B(n123), .C(n124), .A(reg11_4), .Y(r_rxords_ena[4]) );
  NOR3XL U554 ( .A(r_rxords_ena[0]), .B(r_rxords_ena[2]), .C(r_rxords_ena[1]), 
        .Y(n123) );
  NOR3XL U555 ( .A(r_rxords_ena[3]), .B(r_rxords_ena[6]), .C(r_rxords_ena[5]), 
        .Y(n124) );
  ENOX1 U556 ( .A(n125), .B(n176), .C(inst_ofs_plus[0]), .D(n130), .Y(wd18[0])
         );
  INVX1 U557 ( .A(regD3_3), .Y(r_gpio_ie[0]) );
  INVX1 U558 ( .A(r_phyrst[1]), .Y(n394) );
  INVX1 U559 ( .A(n136), .Y(prstz) );
  AOI31X1 U560 ( .A(drstz[1]), .B(n394), .C(n137), .D(atpg_en), .Y(n136) );
  AOI22X1 U561 ( .A(reg27[6]), .B(irq28[6]), .C(reg27[7]), .D(irq28[7]), .Y(
        n147) );
  AND2X1 U562 ( .A(prx_setsta[5]), .B(n369), .Y(set03[5]) );
  NAND4X1 U563 ( .A(n147), .B(n148), .C(n149), .D(n150), .Y(o_intr[2]) );
  AOI22X1 U564 ( .A(reg27[4]), .B(irq28[4]), .C(reg27[5]), .D(irq28[5]), .Y(
        n148) );
  AOI22X1 U565 ( .A(reg27[0]), .B(irq28[0]), .C(reg27[1]), .D(irq28[1]), .Y(
        n150) );
  NOR21XL U566 ( .B(i_goidle), .A(prl_cany0), .Y(set04[1]) );
  XOR2X1 U567 ( .A(N27), .B(rstcnt[2]), .Y(N28) );
  XOR2X1 U568 ( .A(N28), .B(rstcnt[1]), .Y(N29) );
  AND2X1 U569 ( .A(ptx_ack), .B(n369), .Y(set04[0]) );
  XOR2X1 U570 ( .A(N29), .B(rstcnt[0]), .Y(N30) );
  XNOR2XL U571 ( .A(n397), .B(rstcnt[3]), .Y(N27) );
  INVX1 U572 ( .A(rstcnt[4]), .Y(n397) );
  AO22AXL U573 ( .A(reg94[5]), .B(m_scp_sta), .C(s_scp_sta), .D(reg94[5]), .Y(
        setAE[4]) );
  NAND4X1 U574 ( .A(n139), .B(n140), .C(n141), .D(n142), .Y(o_intr[4]) );
  AOI22X1 U575 ( .A(regAF[6]), .B(irqAE[6]), .C(regAF[7]), .D(irqAE[7]), .Y(
        n139) );
  AOI22X1 U576 ( .A(regAF[0]), .B(irqAE[0]), .C(regAF[1]), .D(irqAE[1]), .Y(
        n142) );
  AOI22X1 U577 ( .A(reg27[2]), .B(irq28[2]), .C(reg27[3]), .D(irq28[3]), .Y(
        n149) );
  AOI22X1 U578 ( .A(irqAE[4]), .B(regAF[4]), .C(irqAE[5]), .D(regAF[5]), .Y(
        n140) );
  XNOR2XL U579 ( .A(d_p0[0]), .B(n386), .Y(setDF[0]) );
  XNOR2XL U580 ( .A(d_p0[1]), .B(n388), .Y(setDF[1]) );
  XNOR2XL U581 ( .A(d_p0[2]), .B(n387), .Y(setDF[2]) );
  XNOR2XL U582 ( .A(d_p0[3]), .B(n385), .Y(setDF[3]) );
  XNOR2XL U583 ( .A(d_p0[4]), .B(n384), .Y(setDF[4]) );
  AO22AXL U584 ( .A(reg94[4]), .B(m_ovp_sta), .C(s_ovp_sta), .D(reg94[4]), .Y(
        setAE[2]) );
  XNOR2XL U585 ( .A(d_p0[5]), .B(n383), .Y(setDF[5]) );
  INVX1 U586 ( .A(prl_cany0), .Y(n369) );
  AND2X1 U587 ( .A(prx_setsta[0]), .B(n369), .Y(set03[0]) );
  NAND2X1 U588 ( .A(rstcnt[4]), .B(n121), .Y(n104) );
  INVX1 U589 ( .A(reg25_0_), .Y(r_i2c_ninc) );
  NOR4XL U590 ( .A(rstcnt[0]), .B(rstcnt[1]), .C(rstcnt[2]), .D(rstcnt[3]), 
        .Y(n121) );
  NOR42XL U591 ( .C(n194), .D(r_inst_ofs[10]), .A(r_inst_ofs[8]), .B(n195), 
        .Y(n162) );
  NAND4X1 U592 ( .A(r_inst_ofs[14]), .B(r_inst_ofs[13]), .C(r_inst_ofs[12]), 
        .D(r_inst_ofs[11]), .Y(n195) );
  NOR2X1 U593 ( .A(n16), .B(r_inst_ofs[9]), .Y(n194) );
  AOI22X1 U594 ( .A(regDE[0]), .B(irqDF[0]), .C(regDE[1]), .D(irqDF[1]), .Y(
        n146) );
  AOI22X1 U595 ( .A(regDE[2]), .B(irqDF[2]), .C(regDE[3]), .D(irqDF[3]), .Y(
        n145) );
  AOI22X1 U596 ( .A(irqAE[2]), .B(regAF[2]), .C(regAF[3]), .D(irqAE[3]), .Y(
        n141) );
  OAI32X1 U597 ( .A(n389), .B(r_phyrst[1]), .C(n164), .D(r_phyrst[0]), .E(n394), .Y(n1220) );
  XNOR2XL U598 ( .A(d_p0[6]), .B(n381), .Y(setDF[6]) );
  XNOR2XL U599 ( .A(d_p0[7]), .B(n382), .Y(setDF[7]) );
  INVX1 U600 ( .A(ff_p0[0]), .Y(n386) );
  INVX1 U601 ( .A(ff_p0[2]), .Y(n387) );
  INVX1 U602 ( .A(ff_p0[1]), .Y(n388) );
  INVX1 U603 ( .A(ff_p0[3]), .Y(n385) );
  INVX1 U604 ( .A(ff_p0[5]), .Y(n383) );
  INVX1 U605 ( .A(ff_p0[4]), .Y(n384) );
  INVX1 U606 ( .A(ff_p0[7]), .Y(n382) );
  INVX1 U607 ( .A(ff_p0[6]), .Y(n381) );
  NAND4X1 U608 ( .A(n143), .B(n144), .C(n145), .D(n146), .Y(o_intr[3]) );
  AOI22X1 U609 ( .A(regDE[6]), .B(irqDF[6]), .C(regDE[7]), .D(irqDF[7]), .Y(
        n143) );
  AOI22X1 U610 ( .A(regDE[4]), .B(irqDF[4]), .C(regDE[5]), .D(irqDF[5]), .Y(
        n144) );
  NOR2X1 U611 ( .A(n392), .B(lg_pulse_cnt[2]), .Y(n201) );
  NOR2X1 U612 ( .A(lg_pulse_cnt[1]), .B(lg_pulse_cnt[0]), .Y(n202) );
  NOR2X1 U613 ( .A(n391), .B(lg_pulse_cnt[3]), .Y(n198) );
  INVX1 U614 ( .A(lg_pulse_cnt[4]), .Y(n390) );
  INVX1 U615 ( .A(lg_pulse_len[1]), .Y(n377) );
  INVX1 U616 ( .A(r_first), .Y(n363) );
  INVX1 U617 ( .A(lg_pulse_len[0]), .Y(n378) );
  INVX1 U618 ( .A(r_last), .Y(n380) );
  INVX1 U619 ( .A(r_phyrst[0]), .Y(n389) );
  NAND42X1 U620 ( .C(di_rd_det_clr), .D(dm_fault_clr), .A(n92), .B(n178), .Y(
        aswkup) );
  NOR2X1 U621 ( .A(p0_chg_clr), .B(i_tmrf), .Y(n178) );
  NOR21XL U622 ( .B(n3), .A(n20), .Y(n203) );
  OAI21BX1 U623 ( .C(n203), .B(osc_low_clr), .A(n260), .Y(osc_low_rstz) );
  AOI22X1 U624 ( .A(regDE[1]), .B(n183), .C(regDE[0]), .D(n184), .Y(n182) );
  XNOR2XL U625 ( .A(di_p0[0]), .B(n386), .Y(n184) );
  XNOR2XL U626 ( .A(di_p0[1]), .B(n388), .Y(n183) );
  NAND4X1 U627 ( .A(n179), .B(n180), .C(n181), .D(n182), .Y(as_p0_chg) );
  AOI22X1 U628 ( .A(regDE[7]), .B(n189), .C(regDE[6]), .D(n190), .Y(n179) );
  AOI22X1 U629 ( .A(regDE[5]), .B(n187), .C(regDE[4]), .D(n188), .Y(n180) );
  AOI22X1 U630 ( .A(regDE[3]), .B(n185), .C(regDE[2]), .D(n186), .Y(n181) );
  INVX1 U631 ( .A(sfr_addr[7]), .Y(n262) );
  NOR4XL U632 ( .A(prl_fsm[3]), .B(prl_fsm[2]), .C(prl_fsm[1]), .D(prl_fsm[0]), 
        .Y(n196) );
  INVXL U633 ( .A(n12), .Y(n134) );
  NOR2XL U634 ( .A(n132), .B(n12), .Y(n99) );
  NAND21XL U635 ( .B(n309), .A(n12), .Y(n266) );
  NAND21XL U636 ( .B(n306), .A(n12), .Y(n333) );
endmodule


module regbank_a0_DW_rightsh_2 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n131, n132, n133, n134, n135,
         n136, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n195, n196, n197, n198, n199, n200, n201, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n219, n220, n221, n222, n223, n224, n225, n227, n228, n229,
         n230, n231, n232, n235, n236, n237, n238, n239, n240, n307, n312,
         n314, n315, n316, n317, n318, n491, n492, n497, n498, n503, n504,
         n509, n510, n515, n516, n521, n527, n533, n534, n539, n540, n545,
         n546, n551, n552, n557, n558, n563, n564, n569, n576, n585, n586,
         n589, n590, n593, n594, n597, n598, n601, n602, n605, n606, n609,
         n610, n613, n614, n617, n618, n621, n622, n625, n626, n629, n630,
         n633, n634, n637, n638, n641, n642, n645, n646, n649, n650, n653,
         n654, n657, n658, n661, n662, n665, n666, n669, n670, n673, n674,
         n677, n678, n681, n684, n687, n690, n693, n696, n699, n702, n705,
         n706, n709, n710, n713, n714, n717, n718, n721, n722, n725, n726,
         n729, n730, n733, n734, n737, n740, n743, n746, n749, n752, n755,
         n758, n761, n762, n765, n766, n769, n770, n773, n774, n777, n778,
         n785, n786, n796, n802, n808, n813, n814, n819, n820, n825, n837,
         n843, n844, n849, n850, n855, n856, n862, n868, n873, n879, n880,
         n886, n891, n892, n897, n898, n903, n904, n909, n910, n915, n916,
         n922, n928, n933, n937, n938, n941, n942, n945, n946, n949, n950,
         n953, n954, n957, n958, n961, n962, n965, n966, n969, n970, n973,
         n974, n977, n978, n981, n982, n985, n986, n989, n990, n993, n994,
         n997, n998, n1004, n1010, n1016, n1022, n1028, n1033, n1034, n1040,
         n1045, n1049, n1050, n1053, n1054, n1057, n1058, n1061, n1062, n1065,
         n1066, n1069, n1070, n1073, n1074, n1077, n1078, n1081, n1082, n1085,
         n1086, n1089, n1090, n1093, n1094, n1097, n1098, n1105, n1106, n1113,
         n1114, n1117, n1118, n1121, n1122, n1125, n1126, n1129, n1130, n1133,
         n1134, n1137, n1138, n1141, n1142, n1145, n1146, n1149, n1153, n1154,
         n1157, n1158, n1161, n1162, n1165, n1166, n1169, n1170, n1173, n1174,
         n1177, n1178, n1181, n1182, n1185, n1186, n1189, n1190, n1193, n1194,
         n1197, n1198, n1201, n1202, n1205, n1206, n1209, n1210, n1213, n1214,
         n1217, n1218, n1221, n1222, n1225, n1226, n1229, n1230, n1233, n1234,
         n1237, n1238, n1241, n1244, n1247, n1250, n1253, n1256, n1259, n1262,
         n1269, n1272, n1275, n1278, n1281, n1284, n1287, n1290, n1293, n1296,
         n1299, n1302, n1305, n1308, n1311, n1312, n1315, n1316, n1319, n1320,
         n1323, n1324, n1327, n1328, n1331, n1335, n1336, n1339, n1340, n1343,
         n1344, n1347, n1348, n1351, n1352, n1355, n1356, n1359, n1360, n1363,
         n1364, n1367, n1368, n1371, n1372, n1378, n1383, n1384, n1390, n1396,
         n1402, n1408, n1426, n1431, n1432, n1438, n1444, n1450, n1468, n1471,
         n1472, n1475, n1476, n1479, n1480, n1483, n1484, n1487, n1488, n1491,
         n1492, n1495, n1496, n1499, n1500, n1503, n1504, n1507, n1508, n1511,
         n1512, n1515, n1516, n1519, n1520, n1523, n1527, n1528, n1531, n1535,
         n1536, n1539, n1540, n1543, n1544, n1547, n1548, n1551, n1552, n1555,
         n1556, n1559, n1560, n1563, n1564, n1583, n1586, n1587, n1588, n1590,
         n1599, n1602, n1603, n1604, n1606, n1608, n1610, n1611, n1612, n1614,
         n1615, n1616, n1618, n1619, n1620, n1622, n1624, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1634, n1635, n1636, n1638, n1641, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1666,
         n1667, n1668, n1669, n1671, n1673, n1674, n1675, n1676, n1678, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1689, n1690, n1691,
         n1692, n1694, n1696, n1697, n1698, n1699, n1700, n1702, n1703, n1705,
         n1706, n1707, n1708, n1709, n1710, n1713, n1714, n1715, n1716, n1717,
         n1718, n1721, n1722, n1723, n1724, n1725, n1726, n1729, n1730, n1731,
         n1732, n1733, n1734, n1740, n1741, n1742, n1746, n1747, n1756, n1757,
         n1758, n1761, n1762, n1763, n1776, n1778, n1779, n1780, n1781, n1782,
         n1792, n1794, n1795, n1796, n1797, n1798, n1799, n1802, n1803, n1804,
         n1805, n1806, n1807, n1810, n1811, n1812, n1813, n1814, n1818, n1819,
         n1820, n1821, n1822, n1823, n1826, n1827, n1828, n1829, n1830, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079;

  AO22X1 U500 ( .A(n4013), .B(n491), .C(n492), .D(n3996), .Y(n1830) );
  AO22X1 U510 ( .A(n4009), .B(n497), .C(n498), .D(n3996), .Y(n1829) );
  AO22X1 U514 ( .A(n3777), .B(A[510]), .C(n3824), .D(A[1022]), .Y(n498) );
  AO22X1 U520 ( .A(n4011), .B(n503), .C(n504), .D(n3996), .Y(n1828) );
  AO22X1 U530 ( .A(n4009), .B(n509), .C(n510), .D(n3996), .Y(n1827) );
  AO22X1 U534 ( .A(n3777), .B(A[508]), .C(n3824), .D(A[1020]), .Y(n510) );
  AO22X1 U540 ( .A(n4006), .B(n515), .C(n516), .D(n3996), .Y(n1826) );
  AO22X1 U555 ( .A(n4061), .B(A[250]), .C(n4029), .D(A[762]), .Y(n521) );
  AO22X1 U570 ( .A(n4010), .B(n533), .C(n534), .D(n3996), .Y(n1823) );
  AO22X1 U574 ( .A(n4061), .B(A[504]), .C(n3684), .D(A[1016]), .Y(n534) );
  AO22X1 U575 ( .A(n4061), .B(A[248]), .C(n4041), .D(A[760]), .Y(n533) );
  AO22X1 U580 ( .A(n4005), .B(n539), .C(n540), .D(n3995), .Y(n1822) );
  AO22X1 U590 ( .A(n4010), .B(n545), .C(n546), .D(n3995), .Y(n1821) );
  AO22X1 U600 ( .A(n4011), .B(n551), .C(n552), .D(n3995), .Y(n1820) );
  AO22X1 U610 ( .A(n4010), .B(n557), .C(n558), .D(n3995), .Y(n1819) );
  AO22X1 U614 ( .A(n4062), .B(A[500]), .C(n3766), .D(A[1012]), .Y(n558) );
  AO22X1 U620 ( .A(n4012), .B(n563), .C(n564), .D(n3995), .Y(n1818) );
  NOR2X1 U664 ( .A(n3833), .B(A[239]), .Y(n585) );
  NOR2X1 U672 ( .A(n3833), .B(A[238]), .Y(n589) );
  NOR2X1 U680 ( .A(n4032), .B(A[237]), .Y(n593) );
  NOR2X1 U688 ( .A(n4050), .B(A[236]), .Y(n597) );
  NOR2X1 U696 ( .A(n3801), .B(A[235]), .Y(n601) );
  NOR2X1 U720 ( .A(n4032), .B(A[232]), .Y(n613) );
  NOR2X1 U728 ( .A(n4050), .B(A[231]), .Y(n617) );
  NOR2X1 U736 ( .A(n4075), .B(A[230]), .Y(n621) );
  NOR2X1 U744 ( .A(n3769), .B(A[229]), .Y(n625) );
  NOR2X1 U752 ( .A(n3821), .B(A[228]), .Y(n629) );
  NOR2X1 U760 ( .A(n4075), .B(A[227]), .Y(n633) );
  NOR2X1 U768 ( .A(n4049), .B(A[226]), .Y(n637) );
  NOR2X1 U776 ( .A(n4037), .B(A[225]), .Y(n641) );
  NOR2X1 U792 ( .A(n3781), .B(A[223]), .Y(n649) );
  NOR2X1 U800 ( .A(n3833), .B(A[222]), .Y(n653) );
  NOR2X1 U808 ( .A(n3820), .B(A[221]), .Y(n657) );
  NOR2X1 U816 ( .A(n3821), .B(A[220]), .Y(n661) );
  NOR2X1 U824 ( .A(n3768), .B(A[219]), .Y(n665) );
  NOR2X1 U840 ( .A(n4027), .B(A[217]), .Y(n673) );
  NOR2X1 U1031 ( .A(n3721), .B(A[447]), .Y(n762) );
  NOR2X1 U1039 ( .A(n3805), .B(A[446]), .Y(n766) );
  NOR2X1 U1047 ( .A(n3805), .B(A[445]), .Y(n770) );
  NOR2X1 U1055 ( .A(n3766), .B(A[444]), .Y(n774) );
  NOR2X1 U1063 ( .A(n4050), .B(A[443]), .Y(n778) );
  AO22X1 U1096 ( .A(n3710), .B(A[439]), .C(n3766), .D(A[951]), .Y(n796) );
  AO22X1 U1106 ( .A(n4063), .B(A[438]), .C(n3820), .D(A[950]), .Y(n802) );
  AO22X1 U1116 ( .A(n3710), .B(A[437]), .C(n3820), .D(A[949]), .Y(n808) );
  AO22X1 U1127 ( .A(n4063), .B(A[180]), .C(n3820), .D(A[692]), .Y(n813) );
  AO22X1 U1136 ( .A(n3710), .B(A[435]), .C(n3820), .D(A[947]), .Y(n820) );
  AO22X1 U1167 ( .A(n4064), .B(A[176]), .C(n3830), .D(A[688]), .Y(n837) );
  AO22X1 U1246 ( .A(n4065), .B(A[424]), .C(n3683), .D(A[936]), .Y(n886) );
  AO22X1 U1262 ( .A(n4006), .B(n897), .C(n898), .D(n3992), .Y(n1741) );
  AO22X1 U1272 ( .A(n4014), .B(n903), .C(n904), .D(n3991), .Y(n1740) );
  AO22X1 U1287 ( .A(n4068), .B(A[164]), .C(n3820), .D(A[676]), .Y(n909) );
  AO22X1 U1327 ( .A(n4072), .B(A[160]), .C(n4043), .D(A[672]), .Y(n933) );
  AO22X1 U1464 ( .A(n3710), .B(A[399]), .C(n4050), .D(A[911]), .Y(n1004) );
  AO22X1 U1474 ( .A(n3823), .B(A[398]), .C(n4050), .D(A[910]), .Y(n1010) );
  AO22X1 U1510 ( .A(n4006), .B(n1033), .C(n1034), .D(n3991), .Y(n1713) );
  AO22X1 U1514 ( .A(n4068), .B(A[394]), .C(n3782), .D(A[906]), .Y(n1034) );
  AO22X1 U1535 ( .A(n4066), .B(A[136]), .C(n3830), .D(A[648]), .Y(n1045) );
  NOR2X1 U1543 ( .A(n4045), .B(A[391]), .Y(n1050) );
  NOR2X1 U1544 ( .A(n4045), .B(A[135]), .Y(n1049) );
  NOR2X1 U1551 ( .A(n3801), .B(A[390]), .Y(n1054) );
  NOR2X1 U1559 ( .A(n4040), .B(A[389]), .Y(n1058) );
  NOR2X1 U1567 ( .A(n4040), .B(A[388]), .Y(n1062) );
  NOR2X1 U1575 ( .A(n4040), .B(A[387]), .Y(n1066) );
  NOR2X1 U1583 ( .A(n4040), .B(A[386]), .Y(n1070) );
  NOR2X1 U1584 ( .A(n4040), .B(A[130]), .Y(n1069) );
  NOR2X1 U1591 ( .A(n4031), .B(A[385]), .Y(n1074) );
  NOR2X1 U1599 ( .A(n3684), .B(A[384]), .Y(n1078) );
  NOR2X1 U1600 ( .A(n4039), .B(A[128]), .Y(n1077) );
  NOR2X1 U1607 ( .A(n3793), .B(A[383]), .Y(n1082) );
  NOR2X1 U1615 ( .A(n3769), .B(A[382]), .Y(n1086) );
  NOR2X1 U1623 ( .A(n3818), .B(A[381]), .Y(n1090) );
  NOR2X1 U1631 ( .A(n3824), .B(A[380]), .Y(n1094) );
  NOR2X1 U1639 ( .A(n3768), .B(A[379]), .Y(n1098) );
  NOR2X1 U1655 ( .A(n4038), .B(A[377]), .Y(n1106) );
  NOR2X1 U1671 ( .A(n3818), .B(A[375]), .Y(n1114) );
  NOR2X1 U1679 ( .A(n3833), .B(A[374]), .Y(n1118) );
  NOR2X1 U1687 ( .A(n3818), .B(A[373]), .Y(n1122) );
  NOR2X1 U1695 ( .A(n4033), .B(A[372]), .Y(n1126) );
  NOR2X1 U1703 ( .A(n4033), .B(A[371]), .Y(n1130) );
  NOR2X1 U1735 ( .A(n4028), .B(A[367]), .Y(n1146) );
  NOR2X1 U1751 ( .A(n3833), .B(A[365]), .Y(n1154) );
  NOR2X1 U1759 ( .A(n3758), .B(A[364]), .Y(n1158) );
  NOR2X1 U1767 ( .A(n3833), .B(A[363]), .Y(n1162) );
  NOR2X1 U1799 ( .A(n3833), .B(A[359]), .Y(n1178) );
  NOR2X1 U1815 ( .A(n3833), .B(A[357]), .Y(n1186) );
  NOR2X1 U1823 ( .A(n3833), .B(A[356]), .Y(n1190) );
  NOR2X1 U1831 ( .A(n3808), .B(A[355]), .Y(n1194) );
  NOR2X1 U1871 ( .A(n3758), .B(A[350]), .Y(n1214) );
  NOR2X1 U1879 ( .A(n3808), .B(A[349]), .Y(n1218) );
  NOR2X1 U1887 ( .A(n4030), .B(A[348]), .Y(n1222) );
  NOR2X1 U1895 ( .A(n3768), .B(A[347]), .Y(n1226) );
  NOR2X1 U1903 ( .A(n4050), .B(A[346]), .Y(n1230) );
  NOR2X1 U1911 ( .A(n4039), .B(A[345]), .Y(n1234) );
  NOR21X1 U1920 ( .B(n4039), .A(A[600]), .Y(n1237) );
  NAND21X1 U1938 ( .B(n3989), .A(n1247), .Y(n1660) );
  NAND21X1 U1945 ( .B(n3989), .A(n1250), .Y(n1659) );
  NAND21X1 U1952 ( .B(n3989), .A(n1253), .Y(n1658) );
  NAND21X1 U1959 ( .B(n3989), .A(n1256), .Y(n1657) );
  NAND21X1 U1966 ( .B(n3989), .A(n1259), .Y(n1656) );
  NAND21X1 U1973 ( .B(n3989), .A(n1262), .Y(n1655) );
  NAND21X1 U1980 ( .B(n3989), .A(n3818), .Y(n1654) );
  NAND21X1 U1986 ( .B(n3989), .A(n3818), .Y(n1653) );
  NAND21X1 U1992 ( .B(n3989), .A(n1269), .Y(n1652) );
  NAND21X1 U1999 ( .B(n3673), .A(n1272), .Y(n1651) );
  NAND21X1 U2006 ( .B(n3673), .A(n1275), .Y(n1650) );
  NAND21X1 U2013 ( .B(n3989), .A(n1278), .Y(n1649) );
  NAND21X1 U2020 ( .B(n3672), .A(n1281), .Y(n1648) );
  NAND21X1 U2027 ( .B(n3672), .A(n1284), .Y(n1647) );
  AO22X1 U2222 ( .A(n4068), .B(A[303]), .C(n3824), .D(A[815]), .Y(n1378) );
  AO22X1 U2313 ( .A(n4059), .B(A[38]), .C(n4047), .D(A[550]), .Y(n1431) );
  AO22X1 U2332 ( .A(n4059), .B(A[292]), .C(n4047), .D(A[804]), .Y(n1444) );
  NOR21X1 U2430 ( .B(n4036), .A(A[537]), .Y(n1495) );
  MUX2IX4 U2611 ( .D0(n9), .D1(n1), .S(n3648), .Y(B[0]) );
  INVX16 U2612 ( .A(n3973), .Y(n3648) );
  MUX2IX1 U2613 ( .D0(n957), .D1(n958), .S(n4018), .Y(n1729) );
  MUX2IX1 U2614 ( .D0(n3911), .D1(n3653), .S(n3938), .Y(n139) );
  AOI22CX1 U2615 ( .C(n886), .D(n3992), .A(n3734), .B(n3990), .Y(n3903) );
  MUX2IXL U2616 ( .D0(A[489]), .D1(A[1001]), .S(n3755), .Y(n610) );
  MUX2IX1 U2617 ( .D0(n1069), .D1(n1070), .S(n3977), .Y(n1705) );
  MUX2IX2 U2618 ( .D0(n3764), .D1(n3765), .S(n3965), .Y(n106) );
  INVX2 U2619 ( .A(n3809), .Y(n4065) );
  AOI22X1 U2620 ( .A(n4059), .B(A[290]), .C(n4046), .D(A[802]), .Y(n3759) );
  NOR21X1 U2621 ( .B(n4029), .A(A[521]), .Y(n1559) );
  AO22X1 U2622 ( .A(n4065), .B(A[170]), .C(n4043), .D(A[682]), .Y(n873) );
  AOI22CXL U2623 ( .C(n4046), .D(A[938]), .A(n4077), .B(n3753), .Y(n3905) );
  INVX4 U2624 ( .A(SH[8]), .Y(n4001) );
  AOI22CX1 U2625 ( .C(n4071), .D(A[40]), .A(n3767), .B(n3700), .Y(n3900) );
  MUX2IX2 U2626 ( .D0(n113), .D1(n121), .S(n3964), .Y(n49) );
  MUX2IX1 U2627 ( .D0(n115), .D1(n123), .S(n3966), .Y(n51) );
  NAND2X1 U2628 ( .A(n3655), .B(n3948), .Y(n115) );
  NOR21X2 U2629 ( .B(n4029), .A(A[592]), .Y(n1262) );
  INVX4 U2630 ( .A(n4054), .Y(n4029) );
  INVX4 U2631 ( .A(n4002), .Y(n3981) );
  INVX2 U2632 ( .A(SH[8]), .Y(n4002) );
  MUX2IX4 U2633 ( .D0(n185), .D1(n177), .S(n3756), .Y(n81) );
  MUX2IX2 U2634 ( .D0(n3862), .D1(n3906), .S(n3814), .Y(n185) );
  INVX3 U2635 ( .A(n4059), .Y(n4050) );
  INVX2 U2636 ( .A(n4074), .Y(n4059) );
  MUX2IX4 U2637 ( .D0(n49), .D1(n57), .S(n3747), .Y(n17) );
  NAND2X2 U2638 ( .A(n3744), .B(n3745), .Y(n57) );
  INVX3 U2639 ( .A(n4051), .Y(n4076) );
  INVX2 U2640 ( .A(SH[9]), .Y(n4051) );
  INVX1 U2641 ( .A(A[1009]), .Y(n3712) );
  INVX2 U2642 ( .A(SH[8]), .Y(n3999) );
  NOR2X1 U2643 ( .A(n3808), .B(A[369]), .Y(n1138) );
  INVX1 U2644 ( .A(A[609]), .Y(n3708) );
  NOR2XL U2645 ( .A(n4039), .B(A[353]), .Y(n1202) );
  INVX1 U2646 ( .A(A[681]), .Y(n3697) );
  INVX1 U2647 ( .A(A[425]), .Y(n3772) );
  INVXL U2648 ( .A(n3952), .Y(n3937) );
  INVX2 U2649 ( .A(SH[4]), .Y(n3949) );
  INVX1 U2650 ( .A(A[184]), .Y(n3701) );
  INVX1 U2651 ( .A(A[696]), .Y(n3702) );
  OR2X1 U2652 ( .A(n4039), .B(A[376]), .Y(n3840) );
  INVX1 U2653 ( .A(n3976), .Y(n3839) );
  INVX2 U2654 ( .A(n4003), .Y(n3978) );
  INVX1 U2655 ( .A(A[560]), .Y(n3800) );
  INVX1 U2656 ( .A(A[536]), .Y(n3799) );
  INVX1 U2657 ( .A(A[216]), .Y(n3775) );
  INVX1 U2658 ( .A(n3958), .Y(n4074) );
  INVX2 U2659 ( .A(n4026), .Y(n4058) );
  INVX1 U2660 ( .A(A[505]), .Y(n3729) );
  INVX1 U2661 ( .A(A[761]), .Y(n3707) );
  INVX1 U2662 ( .A(A[497]), .Y(n3711) );
  INVX1 U2663 ( .A(A[753]), .Y(n3693) );
  INVX2 U2664 ( .A(n3767), .Y(n4022) );
  INVX1 U2665 ( .A(n4070), .Y(n4040) );
  INVX1 U2666 ( .A(A[426]), .Y(n3753) );
  MUX2X1 U2667 ( .D0(A[186]), .D1(A[698]), .S(n4023), .Y(n3895) );
  INVX1 U2668 ( .A(A[650]), .Y(n3752) );
  INVX1 U2669 ( .A(A[138]), .Y(n3751) );
  NOR21XL U2670 ( .B(n3842), .A(A[538]), .Y(n1491) );
  INVX1 U2671 ( .A(A[121]), .Y(n3719) );
  INVX1 U2672 ( .A(A[633]), .Y(n3720) );
  INVX1 U2673 ( .A(A[585]), .Y(n3689) );
  NOR21XL U2674 ( .B(n4074), .A(A[601]), .Y(n1233) );
  NOR21XL U2675 ( .B(n4046), .A(A[561]), .Y(n1367) );
  ENOX1 U2676 ( .A(n4037), .B(n3725), .C(n3682), .D(A[929]), .Y(n928) );
  INVX1 U2677 ( .A(A[417]), .Y(n3725) );
  INVX1 U2678 ( .A(A[249]), .Y(n3706) );
  INVX1 U2679 ( .A(A[241]), .Y(n3692) );
  MUX2IX1 U2680 ( .D0(n674), .D1(n673), .S(n4009), .Y(n1792) );
  MUX2IX1 U2681 ( .D0(A[473]), .D1(A[985]), .S(n4036), .Y(n674) );
  AND2X1 U2682 ( .A(n4029), .B(n3723), .Y(n699) );
  INVX1 U2683 ( .A(A[977]), .Y(n3723) );
  AND2X1 U2684 ( .A(n4039), .B(n3704), .Y(n755) );
  INVX1 U2685 ( .A(A[961]), .Y(n3704) );
  AND2X1 U2686 ( .A(n4029), .B(n3727), .Y(n993) );
  INVX1 U2687 ( .A(A[657]), .Y(n3727) );
  EORX1 U2688 ( .A(n1040), .B(n3672), .C(n3760), .D(n3984), .Y(n3774) );
  INVX1 U2689 ( .A(A[393]), .Y(n3822) );
  INVX1 U2690 ( .A(A[296]), .Y(n3797) );
  INVX1 U2691 ( .A(A[808]), .Y(n3798) );
  INVX1 U2692 ( .A(A[552]), .Y(n3700) );
  NOR21XL U2693 ( .B(n3782), .A(A[528]), .Y(n1531) );
  AND2X1 U2694 ( .A(n3755), .B(n3804), .Y(n758) );
  INVX1 U2695 ( .A(A[960]), .Y(n3804) );
  INVX1 U2696 ( .A(A[1008]), .Y(n3685) );
  INVX1 U2697 ( .A(A[496]), .Y(n3740) );
  MUX2IX1 U2698 ( .D0(A[480]), .D1(A[992]), .S(n4039), .Y(n646) );
  INVX1 U2699 ( .A(A[240]), .Y(n3688) );
  INVX1 U2700 ( .A(n4004), .Y(n4015) );
  INVX1 U2701 ( .A(n3947), .Y(n3844) );
  NOR2X1 U2702 ( .A(n3808), .B(A[370]), .Y(n1134) );
  NOR2X1 U2703 ( .A(n4033), .B(A[354]), .Y(n1198) );
  NOR21XL U2704 ( .B(n3670), .A(A[978]), .Y(n696) );
  NOR21XL U2705 ( .B(n4035), .A(A[530]), .Y(n1523) );
  NOR21XL U2706 ( .B(n4029), .A(A[593]), .Y(n1259) );
  AND2X1 U2707 ( .A(n3986), .B(n1305), .Y(n3875) );
  MUX2X1 U2708 ( .D0(n1201), .D1(n1202), .S(n3978), .Y(n3763) );
  MUX2X1 U2709 ( .D0(n1696), .D1(n1680), .S(n3835), .Y(n170) );
  NOR21XL U2710 ( .B(n4034), .A(A[569]), .Y(n1335) );
  MUX2IX1 U2711 ( .D0(n3743), .D1(n3742), .S(n3730), .Y(n122) );
  INVX1 U2712 ( .A(n3675), .Y(n3730) );
  MUX2X1 U2713 ( .D0(n1527), .D1(n1528), .S(n3987), .Y(n3868) );
  INVX1 U2714 ( .A(n3955), .Y(n3757) );
  MUX2X1 U2715 ( .D0(n786), .D1(n785), .S(n3773), .Y(n3783) );
  OR2X1 U2716 ( .A(n4042), .B(A[440]), .Y(n3749) );
  AND2X1 U2717 ( .A(n4036), .B(n3817), .Y(n1141) );
  INVX1 U2718 ( .A(A[624]), .Y(n3817) );
  NOR21XL U2719 ( .B(n4036), .A(A[608]), .Y(n1205) );
  AND2X1 U2720 ( .A(n3986), .B(n1308), .Y(n3874) );
  MUX2X1 U2721 ( .D0(n1647), .D1(n1663), .S(n3940), .Y(n153) );
  MUX2IX1 U2722 ( .D0(n3838), .D1(n3652), .S(n3733), .Y(n169) );
  INVX1 U2723 ( .A(n3940), .Y(n3733) );
  MUX2IX1 U2724 ( .D0(n3840), .D1(n3841), .S(n3839), .Y(n3838) );
  MUX2IX2 U2725 ( .D0(n3811), .D1(n3812), .S(n3810), .Y(n3765) );
  INVX3 U2726 ( .A(n4078), .Y(n4053) );
  INVX1 U2727 ( .A(n4078), .Y(n3827) );
  MUX2IX2 U2728 ( .D0(n153), .D1(n145), .S(n3756), .Y(n65) );
  INVX1 U2729 ( .A(n3958), .Y(n3807) );
  INVXL U2730 ( .A(n4054), .Y(n4032) );
  INVX1 U2731 ( .A(n4076), .Y(n4067) );
  INVX1 U2732 ( .A(n3943), .Y(n3814) );
  INVX1 U2733 ( .A(n3969), .Y(n3968) );
  INVX1 U2734 ( .A(n3948), .Y(n3835) );
  INVX2 U2735 ( .A(n3951), .Y(n3940) );
  INVX6 U2736 ( .A(n3732), .Y(n4036) );
  INVX1 U2737 ( .A(SH[3]), .Y(n3970) );
  INVXL U2738 ( .A(n4016), .Y(n4008) );
  INVX1 U2739 ( .A(n3997), .Y(n3705) );
  INVX1 U2740 ( .A(n3950), .Y(n3944) );
  INVXL U2741 ( .A(n3948), .Y(n3690) );
  INVX1 U2742 ( .A(n3969), .Y(n3964) );
  INVX1 U2743 ( .A(n3953), .Y(n3776) );
  INVX1 U2744 ( .A(n3963), .Y(n3756) );
  INVXL U2745 ( .A(n3844), .Y(n3810) );
  INVXL U2746 ( .A(n3951), .Y(n3703) );
  INVX1 U2747 ( .A(n3790), .Y(n4019) );
  INVX1 U2748 ( .A(n4020), .Y(n4005) );
  INVX1 U2749 ( .A(n4017), .Y(n4006) );
  BUFX8 U2750 ( .A(n3961), .Y(n3732) );
  INVX1 U2751 ( .A(n3813), .Y(n4049) );
  INVX1 U2752 ( .A(n3957), .Y(n3747) );
  INVX1 U2753 ( .A(n3790), .Y(n4020) );
  INVXL U2754 ( .A(n4015), .Y(n4012) );
  INVX1 U2755 ( .A(n3972), .Y(n3971) );
  INVX1 U2756 ( .A(SH[7]), .Y(n3974) );
  INVX1 U2757 ( .A(n3974), .Y(n3973) );
  AOI22X1 U2758 ( .A(n4013), .B(n909), .C(n910), .D(n3673), .Y(n3649) );
  AND2X1 U2759 ( .A(n702), .B(n3988), .Y(n3650) );
  INVX1 U2760 ( .A(n3963), .Y(n3834) );
  AOI22XL U2761 ( .A(n4005), .B(n819), .C(n820), .D(n3992), .Y(n3651) );
  INVXL U2762 ( .A(n3949), .Y(n3946) );
  INVXL U2763 ( .A(n3951), .Y(n3939) );
  INVX1 U2764 ( .A(n3844), .Y(n3686) );
  MUX2X1 U2765 ( .D0(n1173), .D1(n1174), .S(n3978), .Y(n3652) );
  MUX2X1 U2766 ( .D0(n1331), .D1(n3866), .S(n3705), .Y(n3653) );
  MUX2X1 U2767 ( .D0(n637), .D1(n638), .S(n3979), .Y(n3654) );
  MUX2X1 U2768 ( .D0(n1523), .D1(n3873), .S(n3679), .Y(n3655) );
  MUX2X1 U2769 ( .D0(n1555), .D1(n1556), .S(n3984), .Y(n3656) );
  MUX2X1 U2770 ( .D0(n993), .D1(n994), .S(n4018), .Y(n3657) );
  AND2X1 U2771 ( .A(n3987), .B(n752), .Y(n3658) );
  AND2X1 U2772 ( .A(n3988), .B(n755), .Y(n3659) );
  AND2X1 U2773 ( .A(n3716), .B(n3717), .Y(n3660) );
  AND2X1 U2774 ( .A(n758), .B(n3988), .Y(n3661) );
  AOI22X1 U2775 ( .A(n4004), .B(n915), .C(n916), .D(n3991), .Y(n3662) );
  AOI22X1 U2776 ( .A(n4012), .B(n813), .C(n814), .D(n3993), .Y(n3663) );
  AOI22X1 U2777 ( .A(n4012), .B(n1383), .C(n1384), .D(n3994), .Y(n3664) );
  AOI22X1 U2778 ( .A(n4012), .B(n855), .C(n856), .D(n3991), .Y(n3665) );
  INVX1 U2779 ( .A(n3969), .Y(n3967) );
  MUX2X1 U2780 ( .D0(n1507), .D1(n1508), .S(n3681), .Y(n3666) );
  INVX2 U2781 ( .A(n4021), .Y(n3980) );
  INVX3 U2782 ( .A(n3755), .Y(n4054) );
  AOI22X1 U2783 ( .A(n4013), .B(n849), .C(n850), .D(n3993), .Y(n3667) );
  AOI22X1 U2784 ( .A(n4014), .B(n843), .C(n844), .D(n3993), .Y(n3668) );
  AOI22X1 U2785 ( .A(n4007), .B(n1431), .C(n1432), .D(n3994), .Y(n3669) );
  INVX2 U2786 ( .A(n4078), .Y(n4060) );
  INVX8 U2787 ( .A(SH[9]), .Y(n3961) );
  INVX3 U2788 ( .A(SH[9]), .Y(n4052) );
  INVXL U2789 ( .A(n4067), .Y(n3670) );
  INVX1 U2790 ( .A(n3990), .Y(n3671) );
  INVX2 U2791 ( .A(n3671), .Y(n3672) );
  INVXL U2792 ( .A(n3671), .Y(n3673) );
  INVX1 U2793 ( .A(n3956), .Y(n3953) );
  INVX2 U2794 ( .A(n3732), .Y(n4037) );
  INVX2 U2795 ( .A(n3732), .Y(n4027) );
  INVXL U2796 ( .A(n3732), .Y(n4075) );
  INVXL U2797 ( .A(n3937), .Y(n3674) );
  INVXL U2798 ( .A(n3674), .Y(n3675) );
  INVX1 U2799 ( .A(n3674), .Y(n3676) );
  INVX1 U2800 ( .A(n4000), .Y(n3986) );
  INVX1 U2801 ( .A(n4000), .Y(n3985) );
  AND2X1 U2802 ( .A(n3684), .B(n3799), .Y(n1499) );
  AND2X1 U2803 ( .A(n3684), .B(n3708), .Y(n1201) );
  INVX1 U2804 ( .A(n4077), .Y(n3778) );
  INVX1 U2805 ( .A(n3970), .Y(n3963) );
  INVX1 U2806 ( .A(n3970), .Y(n3816) );
  INVXL U2807 ( .A(n3951), .Y(n3945) );
  INVX3 U2808 ( .A(n4053), .Y(n4039) );
  INVX1 U2809 ( .A(n4053), .Y(n3808) );
  INVX1 U2810 ( .A(n4053), .Y(n4033) );
  INVXL U2811 ( .A(n4063), .Y(n3677) );
  NOR21XL U2812 ( .B(n3677), .A(A[714]), .Y(n725) );
  NOR21XL U2813 ( .B(n3677), .A(A[970]), .Y(n726) );
  EORX1 U2814 ( .A(n3677), .B(A[1017]), .C(n3788), .D(n3729), .Y(n3789) );
  NOR21XL U2815 ( .B(n4076), .A(A[713]), .Y(n729) );
  ENOX1 U2816 ( .A(n4073), .B(n3822), .C(n4076), .D(A[905]), .Y(n1040) );
  INVX3 U2817 ( .A(n4076), .Y(n4068) );
  INVX1 U2818 ( .A(n4079), .Y(n4063) );
  INVXL U2819 ( .A(n3986), .Y(n3678) );
  INVXL U2820 ( .A(n3678), .Y(n3679) );
  INVXL U2821 ( .A(n3678), .Y(n3680) );
  INVXL U2822 ( .A(n3678), .Y(n3681) );
  INVX2 U2823 ( .A(n4052), .Y(n3682) );
  INVX2 U2824 ( .A(n4052), .Y(n3683) );
  INVX3 U2825 ( .A(n4052), .Y(n4043) );
  INVX1 U2826 ( .A(n4052), .Y(n4042) );
  INVXL U2827 ( .A(n3961), .Y(n3684) );
  OAI22X1 U2828 ( .A(n4077), .B(n3740), .C(n4052), .D(n3685), .Y(n3815) );
  MUX2BX1 U2829 ( .D0(n1655), .D1(n3874), .S(n3952), .Y(n145) );
  INVXL U2830 ( .A(SH[4]), .Y(n3952) );
  AOI22CX1 U2831 ( .C(n4043), .D(A[752]), .A(n4079), .B(n3688), .Y(n3722) );
  BUFXL U2832 ( .A(n4079), .Y(n3696) );
  MUX2IX1 U2833 ( .D0(n3701), .D1(n3702), .S(n4026), .Y(n3750) );
  INVX6 U2834 ( .A(n3958), .Y(n4026) );
  MUX2IX1 U2835 ( .D0(A[280]), .D1(A[792]), .S(n4046), .Y(n1500) );
  MUX2IX4 U2836 ( .D0(n33), .D1(n41), .S(SH[6]), .Y(n9) );
  AOI22CX1 U2837 ( .C(n3790), .D(n933), .A(n3754), .B(n4000), .Y(n3902) );
  INVX3 U2838 ( .A(n4021), .Y(n3984) );
  INVX1 U2839 ( .A(SH[8]), .Y(n3790) );
  INVX3 U2840 ( .A(n3999), .Y(n3990) );
  MUX2IX2 U2841 ( .D0(n1807), .D1(n1823), .S(n3686), .Y(n3843) );
  MUX2X2 U2842 ( .D0(n3687), .D1(n1703), .S(n3690), .Y(n177) );
  MUX2IXL U2843 ( .D0(n997), .D1(n998), .S(n3978), .Y(n3687) );
  AOI22BX1 U2844 ( .B(n3705), .A(n837), .D(n3960), .C(n4019), .Y(n3959) );
  INVXL U2845 ( .A(n3990), .Y(n4013) );
  MUX2IX1 U2846 ( .D0(n3902), .D1(n3959), .S(n3703), .Y(n193) );
  MUX2IX1 U2847 ( .D0(A[264]), .D1(A[776]), .S(n4034), .Y(n1564) );
  INVX1 U2848 ( .A(n4051), .Y(n4034) );
  INVXL U2849 ( .A(n4051), .Y(n4044) );
  INVX2 U2850 ( .A(n4052), .Y(n4046) );
  INVX1 U2851 ( .A(n4007), .Y(n3826) );
  MUX2IX4 U2852 ( .D0(n73), .D1(n65), .S(n3776), .Y(n25) );
  MUX2IX2 U2853 ( .D0(n169), .D1(n161), .S(n3756), .Y(n73) );
  MUX2IX1 U2854 ( .D0(n122), .D1(n114), .S(n3834), .Y(n50) );
  AND2X1 U2855 ( .A(n4029), .B(n3689), .Y(n1281) );
  INVXL U2856 ( .A(n3950), .Y(n3943) );
  MUX2IX1 U2857 ( .D0(n1632), .D1(n1616), .S(n3690), .Y(n3726) );
  AOI22X1 U2858 ( .A(n576), .B(n3995), .C(n3790), .D(n3691), .Y(n3786) );
  OAI22X1 U2859 ( .A(n3683), .B(n3692), .C(n4051), .D(n3693), .Y(n3691) );
  MUX2IX1 U2860 ( .D0(n58), .D1(n50), .S(n3757), .Y(n18) );
  MUX2IX1 U2861 ( .D0(n98), .D1(n106), .S(n3954), .Y(n42) );
  MUX2IX1 U2862 ( .D0(n18), .D1(n26), .S(SH[6]), .Y(n2) );
  INVXL U2863 ( .A(n3844), .Y(n3694) );
  MUX2IX1 U2864 ( .D0(n42), .D1(n34), .S(n3972), .Y(n10) );
  INVXL U2865 ( .A(n3705), .Y(n3748) );
  INVX1 U2866 ( .A(n4020), .Y(n3773) );
  AOI22CX1 U2867 ( .C(n4009), .D(n527), .A(n3789), .B(n4009), .Y(n3812) );
  MUX2IXL U2868 ( .D0(n227), .D1(n235), .S(n3816), .Y(n107) );
  MUX2IX1 U2869 ( .D0(n3654), .D1(n3914), .S(n3946), .Y(n227) );
  MUX2IX1 U2870 ( .D0(A[185]), .D1(A[697]), .S(n4026), .Y(n785) );
  MUX2IX1 U2871 ( .D0(n3784), .D1(n3783), .S(n3940), .Y(n3771) );
  INVXL U2872 ( .A(SH[6]), .Y(n3972) );
  AOI22CX1 U2873 ( .C(n928), .D(n3992), .A(n3672), .B(n3695), .Y(n3795) );
  AOI22X1 U2874 ( .A(n4058), .B(A[161]), .C(n3682), .D(A[673]), .Y(n3695) );
  INVX4 U2875 ( .A(n3981), .Y(n4004) );
  INVX6 U2876 ( .A(n4079), .Y(n3958) );
  INVX2 U2877 ( .A(n4061), .Y(n4038) );
  NOR2XL U2878 ( .A(n4038), .B(A[361]), .Y(n1170) );
  AO22AX1 U2879 ( .A(n4060), .B(A[169]), .C(n4043), .D(n3697), .Y(n879) );
  EORX1 U2880 ( .A(n4005), .B(n3698), .C(n3699), .D(n3998), .Y(n3794) );
  AO22X1 U2881 ( .A(n4061), .B(A[177]), .C(n3755), .D(A[689]), .Y(n3698) );
  AOI22X1 U2882 ( .A(n3755), .B(A[945]), .C(n3778), .D(A[433]), .Y(n3699) );
  INVXL U2883 ( .A(n3998), .Y(n3993) );
  INVXL U2884 ( .A(n3944), .Y(n3724) );
  MUX2IX4 U2885 ( .D0(n81), .D1(n89), .S(n3747), .Y(n33) );
  MUX2IX2 U2886 ( .D0(n193), .D1(n201), .S(n3816), .Y(n89) );
  AO22XL U2887 ( .A(n4011), .B(n891), .C(n892), .D(n3993), .Y(n1742) );
  INVXL U2888 ( .A(n3942), .Y(n3728) );
  MUX2IX1 U2889 ( .D0(n3875), .D1(n314), .S(n3942), .Y(n146) );
  INVXL U2890 ( .A(n3961), .Y(n3848) );
  INVX1 U2891 ( .A(n4074), .Y(n4071) );
  INVXL U2892 ( .A(n3941), .Y(n3761) );
  MUX2X1 U2893 ( .D0(A[122]), .D1(A[634]), .S(n4046), .Y(n3892) );
  AO22XL U2894 ( .A(n4057), .B(A[397]), .C(n4050), .D(A[909]), .Y(n1016) );
  MUX2X1 U2895 ( .D0(n1583), .D1(n1599), .S(n3675), .Y(n121) );
  INVX4 U2896 ( .A(n3796), .Y(n4021) );
  INVX1 U2897 ( .A(n3958), .Y(n3830) );
  OAI22CXL U2898 ( .C(n3732), .D(n3806), .A(n4060), .B(A[288]), .Y(n1468) );
  MUX2IX1 U2899 ( .D0(n107), .D1(n99), .S(n3957), .Y(n43) );
  MUX2IX1 U2900 ( .D0(n11), .D1(n3), .S(n3974), .Y(B[2]) );
  MUX2IXL U2901 ( .D0(A[921]), .D1(A[409]), .S(n3778), .Y(n962) );
  NOR2X1 U2902 ( .A(n3696), .B(A[441]), .Y(n786) );
  MUX2IX1 U2903 ( .D0(n1776), .D1(n1792), .S(n3703), .Y(n3709) );
  MUX2IX1 U2904 ( .D0(A[265]), .D1(A[777]), .S(n4026), .Y(n1560) );
  INVX1 U2905 ( .A(SH[4]), .Y(n3951) );
  OAI22AX1 U2906 ( .D(n3999), .C(n3779), .A(n4008), .B(n3780), .Y(n1608) );
  INVX2 U2907 ( .A(n4021), .Y(n4018) );
  INVX2 U2908 ( .A(n4003), .Y(n4016) );
  INVX2 U2909 ( .A(SH[8]), .Y(n3997) );
  INVXL U2910 ( .A(n4079), .Y(n4055) );
  OAI22AX1 U2911 ( .D(n4073), .C(n3707), .A(n4037), .B(n3706), .Y(n527) );
  INVX1 U2912 ( .A(n3997), .Y(n3996) );
  INVX1 U2913 ( .A(n3997), .Y(n3994) );
  INVXL U2914 ( .A(n4054), .Y(n4030) );
  MUX2BX1 U2915 ( .D0(n3709), .D1(n210), .S(n3834), .Y(n98) );
  MUX2IX1 U2916 ( .D0(n211), .D1(n219), .S(n3964), .Y(n99) );
  INVXL U2917 ( .A(n4026), .Y(n3710) );
  OAI22AX1 U2918 ( .D(n3682), .C(n3712), .A(n3848), .B(n3711), .Y(n576) );
  NOR21XL U2919 ( .B(n4035), .A(A[607]), .Y(n1209) );
  NOR21XL U2920 ( .B(n4035), .A(A[614]), .Y(n1181) );
  MUX2IX1 U2921 ( .D0(n51), .D1(n59), .S(n3955), .Y(n19) );
  NAND2X1 U2922 ( .A(n3726), .B(n3966), .Y(n3713) );
  NAND2X1 U2923 ( .A(n3660), .B(n3756), .Y(n3714) );
  NAND2X1 U2924 ( .A(n3713), .B(n3714), .Y(n58) );
  NAND2X1 U2925 ( .A(n1608), .B(n3715), .Y(n3716) );
  NAND2X1 U2926 ( .A(n1624), .B(n3676), .Y(n3717) );
  INVXL U2927 ( .A(n3675), .Y(n3715) );
  INVX2 U2928 ( .A(n4060), .Y(n3741) );
  INVX6 U2929 ( .A(n4079), .Y(n4056) );
  INVXL U2930 ( .A(n4075), .Y(n3718) );
  MUX2X1 U2931 ( .D0(n609), .D1(n610), .S(n4019), .Y(n3811) );
  MUX2X1 U2932 ( .D0(n3720), .D1(n3719), .S(n4053), .Y(n1105) );
  NOR21X1 U2933 ( .B(n4043), .A(A[617]), .Y(n1169) );
  INVXL U2934 ( .A(n3777), .Y(n3721) );
  MUX2X1 U2935 ( .D0(A[120]), .D1(A[632]), .S(n4043), .Y(n3841) );
  INVXL U2936 ( .A(n4076), .Y(n4072) );
  INVXL U2937 ( .A(n4052), .Y(n3788) );
  MUX2X1 U2938 ( .D0(n1073), .D1(n1074), .S(n3977), .Y(n3916) );
  AOI22CX1 U2939 ( .C(n3815), .D(n3995), .A(n4015), .B(n3722), .Y(n3731) );
  INVX1 U2940 ( .A(n4015), .Y(n4011) );
  MUX2IXL U2941 ( .D0(A[472]), .D1(A[984]), .S(n4079), .Y(n678) );
  INVX4 U2942 ( .A(n3999), .Y(n3989) );
  INVX4 U2943 ( .A(n3999), .Y(n3988) );
  INVX1 U2944 ( .A(n1656), .Y(n314) );
  MUX2IX1 U2945 ( .D0(n3850), .D1(n3659), .S(n3724), .Y(n210) );
  INVXL U2946 ( .A(n4076), .Y(n4066) );
  MUX2IX2 U2947 ( .D0(n203), .D1(n195), .S(n3834), .Y(n91) );
  INVX2 U2948 ( .A(n4036), .Y(n4069) );
  OAI22AX1 U2949 ( .D(n4027), .C(n3752), .A(n4023), .B(n3751), .Y(n1033) );
  NOR2XL U2950 ( .A(n4038), .B(A[362]), .Y(n1166) );
  INVX1 U2951 ( .A(n4055), .Y(n3782) );
  MUX2IXL U2952 ( .D0(A[920]), .D1(A[408]), .S(n3732), .Y(n966) );
  MUX2X1 U2953 ( .D0(n961), .D1(n962), .S(n3980), .Y(n3849) );
  AOI22X1 U2954 ( .A(n4060), .B(A[34]), .C(n3788), .D(A[546]), .Y(n3910) );
  MUX2X2 U2955 ( .D0(n1559), .D1(n1560), .S(n3975), .Y(n3742) );
  AO22XL U2956 ( .A(n4070), .B(A[295]), .C(n3805), .D(A[807]), .Y(n1426) );
  AO22XL U2957 ( .A(n4070), .B(A[293]), .C(n4047), .D(A[805]), .Y(n1438) );
  AO22XL U2958 ( .A(n4070), .B(A[291]), .C(n4047), .D(A[803]), .Y(n1450) );
  MUX2IX4 U2959 ( .D0(n3843), .D1(n105), .S(n3962), .Y(n41) );
  MUX2IX4 U2960 ( .D0(n225), .D1(n3803), .S(n3776), .Y(n105) );
  MUX2IX1 U2961 ( .D0(A[305]), .D1(A[817]), .S(n4036), .Y(n1368) );
  INVX1 U2962 ( .A(n3796), .Y(n3998) );
  INVX2 U2963 ( .A(n3998), .Y(n3992) );
  MUX2IX1 U2964 ( .D0(n3657), .D1(n3916), .S(n3728), .Y(n178) );
  AND2X1 U2965 ( .A(n3988), .B(n699), .Y(n3850) );
  AOI22X1 U2966 ( .A(n4064), .B(A[434]), .C(n3741), .D(A[946]), .Y(n3913) );
  INVX1 U2967 ( .A(n3949), .Y(n3947) );
  AOI22AX1 U2968 ( .A(n922), .B(n3673), .D(n3908), .C(n4014), .Y(n3907) );
  AO22X1 U2969 ( .A(n4064), .B(A[178]), .C(n4047), .D(A[690]), .Y(n825) );
  INVXL U2970 ( .A(n3944), .Y(n3785) );
  NOR2XL U2971 ( .A(n4027), .B(A[344]), .Y(n1238) );
  MUX2IX1 U2972 ( .D0(n154), .D1(n146), .S(n3969), .Y(n66) );
  MUX2IX1 U2973 ( .D0(n74), .D1(n66), .S(n3776), .Y(n26) );
  INVXL U2974 ( .A(n3718), .Y(n4025) );
  NOR2XL U2975 ( .A(n3741), .B(A[360]), .Y(n1174) );
  MUX2IX4 U2976 ( .D0(n25), .D1(n17), .S(n3972), .Y(n1) );
  MUX2IX1 U2977 ( .D0(n3770), .D1(n3771), .S(n3963), .Y(n90) );
  NOR21XL U2978 ( .B(n4034), .A(A[602]), .Y(n1229) );
  NOR21XL U2979 ( .B(n4034), .A(A[570]), .Y(n1331) );
  MUX2AX2 U2980 ( .D0(n3731), .D1(n1799), .S(n3814), .Y(n225) );
  INVX8 U2981 ( .A(n4056), .Y(n3755) );
  MUX2X1 U2982 ( .D0(n1371), .D1(n1372), .S(n3982), .Y(n3746) );
  INVX3 U2983 ( .A(n4021), .Y(n3979) );
  MUX2IX1 U2984 ( .D0(n3863), .D1(n3903), .S(n3690), .Y(n201) );
  INVX6 U2985 ( .A(n4004), .Y(n3975) );
  AO22XL U2986 ( .A(n3823), .B(A[253]), .C(n3824), .D(A[765]), .Y(n503) );
  AO22XL U2987 ( .A(n3777), .B(A[251]), .C(n3824), .D(A[763]), .Y(n515) );
  AO22XL U2988 ( .A(n4071), .B(A[247]), .C(n4025), .D(A[759]), .Y(n539) );
  AO22XL U2989 ( .A(n4071), .B(A[243]), .C(n3766), .D(A[755]), .Y(n563) );
  MUX2X2 U2990 ( .D0(n3825), .D1(n3746), .S(n3703), .Y(n3831) );
  MUX2IX1 U2991 ( .D0(n1233), .D1(n1234), .S(n3980), .Y(n1664) );
  AO22XL U2992 ( .A(n4069), .B(A[301]), .C(n3824), .D(A[813]), .Y(n1390) );
  AO22XL U2993 ( .A(n4069), .B(A[299]), .C(n4033), .D(A[811]), .Y(n1402) );
  INVX2 U2994 ( .A(n4026), .Y(n4057) );
  MUX2X2 U2995 ( .D0(n1671), .D1(n1687), .S(n3941), .Y(n161) );
  INVX2 U2996 ( .A(n3997), .Y(n3995) );
  INVX1 U2997 ( .A(n3995), .Y(n3899) );
  INVX2 U2998 ( .A(n4003), .Y(n3977) );
  NAND21XL U2999 ( .B(n3988), .A(n1241), .Y(n1662) );
  NAND21XL U3000 ( .B(n3988), .A(n1244), .Y(n1661) );
  INVX1 U3001 ( .A(SH[8]), .Y(n4003) );
  MUX2IX1 U3002 ( .D0(n1205), .D1(n1206), .S(n3979), .Y(n1671) );
  INVX2 U3003 ( .A(n3796), .Y(n4000) );
  AOI22X1 U3004 ( .A(n4065), .B(A[168]), .C(n3683), .D(A[680]), .Y(n3734) );
  MUX2IX1 U3005 ( .D0(A[474]), .D1(A[986]), .S(n4046), .Y(n670) );
  MUX2IX1 U3006 ( .D0(n186), .D1(n178), .S(n3834), .Y(n82) );
  NAND2X1 U3007 ( .A(n217), .B(n3965), .Y(n3735) );
  NAND2X1 U3008 ( .A(n209), .B(n3969), .Y(n3736) );
  NAND2X1 U3009 ( .A(n3735), .B(n3736), .Y(n3803) );
  NAND2X1 U3010 ( .A(n3836), .B(n3737), .Y(n3738) );
  NAND2X1 U3011 ( .A(n3837), .B(n3835), .Y(n3739) );
  NAND2X1 U3012 ( .A(n3738), .B(n3739), .Y(n217) );
  INVX1 U3013 ( .A(n3835), .Y(n3737) );
  MUX2IX1 U3014 ( .D0(n3661), .D1(n3650), .S(n3944), .Y(n209) );
  INVX2 U3015 ( .A(n4016), .Y(n4009) );
  INVX2 U3016 ( .A(n3983), .Y(n3829) );
  MUX2IX1 U3017 ( .D0(n3849), .D1(n3774), .S(n3814), .Y(n186) );
  MUX2X1 U3018 ( .D0(n1495), .D1(n1496), .S(n3983), .Y(n3743) );
  NAND2X1 U3019 ( .A(n3831), .B(n3756), .Y(n3744) );
  NAND2X1 U3020 ( .A(n3832), .B(n3968), .Y(n3745) );
  MUX2IX1 U3021 ( .D0(n170), .D1(n162), .S(n3834), .Y(n74) );
  AO22XL U3022 ( .A(n4058), .B(A[46]), .C(n4045), .D(A[558]), .Y(n1383) );
  AO22XL U3023 ( .A(n4058), .B(A[300]), .C(n3758), .D(A[812]), .Y(n1396) );
  AO22XL U3024 ( .A(n4058), .B(A[298]), .C(n4048), .D(A[810]), .Y(n1408) );
  AOI22AX1 U3025 ( .A(n880), .B(n3705), .D(n4020), .C(n879), .Y(n3784) );
  MUX2IXL U3026 ( .D0(A[313]), .D1(A[825]), .S(n3682), .Y(n1336) );
  NOR21XL U3027 ( .B(n4043), .A(A[616]), .Y(n1173) );
  INVX2 U3028 ( .A(n4078), .Y(n4061) );
  MUX2IX1 U3029 ( .D0(n82), .D1(n90), .S(n3747), .Y(n34) );
  MUX2IX1 U3030 ( .D0(n3749), .D1(n3750), .S(n3748), .Y(n3863) );
  NOR2XL U3031 ( .A(n4075), .B(A[218]), .Y(n669) );
  MUX2IX1 U3032 ( .D0(n3907), .D1(n3912), .S(n3944), .Y(n195) );
  NOR2XL U3033 ( .A(n3842), .B(A[234]), .Y(n605) );
  AO22XL U3034 ( .A(n4062), .B(A[242]), .C(n3682), .D(A[754]), .Y(n569) );
  NOR2XL U3035 ( .A(n3683), .B(A[233]), .Y(n609) );
  NOR21XL U3036 ( .B(n4043), .A(A[664]), .Y(n965) );
  NOR21XL U3037 ( .B(n4042), .A(A[665]), .Y(n961) );
  MUX2IX1 U3038 ( .D0(n187), .D1(n179), .S(n3969), .Y(n83) );
  AO22XL U3039 ( .A(n3718), .B(A[511]), .C(n3824), .D(A[1023]), .Y(n492) );
  MUX2IX1 U3040 ( .D0(A[400]), .D1(A[912]), .S(n3848), .Y(n998) );
  MUX2IX1 U3041 ( .D0(n3795), .D1(n3794), .S(n3810), .Y(n3770) );
  INVX2 U3042 ( .A(n3961), .Y(n4077) );
  INVX3 U3043 ( .A(n4001), .Y(n3796) );
  OR2X1 U3044 ( .A(n4039), .B(A[378]), .Y(n3893) );
  AO22XL U3045 ( .A(n3777), .B(A[175]), .C(n4045), .D(A[687]), .Y(n843) );
  MUX2IX1 U3046 ( .D0(n645), .D1(n646), .S(n3983), .Y(n1799) );
  NOR2XL U3047 ( .A(n4037), .B(A[224]), .Y(n645) );
  AOI22X1 U3048 ( .A(n4068), .B(A[416]), .C(n3807), .D(A[928]), .Y(n3754) );
  MUX2IXL U3049 ( .D0(n3871), .D1(n3898), .S(n3947), .Y(n235) );
  AOI22AX1 U3050 ( .A(n4009), .B(n521), .D(n3872), .C(n3996), .Y(n3898) );
  MUX2IX1 U3051 ( .D0(n91), .D1(n83), .S(n3757), .Y(n35) );
  INVX2 U3052 ( .A(n3949), .Y(n3948) );
  INVXL U3053 ( .A(n3823), .Y(n3758) );
  MUX2IX1 U3054 ( .D0(n67), .D1(n75), .S(n3747), .Y(n27) );
  AOI22AX1 U3055 ( .A(n4011), .B(n569), .D(n3915), .C(n3995), .Y(n3914) );
  AOI22BXL U3056 ( .B(n3759), .A(n3994), .D(n3910), .C(n4008), .Y(n3909) );
  MUX2IXL U3057 ( .D0(A[994]), .D1(A[482]), .S(n4059), .Y(n638) );
  AOI22X1 U3058 ( .A(n4057), .B(A[137]), .C(n4076), .D(A[649]), .Y(n3760) );
  MUX2IX1 U3059 ( .D0(n3762), .D1(n3763), .S(n3761), .Y(n162) );
  MUX2X2 U3060 ( .D0(n1137), .D1(n1138), .S(n3975), .Y(n3762) );
  MUX2IX1 U3061 ( .D0(n3786), .D1(n3787), .S(n3785), .Y(n3764) );
  INVX1 U3062 ( .A(n3777), .Y(n3766) );
  NOR21X1 U3063 ( .B(n4036), .A(A[625]), .Y(n1137) );
  INVXL U3064 ( .A(n4078), .Y(n3767) );
  INVX4 U3065 ( .A(n3961), .Y(n4078) );
  MUX2AX2 U3066 ( .D0(n3904), .D1(n1761), .S(n3944), .Y(n203) );
  INVXL U3067 ( .A(n4061), .Y(n3768) );
  INVXL U3068 ( .A(n4079), .Y(n3828) );
  MUX2IX1 U3069 ( .D0(n1367), .D1(n1368), .S(n3982), .Y(n1624) );
  MUX2IX1 U3070 ( .D0(A[402]), .D1(A[914]), .S(n4022), .Y(n990) );
  MUX2X1 U3071 ( .D0(n1648), .D1(n1664), .S(n3940), .Y(n154) );
  MUX2X1 U3072 ( .D0(n3892), .D1(n3893), .S(n3976), .Y(n1697) );
  MUX2IX1 U3073 ( .D0(n1169), .D1(n1170), .S(n3996), .Y(n1680) );
  INVXL U3074 ( .A(n4068), .Y(n3769) );
  AOI22AX1 U3075 ( .A(n4012), .B(n825), .D(n3913), .C(n3992), .Y(n3912) );
  AOI22X1 U3076 ( .A(n4067), .B(A[162]), .C(n4033), .D(A[674]), .Y(n3908) );
  MUX2IX1 U3077 ( .D0(A[816]), .D1(A[304]), .S(n3827), .Y(n1372) );
  MUX2X1 U3078 ( .D0(n3895), .D1(n3896), .S(n4020), .Y(n1761) );
  MUX2IX1 U3079 ( .D0(A[281]), .D1(A[793]), .S(n3755), .Y(n1496) );
  AO22AX1 U3080 ( .A(n3683), .B(A[937]), .C(n4060), .D(n3772), .Y(n880) );
  MUX2IX1 U3081 ( .D0(A[401]), .D1(A[913]), .S(n3683), .Y(n994) );
  MUX2IXL U3082 ( .D0(A[312]), .D1(A[824]), .S(n3683), .Y(n1340) );
  AO22XL U3083 ( .A(n3823), .B(A[165]), .C(n4028), .D(A[677]), .Y(n903) );
  AO22XL U3084 ( .A(n3823), .B(A[163]), .C(n4028), .D(A[675]), .Y(n915) );
  NOR21XL U3085 ( .B(n4076), .A(A[969]), .Y(n730) );
  INVX3 U3086 ( .A(n4036), .Y(n4070) );
  MUX2IX1 U3087 ( .D0(n1335), .D1(n1336), .S(n3994), .Y(n1632) );
  INVXL U3088 ( .A(n3961), .Y(n4073) );
  MUX2XL U3089 ( .D0(A[272]), .D1(A[784]), .S(n3755), .Y(n3847) );
  MUX2IX1 U3090 ( .D0(A[481]), .D1(A[993]), .S(n4048), .Y(n642) );
  AND2XL U3091 ( .A(n4051), .B(n3775), .Y(n677) );
  AOI22X1 U3092 ( .A(n4060), .B(A[289]), .C(n3788), .D(A[801]), .Y(n3780) );
  AOI22X1 U3093 ( .A(n4058), .B(A[33]), .C(n4046), .D(A[545]), .Y(n3779) );
  AO22XL U3094 ( .A(n4068), .B(A[418]), .C(n3755), .D(A[930]), .Y(n922) );
  INVXL U3095 ( .A(n3848), .Y(n3777) );
  AOI22BX1 U3096 ( .B(n4018), .A(n1045), .D(n3869), .C(n3992), .Y(n3906) );
  INVXL U3097 ( .A(n3823), .Y(n3781) );
  MUX2X1 U3098 ( .D0(n641), .D1(n642), .S(n4018), .Y(n3787) );
  NOR21X1 U3099 ( .B(n4062), .A(A[368]), .Y(n1142) );
  MUX2IX1 U3100 ( .D0(n1141), .D1(n1142), .S(n3975), .Y(n1687) );
  OAI22AX1 U3101 ( .D(n3899), .C(n3791), .A(n3792), .B(n4009), .Y(n1616) );
  AOI22X1 U3102 ( .A(n4070), .B(A[41]), .C(n4048), .D(A[553]), .Y(n3791) );
  AOI22X1 U3103 ( .A(n4069), .B(A[297]), .C(n4073), .D(A[809]), .Y(n3792) );
  INVXL U3104 ( .A(n4071), .Y(n3793) );
  AND2XL U3105 ( .A(n3987), .B(n696), .Y(n3851) );
  MUX2IX1 U3106 ( .D0(n733), .D1(n734), .S(n3981), .Y(n3837) );
  OA22X1 U3107 ( .A(n4046), .B(n3797), .C(n3732), .D(n3798), .Y(n3901) );
  MUX2IX1 U3108 ( .D0(n1499), .D1(n1500), .S(n4019), .Y(n1599) );
  INVXL U3109 ( .A(n3705), .Y(n3846) );
  INVX1 U3110 ( .A(n1531), .Y(n3845) );
  INVXL U3111 ( .A(n4004), .Y(n4017) );
  AND2X2 U3112 ( .A(n4042), .B(n3800), .Y(n1371) );
  BUFXL U3113 ( .A(n3808), .Y(n3801) );
  INVXL U3114 ( .A(n3828), .Y(n3802) );
  INVX2 U3115 ( .A(n4077), .Y(n4064) );
  INVXL U3116 ( .A(n3961), .Y(n4048) );
  MUX2IX1 U3117 ( .D0(n729), .D1(n730), .S(n3982), .Y(n1776) );
  INVX12 U3118 ( .A(n4002), .Y(n3982) );
  INVXL U3119 ( .A(n3710), .Y(n3805) );
  INVX16 U3120 ( .A(A[800]), .Y(n3806) );
  INVX4 U3121 ( .A(n3999), .Y(n3976) );
  INVXL U3122 ( .A(n4051), .Y(n3809) );
  MUX2IX1 U3123 ( .D0(n19), .D1(n27), .S(n3971), .Y(n3) );
  INVXL U3124 ( .A(n3682), .Y(n3813) );
  NOR2XL U3125 ( .A(n4055), .B(A[656]), .Y(n997) );
  INVXL U3126 ( .A(n3710), .Y(n4028) );
  NOR2XL U3127 ( .A(n4061), .B(A[712]), .Y(n733) );
  INVXL U3128 ( .A(n3813), .Y(n3818) );
  AOI22CX1 U3129 ( .C(n1468), .D(n3995), .A(n3819), .B(n3705), .Y(n3825) );
  AOI22X1 U3130 ( .A(n4060), .B(A[32]), .C(n3807), .D(A[544]), .Y(n3819) );
  INVXL U3131 ( .A(n4062), .Y(n3820) );
  INVX1 U3132 ( .A(n4078), .Y(n4062) );
  INVXL U3133 ( .A(n4054), .Y(n3821) );
  NOR2XL U3134 ( .A(n3732), .B(A[968]), .Y(n734) );
  AOI22X1 U3135 ( .A(n4064), .B(A[432]), .C(n3755), .D(A[944]), .Y(n3960) );
  INVXL U3136 ( .A(n4023), .Y(n3823) );
  INVX3 U3137 ( .A(n4064), .Y(n4023) );
  INVXL U3138 ( .A(n3828), .Y(n4031) );
  INVXL U3139 ( .A(n4065), .Y(n3824) );
  OAI22X1 U3140 ( .A(n3900), .B(n3826), .C(n3901), .D(n3899), .Y(n1615) );
  MUX2IX1 U3141 ( .D0(n678), .D1(n677), .S(n3829), .Y(n3836) );
  MUX2IX1 U3142 ( .D0(n1615), .D1(n1631), .S(n3938), .Y(n3832) );
  NOR2XL U3143 ( .A(n4053), .B(A[976]), .Y(n702) );
  INVXL U3144 ( .A(n3823), .Y(n3833) );
  MUX2IX1 U3145 ( .D0(n2), .D1(n10), .S(n3973), .Y(B[1]) );
  INVXL U3146 ( .A(n3823), .Y(n4045) );
  INVXL U3147 ( .A(n3767), .Y(n3842) );
  AOI22AX1 U3148 ( .A(n4013), .B(n873), .D(n3905), .C(n3991), .Y(n3904) );
  MUX2IX1 U3149 ( .D0(n3847), .D1(n3845), .S(n3846), .Y(n3897) );
  AO22XL U3150 ( .A(n4062), .B(A[246]), .C(n4041), .D(A[758]), .Y(n545) );
  AO22XL U3151 ( .A(n4071), .B(A[245]), .C(n4041), .D(A[757]), .Y(n551) );
  NOR21XL U3152 ( .B(n4043), .A(A[520]), .Y(n1563) );
  AO22XL U3153 ( .A(n3718), .B(A[167]), .C(n4075), .D(A[679]), .Y(n891) );
  AO22XL U3154 ( .A(n4068), .B(A[423]), .C(n3682), .D(A[935]), .Y(n892) );
  AO22XL U3155 ( .A(n4067), .B(A[166]), .C(n3683), .D(A[678]), .Y(n897) );
  AO22XL U3156 ( .A(n3718), .B(A[422]), .C(n3682), .D(A[934]), .Y(n898) );
  AO22XL U3157 ( .A(n3718), .B(A[421]), .C(n3683), .D(A[933]), .Y(n904) );
  AO22XL U3158 ( .A(n3710), .B(A[396]), .C(n3801), .D(A[908]), .Y(n1022) );
  AO22XL U3159 ( .A(n4057), .B(A[395]), .C(n3801), .D(A[907]), .Y(n1028) );
  MUX2IX1 U3160 ( .D0(n35), .D1(n43), .S(n3971), .Y(n11) );
  NOR2XL U3161 ( .A(n4039), .B(A[352]), .Y(n1206) );
  AO22XL U3162 ( .A(n4064), .B(A[174]), .C(n4044), .D(A[686]), .Y(n849) );
  AO22XL U3163 ( .A(n4068), .B(A[173]), .C(n4044), .D(A[685]), .Y(n855) );
  AO22XL U3164 ( .A(n4065), .B(A[428]), .C(n4044), .D(A[940]), .Y(n862) );
  AO22XL U3165 ( .A(n4066), .B(A[427]), .C(n4044), .D(A[939]), .Y(n868) );
  INVX8 U3166 ( .A(n3961), .Y(n4079) );
  MUX2X2 U3167 ( .D0(n965), .D1(n966), .S(n3980), .Y(n3862) );
  INVX1 U3168 ( .A(n3950), .Y(n3941) );
  MUX2X1 U3169 ( .D0(n1491), .D1(n1492), .S(n3983), .Y(n3864) );
  INVX2 U3170 ( .A(n4001), .Y(n3983) );
  MUX2X1 U3171 ( .D0(n669), .D1(n670), .S(n3983), .Y(n3870) );
  AOI22X1 U3172 ( .A(n4061), .B(A[506]), .C(n3782), .D(A[1018]), .Y(n3872) );
  MUX2IX1 U3173 ( .D0(n1105), .D1(n1106), .S(n3976), .Y(n1696) );
  AOI22XL U3174 ( .A(n4062), .B(A[498]), .C(n4043), .D(A[1010]), .Y(n3915) );
  AOI22X1 U3175 ( .A(n1408), .B(n3993), .C(n3867), .D(n4007), .Y(n3911) );
  INVXL U3176 ( .A(n4015), .Y(n4010) );
  MUX2IX1 U3177 ( .D0(n3658), .D1(n3851), .S(n3945), .Y(n211) );
  NAND2X1 U3178 ( .A(n3868), .B(n3947), .Y(n114) );
  AO22XL U3179 ( .A(n4058), .B(A[42]), .C(n4048), .D(A[554]), .Y(n3867) );
  MUX2X1 U3180 ( .D0(n725), .D1(n726), .S(n3982), .Y(n3894) );
  OR2X1 U3181 ( .A(n4041), .B(A[442]), .Y(n3896) );
  INVXL U3182 ( .A(n3990), .Y(n4014) );
  INVXL U3183 ( .A(n3828), .Y(n4024) );
  INVXL U3184 ( .A(n4051), .Y(n4041) );
  INVXL U3185 ( .A(n3970), .Y(n3966) );
  INVXL U3186 ( .A(n3970), .Y(n3965) );
  INVXL U3187 ( .A(n3956), .Y(n3955) );
  MUX2IXL U3188 ( .D0(n3852), .D1(n3853), .S(n3945), .Y(n212) );
  MUX2IXL U3189 ( .D0(n3859), .D1(n3857), .S(n3945), .Y(n214) );
  MUX2IXL U3190 ( .D0(n3856), .D1(n3854), .S(n3945), .Y(n213) );
  MUX2IXL U3191 ( .D0(n3858), .D1(n3855), .S(n3686), .Y(n215) );
  MUX2IXL U3192 ( .D0(n3860), .D1(n3861), .S(n3686), .Y(n216) );
  NAND2XL U3193 ( .A(n3897), .B(n3947), .Y(n113) );
  MUX2IX1 U3194 ( .D0(n1197), .D1(n1198), .S(n3978), .Y(n1673) );
  MUX2X1 U3195 ( .D0(n1673), .D1(n1689), .S(n3941), .Y(n163) );
  MUX2IX1 U3196 ( .D0(n3909), .D1(n3865), .S(n3938), .Y(n131) );
  MUX2BX1 U3197 ( .D0(n1641), .D1(n315), .S(n3939), .Y(n147) );
  MUX2IXL U3198 ( .D0(n3894), .D1(n3870), .S(n3944), .Y(n219) );
  MUX2X1 U3199 ( .D0(n1681), .D1(n1697), .S(n3942), .Y(n171) );
  MUX2IXL U3200 ( .D0(n1551), .D1(n1552), .S(n3987), .Y(n1586) );
  AND2XL U3201 ( .A(n3988), .B(n749), .Y(n3852) );
  AND2XL U3202 ( .A(n3988), .B(n693), .Y(n3853) );
  MUX2IXL U3203 ( .D0(n1543), .D1(n1544), .S(n3985), .Y(n1588) );
  AND2XL U3204 ( .A(n3985), .B(n690), .Y(n3854) );
  MUX2BXL U3205 ( .D0(n1685), .D1(n3882), .S(n3942), .Y(n175) );
  MUX2AXL U3206 ( .D0(n3669), .D1(n1629), .S(n3938), .Y(n135) );
  AND2XL U3207 ( .A(n3988), .B(n684), .Y(n3855) );
  AND2XL U3208 ( .A(n3987), .B(n746), .Y(n3856) );
  AND2XL U3209 ( .A(n3985), .B(n687), .Y(n3857) );
  NAND2XL U3210 ( .A(n3985), .B(n1287), .Y(n1646) );
  AND2XL U3211 ( .A(n3988), .B(n740), .Y(n3858) );
  AND2XL U3212 ( .A(n3985), .B(n743), .Y(n3859) );
  AND2XL U3213 ( .A(n3985), .B(n737), .Y(n3860) );
  AND2XL U3214 ( .A(n3985), .B(n681), .Y(n3861) );
  MUX2IXL U3215 ( .D0(A[266]), .D1(A[778]), .S(n4026), .Y(n1556) );
  MUX2XL U3216 ( .D0(n1363), .D1(n1364), .S(n3981), .Y(n3865) );
  MUX2IXL U3217 ( .D0(A[314]), .D1(A[826]), .S(n3682), .Y(n3866) );
  MUX2IXL U3218 ( .D0(A[410]), .D1(A[922]), .S(n4022), .Y(n958) );
  MUX2IX1 U3219 ( .D0(n1237), .D1(n1238), .S(n3979), .Y(n1663) );
  MUX2IX1 U3220 ( .D0(n989), .D1(n990), .S(n3984), .Y(n1721) );
  MUX2IX1 U3221 ( .D0(n1133), .D1(n1134), .S(n3975), .Y(n1689) );
  NOR2XL U3222 ( .A(n4076), .B(A[129]), .Y(n1073) );
  AOI22X1 U3223 ( .A(n4068), .B(A[392]), .C(n4076), .D(A[904]), .Y(n3869) );
  INVXL U3224 ( .A(n1657), .Y(n315) );
  INVXL U3225 ( .A(n1649), .Y(n307) );
  MUX2X1 U3226 ( .D0(n605), .D1(n606), .S(n3994), .Y(n3871) );
  MUX2XL U3227 ( .D0(n1229), .D1(n1230), .S(n3980), .Y(n3891) );
  MUX2IXL U3228 ( .D0(A[274]), .D1(A[786]), .S(n3696), .Y(n3873) );
  NOR2XL U3229 ( .A(n4040), .B(A[131]), .Y(n1065) );
  MUX2XL U3230 ( .D0(n1519), .D1(n1520), .S(n3680), .Y(n3876) );
  AO22XL U3231 ( .A(n3823), .B(A[419]), .C(n4075), .D(A[931]), .Y(n916) );
  AO22XL U3232 ( .A(n4071), .B(A[499]), .C(n3766), .D(A[1011]), .Y(n564) );
  AO22XL U3233 ( .A(n3823), .B(A[507]), .C(n3802), .D(A[1019]), .Y(n516) );
  AND2XL U3234 ( .A(n3987), .B(n1299), .Y(n3877) );
  AO22XL U3235 ( .A(n3813), .B(A[179]), .C(n4045), .D(A[691]), .Y(n819) );
  NOR2XL U3236 ( .A(n4040), .B(A[133]), .Y(n1057) );
  NOR2XL U3237 ( .A(n4040), .B(A[132]), .Y(n1061) );
  MUX2XL U3238 ( .D0(n1515), .D1(n1516), .S(n3680), .Y(n3878) );
  AO22XL U3239 ( .A(n4067), .B(A[420]), .C(n3768), .D(A[932]), .Y(n910) );
  AO22XL U3240 ( .A(n4063), .B(A[436]), .C(n3820), .D(A[948]), .Y(n814) );
  AO22XL U3241 ( .A(n4062), .B(A[244]), .C(n4041), .D(A[756]), .Y(n557) );
  AO22XL U3242 ( .A(n4061), .B(A[252]), .C(n4041), .D(A[764]), .Y(n509) );
  MUX2XL U3243 ( .D0(n1539), .D1(n1540), .S(n3680), .Y(n3879) );
  MUX2XL U3244 ( .D0(n765), .D1(n766), .S(n3981), .Y(n3880) );
  MUX2XL U3245 ( .D0(n761), .D1(n762), .S(n3796), .Y(n3881) );
  MUX2XL U3246 ( .D0(n1085), .D1(n1086), .S(n3977), .Y(n3882) );
  MUX2XL U3247 ( .D0(n769), .D1(n770), .S(n3672), .Y(n3883) );
  MUX2XL U3248 ( .D0(n1315), .D1(n1316), .S(n3984), .Y(n3884) );
  NOR2XL U3249 ( .A(n4040), .B(A[358]), .Y(n1182) );
  NOR2XL U3250 ( .A(n4040), .B(A[134]), .Y(n1053) );
  NOR2XL U3251 ( .A(n3818), .B(A[351]), .Y(n1210) );
  MUX2XL U3252 ( .D0(n1511), .D1(n1512), .S(n3681), .Y(n3885) );
  MUX2XL U3253 ( .D0(n1503), .D1(n1504), .S(n3681), .Y(n3886) );
  MUX2XL U3254 ( .D0(n1117), .D1(n1118), .S(n3976), .Y(n3887) );
  MUX2XL U3255 ( .D0(n1475), .D1(n1476), .S(n3982), .Y(n3888) );
  AO22XL U3256 ( .A(n3777), .B(A[503]), .C(n3805), .D(A[1015]), .Y(n540) );
  AO22XL U3257 ( .A(n3777), .B(A[254]), .C(n3766), .D(A[766]), .Y(n497) );
  AO22XL U3258 ( .A(n3718), .B(A[255]), .C(n3766), .D(A[767]), .Y(n491) );
  AO22XL U3259 ( .A(n3777), .B(A[429]), .C(n4044), .D(A[941]), .Y(n856) );
  AO22XL U3260 ( .A(n4057), .B(A[302]), .C(n3802), .D(A[814]), .Y(n1384) );
  AO22XL U3261 ( .A(n4059), .B(A[294]), .C(n4047), .D(A[806]), .Y(n1432) );
  AO22XL U3262 ( .A(n4071), .B(A[501]), .C(n4041), .D(A[1013]), .Y(n552) );
  AO22XL U3263 ( .A(n4062), .B(A[502]), .C(n4041), .D(A[1014]), .Y(n546) );
  AO22XL U3264 ( .A(n3718), .B(A[509]), .C(n3824), .D(A[1021]), .Y(n504) );
  AND2XL U3265 ( .A(n3987), .B(n1293), .Y(n3889) );
  AND2XL U3266 ( .A(n3985), .B(n1296), .Y(n3890) );
  AO22XL U3267 ( .A(n4064), .B(A[430]), .C(n4044), .D(A[942]), .Y(n850) );
  AO22XL U3268 ( .A(n3718), .B(A[431]), .C(n4045), .D(A[943]), .Y(n844) );
  INVX1 U3269 ( .A(n4000), .Y(n3987) );
  INVX1 U3270 ( .A(n3998), .Y(n3991) );
  INVX1 U3271 ( .A(n4016), .Y(n4007) );
  INVX1 U3272 ( .A(n1654), .Y(n312) );
  INVX1 U3273 ( .A(n3828), .Y(n4035) );
  INVXL U3274 ( .A(n4051), .Y(n4047) );
  INVX1 U3275 ( .A(n3950), .Y(n3942) );
  INVX1 U3276 ( .A(n3951), .Y(n3938) );
  INVX1 U3277 ( .A(n3956), .Y(n3954) );
  NAND2XL U3278 ( .A(n3953), .B(n3963), .Y(n3962) );
  MUX2IXL U3279 ( .D0(n163), .D1(n171), .S(n3966), .Y(n75) );
  INVX1 U3280 ( .A(SH[4]), .Y(n3950) );
  INVX1 U3281 ( .A(SH[5]), .Y(n3956) );
  INVX1 U3282 ( .A(SH[5]), .Y(n3957) );
  INVX1 U3283 ( .A(SH[3]), .Y(n3969) );
  MUX2IXL U3284 ( .D0(n100), .D1(n108), .S(n3954), .Y(n44) );
  MUX2IXL U3285 ( .D0(n212), .D1(n220), .S(n3964), .Y(n100) );
  MUX2IXL U3286 ( .D0(n228), .D1(n236), .S(n3816), .Y(n108) );
  MUX2IXL U3287 ( .D0(n101), .D1(n109), .S(n3955), .Y(n45) );
  MUX2IXL U3288 ( .D0(n213), .D1(n221), .S(n3964), .Y(n101) );
  MUX2IXL U3289 ( .D0(n229), .D1(n237), .S(n3816), .Y(n109) );
  MUX2IXL U3290 ( .D0(n23), .D1(n31), .S(n3971), .Y(n7) );
  MUX2IXL U3291 ( .D0(n71), .D1(n79), .S(n3954), .Y(n31) );
  MUX2IXL U3292 ( .D0(n55), .D1(n63), .S(n3747), .Y(n23) );
  MUX2IXL U3293 ( .D0(n151), .D1(n159), .S(n3967), .Y(n71) );
  MUX2IXL U3294 ( .D0(n102), .D1(n110), .S(n3954), .Y(n46) );
  MUX2IXL U3295 ( .D0(n214), .D1(n222), .S(n3964), .Y(n102) );
  MUX2IXL U3296 ( .D0(n230), .D1(n238), .S(n3816), .Y(n110) );
  MUX2IXL U3297 ( .D0(n103), .D1(n111), .S(n3955), .Y(n47) );
  MUX2IXL U3298 ( .D0(n215), .D1(n223), .S(n3816), .Y(n103) );
  MUX2IXL U3299 ( .D0(n231), .D1(n239), .S(n3816), .Y(n111) );
  MUX2IXL U3300 ( .D0(n104), .D1(n112), .S(n3954), .Y(n48) );
  MUX2IXL U3301 ( .D0(n216), .D1(n224), .S(n3816), .Y(n104) );
  MUX2IXL U3302 ( .D0(n232), .D1(n240), .S(n3816), .Y(n112) );
  NOR21XL U3303 ( .B(n4026), .A(A[962]), .Y(n752) );
  MUX2IX1 U3304 ( .D0(n147), .D1(n155), .S(n3967), .Y(n67) );
  MUX2IX1 U3305 ( .D0(n307), .D1(n3891), .S(n3940), .Y(n155) );
  MUX2X2 U3306 ( .D0(n1705), .D1(n1721), .S(n3941), .Y(n179) );
  MUX2IX1 U3307 ( .D0(n1339), .D1(n1340), .S(n3981), .Y(n1631) );
  MUX2X2 U3308 ( .D0(n1713), .D1(n1729), .S(n3694), .Y(n187) );
  MUX2IX1 U3309 ( .D0(n131), .D1(n139), .S(n3968), .Y(n59) );
  MUX2IX1 U3310 ( .D0(n1563), .D1(n1564), .S(n3984), .Y(n1583) );
  MUX2IXL U3311 ( .D0(n1165), .D1(n1166), .S(n3975), .Y(n1681) );
  MUX2IXL U3312 ( .D0(n3656), .D1(n3864), .S(n3676), .Y(n123) );
  MUX2XL U3313 ( .D0(n1706), .D1(n1722), .S(n3941), .Y(n180) );
  MUX2IXL U3314 ( .D0(n985), .D1(n986), .S(n4018), .Y(n1722) );
  MUX2IXL U3315 ( .D0(n84), .D1(n92), .S(n3955), .Y(n36) );
  MUX2IXL U3316 ( .D0(n196), .D1(n204), .S(n3965), .Y(n92) );
  MUX2IXL U3317 ( .D0(n180), .D1(n188), .S(n3965), .Y(n84) );
  MUX2IXL U3318 ( .D0(n3662), .D1(n3651), .S(n3945), .Y(n196) );
  NOR21XL U3319 ( .B(n4030), .A(A[979]), .Y(n693) );
  MUX2XL U3320 ( .D0(n1802), .D1(n1818), .S(n3945), .Y(n228) );
  MUX2IXL U3321 ( .D0(n633), .D1(n634), .S(n3679), .Y(n1802) );
  MUX2XL U3322 ( .D0(n1610), .D1(n1626), .S(n3938), .Y(n132) );
  MUX2IXL U3323 ( .D0(n1359), .D1(n1360), .S(n3982), .Y(n1626) );
  MUX2XL U3324 ( .D0(n1674), .D1(n1690), .S(n3941), .Y(n164) );
  MUX2IX1 U3325 ( .D0(n1129), .D1(n1130), .S(n3976), .Y(n1690) );
  MUX2IXL U3326 ( .D0(n52), .D1(n60), .S(n3954), .Y(n20) );
  MUX2IXL U3327 ( .D0(n116), .D1(n124), .S(n3965), .Y(n52) );
  MUX2IXL U3328 ( .D0(n132), .D1(n140), .S(n3968), .Y(n60) );
  NAND2XL U3329 ( .A(n3876), .B(n3947), .Y(n116) );
  MUX2XL U3330 ( .D0(n1714), .D1(n1730), .S(n3694), .Y(n188) );
  MUX2IX1 U3331 ( .D0(n953), .D1(n954), .S(n3681), .Y(n1730) );
  MUX2XL U3332 ( .D0(n1746), .D1(n1762), .S(n3945), .Y(n204) );
  MUX2IXL U3333 ( .D0(n777), .D1(n778), .S(n3673), .Y(n1762) );
  MUX2XL U3334 ( .D0(n1778), .D1(n1794), .S(n3945), .Y(n220) );
  MUX2IXL U3335 ( .D0(n721), .D1(n722), .S(n3982), .Y(n1778) );
  MUX2XL U3336 ( .D0(n1618), .D1(n1634), .S(n3938), .Y(n140) );
  MUX2IXL U3337 ( .D0(n1327), .D1(n1328), .S(n3984), .Y(n1634) );
  MUX2XL U3338 ( .D0(n1586), .D1(n1602), .S(n3676), .Y(n124) );
  MUX2XL U3339 ( .D0(n1682), .D1(n1698), .S(n3942), .Y(n172) );
  MUX2IXL U3340 ( .D0(n1161), .D1(n1162), .S(n3975), .Y(n1682) );
  MUX2XL U3341 ( .D0(n1650), .D1(n1666), .S(n3940), .Y(n156) );
  NOR21XL U3342 ( .B(n4037), .A(A[971]), .Y(n722) );
  MUX2XL U3343 ( .D0(n1810), .D1(n1826), .S(n3947), .Y(n236) );
  MUX2IXL U3344 ( .D0(n601), .D1(n602), .S(n3679), .Y(n1810) );
  MUX2IXL U3345 ( .D0(n68), .D1(n76), .S(n3747), .Y(n28) );
  MUX2IXL U3346 ( .D0(n148), .D1(n156), .S(n3967), .Y(n68) );
  MUX2IXL U3347 ( .D0(n164), .D1(n172), .S(n3966), .Y(n76) );
  MUX2IXL U3348 ( .D0(n3877), .D1(n316), .S(n3939), .Y(n148) );
  NOR21XL U3349 ( .B(n3721), .A(A[963]), .Y(n749) );
  MUX2XL U3350 ( .D0(n1707), .D1(n1723), .S(n3694), .Y(n181) );
  MUX2IXL U3351 ( .D0(n981), .D1(n982), .S(n3979), .Y(n1723) );
  MUX2XL U3352 ( .D0(n1803), .D1(n1819), .S(n3946), .Y(n229) );
  MUX2IXL U3353 ( .D0(n629), .D1(n630), .S(n3984), .Y(n1803) );
  MUX2XL U3354 ( .D0(n1611), .D1(n1627), .S(n3938), .Y(n133) );
  MUX2IXL U3355 ( .D0(n1355), .D1(n1356), .S(n3981), .Y(n1627) );
  MUX2IXL U3356 ( .D0(n85), .D1(n93), .S(n3954), .Y(n37) );
  MUX2IXL U3357 ( .D0(n197), .D1(n205), .S(n3964), .Y(n93) );
  MUX2IXL U3358 ( .D0(n181), .D1(n189), .S(n3967), .Y(n85) );
  MUX2IXL U3359 ( .D0(n3649), .D1(n3663), .S(n3939), .Y(n197) );
  MUX2IXL U3360 ( .D0(n53), .D1(n61), .S(n3747), .Y(n21) );
  MUX2IXL U3361 ( .D0(n117), .D1(n125), .S(n3968), .Y(n53) );
  MUX2IXL U3362 ( .D0(n133), .D1(n141), .S(n3968), .Y(n61) );
  NAND2XL U3363 ( .A(n3878), .B(n3948), .Y(n117) );
  MUX2XL U3364 ( .D0(n1715), .D1(n1731), .S(n3694), .Y(n189) );
  MUX2IX1 U3365 ( .D0(n949), .D1(n950), .S(n3681), .Y(n1731) );
  MUX2XL U3366 ( .D0(n1747), .D1(n1763), .S(n3946), .Y(n205) );
  MUX2IXL U3367 ( .D0(n773), .D1(n774), .S(n3673), .Y(n1763) );
  MUX2XL U3368 ( .D0(n1811), .D1(n1827), .S(n3946), .Y(n237) );
  MUX2IXL U3369 ( .D0(n597), .D1(n598), .S(n4018), .Y(n1811) );
  MUX2XL U3370 ( .D0(n1619), .D1(n1635), .S(n3939), .Y(n141) );
  MUX2IXL U3371 ( .D0(n1323), .D1(n1324), .S(n3980), .Y(n1635) );
  MUX2XL U3372 ( .D0(n1683), .D1(n1699), .S(n3942), .Y(n173) );
  MUX2IX1 U3373 ( .D0(n1093), .D1(n1094), .S(n3976), .Y(n1699) );
  MUX2IXL U3374 ( .D0(n69), .D1(n77), .S(n3954), .Y(n29) );
  MUX2IXL U3375 ( .D0(n149), .D1(n157), .S(n3967), .Y(n69) );
  MUX2IXL U3376 ( .D0(n165), .D1(n173), .S(n3966), .Y(n77) );
  MUX2IXL U3377 ( .D0(n3890), .D1(n317), .S(n3939), .Y(n149) );
  NOR21XL U3378 ( .B(n3821), .A(A[980]), .Y(n690) );
  MUX2XL U3379 ( .D0(n1612), .D1(n1628), .S(n3938), .Y(n134) );
  MUX2IXL U3380 ( .D0(n1351), .D1(n1352), .S(n3981), .Y(n1628) );
  MUX2XL U3381 ( .D0(n1676), .D1(n1692), .S(n3941), .Y(n166) );
  MUX2IX1 U3382 ( .D0(n1121), .D1(n1122), .S(n3976), .Y(n1692) );
  MUX2XL U3383 ( .D0(n1708), .D1(n1724), .S(n3694), .Y(n182) );
  MUX2IXL U3384 ( .D0(n977), .D1(n978), .S(n3984), .Y(n1724) );
  MUX2XL U3385 ( .D0(n1740), .D1(n1756), .S(n3686), .Y(n198) );
  MUX2XL U3386 ( .D0(n1804), .D1(n1820), .S(n3686), .Y(n230) );
  MUX2IXL U3387 ( .D0(n625), .D1(n626), .S(n3680), .Y(n1804) );
  MUX2XL U3388 ( .D0(n1675), .D1(n1691), .S(n3941), .Y(n165) );
  MUX2IX1 U3389 ( .D0(n1125), .D1(n1126), .S(n3976), .Y(n1691) );
  MUX2XL U3390 ( .D0(n1709), .D1(n1725), .S(n3694), .Y(n183) );
  MUX2IXL U3391 ( .D0(n973), .D1(n974), .S(n3979), .Y(n1725) );
  MUX2XL U3392 ( .D0(n1741), .D1(n1757), .S(n3945), .Y(n199) );
  MUX2XL U3393 ( .D0(n1805), .D1(n1821), .S(n3676), .Y(n231) );
  MUX2IXL U3394 ( .D0(n621), .D1(n622), .S(n4018), .Y(n1805) );
  MUX2IXL U3395 ( .D0(n54), .D1(n62), .S(n3747), .Y(n22) );
  MUX2IXL U3396 ( .D0(n118), .D1(n126), .S(n3968), .Y(n54) );
  MUX2IXL U3397 ( .D0(n134), .D1(n142), .S(n3968), .Y(n62) );
  NAND2XL U3398 ( .A(n3885), .B(n3948), .Y(n118) );
  MUX2IXL U3399 ( .D0(n86), .D1(n94), .S(n3954), .Y(n38) );
  MUX2IXL U3400 ( .D0(n198), .D1(n206), .S(n3964), .Y(n94) );
  MUX2IXL U3401 ( .D0(n182), .D1(n190), .S(n3967), .Y(n86) );
  MUX2IXL U3402 ( .D0(n3665), .D1(n3883), .S(n3686), .Y(n206) );
  MUX2XL U3403 ( .D0(n1620), .D1(n1636), .S(n3939), .Y(n142) );
  MUX2IXL U3404 ( .D0(n1319), .D1(n1320), .S(n4018), .Y(n1636) );
  MUX2XL U3405 ( .D0(n1588), .D1(n1604), .S(n3676), .Y(n126) );
  MUX2XL U3406 ( .D0(n1684), .D1(n1700), .S(n3942), .Y(n174) );
  MUX2IXL U3407 ( .D0(n1089), .D1(n1090), .S(n3977), .Y(n1700) );
  MUX2XL U3408 ( .D0(n1652), .D1(n1668), .S(n3940), .Y(n158) );
  MUX2XL U3409 ( .D0(n1716), .D1(n1732), .S(n3942), .Y(n190) );
  MUX2IX1 U3410 ( .D0(n945), .D1(n946), .S(n3681), .Y(n1732) );
  MUX2XL U3411 ( .D0(n1780), .D1(n1796), .S(n3946), .Y(n222) );
  MUX2IXL U3412 ( .D0(n713), .D1(n714), .S(n3982), .Y(n1780) );
  MUX2XL U3413 ( .D0(n1779), .D1(n1795), .S(n3946), .Y(n221) );
  MUX2IXL U3414 ( .D0(n717), .D1(n718), .S(n3982), .Y(n1779) );
  MUX2XL U3415 ( .D0(n1587), .D1(n1603), .S(n3676), .Y(n125) );
  MUX2IX1 U3416 ( .D0(n1547), .D1(n1548), .S(n3680), .Y(n1587) );
  MUX2XL U3417 ( .D0(n1651), .D1(n1667), .S(n3940), .Y(n157) );
  MUX2XL U3418 ( .D0(n1717), .D1(n1733), .S(n3686), .Y(n191) );
  MUX2IX1 U3419 ( .D0(n941), .D1(n942), .S(n3680), .Y(n1733) );
  MUX2XL U3420 ( .D0(n1813), .D1(n1829), .S(n3946), .Y(n239) );
  MUX2IXL U3421 ( .D0(n589), .D1(n590), .S(n3680), .Y(n1813) );
  MUX2IXL U3422 ( .D0(n70), .D1(n78), .S(n3955), .Y(n30) );
  MUX2IXL U3423 ( .D0(n150), .D1(n158), .S(n3967), .Y(n70) );
  MUX2IXL U3424 ( .D0(n166), .D1(n174), .S(n3966), .Y(n78) );
  MUX2IXL U3425 ( .D0(n3889), .D1(n318), .S(n3938), .Y(n150) );
  MUX2IXL U3426 ( .D0(n135), .D1(n143), .S(n3967), .Y(n63) );
  MUX2IXL U3427 ( .D0(n3664), .D1(n3884), .S(n3939), .Y(n143) );
  NOR21XL U3428 ( .B(n3766), .A(A[972]), .Y(n718) );
  MUX2XL U3429 ( .D0(n1812), .D1(n1828), .S(n3947), .Y(n238) );
  MUX2IX1 U3430 ( .D0(n593), .D1(n594), .S(n3680), .Y(n1812) );
  MUX2IXL U3431 ( .D0(n167), .D1(n175), .S(n3966), .Y(n79) );
  MUX2IXL U3432 ( .D0(n3931), .D1(n3887), .S(n3941), .Y(n167) );
  MUX2IXL U3433 ( .D0(n87), .D1(n95), .S(n3955), .Y(n39) );
  MUX2IXL U3434 ( .D0(n199), .D1(n207), .S(n3964), .Y(n95) );
  MUX2IXL U3435 ( .D0(n183), .D1(n191), .S(n3966), .Y(n87) );
  MUX2IXL U3436 ( .D0(n3667), .D1(n3880), .S(n3686), .Y(n207) );
  NOR21XL U3437 ( .B(n3721), .A(A[964]), .Y(n746) );
  NOR21XL U3438 ( .B(n3758), .A(A[981]), .Y(n687) );
  NOR21XL U3439 ( .B(n3821), .A(A[982]), .Y(n684) );
  MUX2XL U3440 ( .D0(n1645), .D1(n1661), .S(n3940), .Y(n151) );
  NAND2XL U3441 ( .A(n3985), .B(n1290), .Y(n1645) );
  MUX2XL U3442 ( .D0(n1614), .D1(n1630), .S(n3938), .Y(n136) );
  MUX2IXL U3443 ( .D0(n1343), .D1(n1344), .S(n3981), .Y(n1630) );
  MUX2XL U3444 ( .D0(n1678), .D1(n1694), .S(n3941), .Y(n168) );
  MUX2IX1 U3445 ( .D0(n1113), .D1(n1114), .S(n3976), .Y(n1694) );
  MUX2XL U3446 ( .D0(n1646), .D1(n1662), .S(n3940), .Y(n152) );
  MUX2XL U3447 ( .D0(n1710), .D1(n1726), .S(n3694), .Y(n184) );
  MUX2IXL U3448 ( .D0(n1049), .D1(n1050), .S(n3978), .Y(n1710) );
  MUX2XL U3449 ( .D0(n1742), .D1(n1758), .S(n3694), .Y(n200) );
  MUX2IXL U3450 ( .D0(n56), .D1(n64), .S(n3747), .Y(n24) );
  MUX2IXL U3451 ( .D0(n120), .D1(n128), .S(n3968), .Y(n56) );
  MUX2IXL U3452 ( .D0(n136), .D1(n144), .S(n3967), .Y(n64) );
  NAND2XL U3453 ( .A(n3886), .B(n3947), .Y(n120) );
  MUX2IXL U3454 ( .D0(n88), .D1(n96), .S(n3955), .Y(n40) );
  MUX2IXL U3455 ( .D0(n200), .D1(n208), .S(n3964), .Y(n96) );
  MUX2IXL U3456 ( .D0(n184), .D1(n192), .S(n3966), .Y(n88) );
  MUX2IXL U3457 ( .D0(n3668), .D1(n3881), .S(n3686), .Y(n208) );
  MUX2XL U3458 ( .D0(n1653), .D1(n1669), .S(n3939), .Y(n159) );
  MUX2IX1 U3459 ( .D0(n1213), .D1(n1214), .S(n3681), .Y(n1669) );
  MUX2XL U3460 ( .D0(n1781), .D1(n1797), .S(n3946), .Y(n223) );
  MUX2IXL U3461 ( .D0(n709), .D1(n710), .S(n3981), .Y(n1781) );
  MUX2IXL U3462 ( .D0(n119), .D1(n127), .S(n3968), .Y(n55) );
  NAND2XL U3463 ( .A(n3666), .B(n3948), .Y(n119) );
  MUX2IXL U3464 ( .D0(n3879), .D1(n3888), .S(n3676), .Y(n127) );
  MUX2XL U3465 ( .D0(n1622), .D1(n1638), .S(n3939), .Y(n144) );
  MUX2IXL U3466 ( .D0(n1311), .D1(n1312), .S(n3979), .Y(n1638) );
  MUX2XL U3467 ( .D0(n1590), .D1(n1606), .S(n3676), .Y(n128) );
  MUX2IXL U3468 ( .D0(n1471), .D1(n1472), .S(n3983), .Y(n1606) );
  MUX2XL U3469 ( .D0(n1686), .D1(n1702), .S(n3942), .Y(n176) );
  MUX2IXL U3470 ( .D0(n1081), .D1(n1082), .S(n3977), .Y(n1702) );
  MUX2XL U3471 ( .D0(n1718), .D1(n1734), .S(n3945), .Y(n192) );
  MUX2IX1 U3472 ( .D0(n937), .D1(n938), .S(n3681), .Y(n1734) );
  MUX2XL U3473 ( .D0(n1814), .D1(n1830), .S(n3946), .Y(n240) );
  MUX2IX1 U3474 ( .D0(n585), .D1(n586), .S(n3680), .Y(n1814) );
  MUX2XL U3475 ( .D0(n1782), .D1(n1798), .S(n3946), .Y(n224) );
  MUX2IXL U3476 ( .D0(n705), .D1(n706), .S(n3983), .Y(n1782) );
  MUX2IXL U3477 ( .D0(n72), .D1(n80), .S(n3954), .Y(n32) );
  MUX2IXL U3478 ( .D0(n152), .D1(n160), .S(n3967), .Y(n72) );
  MUX2IXL U3479 ( .D0(n168), .D1(n176), .S(n3966), .Y(n80) );
  MUX2IXL U3480 ( .D0(n312), .D1(n3936), .S(n3939), .Y(n160) );
  MUX2XL U3481 ( .D0(n1806), .D1(n1822), .S(n3947), .Y(n232) );
  MUX2IXL U3482 ( .D0(n617), .D1(n618), .S(n3984), .Y(n1806) );
  NOR21XL U3483 ( .B(n4028), .A(A[973]), .Y(n714) );
  NOR21XL U3484 ( .B(n3818), .A(A[974]), .Y(n710) );
  NOR21XL U3485 ( .B(n3781), .A(A[975]), .Y(n706) );
  NOR21XL U3486 ( .B(n3721), .A(A[965]), .Y(n743) );
  NOR21XL U3487 ( .B(n3721), .A(A[966]), .Y(n740) );
  NOR21XL U3488 ( .B(n3721), .A(A[967]), .Y(n737) );
  NOR21XL U3489 ( .B(n3769), .A(A[983]), .Y(n681) );
  MUX2IXL U3490 ( .D0(n613), .D1(n614), .S(n3986), .Y(n1807) );
  NOR21XL U3491 ( .B(n4029), .A(A[658]), .Y(n989) );
  MUX2IX1 U3492 ( .D0(n1077), .D1(n1078), .S(n3977), .Y(n1703) );
  NOR21XL U3493 ( .B(n4044), .A(A[522]), .Y(n1555) );
  MUX2IXL U3494 ( .D0(A[490]), .D1(A[1002]), .S(n4023), .Y(n606) );
  NOR21XL U3495 ( .B(n4037), .A(A[626]), .Y(n1133) );
  NOR21XL U3496 ( .B(n3755), .A(A[832]), .Y(n1308) );
  NAND2X1 U3497 ( .A(n3987), .B(n1302), .Y(n1641) );
  NOR21XL U3498 ( .B(n3683), .A(A[834]), .Y(n1302) );
  NOR21XL U3499 ( .B(n4047), .A(A[610]), .Y(n1197) );
  NOR21XL U3500 ( .B(n3677), .A(A[666]), .Y(n957) );
  NOR21XL U3501 ( .B(n3682), .A(A[618]), .Y(n1165) );
  NOR21XL U3502 ( .B(n4029), .A(A[584]), .Y(n1284) );
  MUX2IXL U3503 ( .D0(A[273]), .D1(A[785]), .S(n4039), .Y(n1528) );
  NOR21XL U3504 ( .B(n3684), .A(A[529]), .Y(n1527) );
  NOR21XL U3505 ( .B(n4029), .A(A[586]), .Y(n1278) );
  NOR21XL U3506 ( .B(n3808), .A(A[594]), .Y(n1256) );
  MUX2IXL U3507 ( .D0(A[306]), .D1(A[818]), .S(n4027), .Y(n1364) );
  NOR21XL U3508 ( .B(n3696), .A(A[562]), .Y(n1363) );
  MUX2IXL U3509 ( .D0(A[282]), .D1(A[794]), .S(n4026), .Y(n1492) );
  NOR21XL U3510 ( .B(n4042), .A(A[833]), .Y(n1305) );
  MUX2IXL U3511 ( .D0(n1065), .D1(n1066), .S(n3977), .Y(n1706) );
  MUX2IXL U3512 ( .D0(n4), .D1(n12), .S(n3973), .Y(B[3]) );
  MUX2IXL U3513 ( .D0(n20), .D1(n28), .S(SH[6]), .Y(n4) );
  MUX2IXL U3514 ( .D0(n36), .D1(n44), .S(n3971), .Y(n12) );
  AO22AXL U3515 ( .A(n868), .B(n3992), .C(n4014), .D(n3917), .Y(n1746) );
  AOI22XL U3516 ( .A(n4067), .B(A[171]), .C(n4044), .D(A[683]), .Y(n3917) );
  AO22AXL U3517 ( .A(n1450), .B(n3994), .C(n4011), .D(n3918), .Y(n1610) );
  AOI22XL U3518 ( .A(n3718), .B(A[35]), .C(n3820), .D(A[547]), .Y(n3918) );
  MUX2IXL U3519 ( .D0(n1487), .D1(n1488), .S(n3983), .Y(n1602) );
  MUX2IXL U3520 ( .D0(A[283]), .D1(A[795]), .S(n3818), .Y(n1488) );
  NOR21XL U3521 ( .B(n3781), .A(A[539]), .Y(n1487) );
  MUX2IXL U3522 ( .D0(n1193), .D1(n1194), .S(n3978), .Y(n1674) );
  NOR21XL U3523 ( .B(n4049), .A(A[611]), .Y(n1193) );
  MUX2IXL U3524 ( .D0(n1225), .D1(n1226), .S(n3979), .Y(n1666) );
  NOR21XL U3525 ( .B(n3801), .A(A[603]), .Y(n1225) );
  NOR21XL U3526 ( .B(n4035), .A(A[531]), .Y(n1519) );
  MUX2IX1 U3527 ( .D0(A[275]), .D1(A[787]), .S(n4024), .Y(n1520) );
  INVX1 U3528 ( .A(n1658), .Y(n316) );
  NOR21XL U3529 ( .B(n3802), .A(A[595]), .Y(n1253) );
  NOR21XL U3530 ( .B(n3769), .A(A[563]), .Y(n1359) );
  NOR21XL U3531 ( .B(n3821), .A(A[627]), .Y(n1129) );
  NOR21XL U3532 ( .B(n4030), .A(A[659]), .Y(n985) );
  NOR21XL U3533 ( .B(n4027), .A(A[667]), .Y(n953) );
  NOR21XL U3534 ( .B(n4075), .A(A[715]), .Y(n721) );
  NOR21XL U3535 ( .B(n3793), .A(A[571]), .Y(n1327) );
  NOR21XL U3536 ( .B(n4035), .A(A[523]), .Y(n1551) );
  NOR21XL U3537 ( .B(n3821), .A(A[619]), .Y(n1161) );
  MUX2IXL U3538 ( .D0(A[187]), .D1(A[699]), .S(n4023), .Y(n777) );
  MUX2IXL U3539 ( .D0(n1097), .D1(n1098), .S(n3976), .Y(n1698) );
  MUX2IXL U3540 ( .D0(A[123]), .D1(A[635]), .S(n3769), .Y(n1097) );
  MUX2IXL U3541 ( .D0(A[403]), .D1(A[915]), .S(n4022), .Y(n986) );
  MUX2IXL U3542 ( .D0(A[411]), .D1(A[923]), .S(n4022), .Y(n954) );
  MUX2IX1 U3543 ( .D0(A[483]), .D1(A[995]), .S(n4024), .Y(n634) );
  MUX2IXL U3544 ( .D0(A[315]), .D1(A[827]), .S(n3801), .Y(n1328) );
  MUX2IXL U3545 ( .D0(A[307]), .D1(A[819]), .S(n4075), .Y(n1360) );
  MUX2IXL U3546 ( .D0(A[267]), .D1(A[779]), .S(n4028), .Y(n1552) );
  MUX2IXL U3547 ( .D0(n665), .D1(n666), .S(n3673), .Y(n1794) );
  MUX2IXL U3548 ( .D0(A[475]), .D1(A[987]), .S(n4025), .Y(n666) );
  NOR21XL U3549 ( .B(n3821), .A(A[587]), .Y(n1275) );
  AO22AXL U3550 ( .A(n1028), .B(n3673), .C(n4011), .D(n3919), .Y(n1714) );
  AOI22XL U3551 ( .A(n4057), .B(A[139]), .C(n3801), .D(A[651]), .Y(n3919) );
  AO22AXL U3552 ( .A(n1402), .B(n3993), .C(n4005), .D(n3920), .Y(n1618) );
  AOI22XL U3553 ( .A(n4069), .B(A[43]), .C(n4033), .D(A[555]), .Y(n3920) );
  NOR21XL U3554 ( .B(n3769), .A(A[835]), .Y(n1299) );
  AO22AXL U3555 ( .A(n1022), .B(n3673), .C(n4006), .D(n3921), .Y(n1715) );
  AOI22XL U3556 ( .A(n3718), .B(A[140]), .C(n3801), .D(A[652]), .Y(n3921) );
  AO22AXL U3557 ( .A(n862), .B(n3991), .C(n4013), .D(n3922), .Y(n1747) );
  AOI22XL U3558 ( .A(n4065), .B(A[172]), .C(n4044), .D(A[684]), .Y(n3922) );
  AO22AXL U3559 ( .A(n1396), .B(n3994), .C(n4006), .D(n3923), .Y(n1619) );
  AOI22XL U3560 ( .A(n4058), .B(A[44]), .C(n3808), .D(A[556]), .Y(n3923) );
  AO22AXL U3561 ( .A(n1444), .B(n3994), .C(n4008), .D(n3924), .Y(n1611) );
  AOI22XL U3562 ( .A(n4059), .B(A[36]), .C(n4047), .D(A[548]), .Y(n3924) );
  MUX2IXL U3563 ( .D0(n1061), .D1(n1062), .S(n3977), .Y(n1707) );
  MUX2IXL U3564 ( .D0(n1157), .D1(n1158), .S(n3975), .Y(n1683) );
  NOR21XL U3565 ( .B(n4030), .A(A[620]), .Y(n1157) );
  MUX2IXL U3566 ( .D0(n5), .D1(n13), .S(n3973), .Y(B[4]) );
  MUX2IXL U3567 ( .D0(n21), .D1(n29), .S(SH[6]), .Y(n5) );
  MUX2IXL U3568 ( .D0(n37), .D1(n45), .S(n3971), .Y(n13) );
  AO22AXL U3569 ( .A(n1438), .B(n3994), .C(n4014), .D(n3925), .Y(n1612) );
  AOI22XL U3570 ( .A(n4070), .B(A[37]), .C(n4047), .D(A[549]), .Y(n3925) );
  AO22AXL U3571 ( .A(n1016), .B(n3991), .C(n4011), .D(n3926), .Y(n1716) );
  AOI22XL U3572 ( .A(n3828), .B(A[141]), .C(n3801), .D(A[653]), .Y(n3926) );
  AO22AXL U3573 ( .A(n808), .B(n3992), .C(n4005), .D(n3927), .Y(n1756) );
  AOI22XL U3574 ( .A(n3710), .B(A[181]), .C(n3820), .D(A[693]), .Y(n3927) );
  AO22AXL U3575 ( .A(n1010), .B(n3673), .C(n4006), .D(n3928), .Y(n1717) );
  AOI22XL U3576 ( .A(n3710), .B(A[142]), .C(n4050), .D(A[654]), .Y(n3928) );
  AO22AXL U3577 ( .A(n802), .B(n3992), .C(n4011), .D(n3929), .Y(n1757) );
  AOI22XL U3578 ( .A(n4063), .B(A[182]), .C(n4045), .D(A[694]), .Y(n3929) );
  MUX2IXL U3579 ( .D0(n1479), .D1(n1480), .S(n3983), .Y(n1604) );
  MUX2IXL U3580 ( .D0(A[285]), .D1(A[797]), .S(n4025), .Y(n1480) );
  NOR21XL U3581 ( .B(n4030), .A(A[541]), .Y(n1479) );
  MUX2IXL U3582 ( .D0(n661), .D1(n662), .S(n3983), .Y(n1795) );
  MUX2IXL U3583 ( .D0(A[476]), .D1(A[988]), .S(n4025), .Y(n662) );
  MUX2IXL U3584 ( .D0(n1185), .D1(n1186), .S(n3978), .Y(n1676) );
  NOR21XL U3585 ( .B(n4035), .A(A[613]), .Y(n1185) );
  MUX2IXL U3586 ( .D0(n1217), .D1(n1218), .S(n3681), .Y(n1668) );
  NOR21XL U3587 ( .B(n3781), .A(A[605]), .Y(n1217) );
  MUX2IXL U3588 ( .D0(n1057), .D1(n1058), .S(n3977), .Y(n1708) );
  MUX2IXL U3589 ( .D0(n657), .D1(n658), .S(n3979), .Y(n1796) );
  MUX2IXL U3590 ( .D0(A[477]), .D1(A[989]), .S(n4025), .Y(n658) );
  NOR21XL U3591 ( .B(n4035), .A(A[533]), .Y(n1511) );
  MUX2IX1 U3592 ( .D0(A[277]), .D1(A[789]), .S(n4024), .Y(n1512) );
  MUX2IXL U3593 ( .D0(n1483), .D1(n1484), .S(n3982), .Y(n1603) );
  MUX2IXL U3594 ( .D0(A[284]), .D1(A[796]), .S(n4025), .Y(n1484) );
  NOR21XL U3595 ( .B(n3820), .A(A[540]), .Y(n1483) );
  MUX2IXL U3596 ( .D0(n1221), .D1(n1222), .S(n3681), .Y(n1667) );
  NOR21XL U3597 ( .B(n3781), .A(A[604]), .Y(n1221) );
  MUX2IXL U3598 ( .D0(n1053), .D1(n1054), .S(n3977), .Y(n1709) );
  MUX2IX1 U3599 ( .D0(A[276]), .D1(A[788]), .S(n4024), .Y(n1516) );
  NOR21XL U3600 ( .B(n3781), .A(A[532]), .Y(n1515) );
  MUX2IXL U3601 ( .D0(n1153), .D1(n1154), .S(n3975), .Y(n1684) );
  NOR21XL U3602 ( .B(n3821), .A(A[621]), .Y(n1153) );
  INVX1 U3603 ( .A(n1660), .Y(n318) );
  NOR21XL U3604 ( .B(n3802), .A(A[597]), .Y(n1247) );
  INVX1 U3605 ( .A(n1659), .Y(n317) );
  NOR21XL U3606 ( .B(n3802), .A(A[596]), .Y(n1250) );
  NOR21XL U3607 ( .B(n3781), .A(A[629]), .Y(n1121) );
  NOR21XL U3608 ( .B(n4030), .A(A[628]), .Y(n1125) );
  NOR21XL U3609 ( .B(n3793), .A(A[565]), .Y(n1351) );
  NOR21XL U3610 ( .B(n4028), .A(A[525]), .Y(n1543) );
  NOR21XL U3611 ( .B(n3788), .A(A[717]), .Y(n713) );
  NOR21XL U3612 ( .B(n4030), .A(A[660]), .Y(n981) );
  NOR21XL U3613 ( .B(n4049), .A(A[668]), .Y(n949) );
  NOR21XL U3614 ( .B(n3766), .A(A[716]), .Y(n717) );
  NOR21XL U3615 ( .B(n3805), .A(A[564]), .Y(n1355) );
  NOR21XL U3616 ( .B(n3802), .A(A[524]), .Y(n1547) );
  MUX2IXL U3617 ( .D0(A[125]), .D1(A[637]), .S(n4045), .Y(n1089) );
  MUX2IXL U3618 ( .D0(A[188]), .D1(A[700]), .S(n4023), .Y(n773) );
  MUX2IXL U3619 ( .D0(A[124]), .D1(A[636]), .S(n3802), .Y(n1093) );
  MUX2IXL U3620 ( .D0(A[317]), .D1(A[829]), .S(n3768), .Y(n1320) );
  MUX2IXL U3621 ( .D0(A[309]), .D1(A[821]), .S(n4023), .Y(n1352) );
  MUX2IXL U3622 ( .D0(A[269]), .D1(A[781]), .S(n4030), .Y(n1544) );
  MUX2IXL U3623 ( .D0(A[405]), .D1(A[917]), .S(n4022), .Y(n978) );
  MUX2IXL U3624 ( .D0(A[413]), .D1(A[925]), .S(n3768), .Y(n946) );
  MUX2IX1 U3625 ( .D0(A[485]), .D1(A[997]), .S(n4024), .Y(n626) );
  MUX2IXL U3626 ( .D0(A[493]), .D1(A[1005]), .S(n3821), .Y(n594) );
  MUX2IXL U3627 ( .D0(A[404]), .D1(A[916]), .S(n4022), .Y(n982) );
  MUX2IXL U3628 ( .D0(A[412]), .D1(A[924]), .S(n4022), .Y(n950) );
  MUX2IX1 U3629 ( .D0(A[484]), .D1(A[996]), .S(n4024), .Y(n630) );
  MUX2IXL U3630 ( .D0(A[316]), .D1(A[828]), .S(n3768), .Y(n1324) );
  MUX2IXL U3631 ( .D0(A[308]), .D1(A[820]), .S(n4075), .Y(n1356) );
  MUX2IXL U3632 ( .D0(A[268]), .D1(A[780]), .S(n3821), .Y(n1548) );
  MUX2IXL U3633 ( .D0(A[492]), .D1(A[1004]), .S(n3758), .Y(n598) );
  MUX2IXL U3634 ( .D0(n1189), .D1(n1190), .S(n3978), .Y(n1675) );
  NOR21XL U3635 ( .B(n4035), .A(A[612]), .Y(n1189) );
  MUX2IXL U3636 ( .D0(n6), .D1(n14), .S(n3973), .Y(B[5]) );
  MUX2IXL U3637 ( .D0(n38), .D1(n46), .S(n3971), .Y(n14) );
  MUX2IXL U3638 ( .D0(n22), .D1(n30), .S(SH[6]), .Y(n6) );
  NOR21XL U3639 ( .B(n4030), .A(A[588]), .Y(n1272) );
  NOR21XL U3640 ( .B(n4030), .A(A[589]), .Y(n1269) );
  AO22AXL U3641 ( .A(n1390), .B(n3993), .C(n4014), .D(n3930), .Y(n1620) );
  AOI22XL U3642 ( .A(n4069), .B(A[45]), .C(n3833), .D(A[557]), .Y(n3930) );
  MUX2IXL U3643 ( .D0(n7), .D1(n15), .S(n3973), .Y(B[6]) );
  MUX2IXL U3644 ( .D0(n39), .D1(n47), .S(n3971), .Y(n15) );
  MUX2XL U3645 ( .D0(n1181), .D1(n1182), .S(n3978), .Y(n3931) );
  MUX2IXL U3646 ( .D0(A[189]), .D1(A[701]), .S(n4023), .Y(n769) );
  NOR21XL U3647 ( .B(n3769), .A(A[837]), .Y(n1293) );
  NOR21XL U3648 ( .B(n3769), .A(A[836]), .Y(n1296) );
  AO22AXL U3649 ( .A(n1378), .B(n3993), .C(n4014), .D(n3932), .Y(n1622) );
  AOI22XL U3650 ( .A(n4069), .B(A[47]), .C(n3824), .D(A[559]), .Y(n3932) );
  AO22AXL U3651 ( .A(n1004), .B(n3991), .C(n4011), .D(n3933), .Y(n1718) );
  AOI22XL U3652 ( .A(n4061), .B(A[143]), .C(n4050), .D(A[655]), .Y(n3933) );
  AO22AXL U3653 ( .A(n796), .B(n3993), .C(n4012), .D(n3934), .Y(n1758) );
  AOI22XL U3654 ( .A(n3710), .B(A[183]), .C(n3766), .D(A[695]), .Y(n3934) );
  MUX2IXL U3655 ( .D0(n1347), .D1(n1348), .S(n3981), .Y(n1629) );
  MUX2IXL U3656 ( .D0(A[310]), .D1(A[822]), .S(n4023), .Y(n1348) );
  NOR21XL U3657 ( .B(n3793), .A(A[566]), .Y(n1347) );
  NOR21XL U3658 ( .B(n4035), .A(A[534]), .Y(n1507) );
  MUX2IX1 U3659 ( .D0(A[278]), .D1(A[790]), .S(n4024), .Y(n1508) );
  MUX2IXL U3660 ( .D0(n653), .D1(n654), .S(n3980), .Y(n1797) );
  MUX2IXL U3661 ( .D0(A[478]), .D1(A[990]), .S(n4025), .Y(n654) );
  MUX2IXL U3662 ( .D0(n1177), .D1(n1178), .S(n3978), .Y(n1678) );
  NOR21XL U3663 ( .B(n4028), .A(A[615]), .Y(n1177) );
  MUX2IXL U3664 ( .D0(n969), .D1(n970), .S(n4018), .Y(n1726) );
  NOR21XL U3665 ( .B(n4028), .A(A[663]), .Y(n969) );
  MUX2IXL U3666 ( .D0(A[407]), .D1(A[919]), .S(n4026), .Y(n970) );
  MUX2IXL U3667 ( .D0(n649), .D1(n650), .S(n3980), .Y(n1798) );
  MUX2IXL U3668 ( .D0(A[479]), .D1(A[991]), .S(n3818), .Y(n650) );
  MUX2IX1 U3669 ( .D0(A[279]), .D1(A[791]), .S(n4024), .Y(n1504) );
  NOR21XL U3670 ( .B(n3781), .A(A[535]), .Y(n1503) );
  MUX2IXL U3671 ( .D0(n1535), .D1(n1536), .S(n3985), .Y(n1590) );
  MUX2IXL U3672 ( .D0(A[271]), .D1(A[783]), .S(n3805), .Y(n1536) );
  NOR21XL U3673 ( .B(n3781), .A(A[527]), .Y(n1535) );
  MUX2IXL U3674 ( .D0(n1149), .D1(n3777), .S(n3975), .Y(n1685) );
  NOR21XL U3675 ( .B(n3768), .A(A[622]), .Y(n1149) );
  MUX2IXL U3676 ( .D0(n1145), .D1(n1146), .S(n3975), .Y(n1686) );
  NOR21XL U3677 ( .B(n3721), .A(A[623]), .Y(n1145) );
  NOR21XL U3678 ( .B(n3802), .A(A[598]), .Y(n1244) );
  NOR21XL U3679 ( .B(n3768), .A(A[599]), .Y(n1241) );
  NOR21XL U3680 ( .B(n3721), .A(A[838]), .Y(n1290) );
  NOR21XL U3681 ( .B(n3793), .A(A[839]), .Y(n1287) );
  NOR21XL U3682 ( .B(n3802), .A(A[575]), .Y(n1311) );
  NOR21XL U3683 ( .B(n3781), .A(A[543]), .Y(n1471) );
  NOR21XL U3684 ( .B(n4028), .A(A[661]), .Y(n977) );
  NOR21XL U3685 ( .B(n4075), .A(A[669]), .Y(n945) );
  NOR21XL U3686 ( .B(n4045), .A(A[606]), .Y(n1213) );
  NOR21XL U3687 ( .B(n4028), .A(A[662]), .Y(n973) );
  NOR21XL U3688 ( .B(n3721), .A(A[670]), .Y(n941) );
  NOR21XL U3689 ( .B(n3758), .A(A[718]), .Y(n709) );
  NOR21XL U3690 ( .B(n3793), .A(A[567]), .Y(n1343) );
  NOR21XL U3691 ( .B(n3769), .A(A[631]), .Y(n1113) );
  NOR21XL U3692 ( .B(n3758), .A(A[719]), .Y(n705) );
  MUX2IXL U3693 ( .D0(A[190]), .D1(A[702]), .S(n4049), .Y(n765) );
  MUX2IXL U3694 ( .D0(A[127]), .D1(A[639]), .S(n3758), .Y(n1081) );
  MUX2IXL U3695 ( .D0(A[191]), .D1(A[703]), .S(n4044), .Y(n761) );
  MUX2IXL U3696 ( .D0(A[406]), .D1(A[918]), .S(n4022), .Y(n974) );
  MUX2IXL U3697 ( .D0(A[414]), .D1(A[926]), .S(n3805), .Y(n942) );
  MUX2IX1 U3698 ( .D0(A[486]), .D1(A[998]), .S(n4024), .Y(n622) );
  MUX2IXL U3699 ( .D0(A[494]), .D1(A[1006]), .S(n3769), .Y(n590) );
  MUX2IXL U3700 ( .D0(A[319]), .D1(A[831]), .S(n3805), .Y(n1312) );
  MUX2IXL U3701 ( .D0(A[311]), .D1(A[823]), .S(n4023), .Y(n1344) );
  MUX2IXL U3702 ( .D0(A[287]), .D1(A[799]), .S(n4025), .Y(n1472) );
  MUX2IXL U3703 ( .D0(A[415]), .D1(A[927]), .S(n3805), .Y(n938) );
  MUX2IX1 U3704 ( .D0(A[487]), .D1(A[999]), .S(n4024), .Y(n618) );
  MUX2IXL U3705 ( .D0(A[495]), .D1(A[1007]), .S(n3818), .Y(n586) );
  MUX2IXL U3706 ( .D0(n8), .D1(n16), .S(n3973), .Y(B[7]) );
  MUX2IXL U3707 ( .D0(n40), .D1(n48), .S(n3971), .Y(n16) );
  MUX2IXL U3708 ( .D0(n24), .D1(n32), .S(n3971), .Y(n8) );
  AO22AXL U3709 ( .A(n1426), .B(n3994), .C(n4008), .D(n3935), .Y(n1614) );
  AOI22XL U3710 ( .A(n4070), .B(A[39]), .C(n4047), .D(A[551]), .Y(n3935) );
  NOR21XL U3711 ( .B(n4045), .A(A[526]), .Y(n1539) );
  MUX2IXL U3712 ( .D0(A[270]), .D1(A[782]), .S(n3758), .Y(n1540) );
  MUX2IXL U3713 ( .D0(A[318]), .D1(A[830]), .S(n3805), .Y(n1316) );
  NOR21XL U3714 ( .B(n3802), .A(A[574]), .Y(n1315) );
  MUX2IXL U3715 ( .D0(A[286]), .D1(A[798]), .S(n4025), .Y(n1476) );
  NOR21XL U3716 ( .B(n3768), .A(A[542]), .Y(n1475) );
  NOR21XL U3717 ( .B(n3793), .A(A[630]), .Y(n1117) );
  MUX2IXL U3718 ( .D0(A[126]), .D1(A[638]), .S(n4025), .Y(n1085) );
  MUX2XL U3719 ( .D0(n1209), .D1(n1210), .S(n3680), .Y(n3936) );
  NOR21XL U3720 ( .B(n3721), .A(A[671]), .Y(n937) );
  NOR21XL U3721 ( .B(n3793), .A(A[568]), .Y(n1339) );
  NOR21XL U3722 ( .B(n3793), .A(A[573]), .Y(n1319) );
  NOR21XL U3723 ( .B(n3793), .A(A[572]), .Y(n1323) );
  MUX2IXL U3724 ( .D0(A[491]), .D1(A[1003]), .S(n3758), .Y(n602) );
  MUX2IXL U3725 ( .D0(A[488]), .D1(A[1000]), .S(n3741), .Y(n614) );
endmodule


module regbank_a0_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module regbank_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regbank_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regbank_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_50 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10838;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_50 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10838), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10838), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10838), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10838), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10838), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10838), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10838), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10838), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10838), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_51 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10856;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_51 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10856), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10856), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10856), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10856), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10856), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10856), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10856), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10856), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10856), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_52 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10874;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_52 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10874), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10874), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10874), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10874), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10874), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10874), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10874), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10874), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10874), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_53 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10892;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_53 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10892), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10892), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10892), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10892), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10892), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10892), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10892), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10892), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10892), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_54 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10910;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_54 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10910), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10910), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10910), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10910), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10910), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10910), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10910), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10910), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10910), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_0000001f ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10928;

  SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10928), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10928), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10928), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10928), .XR(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10928), .XS(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10928), .XS(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10928), .XS(arstz), .Q(rdat[2]) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10928), .XS(arstz), .Q(rdat[1]) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10928), .XS(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000004 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10946;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10946), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net10946), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10946), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10946), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10946), .XR(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10946), .XS(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10946), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10946), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10946), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_4_00000004 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10964;

  SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10964), .TE(test_se) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10964), .XR(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10964), .XS(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10964), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10964), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH7_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net10982;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10982), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net10982), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net10982), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net10982), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net10982), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net10982), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net10982), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net10982), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_55 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11000;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_55 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11000), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11000), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11000), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11000), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11000), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11000), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11000), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11000), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11000), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_55 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_2 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_2 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[7]), .Y(n3) );
  INVX1 U4 ( .A(set2[0]), .Y(n1) );
  INVX1 U5 ( .A(set2[1]), .Y(n14) );
  INVX1 U6 ( .A(set2[3]), .Y(n15) );
  INVX1 U7 ( .A(set2[4]), .Y(n2) );
  INVX1 U8 ( .A(set2[5]), .Y(n12) );
  INVX1 U9 ( .A(set2[2]), .Y(n13) );
  NAND3X1 U10 ( .A(n16), .B(n3), .C(n12), .Y(n21) );
  NAND4X1 U11 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U12 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U13 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U14 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U15 ( .C(n13), .D(n11), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U16 ( .A(rdat[2]), .Y(n11) );
  AOI211X1 U17 ( .C(n1), .D(n10), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U18 ( .A(rdat[0]), .Y(n10) );
  AOI211X1 U19 ( .C(n14), .D(n9), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U20 ( .A(rdat[1]), .Y(n9) );
  AOI211X1 U21 ( .C(n12), .D(n8), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U22 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U23 ( .C(n2), .D(n7), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U24 ( .A(rdat[4]), .Y(n7) );
  AOI211X1 U25 ( .C(n15), .D(n6), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U26 ( .A(rdat[3]), .Y(n6) );
  AOI211X1 U27 ( .C(n16), .D(n5), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U28 ( .A(rdat[6]), .Y(n5) );
  AOI211X1 U29 ( .C(n3), .D(n4), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U30 ( .A(rdat[7]), .Y(n4) );
  NOR2X1 U31 ( .A(rdat[5]), .B(n12), .Y(irq[5]) );
  NOR2X1 U32 ( .A(rdat[4]), .B(n2), .Y(irq[4]) );
  NOR2X1 U33 ( .A(rdat[3]), .B(n15), .Y(irq[3]) );
  NOR2X1 U34 ( .A(rdat[2]), .B(n13), .Y(irq[2]) );
  NOR2X1 U35 ( .A(rdat[0]), .B(n1), .Y(irq[0]) );
  NOR2X1 U36 ( .A(rdat[7]), .B(n3), .Y(irq[7]) );
  NOR2X1 U37 ( .A(rdat[1]), .B(n14), .Y(irq[1]) );
  NOR2X1 U38 ( .A(rdat[6]), .B(n16), .Y(irq[6]) );
  INVX1 U39 ( .A(set2[6]), .Y(n16) );
endmodule


module glreg_WIDTH8_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11018;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11018), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11018), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11018), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11018), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11018), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11018), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11018), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11018), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11018), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_9 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n10, n2, n1;

  SDFFRQX1 db_cnt_reg_1_ ( .D(n9), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n8), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n10), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n10) );
  NOR3XL U7 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n8) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n2), .Y(n9) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_10 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n10, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n9), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n8), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n10), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n10) );
  NOR3XL U7 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n8) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n2), .Y(n9) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_11 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n10, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n9), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n8), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n10), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n1) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n10) );
  NOR3XL U7 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n8) );
  NOR3XL U8 ( .A(n1), .B(test_so), .C(n2), .Y(n9) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_12 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n9, n10, n11, n1, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n10), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n9), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n11), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n3) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n11) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n3), .Y(o_chg) );
  NOR3XL U6 ( .A(n3), .B(test_so), .C(db_cnt_0_), .Y(n9) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n3), .Y(n10) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_13 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n9, n10, n11, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n10), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n9), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n11), .SIN(d_org_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n11) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n9) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n10) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_14 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n4, n5, n6, n2, n1;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n5), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n6), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n4), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(o_dbc), .B(d_org_0_), .Y(n2) );
  AO22AXL U4 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n4) );
  NOR32XL U5 ( .B(test_so), .C(n1), .A(n2), .Y(o_chg) );
  NOR3XL U6 ( .A(n2), .B(test_so), .C(db_cnt_0_), .Y(n6) );
  NOR3XL U7 ( .A(n1), .B(test_so), .C(n2), .Y(n5) );
  INVX1 U8 ( .A(db_cnt_0_), .Y(n1) );
endmodule


module dbnc_WIDTH2_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n1, n2, n3, n6, n7;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n6), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n2), .B(n7), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n2) );
  INVX1 U6 ( .A(test_so), .Y(n1) );
  AO22AXL U7 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR2X1 U8 ( .A(n7), .B(db_cnt_0_), .Y(n6) );
  OAI32X1 U9 ( .A(n2), .B(test_so), .C(n7), .D(n1), .E(n3), .Y(n8) );
  INVX1 U10 ( .A(n6), .Y(n3) );
endmodule


module dbnc_WIDTH2_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n1, n2, n3, n6, n7;

  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n6), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n2), .B(n7), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n2) );
  INVX1 U6 ( .A(test_so), .Y(n1) );
  AO22AXL U7 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR2X1 U8 ( .A(n7), .B(db_cnt_0_), .Y(n6) );
  OAI32X1 U9 ( .A(n2), .B(test_so), .C(n7), .D(n1), .E(n3), .Y(n8) );
  INVX1 U10 ( .A(n6), .Y(n3) );
endmodule


module dbnc_WIDTH2_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n1, n2, n3, n6, n7;

  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n6), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n2), .B(n7), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n7) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n2) );
  AO22AXL U6 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  INVX1 U7 ( .A(test_so), .Y(n1) );
  NOR2X1 U8 ( .A(n7), .B(db_cnt_0_), .Y(n6) );
  OAI32X1 U9 ( .A(n2), .B(test_so), .C(n7), .D(n1), .E(n3), .Y(n8) );
  INVX1 U10 ( .A(n6), .Y(n3) );
endmodule


module dbnc_WIDTH2_3 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n8, n9, n4, n5, n1, n2, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n8), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n5), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n9), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n2), .B(n4), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n2) );
  INVX1 U6 ( .A(test_so), .Y(n1) );
  AO22AXL U7 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n9) );
  NOR2X1 U8 ( .A(n4), .B(db_cnt_0_), .Y(n5) );
  OAI32X1 U9 ( .A(n2), .B(test_so), .C(n4), .D(n1), .E(n3), .Y(n8) );
  INVX1 U10 ( .A(n5), .Y(n3) );
endmodule


module dbnc_WIDTH2_4 ( o_dbc, o_chg, i_org, clk, rstz, test_si, test_so, 
        test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_0_, n5, n6, n4, n7, n1, n2, n3;

  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(n6), .SIN(db_cnt_0_), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(n7), .SIN(o_dbc), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n5), .SIN(d_org_0_), .SMC(test_se), .C(clk), .XR(
        rstz), .Q(o_dbc) );
  NOR3XL U3 ( .A(n2), .B(n4), .C(n1), .Y(o_chg) );
  XNOR2XL U4 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  INVX1 U5 ( .A(db_cnt_0_), .Y(n2) );
  INVX1 U6 ( .A(test_so), .Y(n1) );
  AO22AXL U7 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n5) );
  NOR2X1 U8 ( .A(n4), .B(db_cnt_0_), .Y(n7) );
  OAI32X1 U9 ( .A(n2), .B(test_so), .C(n4), .D(n1), .E(n3), .Y(n6) );
  INVX1 U10 ( .A(n7), .Y(n3) );
endmodule


module dbnc_WIDTH5_TIMEOUT30 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_3_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N8, N9, N10,
         N17, N18, N19, N20, N21, N22, net11036, n6, n3, n4, n5, n7, n8, n9,
         n1, n2;
  wire   [4:2] add_165_carry;

  HAD1X1 add_165_U1_1_1 ( .A(db_cnt_1_), .B(db_cnt_0_), .CO(add_165_carry[2]), 
        .SO(N8) );
  HAD1X1 add_165_U1_1_2 ( .A(db_cnt_2_), .B(add_165_carry[2]), .CO(
        add_165_carry[3]), .SO(N9) );
  HAD1X1 add_165_U1_1_3 ( .A(db_cnt_3_), .B(add_165_carry[3]), .CO(
        add_165_carry[4]), .SO(N10) );
  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH5_TIMEOUT30 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N17), .ENCLK(net11036), .TE(test_se) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 db_cnt_reg_4_ ( .D(N22), .SIN(db_cnt_3_), .SMC(test_se), .C(
        net11036), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N21), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11036), .XR(rstz), .Q(db_cnt_3_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N20), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11036), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N19), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11036), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N18), .SIN(o_dbc), .SMC(test_se), .C(net11036), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n6), .SIN(d_org_0_), .SMC(test_se), .C(net11036), 
        .XR(rstz), .Q(o_dbc) );
  NOR21XL U3 ( .B(N9), .A(n1), .Y(N20) );
  NOR21XL U4 ( .B(N10), .A(n1), .Y(N21) );
  NOR21XL U5 ( .B(N8), .A(n1), .Y(N19) );
  NOR43XL U6 ( .B(db_cnt_1_), .C(n3), .D(n2), .A(n4), .Y(o_chg) );
  AND3X1 U7 ( .A(test_so), .B(db_cnt_2_), .C(db_cnt_3_), .Y(n3) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n4) );
  INVX1 U9 ( .A(db_cnt_0_), .Y(n2) );
  NOR2X1 U10 ( .A(n5), .B(n1), .Y(N22) );
  XNOR2XL U11 ( .A(test_so), .B(add_165_carry[4]), .Y(n5) );
  AO22AXL U12 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n6) );
  INVX1 U13 ( .A(n7), .Y(n1) );
  AOI31X1 U14 ( .A(n8), .B(db_cnt_3_), .C(test_so), .D(n4), .Y(n7) );
  NOR32XL U15 ( .B(db_cnt_1_), .C(db_cnt_2_), .A(db_cnt_0_), .Y(n8) );
  NOR2X1 U16 ( .A(db_cnt_0_), .B(n1), .Y(N18) );
  NAND41X1 U17 ( .D(db_cnt_1_), .A(n2), .B(n4), .C(n9), .Y(N17) );
  NOR3XL U18 ( .A(db_cnt_2_), .B(test_so), .C(db_cnt_3_), .Y(n9) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH5_TIMEOUT30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_0 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N18, N19,
         net11054, n13, n9, n10, n11, n12, n14, n15, n1, n2, n3, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11054), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11054), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11054), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N18), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11054), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11054), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11054), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n12), .Y(n2) );
  OAI31XL U4 ( .A(n1), .B(n5), .C(n6), .D(n4), .Y(n11) );
  INVX1 U5 ( .A(n14), .Y(n4) );
  NOR2X1 U6 ( .A(n3), .B(n5), .Y(n12) );
  OAI32X1 U7 ( .A(n2), .B(n6), .C(n11), .D(n11), .E(n1), .Y(N19) );
  AOI211X1 U8 ( .C(n3), .D(n5), .A(n11), .B(n12), .Y(N17) );
  INVX1 U9 ( .A(n9), .Y(o_chg) );
  XNOR2XL U10 ( .A(o_dbc), .B(d_org_0_), .Y(n14) );
  NAND4X1 U11 ( .A(n4), .B(n3), .C(db_cnt_1_), .D(n10), .Y(n9) );
  NOR2X1 U12 ( .A(n6), .B(n1), .Y(n10) );
  AO22AXL U13 ( .A(n9), .B(o_dbc), .C(d_org_0_), .D(n9), .Y(n13) );
  OAI33XL U14 ( .A(n11), .B(n12), .C(n6), .D(n2), .E(db_cnt_2_), .F(n11), .Y(
        N18) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  INVX1 U16 ( .A(db_cnt_1_), .Y(n5) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n6) );
  INVX1 U18 ( .A(test_so), .Y(n1) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n11), .Y(N16) );
  NAND3X1 U20 ( .A(n14), .B(n3), .C(n15), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n15) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_1 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N18, N19,
         net11072, n13, n9, n10, n11, n12, n14, n15, n1, n2, n3, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11072), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11072), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11072), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N18), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11072), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11072), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11072), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n12), .Y(n2) );
  OAI31XL U4 ( .A(n1), .B(n5), .C(n6), .D(n4), .Y(n11) );
  INVX1 U5 ( .A(n14), .Y(n4) );
  NOR2X1 U6 ( .A(n3), .B(n5), .Y(n12) );
  OAI32X1 U7 ( .A(n2), .B(n6), .C(n11), .D(n11), .E(n1), .Y(N19) );
  AOI211X1 U8 ( .C(n3), .D(n5), .A(n11), .B(n12), .Y(N17) );
  INVX1 U9 ( .A(n9), .Y(o_chg) );
  XNOR2XL U10 ( .A(o_dbc), .B(d_org_0_), .Y(n14) );
  NAND4X1 U11 ( .A(n4), .B(n3), .C(db_cnt_1_), .D(n10), .Y(n9) );
  NOR2X1 U12 ( .A(n6), .B(n1), .Y(n10) );
  AO22AXL U13 ( .A(n9), .B(o_dbc), .C(d_org_0_), .D(n9), .Y(n13) );
  OAI33XL U14 ( .A(n11), .B(n12), .C(n6), .D(n2), .E(db_cnt_2_), .F(n11), .Y(
        N18) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  INVX1 U16 ( .A(db_cnt_1_), .Y(n5) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n6) );
  INVX1 U18 ( .A(test_so), .Y(n1) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n11), .Y(N16) );
  NAND3X1 U20 ( .A(n14), .B(n3), .C(n15), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n15) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_2 ( o_dbc, o_chg, i_org, clk, rstz, test_si, 
        test_so, test_se );
  input i_org, clk, rstz, test_si, test_se;
  output o_dbc, o_chg, test_so;
  wire   d_org_0_, db_cnt_2_, db_cnt_1_, db_cnt_0_, N15, N16, N17, N18, N19,
         net11090, n13, n9, n10, n11, n12, n14, n15, n1, n2, n3, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11090), .TE(test_se) );
  SDFFRQX1 db_cnt_reg_3_ ( .D(N19), .SIN(db_cnt_2_), .SMC(test_se), .C(
        net11090), .XR(rstz), .Q(test_so) );
  SDFFRQX1 db_cnt_reg_0_ ( .D(N16), .SIN(o_dbc), .SMC(test_se), .C(net11090), 
        .XR(rstz), .Q(db_cnt_0_) );
  SDFFRQX1 db_cnt_reg_2_ ( .D(N18), .SIN(db_cnt_1_), .SMC(test_se), .C(
        net11090), .XR(rstz), .Q(db_cnt_2_) );
  SDFFRQX1 db_cnt_reg_1_ ( .D(N17), .SIN(db_cnt_0_), .SMC(test_se), .C(
        net11090), .XR(rstz), .Q(db_cnt_1_) );
  SDFFRQX1 d_org_reg_0_ ( .D(i_org), .SIN(test_si), .SMC(test_se), .C(clk), 
        .XR(rstz), .Q(d_org_0_) );
  SDFFRQX1 d_org_reg_1_ ( .D(n13), .SIN(d_org_0_), .SMC(test_se), .C(net11090), 
        .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n12), .Y(n2) );
  OAI31XL U4 ( .A(n1), .B(n5), .C(n6), .D(n4), .Y(n11) );
  INVX1 U5 ( .A(n14), .Y(n4) );
  NOR2X1 U6 ( .A(n3), .B(n5), .Y(n12) );
  OAI32X1 U7 ( .A(n2), .B(n6), .C(n11), .D(n11), .E(n1), .Y(N19) );
  AOI211X1 U8 ( .C(n3), .D(n5), .A(n11), .B(n12), .Y(N17) );
  INVX1 U9 ( .A(n9), .Y(o_chg) );
  XNOR2XL U10 ( .A(o_dbc), .B(d_org_0_), .Y(n14) );
  NAND4X1 U11 ( .A(n4), .B(n3), .C(db_cnt_1_), .D(n10), .Y(n9) );
  NOR2X1 U12 ( .A(n6), .B(n1), .Y(n10) );
  AO22AXL U13 ( .A(n9), .B(o_dbc), .C(d_org_0_), .D(n9), .Y(n13) );
  OAI33XL U14 ( .A(n11), .B(n12), .C(n6), .D(n2), .E(db_cnt_2_), .F(n11), .Y(
        N18) );
  INVX1 U15 ( .A(db_cnt_0_), .Y(n3) );
  INVX1 U16 ( .A(db_cnt_1_), .Y(n5) );
  INVX1 U17 ( .A(db_cnt_2_), .Y(n6) );
  INVX1 U18 ( .A(test_so), .Y(n1) );
  NOR2X1 U19 ( .A(db_cnt_0_), .B(n11), .Y(N16) );
  NAND3X1 U20 ( .A(n14), .B(n3), .C(n15), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt_1_), .B(test_so), .C(db_cnt_2_), .Y(n15) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000028 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11108;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11108), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11108), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11108), .XR(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11108), .XS(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11108), .XR(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11108), .XS(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11108), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11108), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11108), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_56 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11126;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_56 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11126), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11126), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11126), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11126), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11126), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11126), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11126), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11126), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11126), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_56 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_57 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11144;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_57 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11144), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11144), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11144), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11144), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11144), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11144), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11144), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11144), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11144), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_57 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_58 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11162;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_58 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11162), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11162), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11162), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11162), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11162), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11162), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11162), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11162), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11162), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_58 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_59 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11180;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_59 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11180), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11180), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11180), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11180), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11180), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11180), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11180), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11180), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11180), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_59 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_60 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11198;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_60 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11198), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11198), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11198), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11198), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11198), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11198), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11198), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11198), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11198), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_60 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_61 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11216;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_61 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11216), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11216), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11216), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11216), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11216), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11216), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11216), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11216), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11216), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_61 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_62 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11234;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_62 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11234), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11234), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11234), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11234), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11234), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11234), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11234), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11234), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11234), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_62 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_63 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11252;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_63 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11252), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11252), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11252), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11252), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11252), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11252), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11252), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11252), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11252), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_63 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11270;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11270), .TE(test_se) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11270), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11270), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11270), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11270), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_64 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11288;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_64 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11288), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11288), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11288), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11288), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11288), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11288), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11288), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11288), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11288), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_64 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_3 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_3 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[0]), .Y(n14) );
  INVX1 U4 ( .A(set2[1]), .Y(n16) );
  INVX1 U5 ( .A(set2[2]), .Y(n15) );
  INVX1 U6 ( .A(set2[3]), .Y(n13) );
  INVX1 U7 ( .A(set2[4]), .Y(n12) );
  NAND3X1 U8 ( .A(n9), .B(n10), .C(n11), .Y(n21) );
  AOI211X1 U9 ( .C(n14), .D(n8), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U10 ( .A(rdat[0]), .Y(n8) );
  AOI211X1 U11 ( .C(n16), .D(n7), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U12 ( .A(rdat[1]), .Y(n7) );
  AOI211X1 U13 ( .C(n15), .D(n6), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U14 ( .A(rdat[2]), .Y(n6) );
  AOI211X1 U15 ( .C(n13), .D(n5), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U16 ( .A(rdat[3]), .Y(n5) );
  AOI211X1 U17 ( .C(n12), .D(n4), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U18 ( .A(rdat[4]), .Y(n4) );
  AOI211X1 U19 ( .C(n11), .D(n3), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U20 ( .A(rdat[5]), .Y(n3) );
  AOI211X1 U21 ( .C(n9), .D(n2), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U22 ( .A(rdat[6]), .Y(n2) );
  AOI211X1 U23 ( .C(n10), .D(n1), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U24 ( .A(rdat[7]), .Y(n1) );
  NAND4X1 U25 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U26 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U27 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U28 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  INVX1 U29 ( .A(set2[5]), .Y(n11) );
  NOR2X1 U30 ( .A(rdat[0]), .B(n14), .Y(irq[0]) );
  NOR2X1 U31 ( .A(rdat[1]), .B(n16), .Y(irq[1]) );
  NOR2X1 U32 ( .A(rdat[2]), .B(n15), .Y(irq[2]) );
  NOR2X1 U33 ( .A(rdat[3]), .B(n13), .Y(irq[3]) );
  INVX1 U34 ( .A(set2[6]), .Y(n9) );
  INVX1 U35 ( .A(set2[7]), .Y(n10) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n12), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n9), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[5]), .B(n11), .Y(irq[5]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n10), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11306;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11306), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11306), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11306), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11306), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11306), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11306), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11306), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11306), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11306), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_65 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11324;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_65 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11324), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11324), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11324), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11324), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11324), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11324), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11324), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11324), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11324), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_65 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_66 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11342;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_66 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11342), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11342), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11342), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11342), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11342), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11342), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11342), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11342), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11342), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_66 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000032 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11360;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11360), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11360), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11360), .XR(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11360), .XS(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11360), .XR(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11360), .XS(arstz), .Q(rdat[4]) );
  SDFFSQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11360), .XS(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11360), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11360), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000098 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11378;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11378), .TE(test_se) );
  SDFFSQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11378), .XS(arstz), .Q(rdat[7]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11378), .XS(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11378), .XR(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11378), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11378), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11378), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11378), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11378), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_000000f0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11396;

  SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11396), .TE(test_se) );
  SDFFSQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11396), .XS(arstz), .Q(rdat[7]) );
  SDFFSQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11396), .XS(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11396), .XS(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11396), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11396), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11396), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11396), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11396), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH1_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH1_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH2_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2, n3, n1;

  SDFFRQX1 mem_reg_1_ ( .D(n3), .SIN(rdat[0]), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XR(
        arstz), .Q(rdat[0]) );
  INVX1 U2 ( .A(we), .Y(n1) );
  AO22XL U3 ( .A(wdat[0]), .B(we), .C(rdat[0]), .D(n1), .Y(n2) );
  AO22XL U4 ( .A(we), .B(wdat[1]), .C(rdat[1]), .D(n1), .Y(n3) );
endmodule


module glreg_WIDTH3 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [2:0] wdat;
  output [2:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11414;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11414), .TE(test_se) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11414), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11414), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11414), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000011 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11432;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11432), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11432), .XR(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11432), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11432), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11432), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11432), .XR(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11432), .XS(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11432), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11432), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000001 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11450;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11450), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11450), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11450), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11450), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11450), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11450), .XR(arstz), .Q(rdat[3]) );
  SDFFSQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11450), .XS(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11450), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11450), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_67 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11468;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_67 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11468), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11468), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11468), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11468), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11468), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11468), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11468), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11468), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11468), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_67 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_4 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_4 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[4]), .Y(n13) );
  INVX1 U4 ( .A(set2[7]), .Y(n12) );
  NAND3X1 U5 ( .A(n11), .B(n12), .C(n10), .Y(n21) );
  INVX1 U6 ( .A(set2[3]), .Y(n14) );
  INVX1 U7 ( .A(set2[0]), .Y(n9) );
  INVX1 U8 ( .A(set2[1]), .Y(n16) );
  INVX1 U9 ( .A(set2[5]), .Y(n10) );
  INVX1 U10 ( .A(set2[6]), .Y(n11) );
  INVX1 U11 ( .A(set2[2]), .Y(n15) );
  NAND4X1 U12 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U13 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U14 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U15 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U16 ( .C(n10), .D(n1), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U17 ( .A(rdat[5]), .Y(n1) );
  AOI211X1 U18 ( .C(n9), .D(n8), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U19 ( .A(rdat[0]), .Y(n8) );
  AOI211X1 U20 ( .C(n15), .D(n7), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U21 ( .A(rdat[2]), .Y(n7) );
  AOI211X1 U22 ( .C(n16), .D(n6), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U23 ( .A(rdat[1]), .Y(n6) );
  AOI211X1 U24 ( .C(n12), .D(n5), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U25 ( .A(rdat[7]), .Y(n5) );
  AOI211X1 U26 ( .C(n13), .D(n4), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U27 ( .A(rdat[4]), .Y(n4) );
  AOI211X1 U28 ( .C(n11), .D(n3), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U29 ( .A(rdat[6]), .Y(n3) );
  AOI211X1 U30 ( .C(n14), .D(n2), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U31 ( .A(rdat[3]), .Y(n2) );
  NOR2X1 U32 ( .A(rdat[7]), .B(n12), .Y(irq[7]) );
  NOR2X1 U33 ( .A(rdat[6]), .B(n11), .Y(irq[6]) );
  NOR2X1 U34 ( .A(rdat[3]), .B(n14), .Y(irq[3]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n15), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n9), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[4]), .B(n13), .Y(irq[4]) );
  NOR2X1 U38 ( .A(rdat[1]), .B(n16), .Y(irq[1]) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n10), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_4 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11486;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11486), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11486), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11486), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11486), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11486), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11486), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11486), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11486), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11486), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_68 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11504;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_68 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11504), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11504), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11504), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11504), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11504), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11504), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11504), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11504), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11504), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_68 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_7_70 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11522;

  SNPS_CLOCK_GATE_HIGH_glreg_7_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11522), .TE(test_se) );
  SDFFSQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11522), .XS(arstz), .Q(rdat[6]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11522), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11522), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11522), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11522), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11522), .XR(arstz), .Q(rdat[2]) );
  SDFFSQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11522), .XS(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_7_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_1_1_0 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n2;

  SDFFSQX1 mem_reg_0_ ( .D(n2), .SIN(test_si), .SMC(test_se), .C(clk), .XS(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_1_1_1 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   n1;

  SDFFSQX1 mem_reg_0_ ( .D(n1), .SIN(test_si), .SMC(test_se), .C(clk), .XS(
        arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n1) );
endmodule


module glreg_6_00000018 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11540;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11540), .TE(test_se) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11540), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11540), .XR(arstz), .Q(rdat[5]) );
  SDFFSQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11540), .XS(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11540), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11540), .XR(arstz), .Q(rdat[1]) );
  SDFFSQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11540), .XS(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_69 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11558;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_69 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11558), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11558), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11558), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11558), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11558), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11558), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11558), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11558), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11558), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_69 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_70 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11576;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11576), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11576), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11576), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11576), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11576), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11576), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11576), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11576), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11576), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_71 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11594;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_71 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11594), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11594), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11594), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11594), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11594), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11594), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11594), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11594), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11594), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_71 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_72 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11612;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_72 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11612), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11612), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11612), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11612), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11612), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11612), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11612), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11612), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11612), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_72 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_73 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11630;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_73 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11630), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11630), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11630), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11630), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11630), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11630), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11630), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11630), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11630), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_73 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_2 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11648;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11648), .TE(test_se) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11648), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11648), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11648), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11648), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11648), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_74 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11666;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_74 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11666), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11666), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11666), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11666), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11666), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11666), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11666), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11666), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11666), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_74 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_75 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11684;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_75 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11684), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11684), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11684), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11684), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11684), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11684), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11684), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11684), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11684), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_75 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_76 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11702;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_76 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11702), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11702), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11702), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11702), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11702), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11702), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11702), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11702), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11702), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_76 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_77 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11720;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_77 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11720), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11720), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11720), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11720), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11720), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11720), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11720), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11720), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11720), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_77 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_5 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_5 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[4]), .Y(n2) );
  NOR3XL U3 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NAND3X1 U4 ( .A(n14), .B(n1), .C(n3), .Y(n21) );
  INVX1 U5 ( .A(set2[3]), .Y(n4) );
  INVX1 U6 ( .A(set2[2]), .Y(n5) );
  INVX1 U7 ( .A(set2[5]), .Y(n3) );
  NAND4X1 U8 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U9 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U10 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  NOR4XL U11 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  INVX1 U12 ( .A(set2[1]), .Y(n16) );
  INVX1 U13 ( .A(set2[6]), .Y(n14) );
  INVX1 U14 ( .A(set2[0]), .Y(n15) );
  INVX1 U15 ( .A(set2[7]), .Y(n1) );
  NOR2X1 U16 ( .A(rdat[4]), .B(n2), .Y(irq[4]) );
  NOR2X1 U17 ( .A(rdat[5]), .B(n3), .Y(irq[5]) );
  AOI211X1 U18 ( .C(n2), .D(n9), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U19 ( .A(rdat[4]), .Y(n9) );
  AOI211X1 U20 ( .C(n3), .D(n8), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U21 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U22 ( .C(n15), .D(n13), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U23 ( .A(rdat[0]), .Y(n13) );
  AOI211X1 U24 ( .C(n16), .D(n12), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U25 ( .A(rdat[1]), .Y(n12) );
  AOI211X1 U26 ( .C(n5), .D(n11), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U27 ( .A(rdat[2]), .Y(n11) );
  AOI211X1 U28 ( .C(n4), .D(n10), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U29 ( .A(rdat[3]), .Y(n10) );
  AOI211X1 U30 ( .C(n1), .D(n7), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U31 ( .A(rdat[7]), .Y(n7) );
  AOI211X1 U32 ( .C(n14), .D(n6), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U33 ( .A(rdat[6]), .Y(n6) );
  NOR2X1 U34 ( .A(rdat[2]), .B(n5), .Y(irq[2]) );
  NOR2X1 U35 ( .A(rdat[3]), .B(n4), .Y(irq[3]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n15), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n14), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[1]), .B(n16), .Y(irq[1]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n1), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_5 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11738;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11738), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11738), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11738), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11738), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11738), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11738), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11738), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11738), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11738), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_6 ( clk, arstz, rst0, set2, clr1, rdat, irq, test_si, test_se
 );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0, test_si, test_se;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_6 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat), .test_si(test_si), .test_se(test_se) );
  INVX1 U2 ( .A(set2[7]), .Y(n2) );
  INVX1 U3 ( .A(set2[3]), .Y(n4) );
  NAND4X1 U4 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U5 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U6 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  NOR3XL U7 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  INVX1 U8 ( .A(set2[1]), .Y(n1) );
  INVX1 U9 ( .A(set2[2]), .Y(n3) );
  INVX1 U10 ( .A(set2[4]), .Y(n6) );
  NOR4XL U11 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NAND3X1 U12 ( .A(n5), .B(n2), .C(n15), .Y(n21) );
  INVX1 U13 ( .A(set2[6]), .Y(n5) );
  INVX1 U14 ( .A(set2[0]), .Y(n16) );
  NOR2X1 U15 ( .A(rdat[0]), .B(n16), .Y(irq[0]) );
  NOR2X1 U16 ( .A(rdat[1]), .B(n1), .Y(irq[1]) );
  NOR2X1 U17 ( .A(rdat[6]), .B(n5), .Y(irq[6]) );
  NOR2X1 U18 ( .A(rdat[7]), .B(n2), .Y(irq[7]) );
  AOI211X1 U19 ( .C(n16), .D(n14), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U20 ( .A(rdat[0]), .Y(n14) );
  AOI211X1 U21 ( .C(n1), .D(n13), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U22 ( .A(rdat[1]), .Y(n13) );
  AOI211X1 U23 ( .C(n3), .D(n12), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U24 ( .A(rdat[2]), .Y(n12) );
  AOI211X1 U25 ( .C(n4), .D(n11), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U26 ( .A(rdat[3]), .Y(n11) );
  AOI211X1 U27 ( .C(n6), .D(n10), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U28 ( .A(rdat[4]), .Y(n10) );
  AOI211X1 U29 ( .C(n15), .D(n9), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U30 ( .A(rdat[5]), .Y(n9) );
  AOI211X1 U31 ( .C(n5), .D(n8), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U32 ( .A(rdat[6]), .Y(n8) );
  AOI211X1 U33 ( .C(n2), .D(n7), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U34 ( .A(rdat[7]), .Y(n7) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n3), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n6), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[3]), .B(n4), .Y(irq[3]) );
  INVX1 U38 ( .A(set2[5]), .Y(n15) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n15), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_6 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11756;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11756), .TE(test_se) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11756), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11756), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11756), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11756), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11756), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11756), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11756), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11756), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_78 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11774;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_78 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11774), .TE(test_se) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11774), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11774), .XR(arstz), .Q(rdat[7]) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11774), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11774), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11774), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11774), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11774), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11774), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_78 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_79 ( clk, arstz, we, wdat, rdat, test_si, test_se );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we, test_si, test_se;
  wire   net11792;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_79 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11792), .TE(test_se) );
  SDFFRQX1 mem_reg_5_ ( .D(wdat[5]), .SIN(rdat[4]), .SMC(test_se), .C(net11792), .XR(arstz), .Q(rdat[5]) );
  SDFFRQX1 mem_reg_4_ ( .D(wdat[4]), .SIN(rdat[3]), .SMC(test_se), .C(net11792), .XR(arstz), .Q(rdat[4]) );
  SDFFRQX1 mem_reg_3_ ( .D(wdat[3]), .SIN(rdat[2]), .SMC(test_se), .C(net11792), .XR(arstz), .Q(rdat[3]) );
  SDFFRQX1 mem_reg_2_ ( .D(wdat[2]), .SIN(rdat[1]), .SMC(test_se), .C(net11792), .XR(arstz), .Q(rdat[2]) );
  SDFFRQX1 mem_reg_1_ ( .D(wdat[1]), .SIN(rdat[0]), .SMC(test_se), .C(net11792), .XR(arstz), .Q(rdat[1]) );
  SDFFRQX1 mem_reg_0_ ( .D(wdat[0]), .SIN(test_si), .SMC(test_se), .C(net11792), .XR(arstz), .Q(rdat[0]) );
  SDFFRQX1 mem_reg_6_ ( .D(wdat[6]), .SIN(rdat[5]), .SMC(test_se), .C(net11792), .XR(arstz), .Q(rdat[6]) );
  SDFFRQX1 mem_reg_7_ ( .D(wdat[7]), .SIN(rdat[6]), .SMC(test_se), .C(net11792), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_79 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ictlr_a0 ( bkpt_ena, bkpt_pc, memaddr_c, memaddr, mcu_psr_c, mcu_psw, 
        hit_ps_c, hit_ps, mempsack, memdatao, o_set_hold, o_bkp_hold, 
        o_ofs_inc, o_inst, d_inst, sfr_psrack, sfr_psofs, sfr_psr, sfr_psw, 
        dw_rst, dw_ena, sfr_wdat, pmem_pgm, pmem_re, pmem_csb, pmem_clk, 
        pmem_a, pmem_q0, pmem_q1, pmem_twlb, wd_twlb, we_twlb, pwrdn_rst, 
        r_pwdn_en, r_multi, r_hold_mcu, clk, srst, test_si3, test_si2, 
        test_si1, test_so2, test_so1, test_se );
  input [14:0] bkpt_pc;
  input [14:0] memaddr_c;
  input [14:0] memaddr;
  input [7:0] memdatao;
  output [7:0] o_inst;
  output [7:0] d_inst;
  input [14:0] sfr_psofs;
  input [7:0] sfr_wdat;
  output [1:0] pmem_clk;
  output [15:0] pmem_a;
  input [7:0] pmem_q0;
  input [7:0] pmem_q1;
  output [1:0] pmem_twlb;
  input [1:0] wd_twlb;
  input bkpt_ena, mcu_psr_c, mcu_psw, hit_ps_c, hit_ps, sfr_psr, sfr_psw,
         dw_rst, dw_ena, we_twlb, pwrdn_rst, r_pwdn_en, r_multi, r_hold_mcu,
         clk, srst, test_si3, test_si2, test_si1, test_se;
  output mempsack, o_set_hold, o_bkp_hold, o_ofs_inc, sfr_psrack, pmem_pgm,
         pmem_re, pmem_csb, test_so2, test_so1;
  wire   N152, N153, N154, c_buf_22__7_, c_buf_22__6_, c_buf_22__5_,
         c_buf_22__4_, c_buf_22__3_, c_buf_22__2_, c_buf_22__1_, c_buf_22__0_,
         c_buf_21__7_, c_buf_21__6_, c_buf_21__5_, c_buf_21__4_, c_buf_21__3_,
         c_buf_21__2_, c_buf_21__1_, c_buf_21__0_, c_buf_20__7_, c_buf_20__6_,
         c_buf_20__5_, c_buf_20__4_, c_buf_20__3_, c_buf_20__2_, c_buf_20__1_,
         c_buf_20__0_, c_buf_19__7_, c_buf_19__6_, c_buf_19__5_, c_buf_19__4_,
         c_buf_19__3_, c_buf_19__2_, c_buf_19__1_, c_buf_19__0_, c_buf_18__7_,
         c_buf_18__6_, c_buf_18__5_, c_buf_18__4_, c_buf_18__3_, c_buf_18__2_,
         c_buf_18__1_, c_buf_18__0_, c_buf_17__7_, c_buf_17__6_, c_buf_17__5_,
         c_buf_17__4_, c_buf_17__3_, c_buf_17__2_, c_buf_17__1_, c_buf_17__0_,
         c_buf_16__7_, c_buf_16__6_, c_buf_16__5_, c_buf_16__4_, c_buf_16__3_,
         c_buf_16__2_, c_buf_16__1_, c_buf_16__0_, wspp_cnt_5_, wspp_cnt_4_,
         wspp_cnt_3_, wspp_cnt_2_, wspp_cnt_1_, wspp_cnt_0_, d_psrd, r_rdy,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617,
         N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628,
         N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639,
         N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650,
         N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661,
         N662, N757, N759, N786, N787, N788, N789, N790, N791, N792, N793,
         N795, N796, N797, N798, N799, N800, N801, N820, N821, N822, N823,
         N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834,
         N835, N836, N837, N838, N839, N840, N842, N843, N844, N845, N846,
         N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863,
         N864, N865, N866, N867, N868, N874, N875, N876, N877, N878, N879,
         N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890,
         N891, N892, N893, N894, N895, N896, N897, N898, N899, un_hold,
         net11818, net11824, net11829, net11834, net11839, net11844, net11849,
         net11854, net11859, net11864, net11869, net11874, net11879, net11884,
         net11889, net11894, net11899, net11904, net11909, net11914, net11919,
         net11924, net11929, net11934, net11939, net11944, net11949, net11954,
         net11959, net11964, n93, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n923, n249, n250, n251, n252, n253, n254,
         n255, n259, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n415, n416, n420, n453, n459, n460, n461, n464, n465, n466,
         n470, n502, n529, n532, n543, n546, n547, n550, n553, n554, n555,
         n556, n557, n558, n575, n576, n577, n578, n579, n589, n590, n591,
         n593, n603, n605, n606, n607, n608, n609, n610, n611, n615, n621,
         n625, n682, n693, n709, n710, n711, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n762, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n256, n257, n258, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n412, n413,
         n414, n417, n418, n419, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n454, n455, n456, n457, n458, n462, n463, n467,
         n468, n469, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n530, n531, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n544, n545, n548, n549, n551, n552,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n592, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n604, n612, n613, n614, n616, n617, n618, n619, n620,
         n622, n623, n624, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n712, n713, n714, n733,
         n734, n748, n749, n759, n760, n761, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951;
  wire   [3:0] d_hold;
  wire   [1:0] dummy;
  wire   [3:0] cs_ft;
  wire   [4:0] c_ptr;
  wire   [14:0] c_adr;
  wire   [14:13] adr_p;
  wire   [7:0] rd_buf;
  wire   [7:0] dbg_01;
  wire   [7:0] dbg_02;
  wire   [7:0] dbg_03;
  wire   [7:0] dbg_04;
  wire   [7:0] dbg_05;
  wire   [7:0] dbg_06;
  wire   [7:0] dbg_07;
  wire   [7:0] dbg_08;
  wire   [7:0] dbg_09;
  wire   [7:0] dbg_0a;
  wire   [7:0] dbg_0b;
  wire   [7:0] dbg_0c;
  wire   [7:0] dbg_0d;
  wire   [7:0] dbg_0e;
  wire   [7:0] dbg_0f;
  wire   [7:0] wr_buf;
  wire   [14:0] pre_1_adr;

  SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 clk_gate_wspp_cnt_reg ( .CLK(clk), .EN(N899), 
        .ENCLK(net11818), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 clk_gate_a_bit_reg ( .CLK(clk), .EN(N898), 
        .ENCLK(net11824), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 clk_gate_adr_p_reg ( .CLK(clk), .EN(N853), 
        .ENCLK(net11829), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 clk_gate_c_buf_reg_23_ ( .CLK(clk), .EN(
        N897), .ENCLK(net11834), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 clk_gate_c_buf_reg_22_ ( .CLK(clk), .EN(
        N896), .ENCLK(net11839), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 clk_gate_c_buf_reg_21_ ( .CLK(clk), .EN(
        N895), .ENCLK(net11844), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 clk_gate_c_buf_reg_20_ ( .CLK(clk), .EN(
        N894), .ENCLK(net11849), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 clk_gate_c_buf_reg_19_ ( .CLK(clk), .EN(
        N893), .ENCLK(net11854), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 clk_gate_c_buf_reg_18_ ( .CLK(clk), .EN(
        N892), .ENCLK(net11859), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 clk_gate_c_buf_reg_17_ ( .CLK(clk), .EN(
        N891), .ENCLK(net11864), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 clk_gate_c_buf_reg_16_ ( .CLK(clk), .EN(
        N890), .ENCLK(net11869), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 clk_gate_c_buf_reg_15_ ( .CLK(clk), .EN(
        N889), .ENCLK(net11874), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 clk_gate_c_buf_reg_14_ ( .CLK(clk), .EN(
        N888), .ENCLK(net11879), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 clk_gate_c_buf_reg_13_ ( .CLK(clk), .EN(
        N887), .ENCLK(net11884), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 clk_gate_c_buf_reg_12_ ( .CLK(clk), .EN(
        N886), .ENCLK(net11889), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 clk_gate_c_buf_reg_11_ ( .CLK(clk), .EN(
        N885), .ENCLK(net11894), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 clk_gate_c_buf_reg_10_ ( .CLK(clk), .EN(
        N884), .ENCLK(net11899), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 clk_gate_c_buf_reg_9_ ( .CLK(clk), .EN(N883), .ENCLK(net11904), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 clk_gate_c_buf_reg_8_ ( .CLK(clk), .EN(N882), .ENCLK(net11909), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 clk_gate_c_buf_reg_7_ ( .CLK(clk), .EN(N881), .ENCLK(net11914), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 clk_gate_c_buf_reg_6_ ( .CLK(clk), .EN(N880), .ENCLK(net11919), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 clk_gate_c_buf_reg_5_ ( .CLK(clk), .EN(N879), 
        .ENCLK(net11924), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 clk_gate_c_buf_reg_4_ ( .CLK(clk), .EN(N878), 
        .ENCLK(net11929), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 clk_gate_c_buf_reg_3_ ( .CLK(clk), .EN(N877), 
        .ENCLK(net11934), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 clk_gate_c_buf_reg_2_ ( .CLK(clk), .EN(N876), 
        .ENCLK(net11939), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 clk_gate_c_buf_reg_1_ ( .CLK(clk), .EN(N875), 
        .ENCLK(net11944), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 clk_gate_c_buf_reg_0_ ( .CLK(clk), .EN(N874), 
        .ENCLK(net11949), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 clk_gate_c_ptr_reg ( .CLK(clk), .EN(n93), 
        .ENCLK(net11954), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 clk_gate_c_adr_reg ( .CLK(clk), .EN(N825), 
        .ENCLK(net11959), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 clk_gate_cs_ft_reg ( .CLK(clk), .EN(N820), 
        .ENCLK(net11964), .TE(test_se) );
  ictlr_a0_DW01_inc_1 add_242 ( .A(c_adr), .SUM({N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431}) );
  ictlr_a0_DW01_inc_2 r492 ( .A({adr_p, pmem_a[15:9], pmem_a[5:0]}), .SUM(
        pre_1_adr) );
  SDFFNQXL ck_n_reg_1_ ( .D(n642), .SIN(pmem_clk[0]), .SMC(test_se), .XC(clk), 
        .Q(pmem_clk[1]) );
  SDFFNQX1 ck_n_reg_0_ ( .D(n641), .SIN(test_si1), .SMC(test_se), .XC(clk), 
        .Q(pmem_clk[0]) );
  SDFFQX2 a_bit_reg_2_ ( .D(N759), .SIN(pmem_a[7]), .SMC(test_se), .C(net11824), .Q(pmem_a[8]) );
  SDFFQX2 a_bit_reg_0_ ( .D(N757), .SIN(test_si2), .SMC(test_se), .C(net11824), 
        .Q(pmem_a[6]) );
  SDFFQX1 wspp_cnt_reg_1_ ( .D(N796), .SIN(wspp_cnt_0_), .SMC(test_se), .C(
        net11818), .Q(wspp_cnt_1_) );
  SDFFQX1 wspp_cnt_reg_2_ ( .D(N797), .SIN(wspp_cnt_1_), .SMC(test_se), .C(
        net11818), .Q(wspp_cnt_2_) );
  SDFFQX1 wspp_cnt_reg_0_ ( .D(N795), .SIN(un_hold), .SMC(test_se), .C(
        net11818), .Q(wspp_cnt_0_) );
  SDFFQX1 d_hold_reg_0_ ( .D(n923), .SIN(cs_ft[3]), .SMC(test_se), .C(clk), 
        .Q(d_hold[0]) );
  SDFFQX1 d_hold_reg_3_ ( .D(N154), .SIN(d_hold[2]), .SMC(test_se), .C(clk), 
        .Q(d_hold[3]) );
  SDFFQX1 dummy_reg_0_ ( .D(n651), .SIN(n24), .SMC(test_se), .C(clk), .Q(
        dummy[0]) );
  SDFFQX1 d_hold_reg_1_ ( .D(N152), .SIN(d_hold[0]), .SMC(test_se), .C(clk), 
        .Q(d_hold[1]) );
  SDFFQX1 d_hold_reg_2_ ( .D(N153), .SIN(d_hold[1]), .SMC(test_se), .C(clk), 
        .Q(d_hold[2]) );
  SDFFQX1 dummy_reg_1_ ( .D(n650), .SIN(dummy[0]), .SMC(test_se), .C(clk), .Q(
        dummy[1]) );
  SDFFQX2 adr_p_reg_4_ ( .D(N858), .SIN(pmem_a[3]), .SMC(test_se), .C(net11829), .Q(pmem_a[4]) );
  SDFFQX2 adr_p_reg_3_ ( .D(N857), .SIN(pmem_a[2]), .SMC(test_se), .C(net11829), .Q(pmem_a[3]) );
  SDFFQX2 adr_p_reg_5_ ( .D(N859), .SIN(pmem_a[4]), .SMC(test_se), .C(net11829), .Q(pmem_a[5]) );
  SDFFQX1 d_psrd_reg ( .D(n649), .SIN(d_hold[3]), .SMC(test_se), .C(net11964), 
        .Q(d_psrd) );
  SDFFQX2 adr_p_reg_2_ ( .D(N856), .SIN(pmem_a[1]), .SMC(test_se), .C(net11829), .Q(pmem_a[2]) );
  SDFFQX2 adr_p_reg_1_ ( .D(N855), .SIN(pmem_a[0]), .SMC(test_se), .C(net11829), .Q(pmem_a[1]) );
  SDFFQX1 c_adr_reg_14_ ( .D(N840), .SIN(c_adr[13]), .SMC(test_se), .C(
        net11959), .Q(c_adr[14]) );
  SDFFQX1 c_adr_reg_13_ ( .D(N839), .SIN(c_adr[12]), .SMC(test_se), .C(
        net11959), .Q(c_adr[13]) );
  SDFFQX1 c_adr_reg_12_ ( .D(N838), .SIN(c_adr[11]), .SMC(test_se), .C(
        net11959), .Q(c_adr[12]) );
  SDFFQX1 c_adr_reg_11_ ( .D(N837), .SIN(c_adr[10]), .SMC(test_se), .C(
        net11959), .Q(c_adr[11]) );
  SDFFQX1 c_adr_reg_10_ ( .D(N836), .SIN(c_adr[9]), .SMC(test_se), .C(net11959), .Q(c_adr[10]) );
  SDFFQX1 c_adr_reg_7_ ( .D(N833), .SIN(c_adr[6]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[7]) );
  SDFFQX1 c_adr_reg_8_ ( .D(N834), .SIN(c_adr[7]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[8]) );
  SDFFQX1 c_adr_reg_9_ ( .D(N835), .SIN(c_adr[8]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[9]) );
  SDFFQX1 c_adr_reg_6_ ( .D(N832), .SIN(c_adr[5]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[6]) );
  SDFFQX1 c_ptr_reg_4_ ( .D(N846), .SIN(c_ptr[3]), .SMC(test_se), .C(net11954), 
        .Q(c_ptr[4]) );
  SDFFQX1 c_adr_reg_5_ ( .D(N831), .SIN(c_adr[4]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[5]) );
  SDFFQX1 c_ptr_reg_3_ ( .D(N845), .SIN(c_ptr[2]), .SMC(test_se), .C(net11954), 
        .Q(c_ptr[3]) );
  SDFFQX1 c_ptr_reg_2_ ( .D(N844), .SIN(c_ptr[1]), .SMC(test_se), .C(net11954), 
        .Q(c_ptr[2]) );
  SDFFQX1 c_ptr_reg_1_ ( .D(N843), .SIN(c_ptr[0]), .SMC(test_se), .C(net11954), 
        .Q(c_ptr[1]) );
  SDFFQX1 c_ptr_reg_0_ ( .D(N842), .SIN(wr_buf[7]), .SMC(test_se), .C(net11954), .Q(c_ptr[0]) );
  SDFFQX1 adr_p_reg_14_ ( .D(N868), .SIN(adr_p[13]), .SMC(test_se), .C(
        net11829), .Q(adr_p[14]) );
  SDFFQX1 adr_p_reg_13_ ( .D(N867), .SIN(pmem_a[14]), .SMC(test_se), .C(
        net11829), .Q(adr_p[13]) );
  SDFFQX2 adr_p_reg_9_ ( .D(N863), .SIN(pmem_a[11]), .SMC(test_se), .C(
        net11829), .Q(pmem_a[12]) );
  SDFFQX1 wspp_cnt_reg_3_ ( .D(N798), .SIN(wspp_cnt_2_), .SMC(test_se), .C(
        net11818), .Q(wspp_cnt_3_) );
  SDFFQX1 wspp_cnt_reg_5_ ( .D(N800), .SIN(wspp_cnt_4_), .SMC(test_se), .C(
        net11818), .Q(wspp_cnt_5_) );
  SDFFQX1 wspp_cnt_reg_6_ ( .D(N801), .SIN(wspp_cnt_5_), .SMC(test_se), .C(
        net11818), .Q(test_so2) );
  SDFFQX1 wspp_cnt_reg_4_ ( .D(N799), .SIN(wspp_cnt_3_), .SMC(test_se), .C(
        net11818), .Q(wspp_cnt_4_) );
  SDFFQX2 adr_p_reg_7_ ( .D(N861), .SIN(pmem_a[9]), .SMC(test_se), .C(net11829), .Q(pmem_a[10]) );
  SDFFQX2 adr_p_reg_10_ ( .D(N864), .SIN(pmem_a[12]), .SMC(test_se), .C(
        net11829), .Q(pmem_a[13]) );
  SDFFQX2 adr_p_reg_11_ ( .D(N865), .SIN(pmem_a[13]), .SMC(test_se), .C(
        net11829), .Q(pmem_a[14]) );
  SDFFQX2 adr_p_reg_12_ ( .D(N866), .SIN(test_si3), .SMC(test_se), .C(net11829), .Q(pmem_a[15]) );
  SDFFNQXL cs_n_reg ( .D(n643), .SIN(pmem_clk[1]), .SMC(test_se), .XC(clk), 
        .Q(test_so1) );
  SDFFQX1 re_p_reg ( .D(n647), .SIN(pmem_twlb[1]), .SMC(test_se), .C(clk), .Q(
        pmem_re) );
  SDFFQX1 pgm_p_reg ( .D(n644), .SIN(dummy[1]), .SMC(test_se), .C(net11964), 
        .Q(pmem_pgm) );
  SDFFQX1 un_hold_reg ( .D(n762), .SIN(pmem_re), .SMC(test_se), .C(clk), .Q(
        un_hold) );
  SDFFQX1 r_rdy_reg ( .D(n648), .SIN(pmem_pgm), .SMC(test_se), .C(clk), .Q(
        r_rdy) );
  SDFFQX1 r_twlb_reg_1_ ( .D(n645), .SIN(pmem_twlb[0]), .SMC(test_se), .C(clk), 
        .Q(pmem_twlb[1]) );
  SDFFQX1 r_twlb_reg_0_ ( .D(n646), .SIN(r_rdy), .SMC(test_se), .C(clk), .Q(
        pmem_twlb[0]) );
  SDFFQX1 c_buf_reg_0__2_ ( .D(N481), .SIN(rd_buf[1]), .SMC(test_se), .C(
        net11949), .Q(rd_buf[2]) );
  SDFFQX1 c_buf_reg_0__1_ ( .D(N480), .SIN(rd_buf[0]), .SMC(test_se), .C(
        net11949), .Q(rd_buf[1]) );
  SDFFQX1 c_buf_reg_0__0_ ( .D(N479), .SIN(c_adr[14]), .SMC(test_se), .C(
        net11949), .Q(rd_buf[0]) );
  SDFFQX1 c_buf_reg_20__2_ ( .D(N641), .SIN(c_buf_20__1_), .SMC(test_se), .C(
        net11849), .Q(c_buf_20__2_) );
  SDFFQX1 c_buf_reg_22__5_ ( .D(N660), .SIN(c_buf_22__4_), .SMC(test_se), .C(
        net11839), .Q(c_buf_22__5_) );
  SDFFQX1 c_buf_reg_22__4_ ( .D(N659), .SIN(c_buf_22__3_), .SMC(test_se), .C(
        net11839), .Q(c_buf_22__4_) );
  SDFFQX1 c_buf_reg_22__3_ ( .D(N658), .SIN(c_buf_22__2_), .SMC(test_se), .C(
        net11839), .Q(c_buf_22__3_) );
  SDFFQX1 c_buf_reg_22__2_ ( .D(N657), .SIN(c_buf_22__1_), .SMC(test_se), .C(
        net11839), .Q(c_buf_22__2_) );
  SDFFQX1 c_buf_reg_22__1_ ( .D(N656), .SIN(c_buf_22__0_), .SMC(test_se), .C(
        net11839), .Q(c_buf_22__1_) );
  SDFFQX1 c_buf_reg_22__0_ ( .D(N655), .SIN(c_buf_21__7_), .SMC(test_se), .C(
        net11839), .Q(c_buf_22__0_) );
  SDFFQX1 c_buf_reg_21__4_ ( .D(N651), .SIN(c_buf_21__3_), .SMC(test_se), .C(
        net11844), .Q(c_buf_21__4_) );
  SDFFQX1 c_buf_reg_21__2_ ( .D(N649), .SIN(c_buf_21__1_), .SMC(test_se), .C(
        net11844), .Q(c_buf_21__2_) );
  SDFFQX1 c_buf_reg_21__1_ ( .D(N648), .SIN(c_buf_21__0_), .SMC(test_se), .C(
        net11844), .Q(c_buf_21__1_) );
  SDFFQX1 c_buf_reg_21__0_ ( .D(N647), .SIN(c_buf_20__7_), .SMC(test_se), .C(
        net11844), .Q(c_buf_21__0_) );
  SDFFQX1 c_buf_reg_20__4_ ( .D(N643), .SIN(c_buf_20__3_), .SMC(test_se), .C(
        net11849), .Q(c_buf_20__4_) );
  SDFFQX1 c_buf_reg_20__3_ ( .D(N642), .SIN(c_buf_20__2_), .SMC(test_se), .C(
        net11849), .Q(c_buf_20__3_) );
  SDFFQX1 c_buf_reg_20__1_ ( .D(N640), .SIN(c_buf_20__0_), .SMC(test_se), .C(
        net11849), .Q(c_buf_20__1_) );
  SDFFQX1 c_buf_reg_20__0_ ( .D(N639), .SIN(c_buf_19__7_), .SMC(test_se), .C(
        net11849), .Q(c_buf_20__0_) );
  SDFFQX1 c_buf_reg_19__5_ ( .D(N636), .SIN(c_buf_19__4_), .SMC(test_se), .C(
        net11854), .Q(c_buf_19__5_) );
  SDFFQX1 c_buf_reg_19__4_ ( .D(N635), .SIN(c_buf_19__3_), .SMC(test_se), .C(
        net11854), .Q(c_buf_19__4_) );
  SDFFQX1 c_buf_reg_19__3_ ( .D(N634), .SIN(c_buf_19__2_), .SMC(test_se), .C(
        net11854), .Q(c_buf_19__3_) );
  SDFFQX1 c_buf_reg_19__2_ ( .D(N633), .SIN(c_buf_19__1_), .SMC(test_se), .C(
        net11854), .Q(c_buf_19__2_) );
  SDFFQX1 c_buf_reg_19__1_ ( .D(N632), .SIN(c_buf_19__0_), .SMC(test_se), .C(
        net11854), .Q(c_buf_19__1_) );
  SDFFQX1 c_buf_reg_19__0_ ( .D(N631), .SIN(c_buf_18__7_), .SMC(test_se), .C(
        net11854), .Q(c_buf_19__0_) );
  SDFFQX1 c_buf_reg_18__4_ ( .D(N627), .SIN(c_buf_18__3_), .SMC(test_se), .C(
        net11859), .Q(c_buf_18__4_) );
  SDFFQX1 c_buf_reg_18__2_ ( .D(N625), .SIN(c_buf_18__1_), .SMC(test_se), .C(
        net11859), .Q(c_buf_18__2_) );
  SDFFQX1 c_buf_reg_18__1_ ( .D(N624), .SIN(c_buf_18__0_), .SMC(test_se), .C(
        net11859), .Q(c_buf_18__1_) );
  SDFFQX1 c_buf_reg_18__0_ ( .D(N623), .SIN(c_buf_17__7_), .SMC(test_se), .C(
        net11859), .Q(c_buf_18__0_) );
  SDFFQX1 c_buf_reg_17__4_ ( .D(N619), .SIN(c_buf_17__3_), .SMC(test_se), .C(
        net11864), .Q(c_buf_17__4_) );
  SDFFQX1 c_buf_reg_17__2_ ( .D(N617), .SIN(c_buf_17__1_), .SMC(test_se), .C(
        net11864), .Q(c_buf_17__2_) );
  SDFFQX1 c_buf_reg_17__1_ ( .D(N616), .SIN(c_buf_17__0_), .SMC(test_se), .C(
        net11864), .Q(c_buf_17__1_) );
  SDFFQX1 c_buf_reg_17__0_ ( .D(N615), .SIN(c_buf_16__7_), .SMC(test_se), .C(
        net11864), .Q(c_buf_17__0_) );
  SDFFQX1 c_buf_reg_16__4_ ( .D(N611), .SIN(c_buf_16__3_), .SMC(test_se), .C(
        net11869), .Q(c_buf_16__4_) );
  SDFFQX1 c_buf_reg_16__2_ ( .D(N609), .SIN(c_buf_16__1_), .SMC(test_se), .C(
        net11869), .Q(c_buf_16__2_) );
  SDFFQX1 c_buf_reg_16__1_ ( .D(N608), .SIN(c_buf_16__0_), .SMC(test_se), .C(
        net11869), .Q(c_buf_16__1_) );
  SDFFQX1 c_buf_reg_16__0_ ( .D(N607), .SIN(dbg_0f[7]), .SMC(test_se), .C(
        net11869), .Q(c_buf_16__0_) );
  SDFFQX1 c_buf_reg_15__4_ ( .D(N603), .SIN(dbg_0f[3]), .SMC(test_se), .C(
        net11874), .Q(dbg_0f[4]) );
  SDFFQX1 c_buf_reg_15__2_ ( .D(N601), .SIN(dbg_0f[1]), .SMC(test_se), .C(
        net11874), .Q(dbg_0f[2]) );
  SDFFQX1 c_buf_reg_15__1_ ( .D(N600), .SIN(dbg_0f[0]), .SMC(test_se), .C(
        net11874), .Q(dbg_0f[1]) );
  SDFFQX1 c_buf_reg_15__0_ ( .D(N599), .SIN(dbg_0e[7]), .SMC(test_se), .C(
        net11874), .Q(dbg_0f[0]) );
  SDFFQX1 c_buf_reg_14__4_ ( .D(N595), .SIN(dbg_0e[3]), .SMC(test_se), .C(
        net11879), .Q(dbg_0e[4]) );
  SDFFQX1 c_buf_reg_14__2_ ( .D(N593), .SIN(dbg_0e[1]), .SMC(test_se), .C(
        net11879), .Q(dbg_0e[2]) );
  SDFFQX1 c_buf_reg_14__1_ ( .D(N592), .SIN(dbg_0e[0]), .SMC(test_se), .C(
        net11879), .Q(dbg_0e[1]) );
  SDFFQX1 c_buf_reg_14__0_ ( .D(N591), .SIN(dbg_0d[7]), .SMC(test_se), .C(
        net11879), .Q(dbg_0e[0]) );
  SDFFQX1 c_buf_reg_13__4_ ( .D(N587), .SIN(dbg_0d[3]), .SMC(test_se), .C(
        net11884), .Q(dbg_0d[4]) );
  SDFFQX1 c_buf_reg_13__2_ ( .D(N585), .SIN(dbg_0d[1]), .SMC(test_se), .C(
        net11884), .Q(dbg_0d[2]) );
  SDFFQX1 c_buf_reg_13__1_ ( .D(N584), .SIN(dbg_0d[0]), .SMC(test_se), .C(
        net11884), .Q(dbg_0d[1]) );
  SDFFQX1 c_buf_reg_13__0_ ( .D(N583), .SIN(dbg_0c[7]), .SMC(test_se), .C(
        net11884), .Q(dbg_0d[0]) );
  SDFFQX1 c_buf_reg_12__4_ ( .D(N579), .SIN(dbg_0c[3]), .SMC(test_se), .C(
        net11889), .Q(dbg_0c[4]) );
  SDFFQX1 c_buf_reg_12__2_ ( .D(N577), .SIN(dbg_0c[1]), .SMC(test_se), .C(
        net11889), .Q(dbg_0c[2]) );
  SDFFQX1 c_buf_reg_12__1_ ( .D(N576), .SIN(dbg_0c[0]), .SMC(test_se), .C(
        net11889), .Q(dbg_0c[1]) );
  SDFFQX1 c_buf_reg_12__0_ ( .D(N575), .SIN(dbg_0b[7]), .SMC(test_se), .C(
        net11889), .Q(dbg_0c[0]) );
  SDFFQX1 c_buf_reg_11__2_ ( .D(N569), .SIN(dbg_0b[1]), .SMC(test_se), .C(
        net11894), .Q(dbg_0b[2]) );
  SDFFQX1 c_buf_reg_10__2_ ( .D(N561), .SIN(dbg_0a[1]), .SMC(test_se), .C(
        net11899), .Q(dbg_0a[2]) );
  SDFFQX1 c_buf_reg_9__2_ ( .D(N553), .SIN(dbg_09[1]), .SMC(test_se), .C(
        net11904), .Q(dbg_09[2]) );
  SDFFQX1 c_buf_reg_8__2_ ( .D(N545), .SIN(dbg_08[1]), .SMC(test_se), .C(
        net11909), .Q(dbg_08[2]) );
  SDFFQX1 c_buf_reg_7__2_ ( .D(N537), .SIN(dbg_07[1]), .SMC(test_se), .C(
        net11914), .Q(dbg_07[2]) );
  SDFFQX1 c_buf_reg_6__2_ ( .D(N529), .SIN(dbg_06[1]), .SMC(test_se), .C(
        net11919), .Q(dbg_06[2]) );
  SDFFQX1 c_buf_reg_5__2_ ( .D(N521), .SIN(dbg_05[1]), .SMC(test_se), .C(
        net11924), .Q(dbg_05[2]) );
  SDFFQX1 c_buf_reg_4__2_ ( .D(N513), .SIN(dbg_04[1]), .SMC(test_se), .C(
        net11929), .Q(dbg_04[2]) );
  SDFFQX1 c_buf_reg_3__2_ ( .D(N505), .SIN(dbg_03[1]), .SMC(test_se), .C(
        net11934), .Q(dbg_03[2]) );
  SDFFQX1 c_buf_reg_2__2_ ( .D(N497), .SIN(dbg_02[1]), .SMC(test_se), .C(
        net11939), .Q(dbg_02[2]) );
  SDFFQX1 c_buf_reg_1__2_ ( .D(N489), .SIN(dbg_01[1]), .SMC(test_se), .C(
        net11944), .Q(dbg_01[2]) );
  SDFFQX1 c_buf_reg_16__3_ ( .D(N610), .SIN(c_buf_16__2_), .SMC(test_se), .C(
        net11869), .Q(c_buf_16__3_) );
  SDFFQX1 c_buf_reg_23__2_ ( .D(N788), .SIN(wr_buf[1]), .SMC(test_se), .C(
        net11834), .Q(wr_buf[2]) );
  SDFFQX1 c_buf_reg_23__4_ ( .D(N790), .SIN(wr_buf[3]), .SMC(test_se), .C(
        net11834), .Q(wr_buf[4]) );
  SDFFQX1 c_buf_reg_23__1_ ( .D(N787), .SIN(wr_buf[0]), .SMC(test_se), .C(
        net11834), .Q(wr_buf[1]) );
  SDFFQX1 c_buf_reg_23__0_ ( .D(N786), .SIN(c_buf_22__7_), .SMC(test_se), .C(
        net11834), .Q(wr_buf[0]) );
  SDFFQX1 cs_ft_reg_1_ ( .D(N822), .SIN(cs_ft[0]), .SMC(test_se), .C(net11964), 
        .Q(cs_ft[1]) );
  SDFFQX1 cs_ft_reg_3_ ( .D(N824), .SIN(cs_ft[2]), .SMC(test_se), .C(net11964), 
        .Q(cs_ft[3]) );
  SDFFQX1 cs_ft_reg_2_ ( .D(N823), .SIN(cs_ft[1]), .SMC(test_se), .C(net11964), 
        .Q(cs_ft[2]) );
  SDFFQX1 cs_ft_reg_0_ ( .D(N821), .SIN(c_ptr[4]), .SMC(test_se), .C(net11964), 
        .Q(cs_ft[0]) );
  SDFFQX1 c_buf_reg_0__6_ ( .D(N485), .SIN(rd_buf[5]), .SMC(test_se), .C(
        net11949), .Q(rd_buf[6]) );
  SDFFQX1 c_buf_reg_0__5_ ( .D(N484), .SIN(rd_buf[4]), .SMC(test_se), .C(
        net11949), .Q(rd_buf[5]) );
  SDFFQX1 c_buf_reg_0__3_ ( .D(N482), .SIN(rd_buf[2]), .SMC(test_se), .C(
        net11949), .Q(rd_buf[3]) );
  SDFFQX1 c_buf_reg_0__4_ ( .D(N483), .SIN(rd_buf[3]), .SMC(test_se), .C(
        net11949), .Q(rd_buf[4]) );
  SDFFQX1 c_buf_reg_0__7_ ( .D(N486), .SIN(rd_buf[6]), .SMC(test_se), .C(
        net11949), .Q(rd_buf[7]) );
  SDFFQX1 c_buf_reg_22__6_ ( .D(N661), .SIN(c_buf_22__5_), .SMC(test_se), .C(
        net11839), .Q(c_buf_22__6_) );
  SDFFQX1 c_buf_reg_21__6_ ( .D(N653), .SIN(c_buf_21__5_), .SMC(test_se), .C(
        net11844), .Q(c_buf_21__6_) );
  SDFFQX1 c_buf_reg_21__5_ ( .D(N652), .SIN(c_buf_21__4_), .SMC(test_se), .C(
        net11844), .Q(c_buf_21__5_) );
  SDFFQX1 c_buf_reg_21__3_ ( .D(N650), .SIN(c_buf_21__2_), .SMC(test_se), .C(
        net11844), .Q(c_buf_21__3_) );
  SDFFQX1 c_buf_reg_20__6_ ( .D(N645), .SIN(c_buf_20__5_), .SMC(test_se), .C(
        net11849), .Q(c_buf_20__6_) );
  SDFFQX1 c_buf_reg_20__5_ ( .D(N644), .SIN(c_buf_20__4_), .SMC(test_se), .C(
        net11849), .Q(c_buf_20__5_) );
  SDFFQX1 c_buf_reg_19__6_ ( .D(N637), .SIN(c_buf_19__5_), .SMC(test_se), .C(
        net11854), .Q(c_buf_19__6_) );
  SDFFQX1 c_buf_reg_18__6_ ( .D(N629), .SIN(c_buf_18__5_), .SMC(test_se), .C(
        net11859), .Q(c_buf_18__6_) );
  SDFFQX1 c_buf_reg_18__5_ ( .D(N628), .SIN(c_buf_18__4_), .SMC(test_se), .C(
        net11859), .Q(c_buf_18__5_) );
  SDFFQX1 c_buf_reg_18__3_ ( .D(N626), .SIN(c_buf_18__2_), .SMC(test_se), .C(
        net11859), .Q(c_buf_18__3_) );
  SDFFQX1 c_buf_reg_17__6_ ( .D(N621), .SIN(c_buf_17__5_), .SMC(test_se), .C(
        net11864), .Q(c_buf_17__6_) );
  SDFFQX1 c_buf_reg_17__5_ ( .D(N620), .SIN(c_buf_17__4_), .SMC(test_se), .C(
        net11864), .Q(c_buf_17__5_) );
  SDFFQX1 c_buf_reg_17__3_ ( .D(N618), .SIN(c_buf_17__2_), .SMC(test_se), .C(
        net11864), .Q(c_buf_17__3_) );
  SDFFQX1 c_buf_reg_16__6_ ( .D(N613), .SIN(c_buf_16__5_), .SMC(test_se), .C(
        net11869), .Q(c_buf_16__6_) );
  SDFFQX1 c_buf_reg_16__5_ ( .D(N612), .SIN(c_buf_16__4_), .SMC(test_se), .C(
        net11869), .Q(c_buf_16__5_) );
  SDFFQX1 c_buf_reg_15__5_ ( .D(N604), .SIN(dbg_0f[4]), .SMC(test_se), .C(
        net11874), .Q(dbg_0f[5]) );
  SDFFQX1 c_buf_reg_14__6_ ( .D(N597), .SIN(dbg_0e[5]), .SMC(test_se), .C(
        net11879), .Q(dbg_0e[6]) );
  SDFFQX1 c_buf_reg_14__5_ ( .D(N596), .SIN(dbg_0e[4]), .SMC(test_se), .C(
        net11879), .Q(dbg_0e[5]) );
  SDFFQX1 c_buf_reg_14__3_ ( .D(N594), .SIN(dbg_0e[2]), .SMC(test_se), .C(
        net11879), .Q(dbg_0e[3]) );
  SDFFQX1 c_buf_reg_13__5_ ( .D(N588), .SIN(dbg_0d[4]), .SMC(test_se), .C(
        net11884), .Q(dbg_0d[5]) );
  SDFFQX1 c_buf_reg_12__5_ ( .D(N580), .SIN(dbg_0c[4]), .SMC(test_se), .C(
        net11889), .Q(dbg_0c[5]) );
  SDFFQX1 c_buf_reg_11__1_ ( .D(N568), .SIN(dbg_0b[0]), .SMC(test_se), .C(
        net11894), .Q(dbg_0b[1]) );
  SDFFQX1 c_buf_reg_10__1_ ( .D(N560), .SIN(dbg_0a[0]), .SMC(test_se), .C(
        net11899), .Q(dbg_0a[1]) );
  SDFFQX1 c_buf_reg_9__4_ ( .D(N555), .SIN(dbg_09[3]), .SMC(test_se), .C(
        net11904), .Q(dbg_09[4]) );
  SDFFQX1 c_buf_reg_9__1_ ( .D(N552), .SIN(dbg_09[0]), .SMC(test_se), .C(
        net11904), .Q(dbg_09[1]) );
  SDFFQX1 c_buf_reg_9__0_ ( .D(N551), .SIN(dbg_08[7]), .SMC(test_se), .C(
        net11904), .Q(dbg_09[0]) );
  SDFFQX1 c_buf_reg_8__1_ ( .D(N544), .SIN(dbg_08[0]), .SMC(test_se), .C(
        net11909), .Q(dbg_08[1]) );
  SDFFQX1 c_buf_reg_7__1_ ( .D(N536), .SIN(dbg_07[0]), .SMC(test_se), .C(
        net11914), .Q(dbg_07[1]) );
  SDFFQX1 c_buf_reg_6__4_ ( .D(N531), .SIN(dbg_06[3]), .SMC(test_se), .C(
        net11919), .Q(dbg_06[4]) );
  SDFFQX1 c_buf_reg_6__1_ ( .D(N528), .SIN(dbg_06[0]), .SMC(test_se), .C(
        net11919), .Q(dbg_06[1]) );
  SDFFQX1 c_buf_reg_5__1_ ( .D(N520), .SIN(dbg_05[0]), .SMC(test_se), .C(
        net11924), .Q(dbg_05[1]) );
  SDFFQX1 c_buf_reg_4__1_ ( .D(N512), .SIN(dbg_04[0]), .SMC(test_se), .C(
        net11929), .Q(dbg_04[1]) );
  SDFFQX1 c_buf_reg_3__1_ ( .D(N504), .SIN(dbg_03[0]), .SMC(test_se), .C(
        net11934), .Q(dbg_03[1]) );
  SDFFQX1 c_buf_reg_2__1_ ( .D(N496), .SIN(dbg_02[0]), .SMC(test_se), .C(
        net11939), .Q(dbg_02[1]) );
  SDFFQX1 c_buf_reg_1__1_ ( .D(N488), .SIN(dbg_01[0]), .SMC(test_se), .C(
        net11944), .Q(dbg_01[1]) );
  SDFFQX1 c_buf_reg_6__0_ ( .D(N527), .SIN(dbg_05[7]), .SMC(test_se), .C(
        net11919), .Q(dbg_06[0]) );
  SDFFQX1 c_buf_reg_15__6_ ( .D(N605), .SIN(dbg_0f[5]), .SMC(test_se), .C(
        net11874), .Q(dbg_0f[6]) );
  SDFFQX1 c_buf_reg_15__3_ ( .D(N602), .SIN(dbg_0f[2]), .SMC(test_se), .C(
        net11874), .Q(dbg_0f[3]) );
  SDFFQX1 c_buf_reg_13__6_ ( .D(N589), .SIN(dbg_0d[5]), .SMC(test_se), .C(
        net11884), .Q(dbg_0d[6]) );
  SDFFQX1 c_buf_reg_13__3_ ( .D(N586), .SIN(dbg_0d[2]), .SMC(test_se), .C(
        net11884), .Q(dbg_0d[3]) );
  SDFFQX1 c_buf_reg_12__6_ ( .D(N581), .SIN(dbg_0c[5]), .SMC(test_se), .C(
        net11889), .Q(dbg_0c[6]) );
  SDFFQX1 c_buf_reg_12__3_ ( .D(N578), .SIN(dbg_0c[2]), .SMC(test_se), .C(
        net11889), .Q(dbg_0c[3]) );
  SDFFQX1 c_buf_reg_11__6_ ( .D(N573), .SIN(dbg_0b[5]), .SMC(test_se), .C(
        net11894), .Q(dbg_0b[6]) );
  SDFFQX1 c_buf_reg_11__5_ ( .D(N572), .SIN(dbg_0b[4]), .SMC(test_se), .C(
        net11894), .Q(dbg_0b[5]) );
  SDFFQX1 c_buf_reg_11__4_ ( .D(N571), .SIN(dbg_0b[3]), .SMC(test_se), .C(
        net11894), .Q(dbg_0b[4]) );
  SDFFQX1 c_buf_reg_11__3_ ( .D(N570), .SIN(dbg_0b[2]), .SMC(test_se), .C(
        net11894), .Q(dbg_0b[3]) );
  SDFFQX1 c_buf_reg_11__0_ ( .D(N567), .SIN(dbg_0a[7]), .SMC(test_se), .C(
        net11894), .Q(dbg_0b[0]) );
  SDFFQX1 c_buf_reg_10__6_ ( .D(N565), .SIN(dbg_0a[5]), .SMC(test_se), .C(
        net11899), .Q(dbg_0a[6]) );
  SDFFQX1 c_buf_reg_10__5_ ( .D(N564), .SIN(dbg_0a[4]), .SMC(test_se), .C(
        net11899), .Q(dbg_0a[5]) );
  SDFFQX1 c_buf_reg_10__4_ ( .D(N563), .SIN(dbg_0a[3]), .SMC(test_se), .C(
        net11899), .Q(dbg_0a[4]) );
  SDFFQX1 c_buf_reg_10__3_ ( .D(N562), .SIN(dbg_0a[2]), .SMC(test_se), .C(
        net11899), .Q(dbg_0a[3]) );
  SDFFQX1 c_buf_reg_10__0_ ( .D(N559), .SIN(dbg_09[7]), .SMC(test_se), .C(
        net11899), .Q(dbg_0a[0]) );
  SDFFQX1 c_buf_reg_9__6_ ( .D(N557), .SIN(dbg_09[5]), .SMC(test_se), .C(
        net11904), .Q(dbg_09[6]) );
  SDFFQX1 c_buf_reg_9__5_ ( .D(N556), .SIN(dbg_09[4]), .SMC(test_se), .C(
        net11904), .Q(dbg_09[5]) );
  SDFFQX1 c_buf_reg_9__3_ ( .D(N554), .SIN(dbg_09[2]), .SMC(test_se), .C(
        net11904), .Q(dbg_09[3]) );
  SDFFQX1 c_buf_reg_8__6_ ( .D(N549), .SIN(dbg_08[5]), .SMC(test_se), .C(
        net11909), .Q(dbg_08[6]) );
  SDFFQX1 c_buf_reg_8__5_ ( .D(N548), .SIN(dbg_08[4]), .SMC(test_se), .C(
        net11909), .Q(dbg_08[5]) );
  SDFFQX1 c_buf_reg_8__4_ ( .D(N547), .SIN(dbg_08[3]), .SMC(test_se), .C(
        net11909), .Q(dbg_08[4]) );
  SDFFQX1 c_buf_reg_8__3_ ( .D(N546), .SIN(dbg_08[2]), .SMC(test_se), .C(
        net11909), .Q(dbg_08[3]) );
  SDFFQX1 c_buf_reg_8__0_ ( .D(N543), .SIN(dbg_07[7]), .SMC(test_se), .C(
        net11909), .Q(dbg_08[0]) );
  SDFFQX1 c_buf_reg_7__6_ ( .D(N541), .SIN(dbg_07[5]), .SMC(test_se), .C(
        net11914), .Q(dbg_07[6]) );
  SDFFQX1 c_buf_reg_7__5_ ( .D(N540), .SIN(dbg_07[4]), .SMC(test_se), .C(
        net11914), .Q(dbg_07[5]) );
  SDFFQX1 c_buf_reg_7__4_ ( .D(N539), .SIN(dbg_07[3]), .SMC(test_se), .C(
        net11914), .Q(dbg_07[4]) );
  SDFFQX1 c_buf_reg_7__3_ ( .D(N538), .SIN(dbg_07[2]), .SMC(test_se), .C(
        net11914), .Q(dbg_07[3]) );
  SDFFQX1 c_buf_reg_7__0_ ( .D(N535), .SIN(dbg_06[7]), .SMC(test_se), .C(
        net11914), .Q(dbg_07[0]) );
  SDFFQX1 c_buf_reg_6__6_ ( .D(N533), .SIN(dbg_06[5]), .SMC(test_se), .C(
        net11919), .Q(dbg_06[6]) );
  SDFFQX1 c_buf_reg_5__6_ ( .D(N525), .SIN(dbg_05[5]), .SMC(test_se), .C(
        net11924), .Q(dbg_05[6]) );
  SDFFQX1 c_buf_reg_4__6_ ( .D(N517), .SIN(dbg_04[5]), .SMC(test_se), .C(
        net11929), .Q(dbg_04[6]) );
  SDFFQX1 c_buf_reg_3__6_ ( .D(N509), .SIN(dbg_03[5]), .SMC(test_se), .C(
        net11934), .Q(dbg_03[6]) );
  SDFFQX1 c_buf_reg_2__6_ ( .D(N501), .SIN(dbg_02[5]), .SMC(test_se), .C(
        net11939), .Q(dbg_02[6]) );
  SDFFQX1 c_buf_reg_1__6_ ( .D(N493), .SIN(dbg_01[5]), .SMC(test_se), .C(
        net11944), .Q(dbg_01[6]) );
  SDFFQX1 c_buf_reg_6__5_ ( .D(N532), .SIN(dbg_06[4]), .SMC(test_se), .C(
        net11919), .Q(dbg_06[5]) );
  SDFFQX1 c_buf_reg_5__5_ ( .D(N524), .SIN(dbg_05[4]), .SMC(test_se), .C(
        net11924), .Q(dbg_05[5]) );
  SDFFQX1 c_buf_reg_4__5_ ( .D(N516), .SIN(dbg_04[4]), .SMC(test_se), .C(
        net11929), .Q(dbg_04[5]) );
  SDFFQX1 c_buf_reg_3__5_ ( .D(N508), .SIN(dbg_03[4]), .SMC(test_se), .C(
        net11934), .Q(dbg_03[5]) );
  SDFFQX1 c_buf_reg_2__5_ ( .D(N500), .SIN(dbg_02[4]), .SMC(test_se), .C(
        net11939), .Q(dbg_02[5]) );
  SDFFQX1 c_buf_reg_1__5_ ( .D(N492), .SIN(dbg_01[4]), .SMC(test_se), .C(
        net11944), .Q(dbg_01[5]) );
  SDFFQX1 c_buf_reg_5__4_ ( .D(N523), .SIN(dbg_05[3]), .SMC(test_se), .C(
        net11924), .Q(dbg_05[4]) );
  SDFFQX1 c_buf_reg_4__4_ ( .D(N515), .SIN(dbg_04[3]), .SMC(test_se), .C(
        net11929), .Q(dbg_04[4]) );
  SDFFQX1 c_buf_reg_3__4_ ( .D(N507), .SIN(dbg_03[3]), .SMC(test_se), .C(
        net11934), .Q(dbg_03[4]) );
  SDFFQX1 c_buf_reg_2__4_ ( .D(N499), .SIN(dbg_02[3]), .SMC(test_se), .C(
        net11939), .Q(dbg_02[4]) );
  SDFFQX1 c_buf_reg_1__4_ ( .D(N491), .SIN(dbg_01[3]), .SMC(test_se), .C(
        net11944), .Q(dbg_01[4]) );
  SDFFQX1 c_buf_reg_6__3_ ( .D(N530), .SIN(dbg_06[2]), .SMC(test_se), .C(
        net11919), .Q(dbg_06[3]) );
  SDFFQX1 c_buf_reg_5__3_ ( .D(N522), .SIN(dbg_05[2]), .SMC(test_se), .C(
        net11924), .Q(dbg_05[3]) );
  SDFFQX1 c_buf_reg_4__3_ ( .D(N514), .SIN(dbg_04[2]), .SMC(test_se), .C(
        net11929), .Q(dbg_04[3]) );
  SDFFQX1 c_buf_reg_3__3_ ( .D(N506), .SIN(dbg_03[2]), .SMC(test_se), .C(
        net11934), .Q(dbg_03[3]) );
  SDFFQX1 c_buf_reg_2__3_ ( .D(N498), .SIN(dbg_02[2]), .SMC(test_se), .C(
        net11939), .Q(dbg_02[3]) );
  SDFFQX1 c_buf_reg_1__3_ ( .D(N490), .SIN(dbg_01[2]), .SMC(test_se), .C(
        net11944), .Q(dbg_01[3]) );
  SDFFQX1 c_buf_reg_5__0_ ( .D(N519), .SIN(dbg_04[7]), .SMC(test_se), .C(
        net11924), .Q(dbg_05[0]) );
  SDFFQX1 c_buf_reg_4__0_ ( .D(N511), .SIN(dbg_03[7]), .SMC(test_se), .C(
        net11929), .Q(dbg_04[0]) );
  SDFFQX1 c_buf_reg_3__0_ ( .D(N503), .SIN(dbg_02[7]), .SMC(test_se), .C(
        net11934), .Q(dbg_03[0]) );
  SDFFQX1 c_buf_reg_2__0_ ( .D(N495), .SIN(dbg_01[7]), .SMC(test_se), .C(
        net11939), .Q(dbg_02[0]) );
  SDFFQX1 c_buf_reg_1__0_ ( .D(N487), .SIN(rd_buf[7]), .SMC(test_se), .C(
        net11944), .Q(dbg_01[0]) );
  SDFFQX1 c_buf_reg_22__7_ ( .D(N662), .SIN(c_buf_22__6_), .SMC(test_se), .C(
        net11839), .Q(c_buf_22__7_) );
  SDFFQX1 c_buf_reg_21__7_ ( .D(N654), .SIN(c_buf_21__6_), .SMC(test_se), .C(
        net11844), .Q(c_buf_21__7_) );
  SDFFQX1 c_buf_reg_20__7_ ( .D(N646), .SIN(c_buf_20__6_), .SMC(test_se), .C(
        net11849), .Q(c_buf_20__7_) );
  SDFFQX1 c_buf_reg_19__7_ ( .D(N638), .SIN(c_buf_19__6_), .SMC(test_se), .C(
        net11854), .Q(c_buf_19__7_) );
  SDFFQX1 c_buf_reg_18__7_ ( .D(N630), .SIN(c_buf_18__6_), .SMC(test_se), .C(
        net11859), .Q(c_buf_18__7_) );
  SDFFQX1 c_buf_reg_17__7_ ( .D(N622), .SIN(c_buf_17__6_), .SMC(test_se), .C(
        net11864), .Q(c_buf_17__7_) );
  SDFFQX1 c_buf_reg_16__7_ ( .D(N614), .SIN(c_buf_16__6_), .SMC(test_se), .C(
        net11869), .Q(c_buf_16__7_) );
  SDFFQX1 c_buf_reg_15__7_ ( .D(N606), .SIN(dbg_0f[6]), .SMC(test_se), .C(
        net11874), .Q(dbg_0f[7]) );
  SDFFQX1 c_buf_reg_14__7_ ( .D(N598), .SIN(dbg_0e[6]), .SMC(test_se), .C(
        net11879), .Q(dbg_0e[7]) );
  SDFFQX1 c_buf_reg_13__7_ ( .D(N590), .SIN(dbg_0d[6]), .SMC(test_se), .C(
        net11884), .Q(dbg_0d[7]) );
  SDFFQX1 c_buf_reg_12__7_ ( .D(N582), .SIN(dbg_0c[6]), .SMC(test_se), .C(
        net11889), .Q(dbg_0c[7]) );
  SDFFQX1 c_buf_reg_11__7_ ( .D(N574), .SIN(dbg_0b[6]), .SMC(test_se), .C(
        net11894), .Q(dbg_0b[7]) );
  SDFFQX1 c_buf_reg_9__7_ ( .D(N558), .SIN(dbg_09[6]), .SMC(test_se), .C(
        net11904), .Q(dbg_09[7]) );
  SDFFQX1 c_buf_reg_8__7_ ( .D(N550), .SIN(dbg_08[6]), .SMC(test_se), .C(
        net11909), .Q(dbg_08[7]) );
  SDFFQX1 c_buf_reg_7__7_ ( .D(N542), .SIN(dbg_07[6]), .SMC(test_se), .C(
        net11914), .Q(dbg_07[7]) );
  SDFFQX1 c_buf_reg_6__7_ ( .D(N534), .SIN(dbg_06[6]), .SMC(test_se), .C(
        net11919), .Q(dbg_06[7]) );
  SDFFQX1 c_buf_reg_5__7_ ( .D(N526), .SIN(dbg_05[6]), .SMC(test_se), .C(
        net11924), .Q(dbg_05[7]) );
  SDFFQX1 c_buf_reg_4__7_ ( .D(N518), .SIN(dbg_04[6]), .SMC(test_se), .C(
        net11929), .Q(dbg_04[7]) );
  SDFFQX1 c_buf_reg_3__7_ ( .D(N510), .SIN(dbg_03[6]), .SMC(test_se), .C(
        net11934), .Q(dbg_03[7]) );
  SDFFQX1 c_buf_reg_2__7_ ( .D(N502), .SIN(dbg_02[6]), .SMC(test_se), .C(
        net11939), .Q(dbg_02[7]) );
  SDFFQX1 c_buf_reg_1__7_ ( .D(N494), .SIN(dbg_01[6]), .SMC(test_se), .C(
        net11944), .Q(dbg_01[7]) );
  SDFFQX1 c_buf_reg_23__3_ ( .D(N789), .SIN(wr_buf[2]), .SMC(test_se), .C(
        net11834), .Q(wr_buf[3]) );
  SDFFQX1 c_buf_reg_23__7_ ( .D(N793), .SIN(wr_buf[6]), .SMC(test_se), .C(
        net11834), .Q(wr_buf[7]) );
  SDFFQX1 c_buf_reg_23__6_ ( .D(N792), .SIN(wr_buf[5]), .SMC(test_se), .C(
        net11834), .Q(wr_buf[6]) );
  SDFFQX1 c_buf_reg_23__5_ ( .D(N791), .SIN(wr_buf[4]), .SMC(test_se), .C(
        net11834), .Q(wr_buf[5]) );
  SDFFQX1 c_buf_reg_10__7_ ( .D(N566), .SIN(dbg_0a[6]), .SMC(test_se), .C(
        net11899), .Q(dbg_0a[7]) );
  SDFFQX1 c_adr_reg_4_ ( .D(N830), .SIN(c_adr[3]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[4]) );
  SDFFQX1 c_adr_reg_2_ ( .D(N828), .SIN(c_adr[1]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[2]) );
  SDFFQX1 c_adr_reg_3_ ( .D(N829), .SIN(c_adr[2]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[3]) );
  SDFFQX2 adr_p_reg_6_ ( .D(N860), .SIN(pmem_a[5]), .SMC(test_se), .C(net11829), .Q(pmem_a[9]) );
  SDFFQX2 adr_p_reg_8_ ( .D(N862), .SIN(pmem_a[10]), .SMC(test_se), .C(
        net11829), .Q(pmem_a[11]) );
  SDFFQX2 adr_p_reg_0_ ( .D(N854), .SIN(pmem_a[8]), .SMC(test_se), .C(net11829), .Q(pmem_a[0]) );
  SDFFQX2 a_bit_reg_1_ ( .D(n939), .SIN(pmem_a[6]), .SMC(test_se), .C(net11824), .Q(pmem_a[7]) );
  SDFFQX1 c_adr_reg_1_ ( .D(N827), .SIN(c_adr[0]), .SMC(test_se), .C(net11959), 
        .Q(c_adr[1]) );
  SDFFQX1 c_adr_reg_0_ ( .D(N826), .SIN(adr_p[14]), .SMC(test_se), .C(net11959), .Q(c_adr[0]) );
  AND2X1 U3 ( .A(c_adr[1]), .B(n477), .Y(n476) );
  INVX1 U4 ( .A(memaddr[1]), .Y(n477) );
  AND2X1 U5 ( .A(memaddr[2]), .B(n876), .Y(n39) );
  NAND5XL U6 ( .A(n537), .B(n536), .C(n535), .D(n534), .E(n533), .Y(o_inst[0])
         );
  NAND5XL U7 ( .A(n629), .B(n628), .C(n627), .D(n626), .E(n624), .Y(o_inst[2])
         );
  NAND5XL U8 ( .A(n810), .B(n809), .C(n808), .D(n807), .E(n806), .Y(o_inst[6])
         );
  OA222X1 U9 ( .A(n834), .B(n791), .C(n832), .D(n790), .E(n830), .F(n789), .Y(
        n807) );
  OA222X1 U10 ( .A(n822), .B(n785), .C(n820), .D(n784), .E(n818), .F(n783), 
        .Y(n809) );
  OA222X1 U11 ( .A(n816), .B(n782), .C(n814), .D(n781), .E(n812), .F(n780), 
        .Y(n810) );
  INVX1 U12 ( .A(n507), .Y(n512) );
  NOR3XL U13 ( .A(n509), .B(n508), .C(n516), .Y(n41) );
  NOR2X1 U14 ( .A(n517), .B(n30), .Y(n29) );
  XOR3X1 U15 ( .A(c_adr[3]), .B(memaddr[3]), .C(n497), .Y(n516) );
  NAND21X1 U16 ( .B(n518), .A(n29), .Y(n849) );
  NAND5XL U17 ( .A(n583), .B(n582), .C(n581), .D(n580), .E(n574), .Y(o_inst[1]) );
  NAND5XL U18 ( .A(n704), .B(n703), .C(n702), .D(n701), .E(n700), .Y(o_inst[4]) );
  NAND5XL U19 ( .A(n779), .B(n778), .C(n777), .D(n776), .E(n775), .Y(o_inst[5]) );
  NAND5XL U20 ( .A(n671), .B(n670), .C(n669), .D(n668), .E(n667), .Y(o_inst[3]) );
  AO21X1 U21 ( .B(n451), .C(n412), .A(n390), .Y(n647) );
  INVX1 U22 ( .A(c_adr[2]), .Y(n876) );
  INVXL U23 ( .A(n236), .Y(n1) );
  INVXL U24 ( .A(n1), .Y(n2) );
  OA21XL U25 ( .B(memaddr_c[4]), .C(n159), .A(n158), .Y(n165) );
  INVX1 U26 ( .A(n290), .Y(n3) );
  INVX1 U27 ( .A(n290), .Y(n4) );
  INVX1 U28 ( .A(n282), .Y(n5) );
  INVX1 U29 ( .A(n282), .Y(n6) );
  INVX1 U30 ( .A(n284), .Y(n7) );
  INVX1 U31 ( .A(n284), .Y(n8) );
  INVX1 U32 ( .A(n239), .Y(n9) );
  INVX1 U33 ( .A(n286), .Y(n10) );
  INVX1 U34 ( .A(n286), .Y(n11) );
  INVX1 U35 ( .A(n235), .Y(n12) );
  INVX1 U36 ( .A(n288), .Y(n13) );
  INVX1 U37 ( .A(n288), .Y(n14) );
  INVX1 U38 ( .A(n444), .Y(n15) );
  INVX1 U39 ( .A(n292), .Y(n16) );
  INVX1 U40 ( .A(n292), .Y(n17) );
  BUFX3 U41 ( .A(n242), .Y(n18) );
  AOI21XL U42 ( .B(memaddr_c[3]), .C(n242), .A(n89), .Y(n57) );
  INVX1 U43 ( .A(n237), .Y(n19) );
  INVX1 U44 ( .A(n294), .Y(n20) );
  INVX1 U45 ( .A(n294), .Y(n21) );
  INVX1 U46 ( .A(n317), .Y(n22) );
  INVX1 U47 ( .A(n228), .Y(n23) );
  INVX1 U48 ( .A(n906), .Y(n24) );
  INVX1 U49 ( .A(n280), .Y(n25) );
  INVX1 U50 ( .A(n280), .Y(n26) );
  INVX1 U51 ( .A(n368), .Y(n27) );
  INVX1 U52 ( .A(n368), .Y(n28) );
  OR2XL U53 ( .A(n492), .B(n522), .Y(n812) );
  INVX3 U54 ( .A(n489), .Y(n496) );
  NAND21X1 U55 ( .B(n517), .A(n508), .Y(n489) );
  NAND21X1 U56 ( .B(n522), .A(n496), .Y(n826) );
  NAND21X1 U57 ( .B(n490), .A(n491), .Y(n523) );
  INVX1 U58 ( .A(n516), .Y(n30) );
  INVXL U59 ( .A(memaddr[2]), .Y(n38) );
  NAND21XL U60 ( .B(n518), .A(n496), .Y(n828) );
  OR2XL U61 ( .A(n492), .B(n518), .Y(n820) );
  NAND2XL U62 ( .A(o_inst[4]), .B(o_inst[3]), .Y(n891) );
  INVXL U63 ( .A(o_inst[5]), .Y(n894) );
  INVXL U64 ( .A(o_inst[6]), .Y(n895) );
  NAND32XL U65 ( .B(n508), .C(n516), .A(n509), .Y(n507) );
  NAND21XL U66 ( .B(n509), .A(n508), .Y(n492) );
  NOR43XL U67 ( .B(n805), .C(n804), .D(n803), .A(n31), .Y(n806) );
  OAI222XL U68 ( .A(n857), .B(n802), .C(n855), .D(n801), .E(n853), .F(n800), 
        .Y(n31) );
  NOR43XL U69 ( .B(n774), .C(n773), .D(n772), .A(n32), .Y(n775) );
  OAI222XL U70 ( .A(n857), .B(n771), .C(n855), .D(n770), .E(n853), .F(n769), 
        .Y(n32) );
  NOR43XL U71 ( .B(n666), .C(n665), .D(n664), .A(n33), .Y(n667) );
  OAI222XL U72 ( .A(n857), .B(n663), .C(n855), .D(n662), .E(n853), .F(n661), 
        .Y(n33) );
  NOR43XL U73 ( .B(n699), .C(n698), .D(n697), .A(n34), .Y(n700) );
  OAI222XL U74 ( .A(n857), .B(n696), .C(n855), .D(n695), .E(n853), .F(n694), 
        .Y(n34) );
  NOR43XL U75 ( .B(n573), .C(n572), .D(n571), .A(n35), .Y(n574) );
  OAI222XL U76 ( .A(n857), .B(n570), .C(n855), .D(n569), .E(n853), .F(n568), 
        .Y(n35) );
  NOR43XL U77 ( .B(n531), .C(n530), .D(n528), .A(n36), .Y(n533) );
  OAI222XL U78 ( .A(n857), .B(n527), .C(n855), .D(n526), .E(n853), .F(n525), 
        .Y(n36) );
  NAND21XL U79 ( .B(n484), .A(n490), .Y(n524) );
  NOR43XL U80 ( .B(n623), .C(n622), .D(n620), .A(n37), .Y(n624) );
  OAI222XL U81 ( .A(n857), .B(n619), .C(n855), .D(n618), .E(n853), .F(n617), 
        .Y(n37) );
  OAI221XL U82 ( .A(n880), .B(n140), .C(n877), .D(n371), .E(n130), .Y(n144) );
  OAI22XL U83 ( .A(c_adr[1]), .B(n477), .C(n483), .D(n476), .Y(n478) );
  NAND21X1 U84 ( .B(memaddr[0]), .A(c_adr[0]), .Y(n482) );
  OAI22CX1 U85 ( .C(n39), .D(n478), .A(n38), .B(c_adr[2]), .Y(n497) );
  XOR3XL U86 ( .A(c_adr[2]), .B(memaddr[2]), .C(n478), .Y(n509) );
  OAI21BBX1 U87 ( .A(n90), .B(n319), .C(n376), .Y(N823) );
  OAI21BBX1 U88 ( .A(n90), .B(n320), .C(n440), .Y(N821) );
  NAND21XL U89 ( .B(n877), .A(c_ptr[0]), .Y(n140) );
  OAI221XL U90 ( .A(n274), .B(n341), .C(memdatao[1]), .D(n277), .E(n273), .Y(
        N787) );
  OAI221XL U91 ( .A(n271), .B(n341), .C(memdatao[2]), .D(n277), .E(n270), .Y(
        N788) );
  NAND21XL U92 ( .B(c_adr[3]), .A(n353), .Y(n147) );
  NAND21XL U93 ( .B(n872), .A(c_ptr[3]), .Y(n117) );
  NAND21XL U94 ( .B(c_adr[4]), .A(n355), .Y(n137) );
  INVXL U95 ( .A(c_adr[4]), .Y(n883) );
  INVX1 U96 ( .A(n368), .Y(n365) );
  INVX1 U97 ( .A(n372), .Y(n343) );
  INVX1 U98 ( .A(n345), .Y(n354) );
  INVX1 U99 ( .A(n416), .Y(n920) );
  INVX1 U100 ( .A(n231), .Y(n229) );
  AOI21X1 U101 ( .B(n430), .C(we_twlb), .A(N853), .Y(n40) );
  NAND21X1 U102 ( .B(n244), .A(n368), .Y(n236) );
  NAND21X1 U103 ( .B(n345), .A(n69), .Y(n368) );
  INVX1 U104 ( .A(n202), .Y(n182) );
  NAND21X1 U105 ( .B(n304), .A(n336), .Y(n372) );
  INVX1 U106 ( .A(n308), .Y(n86) );
  INVX1 U107 ( .A(n87), .Y(n85) );
  INVX1 U108 ( .A(n87), .Y(n84) );
  INVX1 U109 ( .A(n87), .Y(n83) );
  INVX1 U110 ( .A(n87), .Y(n82) );
  INVX1 U111 ( .A(n87), .Y(n81) );
  INVX1 U112 ( .A(n87), .Y(n80) );
  INVX1 U113 ( .A(n308), .Y(n79) );
  INVX1 U114 ( .A(n308), .Y(n78) );
  INVX1 U115 ( .A(n308), .Y(n77) );
  INVX1 U116 ( .A(n308), .Y(n76) );
  INVX1 U117 ( .A(n308), .Y(n75) );
  INVX1 U118 ( .A(n308), .Y(n74) );
  INVX1 U119 ( .A(n308), .Y(n73) );
  INVX1 U120 ( .A(n87), .Y(n72) );
  INVX1 U121 ( .A(n87), .Y(n70) );
  INVX1 U122 ( .A(n87), .Y(n71) );
  INVX1 U123 ( .A(n324), .Y(n451) );
  NAND21X1 U124 ( .B(n88), .A(n444), .Y(n345) );
  NAND21X1 U125 ( .B(n433), .A(n451), .Y(n376) );
  INVX1 U126 ( .A(n412), .Y(n387) );
  INVX1 U127 ( .A(n419), .Y(n327) );
  NOR2X1 U128 ( .A(dw_rst), .B(n91), .Y(n416) );
  INVX1 U129 ( .A(n155), .Y(n159) );
  INVX1 U130 ( .A(n156), .Y(n150) );
  INVX1 U131 ( .A(n92), .Y(n91) );
  NAND21X1 U132 ( .B(n524), .A(n41), .Y(n851) );
  NAND21X1 U133 ( .B(n523), .A(n512), .Y(n845) );
  NAND21X1 U134 ( .B(n522), .A(n512), .Y(n843) );
  NAND21X1 U135 ( .B(n518), .A(n41), .Y(n838) );
  NAND21X1 U136 ( .B(n524), .A(n512), .Y(n841) );
  NAND21X1 U137 ( .B(n522), .A(n41), .Y(n836) );
  NAND21X1 U138 ( .B(n523), .A(n41), .Y(n847) );
  NAND21X1 U139 ( .B(n518), .A(n512), .Y(n839) );
  NAND21X1 U140 ( .B(n491), .A(n490), .Y(n518) );
  NAND21X1 U141 ( .B(n523), .A(n496), .Y(n822) );
  NAND21X1 U142 ( .B(n522), .A(n503), .Y(n834) );
  NAND21X1 U143 ( .B(n522), .A(n29), .Y(n857) );
  OR2X1 U144 ( .A(n492), .B(n524), .Y(n816) );
  NAND21X1 U145 ( .B(n524), .A(n503), .Y(n832) );
  NAND21X1 U146 ( .B(n523), .A(n29), .Y(n855) );
  OR2X1 U147 ( .A(n492), .B(n523), .Y(n814) );
  NAND21X1 U148 ( .B(n524), .A(n496), .Y(n818) );
  NAND21X1 U149 ( .B(n524), .A(n29), .Y(n853) );
  NAND21X1 U150 ( .B(n518), .A(n503), .Y(n830) );
  NAND21X1 U151 ( .B(n523), .A(n503), .Y(n824) );
  INVX1 U152 ( .A(n90), .Y(n88) );
  NAND32X1 U153 ( .B(n225), .C(n388), .A(n342), .Y(n231) );
  NAND32X1 U154 ( .B(n374), .C(n373), .A(n372), .Y(N853) );
  INVX1 U155 ( .A(n438), .Y(n304) );
  NAND5XL U156 ( .A(n218), .B(n217), .C(n216), .D(n215), .E(n214), .Y(n342) );
  INVX1 U157 ( .A(n201), .Y(n216) );
  AND4X1 U158 ( .A(n45), .B(n204), .C(n203), .D(n202), .Y(n215) );
  AND4X1 U159 ( .A(n213), .B(n212), .C(n211), .D(n210), .Y(n214) );
  INVX1 U160 ( .A(n228), .Y(n374) );
  NAND21X1 U161 ( .B(n341), .A(n69), .Y(n228) );
  AND4X1 U162 ( .A(n209), .B(n208), .C(n207), .D(n206), .Y(n210) );
  INVX1 U163 ( .A(n87), .Y(n69) );
  INVX1 U164 ( .A(n303), .Y(n87) );
  INVX1 U165 ( .A(n221), .Y(n244) );
  NAND21X1 U166 ( .B(n910), .A(n181), .Y(n202) );
  NAND21X1 U167 ( .B(n911), .A(n178), .Y(n204) );
  AO21X1 U168 ( .B(n349), .C(n359), .A(n365), .Y(N881) );
  AO21X1 U169 ( .B(n351), .C(n359), .A(n27), .Y(N885) );
  AO21X1 U170 ( .B(n343), .C(n342), .A(n373), .Y(n93) );
  INVX1 U171 ( .A(n370), .Y(n366) );
  INVX1 U172 ( .A(n212), .Y(n169) );
  AO21X1 U173 ( .B(n60), .C(n359), .A(n28), .Y(N889) );
  OAI211X1 U174 ( .C(n420), .D(n388), .A(n385), .B(n467), .Y(n332) );
  INVX1 U175 ( .A(n388), .Y(n389) );
  NAND32X1 U176 ( .B(n325), .C(n324), .A(n426), .Y(n419) );
  NAND2X1 U177 ( .A(n426), .B(n430), .Y(n339) );
  NAND42X1 U178 ( .C(n336), .D(n335), .A(n334), .B(n333), .Y(N820) );
  AOI21BBXL U179 ( .B(n947), .C(n379), .A(n546), .Y(n333) );
  INVX1 U180 ( .A(n339), .Y(n335) );
  NOR43XL U181 ( .B(n898), .C(n387), .D(n15), .A(n332), .Y(n334) );
  INVX1 U182 ( .A(n325), .Y(n433) );
  INVX1 U183 ( .A(n448), .Y(n430) );
  NAND21X1 U184 ( .B(n88), .A(n247), .Y(n324) );
  AO21X1 U185 ( .B(n247), .C(n325), .A(n447), .Y(n412) );
  INVX1 U186 ( .A(n213), .Y(n122) );
  NAND21X1 U187 ( .B(o_ofs_inc), .A(n90), .Y(n447) );
  AO21X1 U188 ( .B(n898), .C(n947), .A(n88), .Y(n326) );
  INVX1 U189 ( .A(n239), .Y(n233) );
  INVX1 U190 ( .A(n235), .Y(n234) );
  INVX1 U191 ( .A(n947), .Y(n896) );
  INVX1 U192 ( .A(n90), .Y(n89) );
  INVX1 U193 ( .A(n413), .Y(n436) );
  NAND21X1 U194 ( .B(n426), .A(n451), .Y(n413) );
  INVX1 U195 ( .A(n375), .Y(n454) );
  INVX1 U196 ( .A(srst), .Y(n92) );
  XOR2X1 U197 ( .A(n139), .B(n62), .Y(n155) );
  XNOR2XL U198 ( .A(n693), .B(n144), .Y(n146) );
  XNOR2XL U199 ( .A(n682), .B(n149), .Y(n156) );
  INVX1 U200 ( .A(n868), .Y(n936) );
  INVX1 U201 ( .A(n135), .Y(n172) );
  INVX1 U202 ( .A(n935), .Y(n746) );
  INVX1 U203 ( .A(n180), .Y(n133) );
  NOR43XL U204 ( .B(o_inst[1]), .C(o_inst[0]), .D(o_inst[2]), .A(n891), .Y(
        n893) );
  INVX1 U205 ( .A(n871), .Y(n718) );
  INVX1 U206 ( .A(n141), .Y(n107) );
  INVX1 U207 ( .A(n224), .Y(n321) );
  INVX1 U208 ( .A(n341), .Y(n444) );
  NOR2X1 U209 ( .A(n918), .B(n91), .Y(n923) );
  INVX1 U210 ( .A(n232), .Y(n336) );
  INVX1 U211 ( .A(n249), .Y(o_ofs_inc) );
  INVX1 U212 ( .A(n317), .Y(n898) );
  NOR2X1 U213 ( .A(n909), .B(n22), .Y(n575) );
  INVX1 U214 ( .A(n420), .Y(n445) );
  OA222X1 U215 ( .A(n834), .B(n759), .C(n832), .D(n749), .E(n830), .F(n748), 
        .Y(n776) );
  OA222X1 U216 ( .A(n822), .B(n713), .C(n820), .D(n712), .E(n818), .F(n708), 
        .Y(n778) );
  OA222X1 U217 ( .A(n816), .B(n707), .C(n814), .D(n706), .E(n812), .F(n705), 
        .Y(n779) );
  AND4X1 U218 ( .A(n861), .B(n860), .C(n859), .D(n858), .Y(n862) );
  OA222X1 U219 ( .A(n857), .B(n856), .C(n855), .D(n854), .E(n853), .F(n852), 
        .Y(n858) );
  OA222X1 U220 ( .A(n950), .B(n839), .C(n838), .D(n837), .E(n836), .F(n835), 
        .Y(n861) );
  OA222X1 U221 ( .A(n845), .B(n844), .C(n843), .D(n842), .E(n841), .F(n840), 
        .Y(n860) );
  OA222X1 U222 ( .A(n942), .B(n839), .C(n838), .D(n793), .E(n836), .F(n792), 
        .Y(n805) );
  OA222X1 U223 ( .A(n845), .B(n796), .C(n843), .D(n795), .E(n841), .F(n794), 
        .Y(n804) );
  OA222X1 U224 ( .A(n943), .B(n839), .C(n838), .D(n761), .E(n836), .F(n760), 
        .Y(n774) );
  OA222X1 U225 ( .A(n845), .B(n765), .C(n843), .D(n764), .E(n841), .F(n763), 
        .Y(n773) );
  NAND5X1 U226 ( .A(n866), .B(n865), .C(n864), .D(n863), .E(n862), .Y(
        o_inst[7]) );
  OA222X1 U227 ( .A(n834), .B(n833), .C(n832), .D(n831), .E(n830), .F(n829), 
        .Y(n863) );
  OA222X1 U228 ( .A(n822), .B(n821), .C(n820), .D(n819), .E(n818), .F(n817), 
        .Y(n865) );
  OA222X1 U229 ( .A(n816), .B(n815), .C(n814), .D(n813), .E(n812), .F(n811), 
        .Y(n866) );
  INVX1 U230 ( .A(n482), .Y(n483) );
  NAND21X1 U231 ( .B(n491), .A(n485), .Y(n522) );
  INVX1 U232 ( .A(n498), .Y(n503) );
  NAND21X1 U233 ( .B(n509), .A(n516), .Y(n498) );
  OA222X1 U234 ( .A(n834), .B(n652), .C(n832), .D(n640), .E(n830), .F(n639), 
        .Y(n668) );
  OA222X1 U235 ( .A(n822), .B(n635), .C(n820), .D(n634), .E(n818), .F(n633), 
        .Y(n670) );
  OA222X1 U236 ( .A(n816), .B(n632), .C(n814), .D(n631), .E(n812), .F(n630), 
        .Y(n671) );
  OA222X1 U237 ( .A(n834), .B(n684), .C(n832), .D(n683), .E(n830), .F(n681), 
        .Y(n701) );
  OA222X1 U238 ( .A(n822), .B(n677), .C(n820), .D(n676), .E(n818), .F(n675), 
        .Y(n703) );
  OA222X1 U239 ( .A(n816), .B(n674), .C(n814), .D(n673), .E(n812), .F(n672), 
        .Y(n704) );
  INVX1 U240 ( .A(n484), .Y(n491) );
  OA222X1 U241 ( .A(n944), .B(n839), .C(n838), .D(n654), .E(n836), .F(n653), 
        .Y(n666) );
  OA222X1 U242 ( .A(n845), .B(n657), .C(n843), .D(n656), .E(n841), .F(n655), 
        .Y(n665) );
  OA222X1 U243 ( .A(n945), .B(n839), .C(n838), .D(n686), .E(n836), .F(n685), 
        .Y(n699) );
  OA222X1 U244 ( .A(n845), .B(n689), .C(n843), .D(n688), .E(n841), .F(n687), 
        .Y(n698) );
  OA222X1 U245 ( .A(n941), .B(n839), .C(n838), .D(n561), .E(n836), .F(n560), 
        .Y(n573) );
  OA222X1 U246 ( .A(n845), .B(n564), .C(n843), .D(n563), .E(n841), .F(n562), 
        .Y(n572) );
  OA222X1 U247 ( .A(n946), .B(n839), .C(n838), .D(n511), .E(n836), .F(n510), 
        .Y(n531) );
  OA222X1 U248 ( .A(n845), .B(n515), .C(n843), .D(n514), .E(n841), .F(n513), 
        .Y(n530) );
  OA222X1 U249 ( .A(n940), .B(n839), .C(n838), .D(n601), .E(n836), .F(n600), 
        .Y(n623) );
  OA222X1 U250 ( .A(n845), .B(n612), .C(n843), .D(n604), .E(n841), .F(n602), 
        .Y(n622) );
  INVX1 U251 ( .A(n485), .Y(n490) );
  OA222X1 U252 ( .A(n834), .B(n559), .C(n832), .D(n552), .E(n830), .F(n551), 
        .Y(n580) );
  OA222X1 U253 ( .A(n822), .B(n544), .C(n820), .D(n542), .E(n818), .F(n541), 
        .Y(n582) );
  OA222X1 U254 ( .A(n816), .B(n540), .C(n814), .D(n539), .E(n812), .F(n538), 
        .Y(n583) );
  OA222X1 U255 ( .A(n834), .B(n506), .C(n832), .D(n505), .E(n830), .F(n504), 
        .Y(n534) );
  OA222X1 U256 ( .A(n822), .B(n495), .C(n820), .D(n494), .E(n818), .F(n493), 
        .Y(n536) );
  OA222X1 U257 ( .A(n816), .B(n488), .C(n814), .D(n487), .E(n812), .F(n486), 
        .Y(n537) );
  OA222X1 U258 ( .A(n834), .B(n599), .C(n832), .D(n598), .E(n830), .F(n597), 
        .Y(n626) );
  OA222X1 U259 ( .A(n822), .B(n592), .C(n820), .D(n588), .E(n818), .F(n587), 
        .Y(n628) );
  OA222X1 U260 ( .A(n816), .B(n586), .C(n814), .D(n585), .E(n812), .F(n584), 
        .Y(n629) );
  INVX1 U261 ( .A(n509), .Y(n517) );
  INVX1 U262 ( .A(n462), .Y(n90) );
  NAND32X1 U263 ( .B(n312), .C(n223), .A(n316), .Y(n249) );
  NAND2X1 U264 ( .A(n42), .B(n873), .Y(n878) );
  OAI22XL U265 ( .A(memaddr_c[2]), .B(n876), .C(memaddr_c[3]), .D(n872), .Y(
        n42) );
  NAND21X1 U266 ( .B(n304), .A(n908), .Y(n388) );
  AND2X1 U267 ( .A(n337), .B(n90), .Y(n43) );
  INVX1 U268 ( .A(n873), .Y(n875) );
  OAI32XL U269 ( .A(n884), .B(memaddr_c[4]), .C(n883), .D(n882), .E(n881), .Y(
        n885) );
  AND2XL U270 ( .A(memaddr_c[4]), .B(n883), .Y(n874) );
  OAI211X1 U271 ( .C(n200), .D(n199), .A(n198), .B(n197), .Y(n438) );
  AND2X1 U272 ( .A(n188), .B(n417), .Y(n199) );
  INVX1 U273 ( .A(n207), .Y(n200) );
  AOI32X1 U274 ( .A(n355), .B(n353), .C(n219), .D(n196), .E(n870), .Y(n197) );
  OAI211X1 U275 ( .C(n341), .D(n340), .A(n339), .B(n338), .Y(n373) );
  AND2X1 U276 ( .A(n43), .B(n421), .Y(n338) );
  INVX1 U277 ( .A(memaddr_c[7]), .Y(n914) );
  NAND21X1 U278 ( .B(n914), .A(n166), .Y(n218) );
  OR2X1 U279 ( .A(n345), .B(n340), .Y(n221) );
  NAND32X1 U280 ( .B(n342), .C(n452), .A(n316), .Y(n441) );
  OA222X1 U281 ( .A(memaddr_c[11]), .B(n178), .C(n177), .D(n176), .E(
        memaddr_c[10]), .F(n175), .Y(n184) );
  NAND21X1 U282 ( .B(n174), .A(n217), .Y(n176) );
  OA222X1 U283 ( .A(memaddr_c[9]), .B(n171), .C(n170), .D(n169), .E(
        memaddr_c[8]), .F(n168), .Y(n177) );
  INVX1 U284 ( .A(n203), .Y(n174) );
  EORX1 U285 ( .A(n218), .B(n44), .C(memaddr_c[7]), .D(n166), .Y(n170) );
  OAI22XL U286 ( .A(n165), .B(n201), .C(memaddr_c[6]), .D(n164), .Y(n44) );
  OAI211X1 U287 ( .C(n188), .D(n417), .A(n187), .B(n206), .Y(n207) );
  AO21X1 U288 ( .B(n68), .C(n186), .A(n185), .Y(n187) );
  OAI32X1 U289 ( .A(n184), .B(n183), .C(n182), .D(memaddr_c[12]), .E(n181), 
        .Y(n185) );
  INVX1 U290 ( .A(n204), .Y(n183) );
  INVX1 U291 ( .A(n120), .Y(n153) );
  INVX1 U292 ( .A(memaddr_c[11]), .Y(n911) );
  NAND2X1 U293 ( .A(memaddr_c[7]), .B(n934), .Y(n615) );
  INVX1 U294 ( .A(n308), .Y(n303) );
  INVX1 U295 ( .A(n621), .Y(n884) );
  NOR3XL U296 ( .A(n901), .B(memaddr_c[10]), .C(n607), .Y(n606) );
  AOI32X1 U297 ( .A(n157), .B(n208), .C(n209), .D(n162), .E(n163), .Y(n158) );
  GEN2XL U298 ( .D(n61), .E(n154), .C(n153), .B(n45), .A(n152), .Y(n157) );
  INVX1 U299 ( .A(n146), .Y(n151) );
  INVX1 U300 ( .A(n227), .Y(n322) );
  OAI211X1 U301 ( .C(n226), .D(n225), .A(n321), .B(n908), .Y(n227) );
  INVX1 U302 ( .A(n441), .Y(n226) );
  INVXL U303 ( .A(memaddr_c[1]), .Y(n154) );
  OA22X1 U304 ( .A(n146), .B(n145), .C(n61), .D(n154), .Y(n45) );
  NAND2X1 U305 ( .A(n175), .B(memaddr_c[10]), .Y(n217) );
  INVX1 U306 ( .A(memaddr_c[8]), .Y(n913) );
  INVX1 U307 ( .A(memaddr_c[9]), .Y(n912) );
  NAND21X1 U308 ( .B(n336), .A(n337), .Y(n242) );
  NAND21X1 U309 ( .B(n913), .A(n168), .Y(n212) );
  NAND21X1 U310 ( .B(n362), .A(n361), .Y(n370) );
  OAI22AX1 U311 ( .D(n164), .C(n887), .A(n163), .B(n162), .Y(n201) );
  OAI21BBX1 U312 ( .A(N441), .B(n23), .C(n46), .Y(N836) );
  AOI21X1 U313 ( .B(memaddr_c[10]), .C(n242), .A(n462), .Y(n46) );
  OAI21BBX1 U314 ( .A(N439), .B(n374), .C(n47), .Y(N834) );
  AOI21X1 U315 ( .B(n18), .C(memaddr_c[8]), .A(n462), .Y(n47) );
  INVX1 U316 ( .A(n280), .Y(n295) );
  NAND21X1 U317 ( .B(n356), .A(n279), .Y(n280) );
  INVX1 U318 ( .A(n292), .Y(n301) );
  NAND21X1 U319 ( .B(n356), .A(n291), .Y(n292) );
  INVX1 U320 ( .A(n288), .Y(n299) );
  NAND21X1 U321 ( .B(n356), .A(n287), .Y(n288) );
  INVX1 U322 ( .A(n284), .Y(n297) );
  NAND21X1 U323 ( .B(n356), .A(n283), .Y(n284) );
  INVX1 U324 ( .A(n282), .Y(n296) );
  NAND21X1 U325 ( .B(n356), .A(n281), .Y(n282) );
  INVX1 U326 ( .A(n290), .Y(n300) );
  NAND21X1 U327 ( .B(n356), .A(n289), .Y(n290) );
  INVX1 U328 ( .A(n294), .Y(n302) );
  NAND21X1 U329 ( .B(n356), .A(n293), .Y(n294) );
  INVX1 U330 ( .A(n286), .Y(n298) );
  NAND21X1 U331 ( .B(n356), .A(n285), .Y(n286) );
  NAND21XL U332 ( .B(n155), .A(memaddr_c[4]), .Y(n208) );
  OAI21BBX1 U333 ( .A(N443), .B(n374), .C(n48), .Y(N838) );
  AOI21X1 U334 ( .B(n18), .C(memaddr_c[12]), .A(n89), .Y(n48) );
  OAI21BBX1 U335 ( .A(N435), .B(n23), .C(n49), .Y(N830) );
  AOI21XL U336 ( .B(memaddr_c[4]), .C(n242), .A(n89), .Y(n49) );
  OAI21BBX1 U337 ( .A(N436), .B(n23), .C(n50), .Y(N831) );
  AOI21XL U338 ( .B(memaddr_c[5]), .C(n242), .A(n89), .Y(n50) );
  OAI21BBX1 U339 ( .A(N442), .B(n374), .C(n51), .Y(N837) );
  AOI21X1 U340 ( .B(n18), .C(memaddr_c[11]), .A(n89), .Y(n51) );
  OAI21BBX1 U341 ( .A(N444), .B(n374), .C(n52), .Y(N839) );
  AOI21X1 U342 ( .B(memaddr_c[13]), .C(n242), .A(n89), .Y(n52) );
  OAI21BBX1 U343 ( .A(N440), .B(n374), .C(n53), .Y(N835) );
  AOI21X1 U344 ( .B(n18), .C(memaddr_c[9]), .A(n462), .Y(n53) );
  OAI21BBX1 U345 ( .A(N438), .B(n374), .C(n54), .Y(N833) );
  AOI21X1 U346 ( .B(n18), .C(memaddr_c[7]), .A(n89), .Y(n54) );
  OAI21BBX1 U347 ( .A(N432), .B(n23), .C(n55), .Y(N827) );
  AOI21XL U348 ( .B(memaddr_c[1]), .C(n18), .A(n89), .Y(n55) );
  OAI21BBX1 U349 ( .A(N433), .B(n23), .C(n56), .Y(N828) );
  AOI21XL U350 ( .B(memaddr_c[2]), .C(n242), .A(n462), .Y(n56) );
  OAI21BBX1 U351 ( .A(N434), .B(n374), .C(n57), .Y(N829) );
  OAI21BBX1 U352 ( .A(N437), .B(n23), .C(n58), .Y(N832) );
  AOI21XL U353 ( .B(memaddr_c[6]), .C(n242), .A(n89), .Y(n58) );
  AO21X1 U354 ( .B(n347), .C(n363), .A(n365), .Y(N874) );
  AO21X1 U355 ( .B(n347), .C(n364), .A(n27), .Y(N875) );
  AO21X1 U356 ( .B(n347), .C(n367), .A(n28), .Y(N876) );
  AO21X1 U357 ( .B(n347), .C(n359), .A(n365), .Y(N877) );
  AO21X1 U358 ( .B(n349), .C(n363), .A(n27), .Y(N878) );
  AO21X1 U359 ( .B(n349), .C(n364), .A(n28), .Y(N879) );
  AO21X1 U360 ( .B(n349), .C(n367), .A(n365), .Y(N880) );
  AO21X1 U361 ( .B(n351), .C(n363), .A(n27), .Y(N882) );
  AO21X1 U362 ( .B(n351), .C(n364), .A(n28), .Y(N883) );
  AO21X1 U363 ( .B(n351), .C(n367), .A(n365), .Y(N884) );
  AO21X1 U364 ( .B(n360), .C(n363), .A(n27), .Y(N890) );
  AO21X1 U365 ( .B(n360), .C(n364), .A(n28), .Y(N891) );
  AO21X1 U366 ( .B(n360), .C(n367), .A(n365), .Y(N892) );
  AO21X1 U367 ( .B(n360), .C(n359), .A(n27), .Y(N893) );
  AO21X1 U368 ( .B(n366), .C(n363), .A(n28), .Y(N894) );
  AO21X1 U369 ( .B(n364), .C(n366), .A(n365), .Y(N895) );
  AO21X1 U370 ( .B(n367), .C(n366), .A(n27), .Y(N896) );
  INVX1 U371 ( .A(n344), .Y(n356) );
  INVX1 U372 ( .A(memaddr_c[12]), .Y(n910) );
  INVXL U373 ( .A(memaddr_c[5]), .Y(n163) );
  INVX1 U374 ( .A(n348), .Y(n349) );
  NAND32X1 U375 ( .B(n362), .C(n352), .A(n353), .Y(n348) );
  INVX1 U376 ( .A(n350), .Y(n351) );
  NAND32X1 U377 ( .B(n353), .C(n352), .A(n362), .Y(n350) );
  OAI211X1 U378 ( .C(n371), .D(n370), .A(n377), .B(n369), .Y(N897) );
  AND2X1 U379 ( .A(n368), .B(n419), .Y(n369) );
  NAND21X1 U380 ( .B(n912), .A(n171), .Y(n203) );
  NAND21X1 U381 ( .B(n68), .A(memaddr_c[13]), .Y(n206) );
  AND4X1 U382 ( .A(n710), .B(n711), .C(n721), .D(n709), .Y(n127) );
  XOR2X1 U383 ( .A(n717), .B(n718), .Y(n710) );
  XNOR2XL U384 ( .A(n715), .B(n716), .Y(n711) );
  XNOR2XL U385 ( .A(n719), .B(n870), .Y(n709) );
  AO21X1 U386 ( .B(n60), .C(n363), .A(n28), .Y(N886) );
  AO21X1 U387 ( .B(n60), .C(n364), .A(n365), .Y(N887) );
  AO21X1 U388 ( .B(n60), .C(n367), .A(n27), .Y(N888) );
  INVX1 U389 ( .A(memaddr_c[14]), .Y(n417) );
  OA21X1 U390 ( .B(n367), .C(n364), .A(n244), .Y(N843) );
  NAND31X1 U391 ( .C(n23), .A(n59), .B(n43), .Y(N825) );
  NAND3X1 U392 ( .A(n343), .B(n906), .C(n342), .Y(n59) );
  INVX1 U393 ( .A(memaddr_c[13]), .Y(n186) );
  NOR5X1 U394 ( .A(n125), .B(n124), .C(n736), .D(n735), .E(n755), .Y(n126) );
  NAND3X1 U395 ( .A(n741), .B(n742), .C(n743), .Y(n735) );
  AOI221XL U396 ( .A(n607), .B(n737), .C(n738), .D(n911), .E(n739), .Y(n736)
         );
  NOR3XL U397 ( .A(n362), .B(n353), .C(n352), .Y(n60) );
  AOI211X1 U398 ( .C(n371), .D(n362), .A(n905), .B(n221), .Y(N844) );
  AND2X1 U399 ( .A(n244), .B(n243), .Y(N842) );
  NOR3XL U400 ( .A(n911), .B(n737), .C(n900), .Y(n739) );
  INVX1 U401 ( .A(n129), .Y(n225) );
  NAND5XL U402 ( .A(n720), .B(n128), .C(n198), .D(n127), .E(n126), .Y(n129) );
  XNOR2XL U403 ( .A(n731), .B(n732), .Y(n720) );
  INVX1 U404 ( .A(n625), .Y(n916) );
  AO21X1 U405 ( .B(sfr_psr), .C(n907), .A(n908), .Y(n325) );
  NAND21X1 U406 ( .B(n331), .A(n433), .Y(n448) );
  XOR2X1 U407 ( .A(n205), .B(memaddr_c[14]), .Y(n211) );
  OAI32X1 U408 ( .A(n446), .B(n445), .C(n444), .D(n443), .E(n442), .Y(n648) );
  NAND32X1 U409 ( .B(n949), .C(n88), .A(n948), .Y(n446) );
  OA21X1 U410 ( .B(n441), .C(n440), .A(n439), .Y(n443) );
  GEN2XL U411 ( .D(n420), .E(n948), .C(n462), .B(n440), .A(n438), .Y(n439) );
  NAND21X1 U412 ( .B(n915), .A(n451), .Y(n235) );
  INVX1 U413 ( .A(n418), .Y(n424) );
  OAI21X1 U414 ( .B(n936), .C(n621), .A(n747), .Y(n742) );
  NAND21X1 U415 ( .B(n869), .A(n621), .Y(n747) );
  XOR2X1 U416 ( .A(n868), .B(n886), .Y(n869) );
  OAI211X1 U417 ( .C(n378), .D(n377), .A(n419), .B(n376), .Y(N898) );
  AND2X1 U418 ( .A(n375), .B(n532), .Y(n378) );
  XOR2XL U419 ( .A(memaddr_c[4]), .B(n62), .Y(n731) );
  OAI31XL U420 ( .A(n420), .B(n908), .C(n529), .D(n948), .Y(n546) );
  INVX1 U421 ( .A(n908), .Y(n442) );
  NAND21X1 U422 ( .B(n314), .A(n313), .Y(n947) );
  NAND21X1 U423 ( .B(n896), .A(n948), .Y(n469) );
  AO21X1 U424 ( .B(n275), .C(n421), .A(n462), .Y(n239) );
  INVX1 U425 ( .A(n453), .Y(n456) );
  NAND32X1 U426 ( .B(n312), .C(n311), .A(n316), .Y(n420) );
  OR2X1 U427 ( .A(n311), .B(n314), .Y(n375) );
  NAND21X1 U428 ( .B(n454), .A(n452), .Y(n471) );
  NAND32X1 U429 ( .B(n316), .C(n311), .A(n312), .Y(n467) );
  NAND21X1 U430 ( .B(n922), .A(n90), .Y(n377) );
  INVX1 U431 ( .A(n459), .Y(n473) );
  NAND21X1 U432 ( .B(n316), .A(n315), .Y(n385) );
  AND2X1 U433 ( .A(n90), .B(n382), .Y(N899) );
  OAI22X1 U434 ( .A(n898), .B(n381), .C(n947), .D(n380), .Y(n382) );
  AND2X1 U435 ( .A(n915), .B(n487), .Y(n381) );
  INVX1 U436 ( .A(n379), .Y(n380) );
  OAI21X1 U437 ( .B(n915), .C(n323), .A(n547), .Y(n426) );
  INVX1 U438 ( .A(hit_ps), .Y(n323) );
  NAND4X1 U439 ( .A(sfr_psw), .B(n907), .C(n930), .D(n929), .Y(n547) );
  ENOX1 U440 ( .A(n249), .B(n906), .C(n906), .D(sfr_psr), .Y(sfr_psrack) );
  INVX1 U441 ( .A(n415), .Y(n919) );
  AO21X1 U442 ( .B(n144), .C(n142), .A(n143), .Y(n149) );
  AO21X1 U443 ( .B(n139), .C(n137), .A(n131), .Y(n160) );
  AO21X1 U444 ( .B(n149), .C(n147), .A(n148), .Y(n139) );
  INVX1 U445 ( .A(n136), .Y(n161) );
  NAND21X1 U446 ( .B(n899), .A(n133), .Y(n179) );
  AO21X1 U447 ( .B(n732), .C(n137), .A(n131), .Y(n868) );
  OR2X1 U448 ( .A(n903), .B(n725), .Y(n935) );
  AO21X1 U449 ( .B(n142), .C(n716), .A(n143), .Y(n871) );
  NAND21X1 U450 ( .B(n934), .A(n161), .Y(n167) );
  OR2X1 U451 ( .A(n902), .B(n167), .Y(n135) );
  NAND21X1 U452 ( .B(n113), .A(n114), .Y(n141) );
  NAND21X1 U453 ( .B(n900), .A(n173), .Y(n180) );
  AO21X1 U454 ( .B(n134), .C(n900), .A(n133), .Y(n178) );
  OAI21BBX1 U455 ( .A(n180), .B(n899), .C(n179), .Y(n181) );
  AO21X1 U456 ( .B(n147), .C(n871), .A(n148), .Y(n732) );
  AO21X1 U457 ( .B(n115), .C(n114), .A(n113), .Y(n716) );
  NAND21X1 U458 ( .B(n148), .A(n147), .Y(n682) );
  NAND21X1 U459 ( .B(n143), .A(n142), .Y(n693) );
  NOR2X1 U460 ( .A(n740), .B(n899), .Y(n754) );
  NOR2X1 U461 ( .A(n727), .B(n901), .Y(n737) );
  INVX1 U462 ( .A(n134), .Y(n173) );
  INVX1 U463 ( .A(n933), .Y(n752) );
  XOR2X1 U464 ( .A(n141), .B(n140), .Y(n61) );
  INVX1 U465 ( .A(n130), .Y(n113) );
  INVX1 U466 ( .A(n115), .Y(n118) );
  INVX1 U467 ( .A(n119), .Y(n121) );
  NAND21X1 U468 ( .B(n118), .A(n140), .Y(n119) );
  AO21X1 U469 ( .B(n899), .C(n740), .A(n754), .Y(n758) );
  INVX1 U470 ( .A(n205), .Y(n188) );
  OAI21X1 U471 ( .B(n901), .C(n727), .A(n728), .Y(n723) );
  INVX1 U472 ( .A(n138), .Y(n131) );
  AND2X1 U473 ( .A(n137), .B(n138), .Y(n62) );
  NAND2X1 U474 ( .A(n901), .B(n727), .Y(n728) );
  OAI21X1 U475 ( .B(n902), .C(n729), .A(n730), .Y(n722) );
  OAI21X1 U476 ( .B(n903), .C(n725), .A(n726), .Y(n724) );
  INVX1 U477 ( .A(n726), .Y(n123) );
  INVX1 U478 ( .A(r_hold_mcu), .Y(n918) );
  NOR2X1 U479 ( .A(n918), .B(n931), .Y(n550) );
  AO21X1 U480 ( .B(n223), .C(n311), .A(n106), .Y(n341) );
  NAND32X1 U481 ( .B(n355), .C(n353), .A(n219), .Y(n224) );
  OR2X1 U482 ( .A(n316), .B(n452), .Y(n232) );
  NAND21X1 U483 ( .B(n906), .A(n336), .Y(n421) );
  INVX1 U484 ( .A(n331), .Y(n247) );
  NAND21X1 U485 ( .B(n454), .A(n383), .Y(n317) );
  INVX1 U486 ( .A(n922), .Y(n897) );
  AND2X1 U487 ( .A(n459), .B(n453), .Y(n63) );
  NAND21X1 U488 ( .B(n915), .A(n247), .Y(n277) );
  INVX1 U489 ( .A(n306), .Y(n905) );
  INVX1 U490 ( .A(n532), .Y(n909) );
  INVX1 U491 ( .A(n470), .Y(n927) );
  INVX1 U492 ( .A(n556), .Y(n926) );
  INVX1 U493 ( .A(n555), .Y(n925) );
  INVX1 U494 ( .A(n558), .Y(n928) );
  NAND2X1 U495 ( .A(n465), .B(n470), .Y(n379) );
  NOR2X1 U496 ( .A(n91), .B(n931), .Y(N152) );
  INVX1 U497 ( .A(n371), .Y(n359) );
  XOR3X1 U498 ( .A(c_adr[4]), .B(memaddr[4]), .C(n481), .Y(n508) );
  OAI22X1 U499 ( .A(memaddr[3]), .B(n872), .C(n480), .D(n479), .Y(n481) );
  AND2X1 U500 ( .A(memaddr[3]), .B(n872), .Y(n479) );
  INVX1 U501 ( .A(n497), .Y(n480) );
  OA222X1 U502 ( .A(n851), .B(n850), .C(n849), .D(n848), .E(n847), .F(n846), 
        .Y(n859) );
  INVX1 U503 ( .A(dbg_06[7]), .Y(n850) );
  INVX1 U504 ( .A(dbg_08[7]), .Y(n848) );
  INVX1 U505 ( .A(dbg_07[7]), .Y(n846) );
  OA222X1 U506 ( .A(n851), .B(n799), .C(n849), .D(n798), .E(n847), .F(n797), 
        .Y(n803) );
  INVX1 U507 ( .A(dbg_06[6]), .Y(n799) );
  INVX1 U508 ( .A(dbg_08[6]), .Y(n798) );
  INVX1 U509 ( .A(dbg_07[6]), .Y(n797) );
  OA222X1 U510 ( .A(n851), .B(n768), .C(n849), .D(n767), .E(n847), .F(n766), 
        .Y(n772) );
  INVX1 U511 ( .A(dbg_06[5]), .Y(n768) );
  INVX1 U512 ( .A(dbg_08[5]), .Y(n767) );
  INVX1 U513 ( .A(dbg_07[5]), .Y(n766) );
  XOR3XL U514 ( .A(c_adr[1]), .B(memaddr[1]), .C(n482), .Y(n484) );
  AO21XL U515 ( .B(memaddr[0]), .C(n877), .A(n483), .Y(n485) );
  OA222X1 U516 ( .A(n828), .B(n827), .C(n826), .D(n825), .E(n824), .F(n823), 
        .Y(n864) );
  INVX1 U517 ( .A(c_buf_16__7_), .Y(n827) );
  INVX1 U518 ( .A(c_buf_17__7_), .Y(n825) );
  INVX1 U519 ( .A(dbg_0f[7]), .Y(n823) );
  OA222X1 U520 ( .A(n828), .B(n788), .C(n826), .D(n787), .E(n824), .F(n786), 
        .Y(n808) );
  INVX1 U521 ( .A(c_buf_16__6_), .Y(n788) );
  INVX1 U522 ( .A(c_buf_17__6_), .Y(n787) );
  INVX1 U523 ( .A(dbg_0f[6]), .Y(n786) );
  OA222X1 U524 ( .A(n828), .B(n734), .C(n826), .D(n733), .E(n824), .F(n714), 
        .Y(n777) );
  INVX1 U525 ( .A(c_buf_16__5_), .Y(n734) );
  INVX1 U526 ( .A(c_buf_17__5_), .Y(n733) );
  INVX1 U527 ( .A(dbg_0f[5]), .Y(n714) );
  OA222X1 U528 ( .A(n828), .B(n549), .C(n826), .D(n548), .E(n824), .F(n545), 
        .Y(n581) );
  INVX1 U529 ( .A(c_buf_16__1_), .Y(n549) );
  INVX1 U530 ( .A(c_buf_17__1_), .Y(n548) );
  INVX1 U531 ( .A(dbg_0f[1]), .Y(n545) );
  OA222X1 U532 ( .A(n828), .B(n638), .C(n826), .D(n637), .E(n824), .F(n636), 
        .Y(n669) );
  INVX1 U533 ( .A(c_buf_16__3_), .Y(n638) );
  INVX1 U534 ( .A(c_buf_17__3_), .Y(n637) );
  INVX1 U535 ( .A(dbg_0f[3]), .Y(n636) );
  OA222X1 U536 ( .A(n828), .B(n501), .C(n826), .D(n500), .E(n824), .F(n499), 
        .Y(n535) );
  INVX1 U537 ( .A(c_buf_16__0_), .Y(n501) );
  INVX1 U538 ( .A(c_buf_17__0_), .Y(n500) );
  INVX1 U539 ( .A(dbg_0f[0]), .Y(n499) );
  OA222X1 U540 ( .A(n828), .B(n680), .C(n826), .D(n679), .E(n824), .F(n678), 
        .Y(n702) );
  INVX1 U541 ( .A(c_buf_16__4_), .Y(n680) );
  INVX1 U542 ( .A(c_buf_17__4_), .Y(n679) );
  INVX1 U543 ( .A(dbg_0f[4]), .Y(n678) );
  OA222X1 U544 ( .A(n828), .B(n596), .C(n826), .D(n595), .E(n824), .F(n594), 
        .Y(n627) );
  INVX1 U545 ( .A(c_buf_16__2_), .Y(n596) );
  INVX1 U546 ( .A(c_buf_17__2_), .Y(n595) );
  INVX1 U547 ( .A(dbg_0f[2]), .Y(n594) );
  OA222X1 U548 ( .A(n851), .B(n660), .C(n849), .D(n659), .E(n847), .F(n658), 
        .Y(n664) );
  INVX1 U549 ( .A(dbg_06[3]), .Y(n660) );
  INVX1 U550 ( .A(dbg_08[3]), .Y(n659) );
  INVX1 U551 ( .A(dbg_07[3]), .Y(n658) );
  OA222X1 U552 ( .A(n851), .B(n692), .C(n849), .D(n691), .E(n847), .F(n690), 
        .Y(n697) );
  INVX1 U553 ( .A(dbg_06[4]), .Y(n692) );
  INVX1 U554 ( .A(dbg_08[4]), .Y(n691) );
  INVX1 U555 ( .A(dbg_07[4]), .Y(n690) );
  OA222X1 U556 ( .A(n851), .B(n567), .C(n849), .D(n566), .E(n847), .F(n565), 
        .Y(n571) );
  INVX1 U557 ( .A(dbg_06[1]), .Y(n567) );
  INVX1 U558 ( .A(dbg_08[1]), .Y(n566) );
  INVX1 U559 ( .A(dbg_07[1]), .Y(n565) );
  OA222X1 U560 ( .A(n851), .B(n521), .C(n849), .D(n520), .E(n847), .F(n519), 
        .Y(n528) );
  INVX1 U561 ( .A(dbg_06[0]), .Y(n521) );
  INVX1 U562 ( .A(dbg_08[0]), .Y(n520) );
  INVX1 U563 ( .A(dbg_07[0]), .Y(n519) );
  OA222X1 U564 ( .A(n851), .B(n616), .C(n849), .D(n614), .E(n847), .F(n613), 
        .Y(n620) );
  INVX1 U565 ( .A(dbg_06[2]), .Y(n616) );
  INVX1 U566 ( .A(dbg_08[2]), .Y(n614) );
  INVX1 U567 ( .A(dbg_07[2]), .Y(n613) );
  NAND21X1 U568 ( .B(pwrdn_rst), .A(n92), .Y(n462) );
  AND2X1 U569 ( .A(n90), .B(n475), .Y(n641) );
  AO21X1 U570 ( .B(n474), .C(n473), .A(n472), .Y(n475) );
  OAI31XL U571 ( .A(n471), .B(n469), .C(n468), .D(n467), .Y(n472) );
  INVX1 U572 ( .A(pmem_clk[0]), .Y(n468) );
  AOI21X1 U573 ( .B(n386), .C(n385), .A(n88), .Y(n643) );
  AOI31X1 U574 ( .A(n249), .B(test_so1), .C(n420), .D(n384), .Y(n386) );
  INVX1 U575 ( .A(n383), .Y(n384) );
  AOI21XL U576 ( .B(n463), .C(n467), .A(n88), .Y(n642) );
  AOI32X1 U577 ( .A(pmem_clk[1]), .B(n458), .C(n457), .D(n474), .E(n456), .Y(
        n463) );
  INVX1 U578 ( .A(n471), .Y(n457) );
  INVX1 U579 ( .A(n469), .Y(n458) );
  INVX1 U580 ( .A(c_adr[3]), .Y(n872) );
  INVXL U581 ( .A(c_adr[0]), .Y(n877) );
  OAI22X1 U582 ( .A(mcu_psw), .B(n949), .C(n249), .D(n915), .Y(mempsack) );
  INVX1 U583 ( .A(dbg_0a[7]), .Y(n852) );
  INVX1 U584 ( .A(rd_buf[3]), .Y(n944) );
  INVX1 U585 ( .A(rd_buf[5]), .Y(n943) );
  INVX1 U586 ( .A(rd_buf[6]), .Y(n942) );
  INVX1 U587 ( .A(rd_buf[7]), .Y(n950) );
  INVX1 U588 ( .A(rd_buf[4]), .Y(n945) );
  INVX1 U589 ( .A(wr_buf[5]), .Y(n706) );
  INVX1 U590 ( .A(wr_buf[6]), .Y(n781) );
  INVX1 U591 ( .A(wr_buf[3]), .Y(n631) );
  INVX1 U592 ( .A(wr_buf[7]), .Y(n813) );
  INVX1 U593 ( .A(dbg_02[1]), .Y(n562) );
  INVX1 U594 ( .A(dbg_05[1]), .Y(n560) );
  INVX1 U595 ( .A(dbg_0a[1]), .Y(n568) );
  INVX1 U596 ( .A(dbg_02[0]), .Y(n513) );
  INVX1 U597 ( .A(dbg_05[0]), .Y(n510) );
  INVX1 U598 ( .A(dbg_0a[0]), .Y(n525) );
  INVX1 U599 ( .A(dbg_02[3]), .Y(n655) );
  INVX1 U600 ( .A(dbg_05[3]), .Y(n653) );
  INVX1 U601 ( .A(dbg_0a[3]), .Y(n661) );
  INVX1 U602 ( .A(dbg_02[4]), .Y(n687) );
  INVX1 U603 ( .A(dbg_05[4]), .Y(n685) );
  INVX1 U604 ( .A(dbg_0a[4]), .Y(n694) );
  INVX1 U605 ( .A(c_buf_21__3_), .Y(n630) );
  INVX1 U606 ( .A(c_buf_18__3_), .Y(n633) );
  INVX1 U607 ( .A(dbg_0c[3]), .Y(n639) );
  INVX1 U608 ( .A(dbg_02[5]), .Y(n763) );
  INVX1 U609 ( .A(dbg_05[5]), .Y(n760) );
  INVX1 U610 ( .A(dbg_0a[5]), .Y(n769) );
  INVX1 U611 ( .A(dbg_02[6]), .Y(n794) );
  INVX1 U612 ( .A(dbg_05[6]), .Y(n792) );
  INVX1 U613 ( .A(dbg_0a[6]), .Y(n800) );
  INVX1 U614 ( .A(dbg_02[7]), .Y(n840) );
  INVX1 U615 ( .A(dbg_05[7]), .Y(n835) );
  INVX1 U616 ( .A(c_buf_21__5_), .Y(n705) );
  INVX1 U617 ( .A(c_buf_18__5_), .Y(n708) );
  INVX1 U618 ( .A(dbg_0c[5]), .Y(n748) );
  INVX1 U619 ( .A(c_buf_21__6_), .Y(n780) );
  INVX1 U620 ( .A(c_buf_18__6_), .Y(n783) );
  INVX1 U621 ( .A(dbg_0c[6]), .Y(n789) );
  INVX1 U622 ( .A(c_buf_21__7_), .Y(n811) );
  INVX1 U623 ( .A(c_buf_18__7_), .Y(n817) );
  INVX1 U624 ( .A(dbg_0c[7]), .Y(n829) );
  INVX1 U625 ( .A(dbg_01[1]), .Y(n563) );
  INVX1 U626 ( .A(dbg_04[1]), .Y(n561) );
  INVX1 U627 ( .A(dbg_0b[1]), .Y(n569) );
  INVX1 U628 ( .A(dbg_01[0]), .Y(n514) );
  INVX1 U629 ( .A(dbg_04[0]), .Y(n511) );
  INVX1 U630 ( .A(dbg_0b[0]), .Y(n526) );
  INVX1 U631 ( .A(dbg_01[3]), .Y(n656) );
  INVX1 U632 ( .A(dbg_04[3]), .Y(n654) );
  INVX1 U633 ( .A(dbg_0b[3]), .Y(n662) );
  INVX1 U634 ( .A(dbg_01[4]), .Y(n688) );
  INVX1 U635 ( .A(dbg_04[4]), .Y(n686) );
  INVX1 U636 ( .A(dbg_0b[4]), .Y(n695) );
  INVX1 U637 ( .A(dbg_0e[3]), .Y(n640) );
  INVX1 U638 ( .A(dbg_01[5]), .Y(n764) );
  INVX1 U639 ( .A(dbg_04[5]), .Y(n761) );
  INVX1 U640 ( .A(dbg_0b[5]), .Y(n770) );
  INVX1 U641 ( .A(dbg_01[6]), .Y(n795) );
  INVX1 U642 ( .A(dbg_04[6]), .Y(n793) );
  INVX1 U643 ( .A(dbg_0b[6]), .Y(n801) );
  INVX1 U644 ( .A(dbg_01[7]), .Y(n842) );
  INVX1 U645 ( .A(dbg_04[7]), .Y(n837) );
  INVX1 U646 ( .A(dbg_0b[7]), .Y(n854) );
  INVX1 U647 ( .A(c_buf_20__5_), .Y(n712) );
  INVX1 U648 ( .A(dbg_0e[5]), .Y(n749) );
  INVX1 U649 ( .A(c_buf_20__6_), .Y(n784) );
  INVX1 U650 ( .A(dbg_0e[6]), .Y(n790) );
  INVX1 U651 ( .A(c_buf_20__7_), .Y(n819) );
  INVX1 U652 ( .A(dbg_0e[7]), .Y(n831) );
  INVX1 U653 ( .A(dbg_03[1]), .Y(n564) );
  INVX1 U654 ( .A(dbg_09[1]), .Y(n570) );
  INVX1 U655 ( .A(dbg_03[0]), .Y(n515) );
  INVX1 U656 ( .A(dbg_09[0]), .Y(n527) );
  INVX1 U657 ( .A(dbg_03[3]), .Y(n657) );
  INVX1 U658 ( .A(dbg_09[3]), .Y(n663) );
  INVX1 U659 ( .A(dbg_03[4]), .Y(n689) );
  INVX1 U660 ( .A(dbg_09[4]), .Y(n696) );
  INVX1 U661 ( .A(dbg_0d[3]), .Y(n652) );
  INVX1 U662 ( .A(dbg_03[5]), .Y(n765) );
  INVX1 U663 ( .A(dbg_09[5]), .Y(n771) );
  INVX1 U664 ( .A(dbg_03[6]), .Y(n796) );
  INVX1 U665 ( .A(dbg_09[6]), .Y(n802) );
  INVX1 U666 ( .A(dbg_03[7]), .Y(n844) );
  INVX1 U667 ( .A(dbg_09[7]), .Y(n856) );
  INVX1 U668 ( .A(dbg_0d[5]), .Y(n759) );
  INVX1 U669 ( .A(c_buf_22__6_), .Y(n782) );
  INVX1 U670 ( .A(c_buf_19__6_), .Y(n785) );
  INVX1 U671 ( .A(dbg_0d[6]), .Y(n791) );
  INVX1 U672 ( .A(c_buf_22__7_), .Y(n815) );
  INVX1 U673 ( .A(c_buf_19__7_), .Y(n821) );
  INVX1 U674 ( .A(dbg_0d[7]), .Y(n833) );
  INVX1 U675 ( .A(n253), .Y(o_bkp_hold) );
  INVX1 U676 ( .A(memaddr[12]), .Y(n924) );
  NAND21X1 U677 ( .B(cs_ft[0]), .A(cs_ft[1]), .Y(n223) );
  XNOR2XL U678 ( .A(memaddr[10]), .B(bkpt_pc[10]), .Y(n408) );
  XNOR2XL U679 ( .A(memaddr[7]), .B(bkpt_pc[7]), .Y(n400) );
  XOR2X1 U680 ( .A(bkpt_pc[8]), .B(memaddr[8]), .Y(n395) );
  XOR2X1 U681 ( .A(bkpt_pc[13]), .B(memaddr[13]), .Y(n403) );
  XOR2X1 U682 ( .A(bkpt_pc[9]), .B(memaddr[9]), .Y(n396) );
  XNOR2XL U683 ( .A(bkpt_pc[12]), .B(n924), .Y(n404) );
  INVX1 U684 ( .A(cs_ft[2]), .Y(n316) );
  NAND2X1 U685 ( .A(n391), .B(n392), .Y(n253) );
  NOR4XL U686 ( .A(n393), .B(n394), .C(n395), .D(n396), .Y(n392) );
  NOR4XL U687 ( .A(n401), .B(n402), .C(n403), .D(n404), .Y(n391) );
  NAND3X1 U688 ( .A(n938), .B(r_rdy), .C(bkpt_ena), .Y(n394) );
  INVX1 U689 ( .A(cs_ft[3]), .Y(n312) );
  INVX1 U690 ( .A(mcu_psw), .Y(n915) );
  NAND4X1 U691 ( .A(n408), .B(n409), .C(n410), .D(n411), .Y(n401) );
  XNOR2XL U692 ( .A(memaddr[0]), .B(bkpt_pc[0]), .Y(n409) );
  XNOR2XL U693 ( .A(memaddr[5]), .B(bkpt_pc[5]), .Y(n410) );
  XNOR2XL U694 ( .A(memaddr[4]), .B(bkpt_pc[4]), .Y(n411) );
  NAND4X1 U695 ( .A(n397), .B(n398), .C(n399), .D(n400), .Y(n393) );
  XNOR2XL U696 ( .A(memaddr[3]), .B(bkpt_pc[3]), .Y(n397) );
  XNOR2XL U697 ( .A(memaddr[1]), .B(bkpt_pc[1]), .Y(n398) );
  XNOR2XL U698 ( .A(memaddr[6]), .B(bkpt_pc[6]), .Y(n399) );
  NAND3X1 U699 ( .A(n405), .B(n406), .C(n407), .Y(n402) );
  XNOR2XL U700 ( .A(memaddr[2]), .B(bkpt_pc[2]), .Y(n406) );
  XNOR2XL U701 ( .A(memaddr[14]), .B(bkpt_pc[14]), .Y(n405) );
  XNOR2XL U702 ( .A(memaddr[11]), .B(bkpt_pc[11]), .Y(n407) );
  INVX1 U703 ( .A(rd_buf[1]), .Y(n941) );
  INVX1 U704 ( .A(rd_buf[2]), .Y(n940) );
  INVX1 U705 ( .A(wr_buf[0]), .Y(n487) );
  INVX1 U706 ( .A(rd_buf[0]), .Y(n946) );
  INVX1 U707 ( .A(wr_buf[1]), .Y(n539) );
  INVX1 U708 ( .A(wr_buf[4]), .Y(n673) );
  INVX1 U709 ( .A(wr_buf[2]), .Y(n585) );
  INVX1 U710 ( .A(c_buf_21__1_), .Y(n538) );
  INVX1 U711 ( .A(c_buf_18__1_), .Y(n541) );
  INVX1 U712 ( .A(dbg_0c[1]), .Y(n551) );
  INVX1 U713 ( .A(c_buf_21__0_), .Y(n486) );
  INVX1 U714 ( .A(c_buf_18__0_), .Y(n493) );
  INVX1 U715 ( .A(dbg_0c[0]), .Y(n504) );
  INVX1 U716 ( .A(dbg_02[2]), .Y(n602) );
  INVX1 U717 ( .A(dbg_05[2]), .Y(n600) );
  INVX1 U718 ( .A(dbg_0a[2]), .Y(n617) );
  INVX1 U719 ( .A(c_buf_21__2_), .Y(n584) );
  INVX1 U720 ( .A(c_buf_18__2_), .Y(n587) );
  INVX1 U721 ( .A(dbg_0c[2]), .Y(n597) );
  INVX1 U722 ( .A(c_buf_21__4_), .Y(n672) );
  INVX1 U723 ( .A(c_buf_18__4_), .Y(n675) );
  INVX1 U724 ( .A(dbg_0c[4]), .Y(n681) );
  INVX1 U725 ( .A(c_buf_20__1_), .Y(n542) );
  INVX1 U726 ( .A(dbg_0e[1]), .Y(n552) );
  INVX1 U727 ( .A(c_buf_20__0_), .Y(n494) );
  INVX1 U728 ( .A(dbg_0e[0]), .Y(n505) );
  INVX1 U729 ( .A(dbg_01[2]), .Y(n604) );
  INVX1 U730 ( .A(dbg_04[2]), .Y(n601) );
  INVX1 U731 ( .A(dbg_0b[2]), .Y(n618) );
  INVX1 U732 ( .A(c_buf_20__2_), .Y(n588) );
  INVX1 U733 ( .A(dbg_0e[2]), .Y(n598) );
  INVX1 U734 ( .A(c_buf_20__3_), .Y(n634) );
  INVX1 U735 ( .A(c_buf_20__4_), .Y(n676) );
  INVX1 U736 ( .A(dbg_0e[4]), .Y(n683) );
  INVX1 U737 ( .A(c_buf_22__1_), .Y(n540) );
  INVX1 U738 ( .A(c_buf_19__1_), .Y(n544) );
  INVX1 U739 ( .A(dbg_0d[1]), .Y(n559) );
  INVX1 U740 ( .A(c_buf_22__0_), .Y(n488) );
  INVX1 U741 ( .A(c_buf_19__0_), .Y(n495) );
  INVX1 U742 ( .A(dbg_0d[0]), .Y(n506) );
  INVX1 U743 ( .A(dbg_03[2]), .Y(n612) );
  INVX1 U744 ( .A(dbg_09[2]), .Y(n619) );
  INVX1 U745 ( .A(c_buf_22__2_), .Y(n586) );
  INVX1 U746 ( .A(c_buf_19__2_), .Y(n592) );
  INVX1 U747 ( .A(dbg_0d[2]), .Y(n599) );
  INVX1 U748 ( .A(c_buf_22__3_), .Y(n632) );
  INVX1 U749 ( .A(c_buf_19__3_), .Y(n635) );
  INVX1 U750 ( .A(c_buf_22__4_), .Y(n674) );
  INVX1 U751 ( .A(c_buf_19__4_), .Y(n677) );
  INVX1 U752 ( .A(dbg_0d[4]), .Y(n684) );
  INVX1 U753 ( .A(c_buf_22__5_), .Y(n707) );
  INVX1 U754 ( .A(c_buf_19__5_), .Y(n713) );
  INVX1 U755 ( .A(r_rdy), .Y(n949) );
  INVX1 U756 ( .A(un_hold), .Y(n938) );
  NAND32X1 U757 ( .B(d_psrd), .C(n341), .A(n229), .Y(n337) );
  AO21X1 U758 ( .B(c_adr[7]), .C(n914), .A(n890), .Y(n611) );
  INVX1 U759 ( .A(n615), .Y(n889) );
  OAI221X1 U760 ( .A(c_adr[6]), .B(n887), .C(n886), .D(n885), .E(n615), .Y(
        n888) );
  AO21X1 U761 ( .B(n437), .C(n436), .A(n435), .Y(n646) );
  AND3X1 U762 ( .A(wd_twlb[0]), .B(we_twlb), .C(n433), .Y(n437) );
  MUX2X1 U763 ( .D0(n434), .D1(pmem_twlb[0]), .S(n40), .Y(n435) );
  AO21X1 U764 ( .B(n432), .C(n436), .A(n431), .Y(n645) );
  AND3X1 U765 ( .A(wd_twlb[1]), .B(we_twlb), .C(n433), .Y(n432) );
  MUX2X1 U766 ( .D0(n434), .D1(pmem_twlb[1]), .S(n40), .Y(n431) );
  AOI221XL U767 ( .A(n608), .B(n609), .C(memaddr_c[10]), .D(n901), .E(n607), 
        .Y(n605) );
  NAND2X1 U768 ( .A(c_adr[9]), .B(n912), .Y(n609) );
  AOI32X1 U769 ( .A(n916), .B(n913), .C(c_adr[8]), .D(n610), .E(n611), .Y(n608) );
  AOI21X1 U770 ( .B(memaddr_c[8]), .C(n902), .A(n625), .Y(n610) );
  OAI22X1 U771 ( .A(memaddr_c[13]), .B(n195), .C(n194), .D(n193), .Y(n196) );
  INVX1 U772 ( .A(c_adr[13]), .Y(n195) );
  OA22X1 U773 ( .A(n603), .B(n192), .C(memaddr_c[12]), .D(n899), .Y(n193) );
  AOI211X1 U774 ( .C(c_adr[11]), .D(n911), .A(n605), .B(n606), .Y(n192) );
  OAI32X1 U775 ( .A(n232), .B(d_psrd), .C(n88), .D(n440), .E(n231), .Y(n414)
         );
  NAND21XL U776 ( .B(c_adr[5]), .A(memaddr_c[5]), .Y(n621) );
  NAND32X1 U777 ( .B(d_psrd), .C(n229), .A(n224), .Y(n340) );
  NAND21X1 U778 ( .B(d_psrd), .A(n322), .Y(n308) );
  NAND2X1 U779 ( .A(n2), .B(pre_1_adr[14]), .Y(n429) );
  OAI211X1 U780 ( .C(pre_1_adr[13]), .D(n429), .A(n428), .B(n427), .Y(n434) );
  AOI33X1 U781 ( .A(n426), .B(n425), .C(n424), .D(sfr_psofs[14]), .E(n423), 
        .F(n422), .Y(n427) );
  NAND32X1 U782 ( .B(memaddr_c[13]), .C(n417), .A(n414), .Y(n428) );
  INVX1 U783 ( .A(sfr_psofs[13]), .Y(n422) );
  NOR2X1 U784 ( .A(n911), .B(c_adr[11]), .Y(n607) );
  OAI211X1 U785 ( .C(n240), .D(n239), .A(n418), .B(n238), .Y(N868) );
  INVX1 U786 ( .A(sfr_psofs[14]), .Y(n240) );
  OA21X1 U787 ( .B(n237), .C(n417), .A(n429), .Y(n238) );
  INVX1 U788 ( .A(n414), .Y(n237) );
  NAND21X1 U789 ( .B(d_psrd), .A(n340), .Y(n344) );
  NAND32X1 U790 ( .B(c_ptr[4]), .C(n345), .A(n344), .Y(n352) );
  AO2222XL U791 ( .A(memaddr[10]), .B(n234), .C(sfr_psofs[10]), .D(n233), .E(
        memaddr_c[10]), .F(n414), .G(pre_1_adr[10]), .H(n2), .Y(N864) );
  INVX1 U792 ( .A(n358), .Y(n360) );
  NAND21X1 U793 ( .B(c_ptr[2]), .A(n361), .Y(n358) );
  AO2222XL U794 ( .A(memaddr[8]), .B(n12), .C(sfr_psofs[8]), .D(n9), .E(n19), 
        .F(memaddr_c[8]), .G(pre_1_adr[8]), .H(n2), .Y(N862) );
  AO2222XL U795 ( .A(memaddr[7]), .B(n234), .C(sfr_psofs[7]), .D(n233), .E(
        n414), .F(memaddr_c[7]), .G(pre_1_adr[7]), .H(n236), .Y(N861) );
  AO2222XL U796 ( .A(memaddr[12]), .B(n234), .C(sfr_psofs[12]), .D(n233), .E(
        n19), .F(memaddr_c[12]), .G(pre_1_adr[12]), .H(n2), .Y(N866) );
  AO2222XL U797 ( .A(memaddr[9]), .B(n234), .C(sfr_psofs[9]), .D(n233), .E(n19), .F(memaddr_c[9]), .G(pre_1_adr[9]), .H(n236), .Y(N863) );
  AO2222XL U798 ( .A(memaddr[11]), .B(n234), .C(sfr_psofs[11]), .D(n233), .E(
        n19), .F(memaddr_c[11]), .G(pre_1_adr[11]), .H(n2), .Y(N865) );
  AO2222XL U799 ( .A(memaddr[13]), .B(n234), .C(sfr_psofs[13]), .D(n233), .E(
        memaddr_c[13]), .F(n414), .G(pre_1_adr[13]), .H(n236), .Y(N867) );
  AO2222XL U800 ( .A(memaddr[5]), .B(n234), .C(sfr_psofs[5]), .D(n233), .E(
        memaddr_c[5]), .F(n414), .G(pre_1_adr[5]), .H(n236), .Y(N859) );
  AO2222XL U801 ( .A(memaddr[4]), .B(n234), .C(sfr_psofs[4]), .D(n233), .E(
        memaddr_c[4]), .F(n414), .G(pre_1_adr[4]), .H(n2), .Y(N858) );
  AO21X1 U802 ( .B(N445), .C(n374), .A(n241), .Y(N840) );
  AO21X1 U803 ( .B(memaddr_c[14]), .C(n242), .A(n89), .Y(n241) );
  AO21X1 U804 ( .B(n86), .C(dbg_01[7]), .A(n295), .Y(N486) );
  AO21X1 U805 ( .B(n86), .C(dbg_02[7]), .A(n25), .Y(N494) );
  AO21X1 U806 ( .B(n85), .C(dbg_03[7]), .A(n26), .Y(N502) );
  AO21X1 U807 ( .B(n84), .C(dbg_04[7]), .A(n295), .Y(N510) );
  AO21X1 U808 ( .B(n83), .C(dbg_05[7]), .A(n25), .Y(N518) );
  AO21X1 U809 ( .B(n82), .C(dbg_06[7]), .A(n26), .Y(N526) );
  AO21X1 U810 ( .B(n82), .C(dbg_07[7]), .A(n295), .Y(N534) );
  AO21X1 U811 ( .B(n81), .C(dbg_08[7]), .A(n25), .Y(N542) );
  AO21X1 U812 ( .B(n80), .C(dbg_09[7]), .A(n26), .Y(N550) );
  AO21X1 U813 ( .B(n79), .C(dbg_0a[7]), .A(n295), .Y(N558) );
  AO21X1 U814 ( .B(n78), .C(dbg_0b[7]), .A(n25), .Y(N566) );
  AO21X1 U815 ( .B(n78), .C(dbg_0c[7]), .A(n26), .Y(N574) );
  AO21X1 U816 ( .B(n77), .C(dbg_0d[7]), .A(n295), .Y(N582) );
  AO21X1 U817 ( .B(n76), .C(dbg_0e[7]), .A(n25), .Y(N590) );
  AO21X1 U818 ( .B(n75), .C(dbg_0f[7]), .A(n26), .Y(N598) );
  AO21X1 U819 ( .B(n74), .C(c_buf_16__7_), .A(n295), .Y(N606) );
  AO21X1 U820 ( .B(n74), .C(c_buf_17__7_), .A(n25), .Y(N614) );
  AO21X1 U821 ( .B(n73), .C(c_buf_18__7_), .A(n26), .Y(N622) );
  AO21X1 U822 ( .B(n72), .C(c_buf_19__7_), .A(n295), .Y(N630) );
  AO21X1 U823 ( .B(n71), .C(c_buf_20__7_), .A(n25), .Y(N638) );
  AO21X1 U824 ( .B(n70), .C(c_buf_21__7_), .A(n26), .Y(N646) );
  AO21X1 U825 ( .B(n70), .C(c_buf_22__7_), .A(n295), .Y(N654) );
  AO21X1 U826 ( .B(n69), .C(wr_buf[7]), .A(n25), .Y(N662) );
  AO21X1 U827 ( .B(n303), .C(dbg_01[0]), .A(n302), .Y(N479) );
  AO21X1 U828 ( .B(n303), .C(dbg_01[4]), .A(n298), .Y(N483) );
  AO21X1 U829 ( .B(n303), .C(dbg_01[3]), .A(n299), .Y(N482) );
  AO21X1 U830 ( .B(n303), .C(dbg_01[5]), .A(n297), .Y(N484) );
  AO21X1 U831 ( .B(n86), .C(dbg_01[6]), .A(n296), .Y(N485) );
  AO21X1 U832 ( .B(n86), .C(dbg_02[0]), .A(n20), .Y(N487) );
  AO21X1 U833 ( .B(n85), .C(dbg_03[0]), .A(n21), .Y(N495) );
  AO21X1 U834 ( .B(n85), .C(dbg_04[0]), .A(n302), .Y(N503) );
  AO21X1 U835 ( .B(n84), .C(dbg_05[0]), .A(n20), .Y(N511) );
  AO21X1 U836 ( .B(n83), .C(dbg_06[0]), .A(n21), .Y(N519) );
  AO21X1 U837 ( .B(n86), .C(dbg_02[3]), .A(n13), .Y(N490) );
  AO21X1 U838 ( .B(n85), .C(dbg_03[3]), .A(n14), .Y(N498) );
  AO21X1 U839 ( .B(n84), .C(dbg_04[3]), .A(n299), .Y(N506) );
  AO21X1 U840 ( .B(n84), .C(dbg_05[3]), .A(n13), .Y(N514) );
  AO21X1 U841 ( .B(n83), .C(dbg_06[3]), .A(n14), .Y(N522) );
  AO21X1 U842 ( .B(n82), .C(dbg_07[3]), .A(n299), .Y(N530) );
  AO21X1 U843 ( .B(n86), .C(dbg_02[4]), .A(n10), .Y(N491) );
  AO21X1 U844 ( .B(n85), .C(dbg_03[4]), .A(n11), .Y(N499) );
  AO21X1 U845 ( .B(n84), .C(dbg_04[4]), .A(n298), .Y(N507) );
  AO21X1 U846 ( .B(n83), .C(dbg_05[4]), .A(n10), .Y(N515) );
  AO21X1 U847 ( .B(n83), .C(dbg_06[4]), .A(n11), .Y(N523) );
  AO21X1 U848 ( .B(n86), .C(dbg_02[5]), .A(n7), .Y(N492) );
  AO21X1 U849 ( .B(n85), .C(dbg_03[5]), .A(n8), .Y(N500) );
  AO21X1 U850 ( .B(n84), .C(dbg_04[5]), .A(n297), .Y(N508) );
  AO21X1 U851 ( .B(n83), .C(dbg_05[5]), .A(n7), .Y(N516) );
  AO21X1 U852 ( .B(n83), .C(dbg_06[5]), .A(n8), .Y(N524) );
  AO21X1 U853 ( .B(n82), .C(dbg_07[5]), .A(n297), .Y(N532) );
  AO21X1 U854 ( .B(n86), .C(dbg_02[6]), .A(n5), .Y(N493) );
  AO21X1 U855 ( .B(n85), .C(dbg_03[6]), .A(n6), .Y(N501) );
  AO21X1 U856 ( .B(n84), .C(dbg_04[6]), .A(n296), .Y(N509) );
  AO21X1 U857 ( .B(n83), .C(dbg_05[6]), .A(n5), .Y(N517) );
  AO21X1 U858 ( .B(n82), .C(dbg_06[6]), .A(n6), .Y(N525) );
  AO21X1 U859 ( .B(n82), .C(dbg_07[6]), .A(n296), .Y(N533) );
  AO21X1 U860 ( .B(n81), .C(dbg_08[0]), .A(n302), .Y(N535) );
  AO21X1 U861 ( .B(n81), .C(dbg_08[3]), .A(n13), .Y(N538) );
  AO21X1 U862 ( .B(n81), .C(dbg_08[4]), .A(n298), .Y(N539) );
  AO21X1 U863 ( .B(n81), .C(dbg_08[5]), .A(n7), .Y(N540) );
  AO21X1 U864 ( .B(n81), .C(dbg_08[6]), .A(n5), .Y(N541) );
  AO21X1 U865 ( .B(n81), .C(dbg_09[0]), .A(n20), .Y(N543) );
  AO21X1 U866 ( .B(n80), .C(dbg_09[3]), .A(n14), .Y(N546) );
  AO21X1 U867 ( .B(n80), .C(dbg_09[4]), .A(n10), .Y(N547) );
  AO21X1 U868 ( .B(n80), .C(dbg_09[5]), .A(n8), .Y(N548) );
  AO21X1 U869 ( .B(n80), .C(dbg_09[6]), .A(n6), .Y(N549) );
  AO21X1 U870 ( .B(n80), .C(dbg_0a[3]), .A(n299), .Y(N554) );
  AO21X1 U871 ( .B(n79), .C(dbg_0a[5]), .A(n297), .Y(N556) );
  AO21X1 U872 ( .B(n79), .C(dbg_0a[6]), .A(n296), .Y(N557) );
  AO21X1 U873 ( .B(n79), .C(dbg_0b[0]), .A(n21), .Y(N559) );
  AO21X1 U874 ( .B(n79), .C(dbg_0b[3]), .A(n13), .Y(N562) );
  AO21X1 U875 ( .B(n79), .C(dbg_0b[4]), .A(n11), .Y(N563) );
  AO21X1 U876 ( .B(n79), .C(dbg_0b[5]), .A(n7), .Y(N564) );
  AO21X1 U877 ( .B(n78), .C(dbg_0b[6]), .A(n5), .Y(N565) );
  AO21X1 U878 ( .B(n78), .C(dbg_0c[0]), .A(n302), .Y(N567) );
  AO21X1 U879 ( .B(n78), .C(dbg_0c[3]), .A(n14), .Y(N570) );
  AO21X1 U880 ( .B(n78), .C(dbg_0c[4]), .A(n298), .Y(N571) );
  AO21X1 U881 ( .B(n78), .C(dbg_0c[5]), .A(n8), .Y(N572) );
  AO21X1 U882 ( .B(n78), .C(dbg_0c[6]), .A(n6), .Y(N573) );
  AO21X1 U883 ( .B(n77), .C(dbg_0d[3]), .A(n299), .Y(N578) );
  AO21X1 U884 ( .B(n77), .C(dbg_0d[6]), .A(n296), .Y(N581) );
  AO21X1 U885 ( .B(n76), .C(dbg_0e[3]), .A(n13), .Y(N586) );
  AO21X1 U886 ( .B(n76), .C(dbg_0e[6]), .A(n5), .Y(N589) );
  AO21X1 U887 ( .B(n75), .C(c_buf_16__3_), .A(n14), .Y(N602) );
  AO21X1 U888 ( .B(n74), .C(c_buf_16__6_), .A(n6), .Y(N605) );
  AO21X1 U889 ( .B(n74), .C(c_buf_17__3_), .A(n299), .Y(N610) );
  AO21X1 U890 ( .B(n303), .C(dbg_01[1]), .A(n301), .Y(N480) );
  AO21X1 U891 ( .B(n303), .C(dbg_01[2]), .A(n300), .Y(N481) );
  AO21X1 U892 ( .B(n82), .C(dbg_07[0]), .A(n20), .Y(N527) );
  AO21X1 U893 ( .B(n86), .C(dbg_02[1]), .A(n16), .Y(N488) );
  AO21X1 U894 ( .B(n85), .C(dbg_03[1]), .A(n17), .Y(N496) );
  AO21X1 U895 ( .B(n85), .C(dbg_04[1]), .A(n301), .Y(N504) );
  AO21X1 U896 ( .B(n84), .C(dbg_05[1]), .A(n16), .Y(N512) );
  AO21X1 U897 ( .B(n83), .C(dbg_06[1]), .A(n17), .Y(N520) );
  AO21X1 U898 ( .B(n82), .C(dbg_07[1]), .A(n301), .Y(N528) );
  AO21X1 U899 ( .B(n86), .C(dbg_02[2]), .A(n3), .Y(N489) );
  AO21X1 U900 ( .B(n85), .C(dbg_03[2]), .A(n4), .Y(N497) );
  AO21X1 U901 ( .B(n84), .C(dbg_04[2]), .A(n300), .Y(N505) );
  AO21X1 U902 ( .B(n84), .C(dbg_05[2]), .A(n3), .Y(N513) );
  AO21X1 U903 ( .B(n83), .C(dbg_06[2]), .A(n4), .Y(N521) );
  AO21X1 U904 ( .B(n82), .C(dbg_07[2]), .A(n300), .Y(N529) );
  AO21X1 U905 ( .B(n82), .C(dbg_07[4]), .A(n10), .Y(N531) );
  AO21X1 U906 ( .B(n81), .C(dbg_08[1]), .A(n16), .Y(N536) );
  AO21X1 U907 ( .B(n81), .C(dbg_08[2]), .A(n3), .Y(N537) );
  AO21X1 U908 ( .B(n81), .C(dbg_09[1]), .A(n17), .Y(N544) );
  AO21X1 U909 ( .B(n80), .C(dbg_09[2]), .A(n4), .Y(N545) );
  AO21X1 U910 ( .B(n80), .C(dbg_0a[0]), .A(n21), .Y(N551) );
  AO21X1 U911 ( .B(n80), .C(dbg_0a[1]), .A(n301), .Y(N552) );
  AO21X1 U912 ( .B(n80), .C(dbg_0a[2]), .A(n300), .Y(N553) );
  AO21X1 U913 ( .B(n79), .C(dbg_0a[4]), .A(n11), .Y(N555) );
  AO21X1 U914 ( .B(n79), .C(dbg_0b[1]), .A(n16), .Y(N560) );
  AO21X1 U915 ( .B(n79), .C(dbg_0b[2]), .A(n3), .Y(N561) );
  AO21X1 U916 ( .B(n78), .C(dbg_0c[1]), .A(n17), .Y(N568) );
  AO21X1 U917 ( .B(n78), .C(dbg_0c[2]), .A(n4), .Y(N569) );
  AO21X1 U918 ( .B(n77), .C(dbg_0d[0]), .A(n302), .Y(N575) );
  AO21X1 U919 ( .B(n77), .C(dbg_0d[1]), .A(n301), .Y(N576) );
  AO21X1 U920 ( .B(n77), .C(dbg_0d[2]), .A(n300), .Y(N577) );
  AO21X1 U921 ( .B(n77), .C(dbg_0d[4]), .A(n298), .Y(N579) );
  AO21X1 U922 ( .B(n77), .C(dbg_0d[5]), .A(n297), .Y(N580) );
  AO21X1 U923 ( .B(n77), .C(dbg_0e[0]), .A(n20), .Y(N583) );
  AO21X1 U924 ( .B(n77), .C(dbg_0e[1]), .A(n16), .Y(N584) );
  AO21X1 U925 ( .B(n76), .C(dbg_0e[2]), .A(n3), .Y(N585) );
  AO21X1 U926 ( .B(n76), .C(dbg_0e[4]), .A(n10), .Y(N587) );
  AO21X1 U927 ( .B(n76), .C(dbg_0e[5]), .A(n7), .Y(N588) );
  AO21X1 U928 ( .B(n76), .C(dbg_0f[0]), .A(n21), .Y(N591) );
  AO21X1 U929 ( .B(n76), .C(dbg_0f[1]), .A(n17), .Y(N592) );
  AO21X1 U930 ( .B(n76), .C(dbg_0f[2]), .A(n4), .Y(N593) );
  AO21X1 U931 ( .B(n76), .C(dbg_0f[3]), .A(n13), .Y(N594) );
  AO21X1 U932 ( .B(n75), .C(dbg_0f[4]), .A(n11), .Y(N595) );
  AO21X1 U933 ( .B(n75), .C(dbg_0f[5]), .A(n8), .Y(N596) );
  AO21X1 U934 ( .B(n75), .C(dbg_0f[6]), .A(n296), .Y(N597) );
  AO21X1 U935 ( .B(n75), .C(c_buf_16__0_), .A(n302), .Y(N599) );
  AO21X1 U936 ( .B(n75), .C(c_buf_16__1_), .A(n301), .Y(N600) );
  AO21X1 U937 ( .B(n75), .C(c_buf_16__2_), .A(n300), .Y(N601) );
  AO21X1 U938 ( .B(n75), .C(c_buf_16__4_), .A(n298), .Y(N603) );
  AO21X1 U939 ( .B(n75), .C(c_buf_16__5_), .A(n297), .Y(N604) );
  AO21X1 U940 ( .B(n74), .C(c_buf_17__0_), .A(n20), .Y(N607) );
  AO21X1 U941 ( .B(n74), .C(c_buf_17__1_), .A(n16), .Y(N608) );
  AO21X1 U942 ( .B(n74), .C(c_buf_17__2_), .A(n3), .Y(N609) );
  AO21X1 U943 ( .B(n74), .C(c_buf_17__4_), .A(n10), .Y(N611) );
  AO21X1 U944 ( .B(n74), .C(c_buf_17__5_), .A(n7), .Y(N612) );
  AO21X1 U945 ( .B(n74), .C(c_buf_17__6_), .A(n5), .Y(N613) );
  AO21X1 U946 ( .B(n73), .C(c_buf_18__0_), .A(n21), .Y(N615) );
  AO21X1 U947 ( .B(n73), .C(c_buf_18__1_), .A(n17), .Y(N616) );
  AO21X1 U948 ( .B(n73), .C(c_buf_18__2_), .A(n4), .Y(N617) );
  AO21X1 U949 ( .B(n73), .C(c_buf_18__3_), .A(n14), .Y(N618) );
  AO21X1 U950 ( .B(n73), .C(c_buf_18__4_), .A(n11), .Y(N619) );
  AO21X1 U951 ( .B(n73), .C(c_buf_18__5_), .A(n8), .Y(N620) );
  AO21X1 U952 ( .B(n73), .C(c_buf_18__6_), .A(n6), .Y(N621) );
  AO21X1 U953 ( .B(n73), .C(c_buf_19__0_), .A(n302), .Y(N623) );
  AO21X1 U954 ( .B(n73), .C(c_buf_19__1_), .A(n301), .Y(N624) );
  AO21X1 U955 ( .B(n72), .C(c_buf_19__2_), .A(n300), .Y(N625) );
  AO21X1 U956 ( .B(n72), .C(c_buf_19__3_), .A(n299), .Y(N626) );
  AO21X1 U957 ( .B(n72), .C(c_buf_19__4_), .A(n298), .Y(N627) );
  AO21X1 U958 ( .B(n72), .C(c_buf_19__5_), .A(n297), .Y(N628) );
  AO21X1 U959 ( .B(n72), .C(c_buf_19__6_), .A(n296), .Y(N629) );
  AO21X1 U960 ( .B(n72), .C(c_buf_20__0_), .A(n20), .Y(N631) );
  AO21X1 U961 ( .B(n72), .C(c_buf_20__1_), .A(n16), .Y(N632) );
  AO21X1 U962 ( .B(n72), .C(c_buf_20__2_), .A(n3), .Y(N633) );
  AO21X1 U963 ( .B(n72), .C(c_buf_20__3_), .A(n13), .Y(N634) );
  AO21X1 U964 ( .B(n71), .C(c_buf_20__4_), .A(n10), .Y(N635) );
  AO21X1 U965 ( .B(n71), .C(c_buf_20__5_), .A(n7), .Y(N636) );
  AO21X1 U966 ( .B(n71), .C(c_buf_20__6_), .A(n5), .Y(N637) );
  AO21X1 U967 ( .B(n71), .C(c_buf_21__0_), .A(n21), .Y(N639) );
  AO21X1 U968 ( .B(n71), .C(c_buf_21__1_), .A(n17), .Y(N640) );
  AO21X1 U969 ( .B(n71), .C(c_buf_21__3_), .A(n14), .Y(N642) );
  AO21X1 U970 ( .B(n71), .C(c_buf_21__4_), .A(n11), .Y(N643) );
  AO21X1 U971 ( .B(n71), .C(c_buf_21__5_), .A(n8), .Y(N644) );
  AO21X1 U972 ( .B(n70), .C(c_buf_21__6_), .A(n6), .Y(N645) );
  AO21X1 U973 ( .B(n70), .C(c_buf_22__0_), .A(n302), .Y(N647) );
  AO21X1 U974 ( .B(n70), .C(c_buf_22__1_), .A(n301), .Y(N648) );
  AO21X1 U975 ( .B(n70), .C(c_buf_22__2_), .A(n4), .Y(N649) );
  AO21X1 U976 ( .B(n70), .C(c_buf_22__3_), .A(n299), .Y(N650) );
  AO21X1 U977 ( .B(n70), .C(c_buf_22__4_), .A(n298), .Y(N651) );
  AO21X1 U978 ( .B(n70), .C(c_buf_22__5_), .A(n297), .Y(N652) );
  AO21X1 U979 ( .B(n70), .C(c_buf_22__6_), .A(n296), .Y(N653) );
  AO21X1 U980 ( .B(n69), .C(wr_buf[0]), .A(n20), .Y(N655) );
  AO21X1 U981 ( .B(n69), .C(wr_buf[1]), .A(n16), .Y(N656) );
  AO21X1 U982 ( .B(n69), .C(wr_buf[2]), .A(n300), .Y(N657) );
  AO21X1 U983 ( .B(n69), .C(wr_buf[3]), .A(n13), .Y(N658) );
  AO21X1 U984 ( .B(n69), .C(wr_buf[4]), .A(n10), .Y(N659) );
  AO21X1 U985 ( .B(n69), .C(wr_buf[5]), .A(n7), .Y(N660) );
  AO21X1 U986 ( .B(n69), .C(wr_buf[6]), .A(n5), .Y(N661) );
  AO21X1 U987 ( .B(n71), .C(c_buf_21__2_), .A(n3), .Y(N641) );
  AO21X1 U988 ( .B(N431), .C(n374), .A(n230), .Y(N826) );
  NOR2X1 U989 ( .A(n912), .B(c_adr[9]), .Y(n625) );
  INVX1 U990 ( .A(n357), .Y(n361) );
  NAND43X1 U991 ( .B(c_ptr[3]), .C(n356), .D(n355), .A(n354), .Y(n357) );
  INVX1 U992 ( .A(n346), .Y(n347) );
  NAND32X1 U993 ( .B(c_ptr[2]), .C(n352), .A(n353), .Y(n346) );
  OAI21X1 U994 ( .B(n310), .C(n88), .A(n309), .Y(N822) );
  AND4X1 U995 ( .A(n948), .B(n467), .C(n421), .D(n305), .Y(n310) );
  GEN2XL U996 ( .D(n356), .E(n308), .C(n307), .B(n388), .A(n345), .Y(n309) );
  AOI221XL U997 ( .A(n897), .B(n909), .C(n454), .D(mcu_psw), .E(n343), .Y(n305) );
  INVX1 U998 ( .A(n867), .Y(n886) );
  NAND21XL U999 ( .B(memaddr_c[5]), .A(c_adr[5]), .Y(n867) );
  NAND21X1 U1000 ( .B(c_adr[14]), .A(memaddr_c[14]), .Y(n870) );
  GEN2XL U1001 ( .D(n330), .E(n329), .C(n24), .B(n354), .A(n328), .Y(N824) );
  NAND21X1 U1002 ( .B(n327), .A(n326), .Y(n328) );
  AND3X1 U1003 ( .A(n321), .B(cs_ft[0]), .C(n388), .Y(n330) );
  AOI21X1 U1004 ( .B(n921), .C(n529), .A(n322), .Y(n329) );
  AND2X1 U1005 ( .A(hit_ps_c), .B(mcu_psr_c), .Y(n908) );
  MUX2X1 U1006 ( .D0(n109), .D1(n194), .S(n754), .Y(n110) );
  AND2X1 U1007 ( .A(c_adr[13]), .B(memaddr_c[13]), .Y(n109) );
  NAND32X1 U1008 ( .B(n896), .C(n332), .A(n318), .Y(n319) );
  AOI32X1 U1009 ( .A(n375), .B(mcu_psw), .C(n317), .D(n897), .E(n532), .Y(n318) );
  OAI31XL U1010 ( .A(n932), .B(memaddr_c[10]), .C(n737), .D(n756), .Y(n755) );
  INVX1 U1011 ( .A(n728), .Y(n932) );
  OAI21BX1 U1012 ( .C(n603), .B(n740), .A(n757), .Y(n756) );
  AOI32X1 U1013 ( .A(c_adr[12]), .B(n740), .C(memaddr_c[12]), .D(n758), .E(
        n910), .Y(n757) );
  OAI31XL U1014 ( .A(n112), .B(memaddr_c[8]), .C(n752), .D(n111), .Y(n125) );
  INVX1 U1015 ( .A(n730), .Y(n112) );
  AO21X1 U1016 ( .B(n753), .C(n186), .A(n110), .Y(n111) );
  OAI21X1 U1017 ( .B(c_adr[13]), .C(n754), .A(n719), .Y(n753) );
  AND2X1 U1018 ( .A(n244), .B(n220), .Y(N846) );
  XOR2X1 U1019 ( .A(n355), .B(n502), .Y(n220) );
  NAND2X1 U1020 ( .A(n905), .B(c_ptr[3]), .Y(n502) );
  AND2X1 U1021 ( .A(n222), .B(n244), .Y(N845) );
  XOR2X1 U1022 ( .A(c_ptr[3]), .B(n905), .Y(n222) );
  MUX2IX1 U1023 ( .D0(n64), .D1(n65), .S(n445), .Y(n390) );
  NAND2X1 U1024 ( .A(pmem_re), .B(n387), .Y(n64) );
  NAND2XL U1025 ( .A(n389), .B(n90), .Y(n65) );
  INVX1 U1026 ( .A(n108), .Y(n194) );
  NAND21X1 U1027 ( .B(c_adr[13]), .A(memaddr_c[13]), .Y(n108) );
  INVX1 U1028 ( .A(n191), .Y(n603) );
  NAND21X1 U1029 ( .B(c_adr[12]), .A(memaddr_c[12]), .Y(n191) );
  NAND21X1 U1030 ( .B(memaddr_c[14]), .A(c_adr[14]), .Y(n198) );
  NOR5X1 U1031 ( .A(c_ptr[3]), .B(n438), .C(n306), .D(n24), .E(n355), .Y(n307)
         );
  OAI22XL U1032 ( .A(n88), .B(n421), .C(mcu_psw), .D(n419), .Y(n423) );
  OAI21X1 U1033 ( .B(n935), .C(n615), .A(n744), .Y(n743) );
  AOI32X1 U1034 ( .A(c_adr[7]), .B(n935), .C(memaddr_c[7]), .D(n745), .E(n914), 
        .Y(n744) );
  OAI21X1 U1035 ( .B(c_adr[7]), .C(n746), .A(n729), .Y(n745) );
  NAND21X1 U1036 ( .B(n235), .A(memaddr[14]), .Y(n418) );
  OAI21X1 U1037 ( .B(n933), .C(n916), .A(n750), .Y(n741) );
  AOI32X1 U1038 ( .A(c_adr[9]), .B(n933), .C(memaddr_c[9]), .D(n751), .E(n912), 
        .Y(n750) );
  OAI21X1 U1039 ( .B(c_adr[9]), .C(n752), .A(n727), .Y(n751) );
  INVX1 U1040 ( .A(test_so1), .Y(pmem_csb) );
  NAND21X1 U1041 ( .B(d_psrd), .A(n354), .Y(n440) );
  MUX2X1 U1042 ( .D0(n451), .D1(pmem_pgm), .S(n450), .Y(n644) );
  AND2X1 U1043 ( .A(n449), .B(n448), .Y(n450) );
  INVX1 U1044 ( .A(n447), .Y(n449) );
  MUX2X1 U1045 ( .D0(n100), .D1(n24), .S(n387), .Y(n649) );
  AND2X1 U1046 ( .A(n451), .B(n442), .Y(n100) );
  MUX2BXL U1047 ( .D0(n904), .D1(n589), .S(adr_p[14]), .Y(n453) );
  NOR2X1 U1048 ( .A(n590), .B(n591), .Y(n589) );
  OR4X1 U1049 ( .A(pmem_a[12]), .B(pmem_a[13]), .C(pmem_a[14]), .D(pmem_a[15]), 
        .Y(n590) );
  NAND42X1 U1050 ( .C(pmem_a[10]), .D(pmem_a[11]), .A(pmem_a[9]), .B(n904), 
        .Y(n591) );
  NAND21X1 U1051 ( .B(n312), .A(cs_ft[2]), .Y(n314) );
  INVX1 U1052 ( .A(n94), .Y(n313) );
  NAND21X1 U1053 ( .B(cs_ft[0]), .A(n102), .Y(n94) );
  AOI21BBXL U1054 ( .B(wspp_cnt_3_), .C(n465), .A(test_so2), .Y(n466) );
  NOR4XL U1055 ( .A(wspp_cnt_3_), .B(wspp_cnt_4_), .C(wspp_cnt_5_), .D(
        test_so2), .Y(n465) );
  XNOR2XL U1056 ( .A(wspp_cnt_5_), .B(wspp_cnt_3_), .Y(n464) );
  NAND32X1 U1057 ( .B(n336), .C(n543), .A(n385), .Y(n320) );
  OAI31XL U1058 ( .A(n922), .B(wr_buf[0]), .C(n909), .D(n947), .Y(n543) );
  INVX1 U1059 ( .A(n455), .Y(n474) );
  OAI31XL U1060 ( .A(pmem_re), .B(n461), .C(n460), .D(n469), .Y(n455) );
  AOI221XL U1061 ( .A(wspp_cnt_5_), .B(n937), .C(n464), .D(test_so2), .E(n465), 
        .Y(n461) );
  OAI21X1 U1062 ( .B(n466), .C(wspp_cnt_4_), .A(r_multi), .Y(n460) );
  AO21X1 U1063 ( .B(adr_p[14]), .C(n246), .A(adr_p[13]), .Y(n459) );
  NAND43X1 U1064 ( .B(n593), .C(pmem_a[10]), .D(pmem_a[12]), .A(n245), .Y(n246) );
  INVX1 U1065 ( .A(pmem_a[11]), .Y(n245) );
  OR4X1 U1066 ( .A(pmem_a[9]), .B(pmem_a[13]), .C(pmem_a[14]), .D(pmem_a[15]), 
        .Y(n593) );
  OR2X1 U1067 ( .A(cs_ft[3]), .B(n223), .Y(n452) );
  NAND32X1 U1068 ( .B(n103), .C(n102), .A(n101), .Y(n948) );
  INVX1 U1069 ( .A(cs_ft[0]), .Y(n103) );
  INVX1 U1070 ( .A(n106), .Y(n101) );
  NAND21X1 U1071 ( .B(cs_ft[2]), .A(n312), .Y(n106) );
  NAND21X1 U1072 ( .B(cs_ft[1]), .A(cs_ft[0]), .Y(n311) );
  INVX1 U1073 ( .A(cs_ft[1]), .Y(n102) );
  INVX1 U1074 ( .A(adr_p[13]), .Y(n904) );
  INVX1 U1075 ( .A(wspp_cnt_4_), .Y(n937) );
  NAND43X1 U1076 ( .B(cs_ft[2]), .C(cs_ft[1]), .D(cs_ft[0]), .A(cs_ft[3]), .Y(
        n383) );
  INVX1 U1077 ( .A(n95), .Y(n315) );
  NAND21X1 U1078 ( .B(cs_ft[3]), .A(n313), .Y(n95) );
  NAND2X1 U1079 ( .A(d_psrd), .B(n950), .Y(d_inst[7]) );
  NOR2X1 U1080 ( .A(n906), .B(n946), .Y(d_inst[0]) );
  NAND2X1 U1081 ( .A(n24), .B(n942), .Y(d_inst[6]) );
  NAND2X1 U1082 ( .A(d_psrd), .B(n941), .Y(d_inst[1]) );
  NAND2X1 U1083 ( .A(d_psrd), .B(n940), .Y(d_inst[2]) );
  NAND2X1 U1084 ( .A(n24), .B(n943), .Y(d_inst[5]) );
  NAND2X1 U1085 ( .A(n24), .B(n944), .Y(d_inst[3]) );
  NOR2X1 U1086 ( .A(n906), .B(n945), .Y(d_inst[4]) );
  NAND3X1 U1087 ( .A(n416), .B(sfr_psw), .C(dw_ena), .Y(n415) );
  OAI33XL U1088 ( .A(n415), .B(dummy[1]), .C(dummy[0]), .D(n930), .E(n919), 
        .F(n920), .Y(n651) );
  OAI33XL U1089 ( .A(n415), .B(dummy[1]), .C(n930), .D(n929), .E(n919), .F(
        n920), .Y(n650) );
  NAND21X1 U1090 ( .B(n243), .A(c_ptr[1]), .Y(n371) );
  XOR2X1 U1091 ( .A(n160), .B(c_adr[5]), .Y(n162) );
  INVX1 U1092 ( .A(c_ptr[0]), .Y(n243) );
  NAND31X1 U1093 ( .C(n903), .A(c_adr[5]), .B(n160), .Y(n136) );
  NAND21X1 U1094 ( .B(n880), .A(c_ptr[1]), .Y(n130) );
  OR2X1 U1095 ( .A(n161), .B(n66), .Y(n164) );
  AOI21X1 U1096 ( .B(c_adr[5]), .C(n160), .A(c_adr[6]), .Y(n66) );
  INVX1 U1097 ( .A(n116), .Y(n143) );
  NAND21XL U1098 ( .B(n876), .A(c_ptr[2]), .Y(n116) );
  INVXL U1099 ( .A(c_adr[1]), .Y(n880) );
  NAND21X1 U1100 ( .B(n936), .A(c_adr[5]), .Y(n725) );
  NAND21X1 U1101 ( .B(n729), .A(c_adr[8]), .Y(n933) );
  OR2X1 U1102 ( .A(n173), .B(n67), .Y(n175) );
  AOI21X1 U1103 ( .B(n172), .C(c_adr[9]), .A(c_adr[10]), .Y(n67) );
  NAND21XL U1104 ( .B(c_adr[0]), .A(n243), .Y(n115) );
  NAND31X1 U1105 ( .C(n901), .A(c_adr[9]), .B(n172), .Y(n134) );
  XOR2X1 U1106 ( .A(n167), .B(c_adr[8]), .Y(n168) );
  XOR2X1 U1107 ( .A(n135), .B(c_adr[9]), .Y(n171) );
  XOR2X1 U1108 ( .A(n136), .B(c_adr[7]), .Y(n166) );
  NAND21XL U1109 ( .B(c_adr[2]), .A(n362), .Y(n142) );
  OR2XL U1110 ( .A(c_adr[1]), .B(c_ptr[1]), .Y(n114) );
  INVX1 U1111 ( .A(c_ptr[3]), .Y(n353) );
  INVX1 U1112 ( .A(c_ptr[2]), .Y(n362) );
  NAND2X1 U1113 ( .A(n746), .B(c_adr[7]), .Y(n729) );
  NAND2X1 U1114 ( .A(n752), .B(c_adr[9]), .Y(n727) );
  OAI221XL U1115 ( .A(n265), .B(n341), .C(memdatao[4]), .D(n277), .E(n264), 
        .Y(N790) );
  INVX1 U1116 ( .A(n285), .Y(n265) );
  OA22X1 U1117 ( .A(sfr_wdat[4]), .B(n275), .C(n898), .D(n706), .Y(n264) );
  NAND2X1 U1118 ( .A(n737), .B(c_adr[11]), .Y(n740) );
  INVX1 U1119 ( .A(n117), .Y(n148) );
  NAND21X1 U1120 ( .B(n883), .A(c_ptr[4]), .Y(n138) );
  XOR2X1 U1121 ( .A(n132), .B(c_adr[14]), .Y(n205) );
  NAND21X1 U1122 ( .B(n179), .A(c_adr[13]), .Y(n132) );
  OAI222XL U1123 ( .A(memdatao[7]), .B(n277), .C(n256), .D(n341), .E(
        sfr_wdat[7]), .F(n275), .Y(N793) );
  INVX1 U1124 ( .A(n279), .Y(n256) );
  INVX1 U1125 ( .A(c_ptr[4]), .Y(n355) );
  OAI221XL U1126 ( .A(n278), .B(n341), .C(memdatao[0]), .D(n277), .E(n276), 
        .Y(N786) );
  INVX1 U1127 ( .A(n293), .Y(n278) );
  OA22X1 U1128 ( .A(sfr_wdat[0]), .B(n275), .C(n898), .D(n539), .Y(n276) );
  INVX1 U1129 ( .A(n291), .Y(n274) );
  OA22X1 U1130 ( .A(sfr_wdat[1]), .B(n275), .C(n898), .D(n585), .Y(n273) );
  OAI221X1 U1131 ( .A(n263), .B(n15), .C(memdatao[5]), .D(n277), .E(n262), .Y(
        N791) );
  INVX1 U1132 ( .A(n283), .Y(n263) );
  OA22X1 U1133 ( .A(sfr_wdat[5]), .B(n275), .C(n898), .D(n781), .Y(n262) );
  OAI221XL U1134 ( .A(n268), .B(n341), .C(memdatao[3]), .D(n277), .E(n267), 
        .Y(N789) );
  INVX1 U1135 ( .A(n287), .Y(n268) );
  OA22X1 U1136 ( .A(sfr_wdat[3]), .B(n275), .C(n898), .D(n673), .Y(n267) );
  OAI221X1 U1137 ( .A(n260), .B(n15), .C(memdatao[6]), .D(n277), .E(n258), .Y(
        N792) );
  INVX1 U1138 ( .A(n281), .Y(n260) );
  OA22X1 U1139 ( .A(sfr_wdat[6]), .B(n275), .C(n898), .D(n813), .Y(n258) );
  INVX1 U1140 ( .A(n289), .Y(n271) );
  OA22X1 U1141 ( .A(sfr_wdat[2]), .B(n275), .C(n898), .D(n631), .Y(n270) );
  OAI21X1 U1142 ( .B(c_adr[11]), .C(n737), .A(n740), .Y(n738) );
  XNOR2XL U1143 ( .A(n179), .B(c_adr[13]), .Y(n68) );
  NAND2X1 U1144 ( .A(n754), .B(c_adr[13]), .Y(n719) );
  INVX1 U1145 ( .A(c_adr[6]), .Y(n903) );
  NAND21X1 U1146 ( .B(c_adr[8]), .A(n729), .Y(n730) );
  NAND21X1 U1147 ( .B(c_adr[6]), .A(n725), .Y(n726) );
  INVX1 U1148 ( .A(c_adr[10]), .Y(n901) );
  INVX1 U1149 ( .A(c_adr[7]), .Y(n934) );
  INVX1 U1150 ( .A(c_adr[8]), .Y(n902) );
  INVX1 U1151 ( .A(c_adr[11]), .Y(n900) );
  AND3XL U1152 ( .A(r_rdy), .B(o_inst[7]), .C(n259), .Y(n892) );
  NOR3XL U1153 ( .A(memaddr[0]), .B(memaddr[11]), .C(memaddr[10]), .Y(n259) );
  OAI31XL U1154 ( .A(n250), .B(n251), .C(n252), .D(n253), .Y(o_set_hold) );
  NAND42X1 U1155 ( .C(memaddr[14]), .D(memaddr[13]), .A(n924), .B(n254), .Y(
        n252) );
  NAND43X1 U1156 ( .B(memaddr[5]), .C(memaddr[6]), .D(memaddr[4]), .A(n255), 
        .Y(n251) );
  NAND42X1 U1157 ( .C(n895), .D(n894), .A(n893), .B(n892), .Y(n250) );
  INVX1 U1158 ( .A(n99), .Y(n907) );
  NAND43X1 U1159 ( .B(n98), .C(n97), .D(n96), .A(n550), .Y(n99) );
  INVX1 U1160 ( .A(d_hold[3]), .Y(n98) );
  INVX1 U1161 ( .A(d_hold[1]), .Y(n97) );
  INVX1 U1162 ( .A(c_adr[12]), .Y(n899) );
  INVX1 U1163 ( .A(n189), .Y(n363) );
  NAND21X1 U1164 ( .B(c_ptr[1]), .A(n243), .Y(n189) );
  INVX1 U1165 ( .A(n190), .Y(n219) );
  NAND21X1 U1166 ( .B(c_ptr[2]), .A(n363), .Y(n190) );
  AOI21X1 U1167 ( .B(hit_ps), .C(mcu_psw), .A(n907), .Y(n529) );
  INVX1 U1168 ( .A(d_psrd), .Y(n906) );
  NAND21X1 U1169 ( .B(cs_ft[2]), .A(n315), .Y(n331) );
  OAI31XL U1170 ( .A(n938), .B(n91), .C(r_rdy), .D(n917), .Y(n762) );
  INVX1 U1171 ( .A(n923), .Y(n917) );
  INVX1 U1172 ( .A(dummy[0]), .Y(n930) );
  INVX1 U1173 ( .A(d_hold[0]), .Y(n931) );
  INVX1 U1174 ( .A(dummy[1]), .Y(n929) );
  INVX1 U1175 ( .A(d_hold[2]), .Y(n96) );
  NAND21X1 U1176 ( .B(mcu_psw), .A(n317), .Y(n922) );
  NAND21X1 U1177 ( .B(n63), .A(n248), .Y(n279) );
  MUX2X1 U1178 ( .D0(pmem_q1[7]), .D1(pmem_q0[7]), .S(n473), .Y(n248) );
  NAND21X1 U1179 ( .B(n63), .A(n272), .Y(n291) );
  MUX2X1 U1180 ( .D0(pmem_q1[1]), .D1(pmem_q0[1]), .S(n473), .Y(n272) );
  NAND21X1 U1181 ( .B(n63), .A(n261), .Y(n283) );
  MUX2X1 U1182 ( .D0(pmem_q1[5]), .D1(pmem_q0[5]), .S(n473), .Y(n261) );
  NAND21X1 U1183 ( .B(n63), .A(n266), .Y(n287) );
  MUX2X1 U1184 ( .D0(pmem_q1[3]), .D1(pmem_q0[3]), .S(n473), .Y(n266) );
  NAND21X1 U1185 ( .B(n63), .A(n257), .Y(n281) );
  MUX2X1 U1186 ( .D0(pmem_q1[6]), .D1(pmem_q0[6]), .S(n473), .Y(n257) );
  NAND21X1 U1187 ( .B(n63), .A(n269), .Y(n289) );
  MUX2X1 U1188 ( .D0(pmem_q1[2]), .D1(pmem_q0[2]), .S(n473), .Y(n269) );
  OAI22X1 U1189 ( .A(pmem_q1[0]), .B(n453), .C(pmem_q0[0]), .D(n459), .Y(n293)
         );
  OAI22X1 U1190 ( .A(pmem_q1[4]), .B(n453), .C(pmem_q0[4]), .D(n459), .Y(n285)
         );
  INVX1 U1191 ( .A(memaddr[13]), .Y(n425) );
  NOR3XL U1192 ( .A(memaddr[7]), .B(memaddr[9]), .C(memaddr[8]), .Y(n255) );
  NOR21XL U1193 ( .B(n575), .A(pmem_a[6]), .Y(N757) );
  NAND21X1 U1194 ( .B(n371), .A(c_ptr[2]), .Y(n306) );
  NAND21X1 U1195 ( .B(mcu_psw), .A(n247), .Y(n275) );
  GEN2XL U1196 ( .D(n575), .E(n951), .C(N757), .B(pmem_a[8]), .A(n576), .Y(
        N759) );
  NOR42XL U1197 ( .C(pmem_a[6]), .D(n575), .A(n951), .B(pmem_a[8]), .Y(n576)
         );
  GEN2XL U1198 ( .D(wspp_cnt_1_), .E(wspp_cnt_0_), .C(n558), .B(n896), .A(n897), .Y(N796) );
  GEN2XL U1199 ( .D(wspp_cnt_2_), .E(n928), .C(n470), .B(n896), .A(n897), .Y(
        N797) );
  GEN2XL U1200 ( .D(wspp_cnt_4_), .E(n926), .C(n555), .B(n896), .A(n897), .Y(
        N799) );
  GEN2XL U1201 ( .D(wspp_cnt_5_), .E(n925), .C(n554), .B(n896), .A(n897), .Y(
        N800) );
  INVX1 U1202 ( .A(n577), .Y(n939) );
  AOI32X1 U1203 ( .A(pmem_a[6]), .B(n951), .C(n575), .D(pmem_a[7]), .E(N757), 
        .Y(n577) );
  NOR2X1 U1204 ( .A(n928), .B(wspp_cnt_2_), .Y(n470) );
  OAI21X1 U1205 ( .B(n553), .C(n947), .A(n922), .Y(N801) );
  XNOR2XL U1206 ( .A(test_so2), .B(n554), .Y(n553) );
  NOR2X1 U1207 ( .A(n927), .B(wspp_cnt_3_), .Y(n556) );
  NOR2X1 U1208 ( .A(wspp_cnt_1_), .B(wspp_cnt_0_), .Y(n558) );
  NOR2X1 U1209 ( .A(n926), .B(wspp_cnt_4_), .Y(n555) );
  NAND2X1 U1210 ( .A(n578), .B(n579), .Y(n532) );
  NOR4XL U1211 ( .A(wr_buf[3]), .B(wr_buf[2]), .C(wr_buf[1]), .D(wr_buf[0]), 
        .Y(n578) );
  NOR4XL U1212 ( .A(wr_buf[7]), .B(wr_buf[6]), .C(wr_buf[5]), .D(wr_buf[4]), 
        .Y(n579) );
  NOR3XL U1213 ( .A(memaddr[1]), .B(memaddr[3]), .C(memaddr[2]), .Y(n254) );
  OAI21X1 U1214 ( .B(wspp_cnt_0_), .C(n947), .A(n922), .Y(N795) );
  NOR2X1 U1215 ( .A(n925), .B(wspp_cnt_5_), .Y(n554) );
  NOR21XL U1216 ( .B(d_hold[1]), .A(n91), .Y(N153) );
  NOR21XL U1217 ( .B(d_hold[2]), .A(n91), .Y(N154) );
  INVX1 U1218 ( .A(pmem_a[7]), .Y(n951) );
  INVX1 U1219 ( .A(n104), .Y(n367) );
  NAND21X1 U1220 ( .B(c_ptr[0]), .A(c_ptr[1]), .Y(n104) );
  INVX1 U1221 ( .A(n105), .Y(n364) );
  NAND21X1 U1222 ( .B(c_ptr[1]), .A(c_ptr[0]), .Y(n105) );
  NOR2X1 U1223 ( .A(n557), .B(n947), .Y(N798) );
  AOI21X1 U1224 ( .B(wspp_cnt_3_), .C(n927), .A(n556), .Y(n557) );
  INVX1 U1225 ( .A(r_pwdn_en), .Y(n921) );
  AO2222XL U1226 ( .A(memaddr[6]), .B(n12), .C(sfr_psofs[6]), .D(n9), .E(
        memaddr_c[6]), .F(n19), .G(pre_1_adr[6]), .H(n236), .Y(N860) );
  OAI32XL U1227 ( .A(n123), .B(memaddr_c[6]), .C(n746), .D(n153), .E(n122), 
        .Y(n124) );
  AOI222XL U1228 ( .A(memaddr_c[8]), .B(n722), .C(memaddr_c[10]), .D(n723), 
        .E(memaddr_c[6]), .F(n724), .Y(n721) );
  OAI31XL U1229 ( .A(memaddr_c[6]), .B(n903), .C(n889), .D(n888), .Y(n890) );
  INVXL U1230 ( .A(memaddr_c[6]), .Y(n887) );
  AO2222XL U1231 ( .A(n234), .B(memaddr[2]), .C(sfr_psofs[2]), .D(n233), .E(
        memaddr_c[2]), .F(n414), .G(pre_1_adr[2]), .H(n236), .Y(N856) );
  XNOR2XL U1232 ( .A(memaddr_c[2]), .B(n693), .Y(n715) );
  GEN2XL U1233 ( .D(memaddr_c[2]), .E(n876), .C(n875), .B(n878), .A(n874), .Y(
        n882) );
  INVXL U1234 ( .A(memaddr_c[2]), .Y(n145) );
  AO2222XL U1235 ( .A(n12), .B(memaddr[0]), .C(sfr_psofs[0]), .D(n9), .E(
        memaddr_c[0]), .F(n19), .G(pre_1_adr[0]), .H(n2), .Y(N854) );
  AO21XL U1236 ( .B(memaddr_c[0]), .C(n242), .A(n88), .Y(n230) );
  NAND21XL U1237 ( .B(n121), .A(memaddr_c[0]), .Y(n213) );
  NAND21XL U1238 ( .B(memaddr_c[0]), .A(n121), .Y(n120) );
  AO2222XL U1239 ( .A(n234), .B(memaddr[3]), .C(sfr_psofs[3]), .D(n233), .E(
        memaddr_c[3]), .F(n414), .G(pre_1_adr[3]), .H(n2), .Y(N857) );
  XNOR2XL U1240 ( .A(memaddr_c[3]), .B(n682), .Y(n717) );
  NAND21XL U1241 ( .B(n156), .A(memaddr_c[3]), .Y(n209) );
  OAI22XL U1242 ( .A(memaddr_c[2]), .B(n151), .C(memaddr_c[3]), .D(n150), .Y(
        n152) );
  NAND21XL U1243 ( .B(c_adr[3]), .A(memaddr_c[3]), .Y(n873) );
  AO2222XL U1244 ( .A(n12), .B(memaddr[1]), .C(sfr_psofs[1]), .D(n9), .E(
        memaddr_c[1]), .F(n414), .G(pre_1_adr[1]), .H(n236), .Y(N855) );
  XOR3XL U1245 ( .A(memaddr_c[1]), .B(n107), .C(n118), .Y(n128) );
  GEN2XL U1246 ( .D(memaddr_c[1]), .E(n880), .C(n879), .B(n878), .A(n884), .Y(
        n881) );
  OA22XL U1247 ( .A(memaddr_c[1]), .B(n880), .C(memaddr_c[0]), .D(n877), .Y(
        n879) );
endmodule


module ictlr_a0_DW01_inc_2 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module ictlr_a0_DW01_inc_1 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  HAD1XL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1XL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  XOR2X1 U1 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  INVXL U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mcu51_a0 ( bclki2c, pc_ini, slp2wakeup, r_hold_mcu, wdt_slow, wdtov, 
        mdubsy, cs_run, t0_intr, clki2c, clkmdu, clkur0, clktm0, clktm1, 
        clkwdt, i2c_autoack, i2c_con_ens1, clkcpu, clkper, reset, ro, port0i, 
        exint_9, exint, clkcpuen, clkperen, port0o, port0ff, rxd0o, txd0, 
        rxd0i, rxd0oe, scli, sdai, sclo, sdao, waitstaten, mempsack, memack, 
        memdatai, memdatao, memaddr, mempswr, mempsrd, memwr, memrd, 
        memdatao_comb, memaddr_comb, mempswr_comb, mempsrd_comb, memwr_comb, 
        memrd_comb, ramdatai, ramdatao, ramaddr, ramwe, ramoe, dbgpo, sfrack, 
        sfrdatai, sfrdatao, sfraddr, sfrwe, sfroe, esfrm_wrdata, esfrm_addr, 
        esfrm_we, esfrm_oe, esfrm_rddata, test_si2, test_si1, test_so1, 
        test_se );
  input [15:0] pc_ini;
  output [1:0] wdtov;
  input [7:0] port0i;
  input [7:0] exint;
  output [7:0] port0o;
  output [7:0] port0ff;
  input [7:0] memdatai;
  output [7:0] memdatao;
  output [15:0] memaddr;
  output [7:0] memdatao_comb;
  output [15:0] memaddr_comb;
  input [7:0] ramdatai;
  output [7:0] ramdatao;
  output [7:0] ramaddr;
  output [31:0] dbgpo;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  output [6:0] sfraddr;
  input [7:0] esfrm_wrdata;
  input [6:0] esfrm_addr;
  output [7:0] esfrm_rddata;
  input bclki2c, slp2wakeup, r_hold_mcu, wdt_slow, clki2c, clkmdu, clkur0,
         clktm0, clktm1, clkwdt, i2c_autoack, clkcpu, clkper, reset, exint_9,
         rxd0i, scli, sdai, mempsack, memack, sfrack, esfrm_we, esfrm_oe,
         test_si2, test_si1, test_se;
  output mdubsy, cs_run, t0_intr, i2c_con_ens1, ro, clkcpuen, clkperen, rxd0o,
         txd0, rxd0oe, sclo, sdao, waitstaten, mempswr, mempsrd, memwr, memrd,
         mempswr_comb, mempsrd_comb, memwr_comb, memrd_comb, ramwe, ramoe,
         sfrwe, sfroe, test_so1;
  wire   n143, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, t0_tf1, t1_tf1, t0_tr1, t1_tr1, stop_flag, idle_flag, sfroe_s,
         sfroe_mcu51_per, sfrwe_s, sfrwe_mcu51_per, newinstr, intcall_int,
         cpu_resume, rmwinstr, pmw, p2sel, gf0, c, ac, ov, f0, f1, p, rsttowdt,
         rsttosrst, rst, int0ff, int1ff, rxd0ff, sdaiff, rsttowdtff,
         rsttosrstff, resetff, smod, ip0wdts, wdt_tm, bd, ie0, it0, ie1, it1,
         iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9, isr_tm, i2c_int,
         i2ccon_o_7, tf1_gate, riti0_gate, iex7_gate, iex2_gate, srstflag,
         int_vect_8b, int_vect_93, int_vect_9b, int_vect_a3, wdts, srst,
         pmuintreq_rev, pmuintreq, t1ov, t0ack, t1ack, isr_irq, int0ack,
         int1ack, iex7ack, iex2ack, iex3ack, iex4ack, iex5ack, iex6ack,
         iex8ack, iex9ack, n11, n144, n145, n142, n141, n140, n139, n138, n137,
         n136, n135, n134, n79, n80, n122, n112, n130, n131, n133, n3, n7, n8,
         n9, n10, n12, n1, n2, n4, n5, n6, n13, n14, n15, n16, n18, n19, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n38,
         n39, n40, n41, n42, n43, n54, n55, n56, n57, n58, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n70, n71, n73, n74, n75, n77, n78, n81, n90,
         n91, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5;
  wire   [13:0] timer_1ms;
  wire   [5:0] ien2;
  wire   [6:0] ramsfraddr;
  wire   [4:0] intvect_int;
  wire   [7:0] ckcon;
  wire   [7:0] dph;
  wire   [7:0] dpl;
  wire   [3:0] dps;
  wire   [7:0] p2;
  wire   [5:0] dpc;
  wire   [7:0] sp;
  wire   [7:0] acc_s;
  wire   [7:0] b;
  wire   [1:0] rs;
  wire   [7:0] arcon;
  wire   [7:0] md0;
  wire   [7:0] md1;
  wire   [7:0] md2;
  wire   [7:0] md3;
  wire   [7:0] md4;
  wire   [7:0] md5;
  wire   [3:0] t0_tmod;
  wire   [7:0] tl0;
  wire   [7:0] th0;
  wire   [3:0] t1_tmod;
  wire   [7:0] tl1;
  wire   [7:0] th1;
  wire   [7:0] wdtrel;
  wire   [6:5] t2con;
  wire   [7:0] s0con;
  wire   [7:0] s0buf;
  wire   [7:0] s0rell;
  wire   [7:0] s0relh;
  wire   [7:0] ien0;
  wire   [5:0] ien1;
  wire   [5:0] ip0;
  wire   [5:0] ip1;
  wire   [7:0] i2cdat_o;
  wire   [7:0] i2cadr_o;
  wire   [5:0] i2ccon_o;
  wire   [7:0] i2csta_o;
  wire   [3:0] isreg;

  INVX1 U52 ( .A(n80), .Y(n79) );
  INVX1 U53 ( .A(reset), .Y(n80) );
  INVX8 U50 ( .A(n80), .Y(n3) );
  mcu51_cpu_a0 u_cpu ( .clkcpu(clkcpu), .rst(n92), .mempsack(mempsack), 
        .memack(memack), .memdatai(memdatai), .memaddr(memaddr), .mempsrd(
        mempsrd), .mempswr(mempswr), .memrd(memrd), .memwr(memwr), 
        .memaddr_comb(memaddr_comb), .mempsrd_comb(mempsrd_comb), 
        .mempswr_comb(mempswr_comb), .memrd_comb(memrd_comb), .memwr_comb(
        memwr_comb), .cpu_hold(r_hold_mcu), .cpu_resume(cpu_resume), .irq(
        dbgpo[20]), .intvect(intvect_int), .intcall(intcall_int), .retiinstr(
        dbgpo[21]), .newinstr(newinstr), .rmwinstr(rmwinstr), .waitstaten(
        waitstaten), .ramdatai(ramdatai), .sfrdatai({esfrm_rddata[7:3], n143, 
        n144, n145}), .ramsfraddr({SYNOPSYS_UNCONNECTED_1, ramsfraddr}), 
        .ramdatao(memdatao), .ramoe(), .ramwe(), .sfroe(sfroe_s), .sfrwe(
        sfrwe_s), .sfroe_r(), .sfrwe_r(), .sfroe_comb_s(), .sfrwe_comb_s(), 
        .pc_o(dbgpo[15:0]), .pc_ini(pc_ini), .cs_run(cs_run), .instr(
        dbgpo[31:24]), .codefetch_s(), .sfrack(sfrack), .ramsfraddr_comb(
        ramaddr), .ramdatao_comb(ramdatao), .ramoe_comb(ramoe), .ramwe_comb(
        ramwe), .ckcon(ckcon), .pmw(pmw), .p2sel(p2sel), .gf0(gf0), .stop(
        stop_flag), .idle(idle_flag), .acc(acc_s), .b(b), .rs(rs), .c(c), .ac(
        ac), .ov(ov), .p(p), .f0(f0), .f1(f1), .dph(dph), .dpl(dpl), .dps(dps), 
        .dpc(dpc), .p2(p2), .sp(sp), .test_si(timer_1ms[13]), .test_so(n133), 
        .test_se(test_se) );
  syncneg_a0 u_syncneg ( .clk(clkper), .reset(n79), .rsttowdt(rsttowdt), 
        .rsttosrst(rsttosrst), .rst(rst), .int0(exint[0]), .int1(exint[1]), 
        .port0i(port0i), .rxd0i(rxd0i), .sdai(sdai), .int0ff(int0ff), .int1ff(
        int1ff), .port0ff(port0ff), .t0ff(), .t1ff(), .rxd0ff(rxd0ff), 
        .sdaiff(sdaiff), .rsttowdtff(rsttowdtff), .rsttosrstff(rsttosrstff), 
        .rstff(n122), .resetff(resetff), .test_si(srstflag), .test_se(test_se)
         );
  sfrmux_a0 u_sfrmux ( .isfrwait(n13), .sfraddr({sfraddr[6], n62, n43, n70, 
        n42, n29, n65}), .c(c), .ac(ac), .f0(f0), .rs(rs), .ov(ov), .f1(f1), 
        .p(p), .acc(acc_s), .b(b), .dpl(dpl), .dph(dph), .dps(dps), .dpc(dpc), 
        .p2(p2), .sp(sp), .smod(smod), .pmw(pmw), .p2sel(p2sel), .gf0(gf0), 
        .stop(stop_flag), .idle(idle_flag), .ckcon(ckcon), .port0(port0o), 
        .port0ff(port0ff), .rmwinstr(rmwinstr), .arcon(arcon), .md0(md0), 
        .md1(md1), .md2(md2), .md3(md3), .md4(md4), .md5(md5), .t0_tmod(
        t0_tmod), .t0_tf0(dbgpo[17]), .t0_tf1(t0_tf1), .t0_tr0(dbgpo[16]), 
        .t0_tr1(t0_tr1), .tl0(tl0), .th0(th0), .t1_tmod(t1_tmod), .t1_tf1(
        t1_tf1), .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1), .wdtrel(wdtrel), 
        .ip0wdts(ip0wdts), .wdt_tm(wdt_tm), .t2con({1'b0, t2con, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .s0con(s0con), .s0buf(s0buf), .s0rell(s0rell), 
        .s0relh(s0relh), .bd(bd), .ie0(ie0), .it0(it0), .ie1(ie1), .it1(it1), 
        .iex2(iex2), .iex3(iex3), .iex4(iex4), .iex5(iex5), .iex6(iex6), 
        .iex7(iex7), .iex8(iex8), .iex9(iex9), .iex10(1'b0), .iex11(1'b0), 
        .iex12(1'b0), .ien0({ien0[7], 1'b0, ien0[5:0]}), .ien1(ien1), .ien2(
        ien2), .ip0(ip0), .ip1(ip1), .isr_tm(isr_tm), .i2c_int(i2c_int), 
        .i2cdat_o(i2cdat_o), .i2cadr_o(i2cadr_o), .i2ccon_o({i2ccon_o_7, 
        i2c_con_ens1, i2ccon_o}), .i2csta_o({i2csta_o[7:3], 1'b0, 1'b0, 1'b0}), 
        .sfrdatai(sfrdatai), .tf1_gate(tf1_gate), .riti0_gate(riti0_gate), 
        .iex7_gate(iex7_gate), .iex2_gate(iex2_gate), .srstflag(srstflag), 
        .int_vect_8b(int_vect_8b), .int_vect_93(int_vect_93), .int_vect_9b(
        int_vect_9b), .int_vect_a3(int_vect_a3), .ext_sfr_sel(), .sfrdatao({
        esfrm_rddata[7:3], n143, n144, n145}) );
  pmurstctrl_a0 u_pmurstctrl ( .resetff(resetff), .wdts(wdts), .srst(srst), 
        .pmuintreq(pmuintreq_rev), .stop(stop_flag), .idle(idle_flag), 
        .clkcpu_en(clkcpuen), .clkper_en(clkperen), .cpu_resume(cpu_resume), 
        .rsttowdt(rsttowdt), .rsttosrst(rsttosrst), .rst(rst) );
  wakeupctrl_a0 u_wakeupctrl ( .irq(dbgpo[20]), .int0ff(exint[0]), .int1ff(
        exint[1]), .it0(it0), .it1(it1), .isreg(isreg), .intprior0({ip0[2], 
        ip0[0]}), .intprior1({ip1[2], ip1[0]}), .eal(ien0[7]), .eint0(ien0[0]), 
        .eint1(ien0[2]), .pmuintreq(pmuintreq) );
  mdu_a0 u_mdu ( .clkper(clkmdu), .rst(ro), .mdubsy(mdubsy), .sfrdatai({
        sfrdatao[7], n135, n136, sfrdatao[4:0]}), .sfraddr({n60, n75, n73, n71, 
        n1, n5, n68}), .sfrwe(n40), .sfroe(sfroe_mcu51_per), .arcon(arcon), 
        .md0(md0), .md1(md1), .md2(md2), .md3(md3), .md4(md4), .md5(md5), 
        .test_si(isr_tm), .test_so(n130), .test_se(test_se) );
  ports_a0 u_ports ( .clkper(clkper), .rst(dbgpo[22]), .port0(port0o), 
        .sfrdatai({sfrdatao[7], n135, sfrdatao[5], n137, n138, sfrdatao[2], 
        n140, sfrdatao[0]}), .sfraddr({n81, n75, n73, n26, n56, n5, sfraddr[0]}), .sfrwe(sfrwe_mcu51_per), .test_si(n130), .test_se(test_se) );
  serial0_a0 u_serial0 ( .t_shift_clk(), .r_shift_clk(), .clkper(clkur0), 
        .rst(n92), .newinstr(newinstr), .rxd0ff(rxd0ff), .t1ov(t1ov), .rxd0o(
        rxd0o), .rxd0oe(rxd0oe), .txd0(txd0), .sfrdatai({n134, sfrdatao[6], 
        n136, sfrdatao[4:3], n139, sfrdatao[1], n141}), .sfraddr({n81, n77, 
        sfraddr[4], n26, n56, n5, n67}), .sfrwe(n41), .s0con(s0con), .s0buf(
        s0buf), .s0rell(s0rell), .s0relh(s0relh), .smod(smod), .bd(bd), 
        .test_si(port0o[7]), .test_se(test_se) );
  timer0_a0 u_timer0 ( .clkper(clktm0), .rst(n90), .newinstr(newinstr), .t0ff(
        1'b0), .t0ack(t0ack), .t1ack(t1ack), .int0ff(int0ff), .t0_tf0(
        dbgpo[17]), .t0_tf1(t0_tf1), .sfrdatai({sfrdatao[7:1], n141}), 
        .sfraddr({n81, n75, n73, n71, sfraddr[2], n4, n68}), .sfrwe(n41), 
        .t0_tmod(t0_tmod), .t0_tr0(dbgpo[16]), .t0_tr1(t0_tr1), .tl0(tl0), 
        .th0(th0), .test_si(sdaiff), .test_se(test_se) );
  timer1_a0 u_timer1 ( .clkper(clktm1), .rst(ro), .newinstr(newinstr), .t1ff(
        1'b0), .t1ack(t1ack), .int1ff(int1ff), .t1_tf1(t1_tf1), .t1ov(t1ov), 
        .sfrdatai({n134, sfrdatao[6], n136, sfrdatao[4:3], n139, sfrdatao[1], 
        n141}), .sfraddr({n60, n75, n73, n71, n1, n4, n66}), .sfrwe(n40), 
        .t1_tmod(t1_tmod), .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1), .test_si(
        tl0[7]), .test_se(test_se) );
  watchdog_a0 u_watchdog ( .wdt_slow(wdt_slow), .clkwdt(clkwdt), .clkper(
        clkper), .resetff(rsttowdtff), .newinstr(newinstr), .wdts_s(wdtov), 
        .wdts(wdts), .ip0wdts(ip0wdts), .wdt_tm(wdt_tm), .sfrdatai({
        sfrdatao[7:5], n137, n138, sfrdatao[2], n140, sfrdatao[0]}), .sfraddr(
        {n81, n77, n73, n71, sfraddr[2:1], n68}), .sfrwe(sfrwe_mcu51_per), 
        .wdtrel(wdtrel), .test_si(tl1[7]), .test_se(test_se) );
  isr_a0 u_isr ( .clkper(clkper), .rst(n91), .intcall(intcall_int), 
        .retiinstr(dbgpo[21]), .int_vect_03(ie0), .int_vect_0b(dbgpo[17]), 
        .t0ff(1'b0), .int_vect_13(ie1), .int_vect_1b(tf1_gate), .t1ff(1'b0), 
        .int_vect_23(riti0_gate), .i2c_int(i2c_int), .rxd0ff(rxd0ff), 
        .int_vect_43(iex7_gate), .sdaiff(sdaiff), .int_vect_4b(iex2_gate), 
        .int_vect_53(iex3), .int_vect_5b(iex4), .int_vect_63(iex5), 
        .int_vect_6b(iex6), .int_vect_8b(int_vect_8b), .int_vect_93(
        int_vect_93), .int_vect_9b(int_vect_9b), .int_vect_a3(int_vect_a3), 
        .int_vect_ab(1'b0), .irq(isr_irq), .intvect(intvect_int), .int_ack_03(
        int0ack), .int_ack_0b(t0ack), .int_ack_13(int1ack), .int_ack_1b(t1ack), 
        .int_ack_43(iex7ack), .int_ack_4b(iex2ack), .int_ack_53(iex3ack), 
        .int_ack_5b(iex4ack), .int_ack_63(iex5ack), .int_ack_6b(iex6ack), 
        .int_ack_8b(iex8ack), .int_ack_93(iex9ack), .int_ack_9b(), 
        .int_ack_a3(), .int_ack_ab(), .is_reg(isreg), .ip0(ip0), .ip1(ip1), 
        .ien0({ien0[7], SYNOPSYS_UNCONNECTED_2, ien0[5:0]}), .ien1(ien1), 
        .ien2(ien2), .isr_tm(isr_tm), .sfraddr({n81, n75, n24, n26, n56, n2, 
        n67}), .sfrdatai({sfrdatao[7], n135, sfrdatao[5], n137, sfrdatao[3:0]}), .sfrwe(n41), .test_si(n131), .test_se(test_se) );
  extint_a0 u_extint ( .clkper(clkper), .rst(ro), .newinstr(newinstr), 
        .int0ff(int0ff), .int0ack(int0ack), .int1ff(int1ff), .int1ack(int1ack), 
        .int2ff(exint[2]), .iex2ack(iex2ack), .int3ff(exint[3]), .iex3ack(
        iex3ack), .int4ff(exint[4]), .iex4ack(iex4ack), .int5ff(exint[5]), 
        .iex5ack(iex5ack), .int6ff(exint[6]), .iex6ack(iex6ack), .int7ff(
        exint[7]), .iex7ack(iex7ack), .int8ff(n11), .iex8ack(iex8ack), 
        .int9ff(exint_9), .iex9ack(iex9ack), .ie0(ie0), .it0(it0), .ie1(ie1), 
        .it1(it1), .i2fr(t2con[5]), .iex2(iex2), .i3fr(t2con[6]), .iex3(iex3), 
        .iex4(iex4), .iex5(iex5), .iex6(iex6), .iex7(iex7), .iex8(iex8), 
        .iex9(iex9), .iex10(), .iex11(), .iex12(), .sfraddr({n60, n77, 
        sfraddr[4], n71, n1, n2, n66}), .sfrdatai({sfrdatao[7], n135, n136, 
        n137, sfrdatao[3], n139, n140, n141}), .sfrwe(n41), .test_si(n133), 
        .test_se(test_se) );
  i2c_a0 u_i2c ( .clk(clki2c), .rst(n90), .bclksel(bclki2c), .scli(scli), 
        .sdai(sdai), .sclo(sclo), .sdao(sdao), .intack(i2c_autoack), .si(
        i2c_int), .sfrwe(n40), .sfraddr({n81, n75, n73, n71, n56, n2, n68}), 
        .sfrdatai({sfrdatao[7], n135, sfrdatao[5:4], n138, n139, n140, 
        sfrdatao[0]}), .i2cdat_o(i2cdat_o), .i2cadr_o(i2cadr_o), .i2ccon_o({
        i2ccon_o_7, i2c_con_ens1, i2ccon_o}), .i2csta_o({i2csta_o[7:3], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5}), .test_si2(test_si2), .test_si1(it1), .test_so2(n131), .test_so1(test_so1), 
        .test_se(test_se) );
  softrstctrl_a0 u_softrstctrl ( .clkcpu(clkcpu), .resetff(rsttosrstff), 
        .newinstr(newinstr), .srstreq(srst), .srstflag(srstflag), .sfrdatai({
        sfrdatao[7], n135, sfrdatao[5], n137, n138, sfrdatao[2], n140, 
        sfrdatao[0]}), .sfraddr({n60, n75, n73, n26, n56, n4, n68}), .sfrwe(
        n41), .test_si(txd0), .test_se(test_se) );
  mcu51_a0_DW01_inc_0 add_268 ( .A(timer_1ms), .SUM({N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7}) );
  SDFFQX1 timer_1ms_reg_9_ ( .D(N30), .SIN(timer_1ms[8]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[9]) );
  SDFFQX1 timer_1ms_reg_13_ ( .D(N34), .SIN(timer_1ms[12]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[13]) );
  SDFFQX1 timer_1ms_reg_12_ ( .D(N33), .SIN(timer_1ms[11]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[12]) );
  SDFFQX1 timer_1ms_reg_8_ ( .D(N29), .SIN(timer_1ms[7]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[8]) );
  SDFFQX1 timer_1ms_reg_10_ ( .D(N31), .SIN(timer_1ms[9]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[10]) );
  SDFFQX1 timer_1ms_reg_6_ ( .D(N27), .SIN(timer_1ms[5]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[6]) );
  SDFFQX1 timer_1ms_reg_11_ ( .D(N32), .SIN(timer_1ms[10]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[11]) );
  SDFFQX1 timer_1ms_reg_7_ ( .D(N28), .SIN(timer_1ms[6]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[7]) );
  SDFFQX1 timer_1ms_reg_5_ ( .D(N26), .SIN(timer_1ms[4]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[5]) );
  SDFFQX1 timer_1ms_reg_4_ ( .D(N25), .SIN(timer_1ms[3]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[4]) );
  SDFFQX1 timer_1ms_reg_3_ ( .D(N24), .SIN(timer_1ms[2]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[3]) );
  SDFFQX1 timer_1ms_reg_2_ ( .D(N23), .SIN(timer_1ms[1]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[2]) );
  SDFFQX1 timer_1ms_reg_1_ ( .D(N22), .SIN(timer_1ms[0]), .SMC(test_se), .C(
        clkper), .Q(timer_1ms[1]) );
  SDFFQX1 timer_1ms_reg_0_ ( .D(N21), .SIN(test_si1), .SMC(test_se), .C(clkper), .Q(timer_1ms[0]) );
  MUX2IX2 U3 ( .D0(ramsfraddr[0]), .D1(esfrm_addr[0]), .S(n112), .Y(n61) );
  INVX2 U4 ( .A(n112), .Y(n19) );
  INVX4 U5 ( .A(esfrm_we), .Y(n118) );
  INVX6 U6 ( .A(n78), .Y(sfraddr[5]) );
  NAND21X2 U7 ( .B(esfrm_oe), .A(n118), .Y(n23) );
  INVX6 U8 ( .A(n98), .Y(n62) );
  MUX2IX4 U9 ( .D0(ramsfraddr[5]), .D1(esfrm_addr[5]), .S(n23), .Y(n98) );
  BUFX3 U10 ( .A(n142), .Y(n29) );
  INVX6 U11 ( .A(n35), .Y(sfraddr[6]) );
  AND2X1 U12 ( .A(ramsfraddr[6]), .B(n99), .Y(n25) );
  INVX2 U13 ( .A(esfrm_oe), .Y(n99) );
  INVX1 U14 ( .A(ramsfraddr[4]), .Y(n28) );
  INVX4 U15 ( .A(n62), .Y(n78) );
  INVX1 U16 ( .A(n99), .Y(n18) );
  INVX2 U17 ( .A(n55), .Y(sfraddr[1]) );
  INVX1 U18 ( .A(n118), .Y(n6) );
  INVX1 U19 ( .A(n14), .Y(sfraddr[0]) );
  INVXL U20 ( .A(n57), .Y(n1) );
  INVXL U21 ( .A(n54), .Y(n2) );
  INVXL U22 ( .A(n54), .Y(n4) );
  INVXL U23 ( .A(n54), .Y(n5) );
  MUX2X2 U24 ( .D0(ramsfraddr[2]), .D1(esfrm_addr[2]), .S(n22), .Y(n42) );
  INVX3 U25 ( .A(n58), .Y(n70) );
  BUFXL U26 ( .A(n22), .Y(n13) );
  INVXL U27 ( .A(esfrm_addr[4]), .Y(n27) );
  INVXL U28 ( .A(n65), .Y(n14) );
  INVX3 U29 ( .A(n61), .Y(n65) );
  NAND2X1 U30 ( .A(esfrm_addr[6]), .B(n18), .Y(n30) );
  NAND2X1 U31 ( .A(esfrm_addr[6]), .B(n6), .Y(n32) );
  NAND21X2 U32 ( .B(esfrm_oe), .A(n118), .Y(n22) );
  NAND21X2 U33 ( .B(esfrm_oe), .A(n118), .Y(n112) );
  BUFXL U34 ( .A(n35), .Y(n15) );
  INVXL U35 ( .A(sfraddr[0]), .Y(n16) );
  MUX2IX2 U36 ( .D0(ramsfraddr[1]), .D1(esfrm_addr[1]), .S(n22), .Y(n97) );
  BUFXL U37 ( .A(n70), .Y(sfraddr[3]) );
  NAND2X1 U38 ( .A(n118), .B(n25), .Y(n31) );
  BUFXL U39 ( .A(n42), .Y(sfraddr[2]) );
  MUX2IX2 U40 ( .D0(n28), .D1(n27), .S(n23), .Y(n43) );
  INVX1 U41 ( .A(n26), .Y(n21) );
  BUFXL U42 ( .A(n43), .Y(n24) );
  MUX2IX2 U43 ( .D0(esfrm_addr[3]), .D1(ramsfraddr[3]), .S(n19), .Y(n58) );
  BUFXL U44 ( .A(sfraddr[3]), .Y(n26) );
  INVXL U45 ( .A(n78), .Y(n75) );
  INVXL U46 ( .A(n78), .Y(n77) );
  INVXL U47 ( .A(sfraddr[1]), .Y(n54) );
  INVXL U48 ( .A(n15), .Y(n81) );
  AND3X4 U49 ( .A(n31), .B(n30), .C(n32), .Y(n35) );
  BUFXL U51 ( .A(n144), .Y(esfrm_rddata[1]) );
  INVXL U54 ( .A(sfraddr[2]), .Y(n57) );
  BUFXL U55 ( .A(n118), .Y(n34) );
  INVX3 U56 ( .A(n97), .Y(n142) );
  INVX1 U57 ( .A(n142), .Y(n55) );
  BUFXL U58 ( .A(n145), .Y(esfrm_rddata[0]) );
  BUFXL U59 ( .A(n143), .Y(esfrm_rddata[2]) );
  INVXL U60 ( .A(n13), .Y(n38) );
  INVX1 U61 ( .A(sfrwe_mcu51_per), .Y(n39) );
  INVX1 U62 ( .A(n39), .Y(n40) );
  INVX1 U63 ( .A(n39), .Y(n41) );
  INVXL U64 ( .A(n74), .Y(n73) );
  INVXL U65 ( .A(n57), .Y(n56) );
  INVXL U66 ( .A(n74), .Y(sfraddr[4]) );
  INVXL U67 ( .A(n24), .Y(n74) );
  INVXL U68 ( .A(memdatao[0]), .Y(n115) );
  INVXL U69 ( .A(memdatao[1]), .Y(n113) );
  INVXL U70 ( .A(memdatao[2]), .Y(n110) );
  BUFX3 U71 ( .A(ramdatao[2]), .Y(memdatao_comb[2]) );
  BUFX3 U72 ( .A(ramdatao[4]), .Y(memdatao_comb[4]) );
  BUFX3 U73 ( .A(ramdatao[5]), .Y(memdatao_comb[5]) );
  BUFX3 U74 ( .A(ramdatao[6]), .Y(memdatao_comb[6]) );
  BUFX3 U75 ( .A(ramdatao[7]), .Y(memdatao_comb[7]) );
  INVX1 U76 ( .A(n95), .Y(ro) );
  INVX1 U77 ( .A(n107), .Y(sfrdatao[4]) );
  INVX1 U78 ( .A(n109), .Y(sfrdatao[3]) );
  INVX1 U79 ( .A(n116), .Y(sfrdatao[0]) );
  INVX1 U80 ( .A(n95), .Y(dbgpo[22]) );
  INVX1 U81 ( .A(n101), .Y(sfrdatao[7]) );
  INVX1 U82 ( .A(n103), .Y(sfrdatao[6]) );
  INVX1 U83 ( .A(n114), .Y(sfrdatao[1]) );
  INVX1 U84 ( .A(n105), .Y(sfrdatao[5]) );
  INVX1 U85 ( .A(n111), .Y(sfrdatao[2]) );
  NAND21XL U86 ( .B(n18), .A(n121), .Y(sfroe_mcu51_per) );
  INVXL U87 ( .A(n21), .Y(n71) );
  NOR21XL U88 ( .B(N19), .A(n63), .Y(N33) );
  INVX1 U89 ( .A(n95), .Y(n92) );
  INVX1 U90 ( .A(n96), .Y(n90) );
  NOR21XL U91 ( .B(N18), .A(n64), .Y(N32) );
  NOR21XL U92 ( .B(N17), .A(n63), .Y(N31) );
  NOR21XL U93 ( .B(N16), .A(n64), .Y(N30) );
  INVX1 U94 ( .A(n96), .Y(n91) );
  NOR21XL U95 ( .B(N8), .A(n64), .Y(N22) );
  NOR21XL U96 ( .B(N9), .A(n63), .Y(N23) );
  NOR21XL U97 ( .B(N10), .A(n64), .Y(N24) );
  NOR21XL U98 ( .B(N11), .A(n63), .Y(N25) );
  NOR21XL U99 ( .B(N14), .A(n64), .Y(N28) );
  NOR21XL U100 ( .B(N13), .A(n63), .Y(N27) );
  NOR21XL U101 ( .B(N12), .A(n64), .Y(N26) );
  NOR21XL U102 ( .B(N15), .A(n63), .Y(N29) );
  BUFX3 U103 ( .A(n7), .Y(n63) );
  BUFX3 U104 ( .A(n7), .Y(n64) );
  BUFX3 U105 ( .A(ramdatao[0]), .Y(memdatao_comb[0]) );
  BUFX3 U106 ( .A(ramdatao[1]), .Y(memdatao_comb[1]) );
  BUFX3 U107 ( .A(ramdatao[3]), .Y(memdatao_comb[3]) );
  BUFX3 U108 ( .A(rxd0i), .Y(dbgpo[23]) );
  INVX1 U109 ( .A(n117), .Y(n120) );
  OR2X1 U110 ( .A(pmuintreq), .B(slp2wakeup), .Y(pmuintreq_rev) );
  INVX1 U111 ( .A(n122), .Y(n95) );
  INVX1 U112 ( .A(n107), .Y(n137) );
  INVXL U113 ( .A(memdatao[4]), .Y(n106) );
  INVX1 U114 ( .A(n109), .Y(n138) );
  INVXL U115 ( .A(memdatao[3]), .Y(n108) );
  INVX1 U116 ( .A(n116), .Y(n141) );
  NOR21XL U117 ( .B(isr_irq), .A(r_hold_mcu), .Y(dbgpo[20]) );
  OR2X1 U118 ( .A(t0_tf1), .B(t1_tf1), .Y(dbgpo[19]) );
  OR2X1 U119 ( .A(t0_tr1), .B(t1_tr1), .Y(dbgpo[18]) );
  INVX1 U120 ( .A(n101), .Y(n134) );
  INVX1 U121 ( .A(memdatao[7]), .Y(n100) );
  INVX1 U122 ( .A(n114), .Y(n140) );
  INVX1 U123 ( .A(n105), .Y(n136) );
  INVX1 U124 ( .A(memdatao[5]), .Y(n104) );
  INVX1 U125 ( .A(n103), .Y(n135) );
  INVX1 U126 ( .A(memdatao[6]), .Y(n102) );
  INVX1 U127 ( .A(n111), .Y(n139) );
  AO21XL U128 ( .B(sfroe_s), .C(n119), .A(n18), .Y(sfroe) );
  INVX1 U129 ( .A(sfroe_s), .Y(n121) );
  NOR21XL U130 ( .B(N20), .A(n64), .Y(N34) );
  INVX1 U131 ( .A(n122), .Y(n96) );
  NAND32X1 U132 ( .B(n11), .C(n3), .A(ien2[1]), .Y(n7) );
  NOR21XL U133 ( .B(N7), .A(n63), .Y(N21) );
  NAND43X1 U134 ( .B(timer_1ms[8]), .C(timer_1ms[5]), .D(timer_1ms[12]), .A(
        timer_1ms[0]), .Y(n10) );
  NOR4XL U135 ( .A(n8), .B(n9), .C(n10), .D(n12), .Y(n11) );
  NAND4X1 U136 ( .A(timer_1ms[4]), .B(timer_1ms[3]), .C(timer_1ms[2]), .D(
        timer_1ms[1]), .Y(n8) );
  NAND3X1 U137 ( .A(timer_1ms[7]), .B(timer_1ms[6]), .C(timer_1ms[9]), .Y(n9)
         );
  NAND3X1 U138 ( .A(timer_1ms[11]), .B(timer_1ms[10]), .C(timer_1ms[13]), .Y(
        n12) );
  AND2X1 U139 ( .A(ien0[0]), .B(dbgpo[17]), .Y(t0_intr) );
  INVXL U140 ( .A(n15), .Y(n60) );
  INVXL U141 ( .A(n16), .Y(n68) );
  INVXL U142 ( .A(n16), .Y(n67) );
  INVXL U143 ( .A(n16), .Y(n66) );
  MUX2AXL U153 ( .D0(esfrm_wrdata[6]), .D1(n102), .S(n38), .Y(n103) );
  MUX2AXL U154 ( .D0(esfrm_wrdata[2]), .D1(n110), .S(n38), .Y(n111) );
  MUX2AXL U155 ( .D0(esfrm_wrdata[5]), .D1(n104), .S(n38), .Y(n105) );
  MUX2AXL U156 ( .D0(esfrm_wrdata[7]), .D1(n100), .S(n38), .Y(n101) );
  MUX2AXL U157 ( .D0(esfrm_wrdata[1]), .D1(n113), .S(n38), .Y(n114) );
  MUX2AXL U158 ( .D0(esfrm_wrdata[4]), .D1(n106), .S(n38), .Y(n107) );
  MUX2AXL U159 ( .D0(esfrm_wrdata[3]), .D1(n108), .S(n38), .Y(n109) );
  MUX2AXL U160 ( .D0(esfrm_wrdata[0]), .D1(n115), .S(n38), .Y(n116) );
  NAND21XL U161 ( .B(n13), .A(sfrwe_s), .Y(n117) );
  AO21XL U162 ( .B(n120), .C(n119), .A(n6), .Y(sfrwe) );
  NAND21XL U163 ( .B(n120), .A(n34), .Y(sfrwe_mcu51_per) );
  INVX8 U164 ( .A(n3), .Y(n119) );
endmodule


module mcu51_a0_DW01_inc_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;

  wire   [13:2] carry;

  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module softrstctrl_a0 ( clkcpu, resetff, newinstr, srstreq, srstflag, sfrdatai, 
        sfraddr, sfrwe, test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkcpu, resetff, newinstr, sfrwe, test_si, test_se;
  output srstreq, srstflag;
  wire   srst_ff0, srst_ff1, N37, N38, N41, net11981, n24, n25, n26, n27, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n28, n29,
         n30, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [3:0] srst_count;

  SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 clk_gate_srst_count_reg ( .CLK(clkcpu), 
        .EN(N37), .ENCLK(net11981), .TE(test_se) );
  SDFFQX1 srst_ff1_reg ( .D(n24), .SIN(srst_ff0), .SMC(test_se), .C(clkcpu), 
        .Q(srst_ff1) );
  SDFFQX1 srst_count_reg_1_ ( .D(n6), .SIN(srst_count[0]), .SMC(test_se), .C(
        net11981), .Q(srst_count[1]) );
  SDFFQX1 srst_count_reg_3_ ( .D(N41), .SIN(srst_count[2]), .SMC(test_se), .C(
        net11981), .Q(srst_count[3]) );
  SDFFQX1 srst_ff0_reg ( .D(n26), .SIN(srst_count[3]), .SMC(test_se), .C(
        clkcpu), .Q(srst_ff0) );
  SDFFQX1 srst_count_reg_0_ ( .D(N38), .SIN(test_si), .SMC(test_se), .C(
        net11981), .Q(srst_count[0]) );
  SDFFQX1 srst_count_reg_2_ ( .D(n4), .SIN(srst_count[1]), .SMC(test_se), .C(
        net11981), .Q(srst_count[2]) );
  SDFFQX1 srst_r_reg ( .D(n27), .SIN(srst_ff1), .SMC(test_se), .C(clkcpu), .Q(
        srstreq) );
  SDFFQX1 srstflag_reg ( .D(n25), .SIN(srstreq), .SMC(test_se), .C(clkcpu), 
        .Q(srstflag) );
  INVX1 U3 ( .A(n15), .Y(n2) );
  NAND42X1 U4 ( .C(sfraddr[3]), .D(n20), .A(sfraddr[0]), .B(n21), .Y(n15) );
  NAND2XL U5 ( .A(sfraddr[2]), .B(sfraddr[1]), .Y(n20) );
  AND4X1 U6 ( .A(sfrwe), .B(sfraddr[6]), .C(sfraddr[5]), .D(sfraddr[4]), .Y(
        n21) );
  NAND2X1 U7 ( .A(sfrdatai[0]), .B(n2), .Y(n12) );
  INVX1 U8 ( .A(newinstr), .Y(n3) );
  NOR2X1 U9 ( .A(n16), .B(n5), .Y(n22) );
  INVX1 U10 ( .A(n28), .Y(n5) );
  INVX1 U11 ( .A(n16), .Y(n9) );
  NAND2X1 U12 ( .A(n10), .B(n16), .Y(N37) );
  NOR2X1 U13 ( .A(resetff), .B(n18), .Y(n24) );
  AOI22AXL U14 ( .A(srst_ff0), .B(n2), .D(n19), .C(n8), .Y(n18) );
  AOI32X1 U15 ( .A(srst_ff1), .B(n3), .C(n15), .D(srst_ff0), .E(newinstr), .Y(
        n19) );
  NOR2X1 U16 ( .A(resetff), .B(n11), .Y(n27) );
  AOI32X1 U17 ( .A(n12), .B(n13), .C(srstreq), .D(srst_ff1), .E(n1), .Y(n11)
         );
  NAND3X1 U18 ( .A(srst_count[2]), .B(n5), .C(srst_count[3]), .Y(n13) );
  INVX1 U19 ( .A(n12), .Y(n1) );
  NAND2X1 U20 ( .A(n16), .B(n17), .Y(n25) );
  OAI211X1 U21 ( .C(sfrdatai[0]), .D(n15), .A(n10), .B(srstflag), .Y(n17) );
  AOI21X1 U22 ( .B(n12), .C(n14), .A(resetff), .Y(n26) );
  NAND4X1 U23 ( .A(srst_ff0), .B(n15), .C(n3), .D(n8), .Y(n14) );
  GEN2XL U24 ( .D(n9), .E(n7), .C(n22), .B(srst_count[3]), .A(n23), .Y(N41) );
  NOR4XL U25 ( .A(srst_count[3]), .B(n28), .C(n7), .D(n16), .Y(n23) );
  NAND2X1 U26 ( .A(srstreq), .B(n10), .Y(n16) );
  NAND2X1 U27 ( .A(srst_count[1]), .B(srst_count[0]), .Y(n28) );
  INVX1 U28 ( .A(resetff), .Y(n10) );
  INVX1 U29 ( .A(srst_count[2]), .Y(n7) );
  INVX1 U30 ( .A(srstreq), .Y(n8) );
  INVX1 U31 ( .A(n30), .Y(n6) );
  OAI211X1 U32 ( .C(srst_count[0]), .D(srst_count[1]), .A(n9), .B(n28), .Y(n30) );
  INVX1 U33 ( .A(n29), .Y(n4) );
  AOI32X1 U34 ( .A(n9), .B(n7), .C(n5), .D(srst_count[2]), .E(n22), .Y(n29) );
  NOR2X1 U35 ( .A(srst_count[0]), .B(n16), .Y(N38) );
endmodule


module SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2c_a0 ( clk, rst, bclksel, scli, sdai, sclo, sdao, intack, si, sfrwe, 
        sfraddr, sfrdatai, i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o, test_si2, 
        test_si1, test_so2, test_so1, test_se );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  output [7:0] i2cdat_o;
  output [7:0] i2cadr_o;
  output [7:0] i2ccon_o;
  output [7:0] i2csta_o;
  input clk, rst, bclksel, scli, sdai, intack, sfrwe, test_si2, test_si1,
         test_se;
  output sclo, sdao, si, test_so2, test_so1;
  wire   scli_ff, N180, sdai_ff, N181, sclo_int, adrcomp, adrcompen, nedetect,
         ack_bit, bsd7, pedetect, N225, N226, N227, N232, N233, N234, sclint,
         ack, sdaint, bsd7_tmp, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N332, N333, N335, N336, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N406, N407, N408, N409, N410, N412, N413, N414,
         N431, N432, N433, N468, N469, N470, N471, N491, N492, N493, N494,
         N495, busfree, N510, N511, rst_delay, clk_count1_ov, N653, N654, N655,
         N656, N657, clk_count2_ov, N685, N686, N687, N688, N689, N690, clkint,
         clkint_ff, N700, N746, N747, N748, N749, N1022, N1023, N1024, N1025,
         N1026, N1027, N1063, N1064, N1065, sclscl, starto_en, N1124, N1125,
         N1126, net12020, net12026, net12031, net12036, net12041, net12046,
         net12051, net12056, net12061, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n7,
         n8, n9, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n280, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452;
  wire   [2:0] fsmmod;
  wire   [4:0] fsmsta;
  wire   [3:0] framesync;
  wire   [2:0] fsmdet;
  wire   [2:0] setup_counter_r;
  wire   [2:0] scli_ff_reg0;
  wire   [2:0] sdai_ff_reg0;
  wire   [2:0] indelay;
  wire   [2:0] fsmsync;
  wire   [1:0] bclkcnt;
  wire   [3:0] clk_count1;
  wire   [3:0] clk_count2;

  SNPS_CLOCK_GATE_HIGH_i2c_a0_0 clk_gate_i2ccon_reg ( .CLK(clk), .EN(n28), 
        .ENCLK(net12020), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_8 clk_gate_i2cdat_reg ( .CLK(clk), .EN(N296), 
        .ENCLK(net12026), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_7 clk_gate_setup_counter_r_reg ( .CLK(clk), .EN(
        N332), .ENCLK(net12031), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_6 clk_gate_i2cadr_reg ( .CLK(clk), .EN(N342), 
        .ENCLK(net12036), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_5 clk_gate_indelay_reg ( .CLK(clk), .EN(N468), 
        .ENCLK(net12041), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_4 clk_gate_framesync_reg ( .CLK(clk), .EN(N491), 
        .ENCLK(net12046), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_3 clk_gate_clk_count1_reg ( .CLK(clk), .EN(N653), 
        .ENCLK(net12051), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_2 clk_gate_clk_count2_reg ( .CLK(clk), .EN(N689), 
        .ENCLK(net12056), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_1 clk_gate_fsmsta_reg ( .CLK(clk), .EN(N1022), 
        .ENCLK(net12061), .TE(test_se) );
  SDFFQX1 scli_ff_reg ( .D(N180), .SIN(rst_delay), .SMC(test_se), .C(clk), .Q(
        scli_ff) );
  SDFFQX1 sdai_ff_reg ( .D(N181), .SIN(sclscl), .SMC(test_se), .C(clk), .Q(
        sdai_ff) );
  SDFFQX1 clk_count2_ov_reg ( .D(N690), .SIN(clk_count1[3]), .SMC(test_se), 
        .C(clk), .Q(clk_count2_ov) );
  SDFFQX1 sdai_ff_reg_reg_2_ ( .D(N433), .SIN(sdai_ff_reg0[1]), .SMC(test_se), 
        .C(clk), .Q(sdai_ff_reg0[2]) );
  SDFFQX1 sdai_ff_reg_reg_1_ ( .D(N432), .SIN(sdai_ff_reg0[0]), .SMC(test_se), 
        .C(clk), .Q(sdai_ff_reg0[1]) );
  SDFFQX1 rst_delay_reg ( .D(n23), .SIN(pedetect), .SMC(test_se), .C(clk), .Q(
        rst_delay) );
  SDFFQX1 clk_count1_ov_reg ( .D(n505), .SIN(busfree), .SMC(test_se), .C(clk), 
        .Q(clk_count1_ov) );
  SDFFQX1 ack_bit_reg ( .D(n494), .SIN(test_si1), .SMC(test_se), .C(net12020), 
        .Q(ack_bit) );
  SDFFQX1 clk_count2_reg_3_ ( .D(N688), .SIN(clk_count2[2]), .SMC(test_se), 
        .C(net12056), .Q(clk_count2[3]) );
  SDFFQX1 sdai_ff_reg_reg_0_ ( .D(N431), .SIN(sdai_ff), .SMC(test_se), .C(clk), 
        .Q(sdai_ff_reg0[0]) );
  SDFFQX1 sclscl_reg ( .D(n46), .SIN(sclo_int), .SMC(test_se), .C(clk), .Q(
        sclscl) );
  SDFFQX1 clk_count2_reg_2_ ( .D(N687), .SIN(clk_count2[1]), .SMC(test_se), 
        .C(net12056), .Q(clk_count2[2]) );
  SDFFQX1 setup_counter_r_reg_2_ ( .D(N335), .SIN(setup_counter_r[1]), .SMC(
        test_se), .C(net12031), .Q(setup_counter_r[2]) );
  SDFFQX1 bsd7_reg ( .D(n491), .SIN(bclkcnt[1]), .SMC(test_se), .C(clk), .Q(
        bsd7) );
  SDFFQX1 clk_count2_reg_1_ ( .D(N686), .SIN(clk_count2[0]), .SMC(test_se), 
        .C(net12056), .Q(clk_count2[1]) );
  SDFFQX1 clk_count2_reg_0_ ( .D(N685), .SIN(clk_count2_ov), .SMC(test_se), 
        .C(net12056), .Q(clk_count2[0]) );
  SDFFQX1 starto_en_reg ( .D(n490), .SIN(setup_counter_r[2]), .SMC(test_se), 
        .C(clk), .Q(starto_en) );
  SDFFQX1 bclkcnt_reg_1_ ( .D(N511), .SIN(bclkcnt[0]), .SMC(test_se), .C(clk), 
        .Q(bclkcnt[1]) );
  SDFFQX1 indelay_reg_2_ ( .D(N471), .SIN(indelay[1]), .SMC(test_se), .C(
        net12041), .Q(indelay[2]) );
  SDFFQX1 bclkcnt_reg_0_ ( .D(N510), .SIN(adrcompen), .SMC(test_se), .C(clk), 
        .Q(bclkcnt[0]) );
  SDFFQX1 clkint_ff_reg ( .D(N700), .SIN(clk_count2[3]), .SMC(test_se), .C(clk), .Q(clkint_ff) );
  SDFFQX1 setup_counter_r_reg_0_ ( .D(N333), .SIN(sdao), .SMC(test_se), .C(
        net12031), .Q(setup_counter_r[0]) );
  SDFFQX1 write_data_r_reg ( .D(n500), .SIN(test_si2), .SMC(test_se), .C(clk), 
        .Q(test_so2) );
  SDFFQX1 busfree_reg ( .D(n506), .SIN(bsd7_tmp), .SMC(test_se), .C(clk), .Q(
        busfree) );
  SDFFQX1 bsd7_tmp_reg ( .D(n492), .SIN(bsd7), .SMC(test_se), .C(clk), .Q(
        bsd7_tmp) );
  SDFFQX1 clkint_reg ( .D(n504), .SIN(clkint_ff), .SMC(test_se), .C(clk), .Q(
        clkint) );
  SDFFQX1 scli_ff_reg_reg_1_ ( .D(N413), .SIN(scli_ff_reg0[0]), .SMC(test_se), 
        .C(clk), .Q(scli_ff_reg0[1]) );
  SDFFQX1 scli_ff_reg_reg_0_ ( .D(N412), .SIN(scli_ff), .SMC(test_se), .C(clk), 
        .Q(scli_ff_reg0[0]) );
  SDFFQX1 indelay_reg_1_ ( .D(N470), .SIN(indelay[0]), .SMC(test_se), .C(
        net12041), .Q(indelay[1]) );
  SDFFQX1 setup_counter_r_reg_1_ ( .D(n36), .SIN(setup_counter_r[0]), .SMC(
        test_se), .C(net12031), .Q(setup_counter_r[1]) );
  SDFFQX1 scli_ff_reg_reg_2_ ( .D(N414), .SIN(scli_ff_reg0[1]), .SMC(test_se), 
        .C(clk), .Q(scli_ff_reg0[2]) );
  SDFFQX1 fsmsync_reg_1_ ( .D(N747), .SIN(fsmsync[0]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[1]) );
  SDFFQX1 indelay_reg_0_ ( .D(N469), .SIN(i2csta_o[7]), .SMC(test_se), .C(
        net12041), .Q(indelay[0]) );
  SDFFQX1 fsmsync_reg_0_ ( .D(N746), .SIN(fsmsta[4]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[0]) );
  SDFFQX1 fsmsync_reg_2_ ( .D(N748), .SIN(fsmsync[1]), .SMC(test_se), .C(clk), 
        .Q(fsmsync[2]) );
  SDFFQX1 pedetect_reg ( .D(n497), .SIN(nedetect), .SMC(test_se), .C(clk), .Q(
        pedetect) );
  SDFFQX1 nedetect_reg ( .D(n498), .SIN(indelay[2]), .SMC(test_se), .C(clk), 
        .Q(nedetect) );
  SDFFQX1 clk_count1_reg_2_ ( .D(N656), .SIN(clk_count1[1]), .SMC(test_se), 
        .C(net12051), .Q(clk_count1[2]) );
  SDFFQX1 fsmdet_reg_0_ ( .D(N1063), .SIN(framesync[3]), .SMC(test_se), .C(clk), .Q(fsmdet[0]) );
  SDFFQX1 adrcomp_reg ( .D(n501), .SIN(ack), .SMC(test_se), .C(clk), .Q(
        adrcomp) );
  SDFFQX1 adrcompen_reg ( .D(n496), .SIN(adrcomp), .SMC(test_se), .C(clk), .Q(
        adrcompen) );
  SDFFQX1 clk_count1_reg_1_ ( .D(N655), .SIN(clk_count1[0]), .SMC(test_se), 
        .C(net12051), .Q(clk_count1[1]) );
  SDFFQX1 fsmdet_reg_1_ ( .D(N1064), .SIN(fsmdet[0]), .SMC(test_se), .C(clk), 
        .Q(fsmdet[1]) );
  SDFFQX1 ack_reg ( .D(n493), .SIN(ack_bit), .SMC(test_se), .C(clk), .Q(ack)
         );
  SDFFQX1 fsmdet_reg_2_ ( .D(N1065), .SIN(fsmdet[1]), .SMC(test_se), .C(clk), 
        .Q(fsmdet[2]) );
  SDFFQX1 clk_count1_reg_0_ ( .D(N654), .SIN(clk_count1_ov), .SMC(test_se), 
        .C(net12051), .Q(clk_count1[0]) );
  SDFFQX1 sdaint_reg ( .D(n507), .SIN(sdai_ff_reg0[2]), .SMC(test_se), .C(clk), 
        .Q(sdaint) );
  SDFFQX1 clk_count1_reg_3_ ( .D(N657), .SIN(clk_count1[2]), .SMC(test_se), 
        .C(net12051), .Q(clk_count1[3]) );
  SDFFQX1 sclint_reg ( .D(n499), .SIN(scli_ff_reg0[2]), .SMC(test_se), .C(clk), 
        .Q(sclint) );
  SDFFQX1 fsmmod_reg_0_ ( .D(N1124), .SIN(fsmdet[2]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[0]) );
  SDFFQX1 fsmmod_reg_1_ ( .D(N1125), .SIN(fsmmod[0]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[1]) );
  SDFFQX1 fsmmod_reg_2_ ( .D(N1126), .SIN(fsmmod[1]), .SMC(test_se), .C(clk), 
        .Q(fsmmod[2]) );
  SDFFQX1 framesync_reg_3_ ( .D(N495), .SIN(framesync[2]), .SMC(test_se), .C(
        net12046), .Q(framesync[3]) );
  SDFFQX1 framesync_reg_1_ ( .D(N493), .SIN(framesync[0]), .SMC(test_se), .C(
        net12046), .Q(framesync[1]) );
  SDFFQX1 framesync_reg_2_ ( .D(N494), .SIN(framesync[1]), .SMC(test_se), .C(
        net12046), .Q(framesync[2]) );
  SDFFQX1 framesync_reg_0_ ( .D(N492), .SIN(clkint), .SMC(test_se), .C(
        net12046), .Q(framesync[0]) );
  SDFFQX1 fsmsta_reg_2_ ( .D(N1025), .SIN(fsmsta[1]), .SMC(test_se), .C(
        net12061), .Q(fsmsta[2]) );
  SDFFQX1 fsmsta_reg_1_ ( .D(N1024), .SIN(fsmsta[0]), .SMC(test_se), .C(
        net12061), .Q(fsmsta[1]) );
  SDFFQX1 fsmsta_reg_0_ ( .D(N1023), .SIN(fsmmod[2]), .SMC(test_se), .C(
        net12061), .Q(fsmsta[0]) );
  SDFFQX1 fsmsta_reg_4_ ( .D(N1027), .SIN(fsmsta[3]), .SMC(test_se), .C(
        net12061), .Q(fsmsta[4]) );
  SDFFQX1 fsmsta_reg_3_ ( .D(N1026), .SIN(fsmsta[2]), .SMC(test_se), .C(
        net12061), .Q(fsmsta[3]) );
  SDFFQX1 i2csta_reg_4_ ( .D(N410), .SIN(i2csta_o[6]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[7]) );
  SDFFQX1 i2cdat_reg_7_ ( .D(N304), .SIN(i2cdat_o[6]), .SMC(test_se), .C(
        net12026), .Q(i2cdat_o[7]) );
  SDFFQX1 i2cadr_reg_7_ ( .D(N350), .SIN(i2cadr_o[6]), .SMC(test_se), .C(
        net12036), .Q(i2cadr_o[7]) );
  SDFFQX1 i2cdat_reg_6_ ( .D(N303), .SIN(i2cdat_o[5]), .SMC(test_se), .C(
        net12026), .Q(i2cdat_o[6]) );
  SDFFQX1 i2ccon_reg_7_ ( .D(N234), .SIN(i2ccon_o[6]), .SMC(test_se), .C(
        net12020), .Q(i2ccon_o[7]) );
  SDFFQX1 i2csta_reg_3_ ( .D(N409), .SIN(i2csta_o[5]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[6]) );
  SDFFQX1 i2csta_reg_2_ ( .D(N408), .SIN(i2csta_o[4]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[5]) );
  SDFFQX1 i2cadr_reg_6_ ( .D(N349), .SIN(i2cadr_o[5]), .SMC(test_se), .C(
        net12036), .Q(i2cadr_o[6]) );
  SDFFQX1 i2cdat_reg_5_ ( .D(N302), .SIN(i2cdat_o[4]), .SMC(test_se), .C(
        net12026), .Q(i2cdat_o[5]) );
  SDFFQX1 i2cdat_reg_4_ ( .D(N301), .SIN(i2cdat_o[3]), .SMC(test_se), .C(
        net12026), .Q(i2cdat_o[4]) );
  SDFFQX1 i2ccon_reg_5_ ( .D(N232), .SIN(i2ccon_o[4]), .SMC(test_se), .C(
        net12020), .Q(i2ccon_o[5]) );
  SDFFQX1 i2ccon_reg_6_ ( .D(N233), .SIN(i2ccon_o[5]), .SMC(test_se), .C(
        net12020), .Q(i2ccon_o[6]) );
  SDFFQX1 i2csta_reg_1_ ( .D(N407), .SIN(i2csta_o[3]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[4]) );
  SDFFQX1 i2cadr_reg_4_ ( .D(N347), .SIN(i2cadr_o[3]), .SMC(test_se), .C(
        net12036), .Q(i2cadr_o[4]) );
  SDFFQX1 i2cadr_reg_5_ ( .D(N348), .SIN(i2cadr_o[4]), .SMC(test_se), .C(
        net12036), .Q(i2cadr_o[5]) );
  SDFFQX1 i2ccon_reg_4_ ( .D(n503), .SIN(i2ccon_o[3]), .SMC(test_se), .C(clk), 
        .Q(i2ccon_o[4]) );
  SDFFQX1 i2cdat_reg_3_ ( .D(N300), .SIN(i2cdat_o[2]), .SMC(test_se), .C(
        net12026), .Q(i2cdat_o[3]) );
  SDFFQX1 i2csta_reg_0_ ( .D(N406), .SIN(i2cdat_o[7]), .SMC(test_se), .C(clk), 
        .Q(i2csta_o[3]) );
  SDFFQX1 i2cadr_reg_3_ ( .D(N346), .SIN(i2cadr_o[2]), .SMC(test_se), .C(
        net12036), .Q(i2cadr_o[3]) );
  SDFFQX1 i2ccon_reg_3_ ( .D(n495), .SIN(i2ccon_o[2]), .SMC(test_se), .C(clk), 
        .Q(i2ccon_o[3]) );
  SDFFQX1 sclo_int_reg ( .D(N749), .SIN(sclint), .SMC(test_se), .C(clk), .Q(
        sclo_int) );
  SDFFQX1 wait_for_setup_r_reg ( .D(N336), .SIN(starto_en), .SMC(test_se), .C(
        clk), .Q(test_so1) );
  SDFFQX1 sdao_int_reg ( .D(n502), .SIN(sdaint), .SMC(test_se), .C(clk), .Q(
        sdao) );
  SDFFQX1 i2cadr_reg_1_ ( .D(N344), .SIN(i2cadr_o[0]), .SMC(test_se), .C(
        net12036), .Q(i2cadr_o[1]) );
  SDFFQX1 i2ccon_reg_1_ ( .D(N226), .SIN(i2ccon_o[0]), .SMC(test_se), .C(
        net12020), .Q(i2ccon_o[1]) );
  SDFFQX1 i2cdat_reg_1_ ( .D(N298), .SIN(i2cdat_o[0]), .SMC(test_se), .C(
        net12026), .Q(i2cdat_o[1]) );
  SDFFQX1 i2cadr_reg_2_ ( .D(N345), .SIN(i2cadr_o[1]), .SMC(test_se), .C(
        net12036), .Q(i2cadr_o[2]) );
  SDFFQX1 i2ccon_reg_2_ ( .D(N227), .SIN(i2ccon_o[1]), .SMC(test_se), .C(
        net12020), .Q(i2ccon_o[2]) );
  SDFFQX1 i2ccon_reg_0_ ( .D(N225), .SIN(i2cadr_o[7]), .SMC(test_se), .C(
        net12020), .Q(i2ccon_o[0]) );
  SDFFQX1 i2cdat_reg_0_ ( .D(N297), .SIN(i2ccon_o[7]), .SMC(test_se), .C(
        net12026), .Q(i2cdat_o[0]) );
  SDFFQX1 i2cdat_reg_2_ ( .D(N299), .SIN(i2cdat_o[1]), .SMC(test_se), .C(
        net12026), .Q(i2cdat_o[2]) );
  SDFFQX1 i2cadr_reg_0_ ( .D(N343), .SIN(fsmsync[2]), .SMC(test_se), .C(
        net12036), .Q(i2cadr_o[0]) );
  INVX1 U3 ( .A(1'b1), .Y(i2csta_o[0]) );
  INVX1 U5 ( .A(1'b1), .Y(i2csta_o[1]) );
  INVX1 U7 ( .A(1'b1), .Y(i2csta_o[2]) );
  INVX1 U9 ( .A(n10), .Y(n7) );
  INVX1 U10 ( .A(fsmsta[1]), .Y(n8) );
  INVX1 U11 ( .A(si), .Y(n9) );
  BUFX3 U12 ( .A(n92), .Y(n10) );
  INVX1 U13 ( .A(n129), .Y(n28) );
  NOR2X1 U14 ( .A(n21), .B(n171), .Y(n129) );
  AOI21X1 U15 ( .B(n31), .C(n86), .A(n318), .Y(n208) );
  INVX1 U16 ( .A(n212), .Y(n31) );
  NAND2X1 U17 ( .A(n171), .B(n24), .Y(n126) );
  NOR2X1 U18 ( .A(n16), .B(n126), .Y(n192) );
  OAI21X1 U19 ( .B(n310), .C(n13), .A(n25), .Y(N343) );
  OAI21X1 U20 ( .B(n16), .C(n310), .A(n25), .Y(N346) );
  OAI21X1 U21 ( .B(n20), .C(n310), .A(n25), .Y(N350) );
  NOR2X1 U22 ( .A(n310), .B(n17), .Y(N347) );
  NOR2X1 U23 ( .A(n310), .B(n14), .Y(N344) );
  NOR2X1 U24 ( .A(n310), .B(n15), .Y(N345) );
  NOR2X1 U25 ( .A(n310), .B(n18), .Y(N348) );
  NOR2X1 U26 ( .A(n310), .B(n19), .Y(N349) );
  NAND2X1 U27 ( .A(n25), .B(n310), .Y(N342) );
  NOR2X1 U28 ( .A(n22), .B(n19), .Y(N233) );
  NOR2X1 U29 ( .A(n22), .B(n18), .Y(N232) );
  NOR2X1 U30 ( .A(n22), .B(n20), .Y(N234) );
  NOR2X1 U31 ( .A(n21), .B(n13), .Y(N225) );
  NOR2X1 U32 ( .A(n22), .B(n14), .Y(N226) );
  NOR2X1 U33 ( .A(n21), .B(n15), .Y(N227) );
  INVX1 U34 ( .A(n27), .Y(n22) );
  NOR2X1 U35 ( .A(n88), .B(n86), .Y(n217) );
  INVX1 U36 ( .A(n407), .Y(n104) );
  INVX1 U37 ( .A(n204), .Y(n88) );
  INVX1 U38 ( .A(n26), .Y(n21) );
  INVX1 U39 ( .A(n26), .Y(n23) );
  INVX1 U40 ( .A(n421), .Y(n60) );
  INVX1 U41 ( .A(n432), .Y(n78) );
  OR2X1 U42 ( .A(sdai), .B(n23), .Y(N181) );
  NOR42XL U43 ( .C(sfraddr[1]), .D(n312), .A(sfraddr[0]), .B(sfraddr[2]), .Y(
        n212) );
  NOR42XL U44 ( .C(sfraddr[2]), .D(n312), .A(sfraddr[0]), .B(sfraddr[1]), .Y(
        n171) );
  NOR42XL U45 ( .C(sfraddr[4]), .D(sfraddr[3]), .A(sfraddr[5]), .B(n328), .Y(
        n312) );
  NAND2X1 U46 ( .A(sfrwe), .B(sfraddr[6]), .Y(n328) );
  AOI21X1 U47 ( .B(n175), .C(n204), .A(n174), .Y(n318) );
  INVX1 U48 ( .A(n174), .Y(n30) );
  NAND4X1 U49 ( .A(sfraddr[0]), .B(sfraddr[1]), .C(n311), .D(n312), .Y(n310)
         );
  NOR2XL U50 ( .A(sfraddr[2]), .B(n21), .Y(n311) );
  INVX1 U51 ( .A(sfrdatai[6]), .Y(n19) );
  INVX1 U52 ( .A(sfrdatai[7]), .Y(n20) );
  INVX1 U53 ( .A(sfrdatai[4]), .Y(n17) );
  INVX1 U54 ( .A(sfrdatai[5]), .Y(n18) );
  INVX1 U55 ( .A(sfrdatai[2]), .Y(n15) );
  INVX1 U56 ( .A(sfrdatai[1]), .Y(n14) );
  INVX1 U57 ( .A(sfrdatai[0]), .Y(n13) );
  INVX1 U58 ( .A(sfrdatai[3]), .Y(n16) );
  AOI21X1 U59 ( .B(n105), .C(n436), .A(n417), .Y(n398) );
  INVX1 U60 ( .A(n327), .Y(n436) );
  INVX1 U61 ( .A(n324), .Y(n103) );
  NAND2X1 U62 ( .A(n105), .B(n440), .Y(n407) );
  NAND2X1 U63 ( .A(n323), .B(n147), .Y(n204) );
  INVX1 U64 ( .A(n150), .Y(n77) );
  INVX1 U65 ( .A(n173), .Y(n86) );
  NAND2X1 U66 ( .A(n145), .B(n92), .Y(n376) );
  INVX1 U67 ( .A(rst), .Y(n27) );
  NAND2X1 U68 ( .A(n379), .B(n383), .Y(n405) );
  INVX1 U69 ( .A(n175), .Y(n87) );
  INVX1 U70 ( .A(n187), .Y(n89) );
  INVX1 U71 ( .A(n196), .Y(n69) );
  NOR21XL U72 ( .B(n137), .A(n138), .Y(n133) );
  NAND42X1 U73 ( .C(n152), .D(n104), .A(n363), .B(n325), .Y(n356) );
  OAI21X1 U74 ( .B(n364), .C(n362), .A(n10), .Y(n363) );
  NAND2X1 U75 ( .A(n195), .B(n26), .Y(n432) );
  NAND3X1 U76 ( .A(n78), .B(n434), .C(n435), .Y(n421) );
  AND3X1 U77 ( .A(n380), .B(n325), .C(n384), .Y(n409) );
  NOR4XL U78 ( .A(n432), .B(n198), .C(n69), .D(n434), .Y(n370) );
  NAND2X1 U79 ( .A(n425), .B(n280), .Y(n380) );
  INVX1 U80 ( .A(rst), .Y(n26) );
  INVX1 U81 ( .A(n434), .Y(n85) );
  NOR2X1 U82 ( .A(n385), .B(n99), .Y(n359) );
  NAND2X1 U83 ( .A(n379), .B(n380), .Y(n364) );
  INVX1 U84 ( .A(n154), .Y(n101) );
  INVX1 U85 ( .A(n368), .Y(n59) );
  INVX1 U86 ( .A(n125), .Y(n58) );
  INVX1 U87 ( .A(n392), .Y(n99) );
  INVX1 U88 ( .A(n250), .Y(n76) );
  INVX1 U89 ( .A(n309), .Y(n98) );
  INVX1 U90 ( .A(n116), .Y(n73) );
  NAND42X1 U91 ( .C(n370), .D(n368), .A(n421), .B(n431), .Y(N1022) );
  NOR2X1 U92 ( .A(n34), .B(n432), .Y(n431) );
  NAND2X1 U93 ( .A(n442), .B(n309), .Y(n229) );
  INVX1 U94 ( .A(rst), .Y(n24) );
  INVX1 U95 ( .A(n296), .Y(n62) );
  INVX1 U96 ( .A(n282), .Y(n35) );
  INVX1 U97 ( .A(n335), .Y(n32) );
  NAND2X1 U98 ( .A(n25), .B(n250), .Y(n233) );
  INVX1 U99 ( .A(rst), .Y(n25) );
  NAND2X1 U100 ( .A(n62), .B(n47), .Y(N468) );
  OR2X1 U101 ( .A(scli), .B(n23), .Y(N180) );
  OAI21X1 U102 ( .B(n210), .C(n52), .A(n211), .Y(n492) );
  GEN2XL U103 ( .D(n20), .E(n174), .C(n175), .B(n24), .A(n29), .Y(n211) );
  INVX1 U104 ( .A(n210), .Y(n29) );
  OAI21BBX1 U105 ( .A(n212), .B(n209), .C(n213), .Y(n210) );
  NAND2X1 U106 ( .A(n33), .B(n31), .Y(n174) );
  AOI32X1 U107 ( .A(n212), .B(n33), .C(n87), .D(n209), .E(n31), .Y(n219) );
  OAI22X1 U108 ( .A(n167), .B(n14), .C(n208), .D(n449), .Y(N298) );
  OAI22X1 U109 ( .A(n167), .B(n16), .C(n208), .D(n450), .Y(N300) );
  OAI22X1 U110 ( .A(n167), .B(n15), .C(n208), .D(n452), .Y(N299) );
  OAI22X1 U111 ( .A(n167), .B(n13), .C(n208), .D(n84), .Y(N297) );
  OAI21X1 U112 ( .B(n84), .C(n205), .A(n206), .Y(n493) );
  OAI21BBX1 U113 ( .A(n82), .B(n207), .C(n205), .Y(n206) );
  OAI21X1 U114 ( .B(n208), .C(n66), .A(n207), .Y(n205) );
  NOR2X1 U115 ( .A(n21), .B(n209), .Y(n207) );
  OAI211X1 U116 ( .C(n322), .D(n66), .A(n26), .B(n31), .Y(N296) );
  NOR2X1 U117 ( .A(n86), .B(n318), .Y(n322) );
  INVX1 U118 ( .A(n186), .Y(n92) );
  NAND3X1 U119 ( .A(n441), .B(n443), .C(n438), .Y(n327) );
  NAND3X1 U120 ( .A(n430), .B(n378), .C(n398), .Y(n416) );
  NAND3X1 U121 ( .A(n444), .B(n441), .C(n424), .Y(n430) );
  NAND2X1 U122 ( .A(n424), .B(n105), .Y(n324) );
  AND2X1 U123 ( .A(n307), .B(n436), .Y(n417) );
  OAI221X1 U124 ( .A(n399), .B(n59), .C(n70), .D(n365), .E(n400), .Y(N1024) );
  AOI31X1 U125 ( .A(n156), .B(n84), .C(n60), .D(n370), .Y(n400) );
  NOR4XL U126 ( .A(n401), .B(n402), .C(n391), .D(n403), .Y(n399) );
  ENOX1 U127 ( .A(n409), .B(n360), .C(n376), .D(n101), .Y(n402) );
  NAND2X1 U128 ( .A(n436), .B(n444), .Y(n294) );
  INVX1 U129 ( .A(n230), .Y(n105) );
  NAND2X1 U130 ( .A(n103), .B(n441), .Y(n383) );
  OAI211X1 U131 ( .C(n418), .D(n59), .A(n366), .B(n419), .Y(N1023) );
  NOR2X1 U132 ( .A(n420), .B(n34), .Y(n419) );
  NOR4XL U133 ( .A(n422), .B(n403), .C(n423), .D(n357), .Y(n418) );
  AOI21X1 U134 ( .B(n409), .C(n383), .A(n91), .Y(n423) );
  NAND31X1 U135 ( .C(n334), .A(n146), .B(n340), .Y(n150) );
  NAND31X1 U136 ( .C(n303), .A(n280), .B(n438), .Y(n384) );
  NAND32X1 U137 ( .B(n140), .C(n147), .A(n323), .Y(n173) );
  NOR2X1 U138 ( .A(n22), .B(n188), .Y(n187) );
  NAND2X1 U139 ( .A(n323), .B(n140), .Y(n175) );
  OAI211X1 U140 ( .C(n98), .D(n303), .A(n324), .B(n325), .Y(n147) );
  NOR2X1 U141 ( .A(n89), .B(n445), .Y(n323) );
  AOI21X1 U142 ( .B(n97), .C(n90), .A(n92), .Y(n198) );
  NAND2X1 U143 ( .A(n77), .B(n70), .Y(n196) );
  OAI32X1 U144 ( .A(n154), .B(n156), .C(n448), .D(n186), .E(n294), .Y(n413) );
  NOR2X1 U145 ( .A(n437), .B(n441), .Y(n425) );
  NOR3XL U146 ( .A(n186), .B(n84), .C(n294), .Y(n382) );
  NOR2X1 U147 ( .A(n79), .B(n83), .Y(n244) );
  NAND3X1 U148 ( .A(n440), .B(n438), .C(n280), .Y(n325) );
  NAND2X1 U149 ( .A(n425), .B(n307), .Y(n379) );
  OAI21X1 U150 ( .B(n386), .C(n59), .A(n387), .Y(N1025) );
  OAI21BBX1 U151 ( .A(n156), .B(n84), .C(n60), .Y(n387) );
  NOR41XL U152 ( .D(n388), .A(n389), .B(n390), .C(n391), .Y(n386) );
  NOR2X1 U153 ( .A(n10), .B(n380), .Y(n390) );
  NOR2X1 U154 ( .A(n175), .B(n33), .Y(n209) );
  AOI211X1 U155 ( .C(n385), .D(n393), .A(n394), .B(n395), .Y(n388) );
  AOI21X1 U156 ( .B(n361), .C(n186), .A(n398), .Y(n394) );
  OAI211X1 U157 ( .C(n396), .D(n437), .A(n397), .B(n154), .Y(n395) );
  NAND2X1 U158 ( .A(n441), .B(n444), .Y(n396) );
  NAND4X1 U159 ( .A(n407), .B(n397), .C(n426), .D(n427), .Y(n403) );
  NAND4X1 U160 ( .A(n436), .B(n105), .C(n361), .D(n186), .Y(n426) );
  AOI22X1 U161 ( .A(n99), .B(n393), .C(n385), .D(n360), .Y(n427) );
  NOR2X1 U162 ( .A(n244), .B(n143), .Y(n340) );
  INVX1 U163 ( .A(n292), .Y(n280) );
  NAND2X1 U164 ( .A(n382), .B(n82), .Y(n397) );
  INVX1 U165 ( .A(n301), .Y(n440) );
  INVX1 U166 ( .A(n424), .Y(n437) );
  NOR2X1 U167 ( .A(n274), .B(n21), .Y(n125) );
  NAND32X1 U168 ( .B(n143), .C(n23), .A(n144), .Y(n135) );
  AOI21X1 U169 ( .B(n76), .C(n70), .A(n445), .Y(n144) );
  NOR4XL U170 ( .A(n432), .B(n66), .C(n85), .D(n435), .Y(n368) );
  NOR2X1 U171 ( .A(n188), .B(n278), .Y(n434) );
  AND3X1 U172 ( .A(n188), .B(n244), .C(n80), .Y(n420) );
  NAND2X1 U173 ( .A(n438), .B(n100), .Y(n309) );
  NAND3X1 U174 ( .A(n424), .B(n441), .C(n307), .Y(n154) );
  NOR2X1 U175 ( .A(n75), .B(n272), .Y(n116) );
  NAND3X1 U176 ( .A(n79), .B(n83), .C(n80), .Y(n250) );
  OAI31XL U177 ( .A(n376), .B(n84), .C(n154), .D(n229), .Y(n357) );
  NAND3X1 U178 ( .A(n100), .B(n444), .C(n425), .Y(n392) );
  AOI21X1 U179 ( .B(n188), .C(n341), .A(n420), .Y(n195) );
  NOR2X1 U180 ( .A(n445), .B(n21), .Y(n170) );
  AOI211X1 U181 ( .C(n154), .D(n150), .A(n155), .B(n61), .Y(n153) );
  OAI21X1 U182 ( .B(n156), .C(n84), .A(n157), .Y(n155) );
  OAI22X1 U183 ( .A(n156), .B(n448), .C(n158), .D(n159), .Y(n157) );
  NAND3X1 U184 ( .A(n160), .B(n161), .C(n162), .Y(n159) );
  OAI21X1 U185 ( .B(n141), .C(n92), .A(n147), .Y(n137) );
  OAI21X1 U186 ( .B(n272), .C(n65), .A(n73), .Y(n123) );
  AOI21X1 U187 ( .B(n84), .C(n60), .A(n23), .Y(n366) );
  NOR3XL U188 ( .A(n66), .B(n101), .C(n376), .Y(n435) );
  NOR2X1 U189 ( .A(n65), .B(n75), .Y(n266) );
  NOR2X1 U190 ( .A(n96), .B(n351), .Y(n278) );
  OAI21BBX1 U191 ( .A(n384), .B(n359), .C(n360), .Y(n371) );
  OAI21X1 U192 ( .B(n7), .C(n383), .A(n384), .Y(n381) );
  OAI31XL U193 ( .A(n38), .B(n314), .C(n37), .D(n313), .Y(N335) );
  AOI211X1 U194 ( .C(n51), .D(n48), .A(n256), .B(n261), .Y(N686) );
  AOI211X1 U195 ( .C(n65), .D(n75), .A(n264), .B(n266), .Y(N655) );
  NOR2X1 U196 ( .A(n303), .B(n230), .Y(n385) );
  INVX1 U197 ( .A(n316), .Y(n37) );
  NAND2X1 U198 ( .A(n188), .B(n170), .Y(n172) );
  NOR2X1 U199 ( .A(n61), .B(n70), .Y(n145) );
  AOI31X1 U200 ( .A(n303), .B(n301), .C(n308), .D(n444), .Y(n415) );
  NOR2X1 U201 ( .A(n408), .B(n186), .Y(n374) );
  NAND2X1 U202 ( .A(n377), .B(n378), .Y(n362) );
  INVX1 U203 ( .A(n365), .Y(n34) );
  NAND2X1 U204 ( .A(n125), .B(n64), .Y(N700) );
  NAND2X1 U205 ( .A(n125), .B(n40), .Y(N689) );
  INVX1 U206 ( .A(n237), .Y(n93) );
  INVX1 U207 ( .A(n378), .Y(n439) );
  INVX1 U208 ( .A(n200), .Y(n90) );
  INVX1 U209 ( .A(n360), .Y(n91) );
  INVX1 U210 ( .A(n361), .Y(n81) );
  NAND21X1 U211 ( .B(n145), .A(n146), .Y(n138) );
  NAND3X1 U212 ( .A(n67), .B(n27), .C(n226), .Y(n296) );
  NOR2X1 U213 ( .A(n254), .B(n237), .Y(n335) );
  NOR2X1 U214 ( .A(n291), .B(n10), .Y(n282) );
  NAND2X1 U215 ( .A(n130), .B(n56), .Y(n113) );
  NOR2X1 U216 ( .A(n33), .B(n21), .Y(n298) );
  NOR2X1 U217 ( .A(n63), .B(n68), .Y(n226) );
  OAI22X1 U218 ( .A(n91), .B(n392), .C(n374), .D(n378), .Y(n389) );
  NAND2X1 U219 ( .A(n447), .B(n33), .Y(n239) );
  OAI21X1 U220 ( .B(n33), .C(n57), .A(n68), .Y(n247) );
  NOR2X1 U221 ( .A(n309), .B(n443), .Y(n152) );
  OAI21X1 U222 ( .B(n442), .C(n305), .A(n298), .Y(N408) );
  XNOR2XL U223 ( .A(n230), .B(n438), .Y(n305) );
  OAI21X1 U224 ( .B(n447), .C(n237), .A(n9), .Y(n235) );
  OAI31XL U225 ( .A(n66), .B(n180), .C(n176), .D(n181), .Y(n497) );
  NAND4X1 U226 ( .A(n26), .B(n71), .C(n177), .D(n182), .Y(n181) );
  NOR3XL U227 ( .A(n44), .B(n50), .C(n49), .Y(n182) );
  AOI21X1 U228 ( .B(n230), .C(n438), .A(n441), .Y(n228) );
  AOI21X1 U229 ( .B(n71), .C(n52), .A(n33), .Y(n218) );
  OAI211X1 U230 ( .C(n139), .D(n97), .A(n140), .B(n41), .Y(n134) );
  INVX1 U231 ( .A(n177), .Y(n43) );
  NOR2X1 U232 ( .A(n446), .B(n451), .Y(n115) );
  NOR2X1 U233 ( .A(n74), .B(n273), .Y(n121) );
  NAND2X1 U234 ( .A(n273), .B(n74), .Y(n119) );
  NAND4X1 U235 ( .A(n298), .B(n299), .C(n300), .D(n301), .Y(N410) );
  NAND2X1 U236 ( .A(n152), .B(n444), .Y(n299) );
  NAND2X1 U237 ( .A(n49), .B(n24), .Y(N414) );
  NAND2X1 U238 ( .A(n50), .B(n25), .Y(N413) );
  INVX1 U239 ( .A(n221), .Y(n56) );
  INVX1 U240 ( .A(n246), .Y(n57) );
  INVX1 U241 ( .A(n251), .Y(n47) );
  INVX1 U242 ( .A(n308), .Y(n442) );
  NAND2X1 U243 ( .A(n37), .B(n313), .Y(N336) );
  NAND2X1 U244 ( .A(n298), .B(n306), .Y(N407) );
  OAI21X1 U245 ( .B(n307), .C(n280), .A(n308), .Y(n306) );
  INVX1 U246 ( .A(n270), .Y(n451) );
  INVX1 U247 ( .A(n285), .Y(n94) );
  NOR2X1 U248 ( .A(n96), .B(n95), .Y(n350) );
  NOR2X1 U249 ( .A(n51), .B(n48), .Y(n261) );
  NAND2X1 U250 ( .A(n68), .B(n63), .Y(n225) );
  OAI21AX1 U251 ( .B(n71), .C(n43), .A(n176), .Y(n499) );
  NAND2X1 U252 ( .A(n221), .B(n57), .Y(n336) );
  NAND4X1 U253 ( .A(n289), .B(n187), .C(n291), .D(n237), .Y(N491) );
  NOR21XL U254 ( .B(sclo_int), .A(test_so1), .Y(sclo) );
  NOR32XL U255 ( .B(n172), .C(n220), .A(n21), .Y(n213) );
  NAND4X1 U256 ( .A(n30), .B(n87), .C(nedetect), .D(n66), .Y(n220) );
  OAI22AX1 U257 ( .D(i2cdat_o[4]), .C(n208), .A(n167), .B(n18), .Y(N302) );
  OAI22AX1 U258 ( .D(i2cdat_o[3]), .C(n208), .A(n167), .B(n17), .Y(N301) );
  OAI22AX1 U259 ( .D(i2cdat_o[5]), .C(n208), .A(n167), .B(n19), .Y(N303) );
  OAI22AX1 U260 ( .D(i2cdat_o[6]), .C(n208), .A(n167), .B(n20), .Y(N304) );
  ENOX1 U261 ( .A(n189), .B(n190), .C(i2ccon_o[3]), .D(n189), .Y(n495) );
  AOI21X1 U262 ( .B(n191), .C(n129), .A(n192), .Y(n190) );
  AOI21BBXL U263 ( .B(n193), .C(n192), .A(n191), .Y(n189) );
  AOI21X1 U264 ( .B(n194), .C(n195), .A(n445), .Y(n191) );
  ENOX1 U265 ( .A(n126), .B(n127), .C(n127), .D(i2ccon_o[4]), .Y(n503) );
  OAI21X1 U266 ( .B(sfrdatai[4]), .C(n126), .A(n128), .Y(n127) );
  NAND4X1 U267 ( .A(i2ccon_o[6]), .B(n112), .C(n113), .D(n129), .Y(n128) );
  ENOX1 U268 ( .A(n214), .B(n41), .C(n215), .D(n214), .Y(n491) );
  OAI211X1 U269 ( .C(n216), .D(n175), .A(n24), .B(n217), .Y(n215) );
  NAND3X1 U270 ( .A(n213), .B(n217), .C(n219), .Y(n214) );
  AOI221XL U271 ( .A(i2cdat_o[7]), .B(n30), .C(sfrdatai[7]), .D(n212), .E(n218), .Y(n216) );
  NOR2X1 U272 ( .A(intack), .B(n28), .Y(n193) );
  AND4X1 U273 ( .A(n319), .B(n320), .C(n321), .D(n172), .Y(n167) );
  NAND2X1 U274 ( .A(n25), .B(n445), .Y(n320) );
  OAI21X1 U275 ( .B(n87), .C(n88), .A(i2ccon_o[3]), .Y(n319) );
  OAI21BBX1 U276 ( .A(n175), .B(n217), .C(n212), .Y(n321) );
  OAI22X1 U277 ( .A(n167), .B(n31), .C(n168), .D(n169), .Y(n500) );
  NAND3X1 U278 ( .A(n170), .B(n171), .C(test_so2), .Y(n169) );
  NAND4X1 U279 ( .A(n172), .B(n173), .C(n174), .D(n175), .Y(n168) );
  ENOX1 U280 ( .A(n201), .B(n202), .C(n202), .D(ack_bit), .Y(n494) );
  NOR2X1 U281 ( .A(n21), .B(sfrdatai[2]), .Y(n201) );
  NAND2X1 U282 ( .A(n28), .B(n203), .Y(n202) );
  OAI21X1 U283 ( .B(n33), .C(n204), .A(n24), .Y(n203) );
  BUFX3 U284 ( .A(i2ccon_o[3]), .Y(si) );
  NAND2X1 U285 ( .A(framesync[3]), .B(n200), .Y(n186) );
  NOR3XL U286 ( .A(framesync[1]), .B(framesync[2]), .C(framesync[0]), .Y(n200)
         );
  NOR2X1 U287 ( .A(n438), .B(fsmsta[4]), .Y(n424) );
  INVX1 U288 ( .A(fsmsta[3]), .Y(n441) );
  OAI221X1 U289 ( .A(n374), .B(n377), .C(n91), .D(n300), .E(n404), .Y(n391) );
  AOI222XL U290 ( .A(n405), .B(n186), .C(n104), .D(fsmsta[2]), .E(n81), .F(
        n406), .Y(n404) );
  OAI221X1 U291 ( .A(n186), .B(n384), .C(n92), .D(n294), .E(n383), .Y(n406) );
  NAND2X1 U292 ( .A(fsmsta[0]), .B(fsmsta[1]), .Y(n230) );
  INVX1 U293 ( .A(fsmsta[2]), .Y(n438) );
  OAI21BX1 U294 ( .C(n393), .B(n379), .A(n428), .Y(n422) );
  AOI33X1 U295 ( .A(sdaint), .B(n429), .C(n92), .D(n361), .E(n7), .F(n280), 
        .Y(n428) );
  OAI211X1 U296 ( .C(ack), .D(n294), .A(n377), .B(n102), .Y(n429) );
  INVX1 U297 ( .A(n416), .Y(n102) );
  INVX1 U298 ( .A(fsmsta[4]), .Y(n443) );
  AOI21X1 U299 ( .B(n80), .C(fsmmod[2]), .A(n341), .Y(n146) );
  INVX1 U300 ( .A(fsmsta[1]), .Y(n444) );
  NAND3X1 U301 ( .A(n440), .B(n444), .C(fsmsta[2]), .Y(n378) );
  NAND2X1 U302 ( .A(n92), .B(sdao), .Y(n360) );
  NAND2X1 U303 ( .A(fsmsta[4]), .B(n441), .Y(n301) );
  NOR3XL U304 ( .A(n80), .B(fsmmod[2]), .C(n79), .Y(n143) );
  NOR2X1 U305 ( .A(n444), .B(fsmsta[0]), .Y(n307) );
  NAND2X1 U306 ( .A(fsmsta[0]), .B(n8), .Y(n292) );
  NOR3XL U307 ( .A(fsmmod[0]), .B(fsmmod[2]), .C(n79), .Y(n334) );
  NOR3XL U308 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(n80), .Y(n341) );
  OAI211X1 U309 ( .C(n10), .D(n410), .A(n411), .B(n412), .Y(n401) );
  AOI32X1 U310 ( .A(n92), .B(n408), .C(n439), .D(n415), .E(n98), .Y(n411) );
  AOI22X1 U311 ( .A(n413), .B(n84), .C(sdao), .D(n405), .Y(n412) );
  AOI21X1 U312 ( .B(n81), .C(n416), .A(n417), .Y(n410) );
  NAND2X1 U313 ( .A(fsmsta[3]), .B(n443), .Y(n303) );
  AOI221XL U314 ( .A(n364), .B(n186), .C(n374), .D(n362), .E(n375), .Y(n373)
         );
  OAI22X1 U315 ( .A(ack), .B(n376), .C(n441), .D(n309), .Y(n375) );
  INVX1 U316 ( .A(fsmmod[0]), .Y(n80) );
  AOI32X1 U317 ( .A(pedetect), .B(n196), .C(n92), .D(n197), .E(n85), .Y(n194)
         );
  OAI22X1 U318 ( .A(n69), .B(n198), .C(n199), .D(n70), .Y(n197) );
  NOR2X1 U319 ( .A(n93), .B(n200), .Y(n199) );
  NAND3X1 U320 ( .A(fsmsta[2]), .B(n440), .C(n307), .Y(n377) );
  INVX1 U321 ( .A(fsmmod[2]), .Y(n83) );
  INVX1 U322 ( .A(fsmmod[1]), .Y(n79) );
  OAI211X1 U323 ( .C(adrcomp), .D(n365), .A(n366), .B(n367), .Y(N1026) );
  AOI21X1 U324 ( .B(n368), .C(n369), .A(n370), .Y(n367) );
  NAND4X1 U325 ( .A(n371), .B(n229), .C(n372), .D(n373), .Y(n369) );
  AOI22X1 U326 ( .A(n381), .B(n361), .C(n382), .D(sdaint), .Y(n372) );
  AND3X1 U327 ( .A(fsmdet[0]), .B(n96), .C(fsmdet[1]), .Y(n188) );
  GEN2XL U328 ( .D(framesync[3]), .E(n281), .C(n141), .B(n282), .A(n283), .Y(
        N495) );
  AO2222XL U329 ( .A(n121), .B(n451), .C(i2ccon_o[1]), .D(n122), .E(
        i2ccon_o[0]), .F(n123), .G(clk_count1[0]), .H(n116), .Y(n117) );
  XNOR2XL U330 ( .A(i2cdat_o[0]), .B(i2cadr_o[1]), .Y(n165) );
  NAND21X1 U331 ( .B(i2ccon_o[2]), .A(n82), .Y(n408) );
  XNOR2XL U332 ( .A(i2cdat_o[5]), .B(i2cadr_o[6]), .Y(n160) );
  XNOR2XL U333 ( .A(i2cdat_o[2]), .B(i2cadr_o[3]), .Y(n161) );
  XNOR2XL U334 ( .A(i2cdat_o[3]), .B(i2cadr_o[4]), .Y(n162) );
  AOI21X1 U335 ( .B(n77), .C(i2ccon_o[4]), .A(n278), .Y(n112) );
  NAND2X1 U336 ( .A(n139), .B(framesync[3]), .Y(n237) );
  OAI31XL U337 ( .A(n326), .B(fsmsta[3]), .C(n105), .D(n327), .Y(n140) );
  OAI21X1 U338 ( .B(fsmsta[4]), .C(n444), .A(fsmsta[2]), .Y(n326) );
  NAND2X1 U339 ( .A(sdao), .B(n82), .Y(n361) );
  AOI21X1 U340 ( .B(n71), .C(i2ccon_o[3]), .A(n278), .Y(n289) );
  INVX1 U341 ( .A(sdaint), .Y(n82) );
  NOR31X1 U342 ( .C(framesync[0]), .A(framesync[1]), .B(framesync[2]), .Y(n139) );
  NAND3X1 U343 ( .A(n433), .B(n85), .C(n78), .Y(n365) );
  OAI32X1 U344 ( .A(n90), .B(i2ccon_o[3]), .C(framesync[3]), .D(i2ccon_o[3]), 
        .E(n237), .Y(n433) );
  OAI211X1 U345 ( .C(sclint), .D(n276), .A(n277), .B(n112), .Y(n274) );
  OAI21X1 U346 ( .B(fsmsync[0]), .C(fsmsync[2]), .A(n63), .Y(n277) );
  AOI22AXL U347 ( .A(n130), .B(sclo_int), .D(n107), .C(busfree), .Y(n276) );
  NAND2X1 U348 ( .A(fsmsta[3]), .B(fsmsta[4]), .Y(n308) );
  NOR3XL U349 ( .A(n80), .B(fsmmod[1]), .C(n83), .Y(n107) );
  OAI33XL U350 ( .A(n39), .B(n23), .C(n40), .D(n58), .E(rst_delay), .F(n114), 
        .Y(n505) );
  INVX1 U351 ( .A(rst_delay), .Y(n39) );
  AOI221XL U352 ( .A(n115), .B(n116), .C(n117), .D(n446), .E(n118), .Y(n114)
         );
  NOR43XL U353 ( .B(n119), .C(n120), .D(n451), .A(n446), .Y(n118) );
  INVX1 U354 ( .A(sclint), .Y(n71) );
  OAI32X1 U355 ( .A(n225), .B(n22), .C(n67), .D(clk_count2[0]), .E(n58), .Y(
        N685) );
  NAND2X1 U356 ( .A(sclint), .B(n26), .Y(n178) );
  NAND2X1 U357 ( .A(clk_count1_ov), .B(n125), .Y(n256) );
  INVX1 U358 ( .A(ack), .Y(n84) );
  NAND4X1 U359 ( .A(n452), .B(n450), .C(n449), .D(n414), .Y(n156) );
  NOR4XL U360 ( .A(i2cdat_o[6]), .B(i2cdat_o[5]), .C(i2cdat_o[4]), .D(
        i2cdat_o[3]), .Y(n414) );
  NAND2X1 U361 ( .A(n125), .B(n268), .Y(n264) );
  OAI211X1 U362 ( .C(i2ccon_o[7]), .D(n121), .A(n119), .B(n269), .Y(n268) );
  AOI32X1 U363 ( .A(n270), .B(n446), .C(n271), .D(n115), .E(n73), .Y(n269) );
  AOI22X1 U364 ( .A(i2ccon_o[0]), .B(n123), .C(i2ccon_o[1]), .D(n122), .Y(n271) );
  NAND3X1 U365 ( .A(nedetect), .B(n237), .C(n289), .Y(n291) );
  INVX1 U366 ( .A(adrcomp), .Y(n70) );
  OAI211X1 U367 ( .C(n287), .D(n288), .A(n187), .B(n289), .Y(n283) );
  AOI21X1 U368 ( .B(i2ccon_o[5]), .C(n294), .A(n239), .Y(n287) );
  AOI22AXL U369 ( .A(n93), .B(n290), .D(n291), .C(n92), .Y(n288) );
  OAI211X1 U370 ( .C(fsmsta[0]), .D(n438), .A(n292), .B(n293), .Y(n290) );
  OAI21X1 U371 ( .B(n110), .C(n89), .A(n25), .Y(n506) );
  AOI211X1 U372 ( .C(sclint), .D(n55), .A(n111), .B(busfree), .Y(n110) );
  INVX1 U373 ( .A(n113), .Y(n55) );
  NAND2X1 U374 ( .A(i2ccon_o[6]), .B(n112), .Y(n111) );
  OAI21X1 U375 ( .B(rst_delay), .C(n275), .A(n26), .Y(N653) );
  NOR4XL U376 ( .A(n120), .B(n274), .C(n270), .D(n446), .Y(n275) );
  AOI211X1 U377 ( .C(n70), .D(n148), .A(n149), .B(n85), .Y(n501) );
  OAI211X1 U378 ( .C(n150), .D(n447), .A(n151), .B(n24), .Y(n149) );
  NAND4X1 U379 ( .A(nedetect), .B(n141), .C(i2ccon_o[2]), .D(n153), .Y(n148)
         );
  OAI31XL U380 ( .A(n101), .B(n152), .C(n104), .D(i2ccon_o[3]), .Y(n151) );
  OAI21BBX1 U381 ( .A(clk_count1[3]), .B(n266), .C(n272), .Y(n122) );
  AOI21X1 U382 ( .B(fsmsta[3]), .C(fsmsta[1]), .A(n443), .Y(n293) );
  NOR3XL U383 ( .A(n137), .B(ack_bit), .C(n138), .Y(n136) );
  NAND2X1 U384 ( .A(fsmdet[0]), .B(n95), .Y(n351) );
  NAND2X1 U385 ( .A(clk_count1[3]), .B(clk_count1[2]), .Y(n272) );
  INVX1 U386 ( .A(fsmsta[0]), .Y(n100) );
  ENOX1 U387 ( .A(n131), .B(n132), .C(n131), .D(sdao), .Y(n502) );
  AOI211X1 U388 ( .C(n141), .D(nedetect), .A(n133), .B(n142), .Y(n131) );
  AOI211X1 U389 ( .C(n133), .D(n134), .A(n135), .B(n136), .Y(n132) );
  OR2X1 U390 ( .A(n138), .B(n135), .Y(n142) );
  ENOX1 U391 ( .A(n267), .B(n264), .C(n25), .D(n238), .Y(N656) );
  XNOR2XL U392 ( .A(n266), .B(clk_count1[2]), .Y(n267) );
  INVX1 U393 ( .A(fsmdet[2]), .Y(n96) );
  INVX1 U394 ( .A(fsmdet[1]), .Y(n95) );
  OAI211X1 U395 ( .C(n354), .D(n59), .A(n24), .B(n355), .Y(N1027) );
  AOI22X1 U396 ( .A(n60), .B(ack), .C(n78), .D(n85), .Y(n355) );
  NOR3XL U397 ( .A(n356), .B(n357), .C(n358), .Y(n354) );
  ENOX1 U398 ( .A(n359), .B(n360), .C(n361), .D(n362), .Y(n358) );
  NOR2X1 U399 ( .A(n186), .B(sdao), .Y(n393) );
  NAND2X1 U400 ( .A(n103), .B(fsmsta[3]), .Y(n300) );
  OAI21AX1 U401 ( .B(framesync[0]), .C(n35), .A(n283), .Y(N492) );
  INVX1 U402 ( .A(clk_count1[1]), .Y(n75) );
  INVX1 U403 ( .A(clk_count1[0]), .Y(n65) );
  INVX1 U404 ( .A(i2cdat_o[1]), .Y(n452) );
  NOR2X1 U405 ( .A(n37), .B(setup_counter_r[0]), .Y(N333) );
  INVX1 U406 ( .A(framesync[3]), .Y(n97) );
  NAND4X1 U407 ( .A(n163), .B(n164), .C(n165), .D(n166), .Y(n158) );
  XNOR2XL U408 ( .A(i2cdat_o[6]), .B(i2cadr_o[7]), .Y(n164) );
  XNOR2XL U409 ( .A(i2cdat_o[1]), .B(i2cadr_o[2]), .Y(n163) );
  XNOR2XL U410 ( .A(i2cdat_o[4]), .B(i2cadr_o[5]), .Y(n166) );
  INVX1 U411 ( .A(i2cdat_o[0]), .Y(n449) );
  INVX1 U412 ( .A(i2cdat_o[2]), .Y(n450) );
  AOI22AXL U413 ( .A(n38), .B(n314), .D(n317), .C(n178), .Y(n316) );
  NOR2X1 U414 ( .A(n22), .B(test_so2), .Y(n317) );
  INVX1 U415 ( .A(adrcompen), .Y(n61) );
  NAND2X1 U416 ( .A(n124), .B(n125), .Y(n504) );
  XNOR2XL U417 ( .A(clkint), .B(clk_count2_ov), .Y(n124) );
  NOR2X1 U418 ( .A(n263), .B(n264), .Y(N657) );
  XNOR2XL U419 ( .A(clk_count1[3]), .B(n265), .Y(n263) );
  AND2X1 U420 ( .A(clk_count1[2]), .B(n266), .Y(n265) );
  NOR2X1 U421 ( .A(clk_count1[0]), .B(n264), .Y(N654) );
  NOR2X1 U422 ( .A(n262), .B(n256), .Y(N687) );
  XNOR2XL U423 ( .A(n261), .B(clk_count2[2]), .Y(n262) );
  NOR2X1 U424 ( .A(n259), .B(n256), .Y(N688) );
  XNOR2XL U425 ( .A(clk_count2[3]), .B(n260), .Y(n259) );
  AND2X1 U426 ( .A(clk_count2[2]), .B(n261), .Y(n260) );
  NOR2X1 U427 ( .A(n255), .B(n256), .Y(N690) );
  AOI22X1 U428 ( .A(clk_count2[0]), .B(n257), .C(i2ccon_o[7]), .D(i2ccon_o[1]), 
        .Y(n255) );
  ENOX1 U429 ( .A(n258), .B(n48), .C(i2ccon_o[0]), .D(i2ccon_o[7]), .Y(n257)
         );
  AOI21X1 U430 ( .B(clk_count2[3]), .C(clk_count2[2]), .A(n446), .Y(n258) );
  INVX1 U431 ( .A(n315), .Y(n36) );
  AOI32X1 U432 ( .A(setup_counter_r[1]), .B(n316), .C(setup_counter_r[0]), .D(
        n42), .E(N333), .Y(n315) );
  INVX1 U433 ( .A(setup_counter_r[1]), .Y(n42) );
  AOI31X1 U434 ( .A(n50), .B(n44), .C(n49), .D(test_so1), .Y(n177) );
  NAND31X1 U435 ( .C(n278), .A(n345), .B(n170), .Y(n332) );
  NAND3X1 U436 ( .A(n10), .B(pedetect), .C(n101), .Y(n345) );
  NOR21XL U437 ( .B(bclkcnt[1]), .A(n11), .Y(n120) );
  XNOR2XL U438 ( .A(bclksel), .B(bclkcnt[0]), .Y(n11) );
  INVX1 U439 ( .A(i2ccon_o[3]), .Y(n33) );
  NAND2X1 U440 ( .A(clkint_ff), .B(n64), .Y(n221) );
  NOR2X1 U441 ( .A(n64), .B(clkint_ff), .Y(n246) );
  NAND2X1 U442 ( .A(i2ccon_o[1]), .B(i2ccon_o[0]), .Y(n270) );
  NAND3X1 U443 ( .A(indelay[1]), .B(n54), .C(indelay[2]), .Y(n251) );
  NAND2X1 U444 ( .A(framesync[1]), .B(framesync[0]), .Y(n285) );
  NOR3XL U445 ( .A(clk_count1[1]), .B(clk_count1[2]), .C(clk_count1[0]), .Y(
        n273) );
  INVX1 U446 ( .A(i2ccon_o[7]), .Y(n446) );
  NOR3XL U447 ( .A(fsmmod[0]), .B(fsmmod[1]), .C(n83), .Y(n130) );
  INVX1 U448 ( .A(fsmsync[0]), .Y(n68) );
  INVX1 U449 ( .A(pedetect), .Y(n66) );
  INVX1 U450 ( .A(i2ccon_o[6]), .Y(n445) );
  NOR2X1 U451 ( .A(n281), .B(framesync[3]), .Y(n141) );
  INVX1 U452 ( .A(fsmsync[1]), .Y(n63) );
  OAI221X1 U453 ( .A(fsmsta[1]), .B(n309), .C(fsmsta[0]), .D(n442), .E(n298), 
        .Y(N406) );
  AOI31X1 U454 ( .A(scli_ff_reg0[2]), .B(N414), .C(N413), .D(n43), .Y(n180) );
  OAI21X1 U455 ( .B(n35), .C(n286), .A(n187), .Y(N493) );
  OAI21X1 U456 ( .B(framesync[1]), .C(framesync[0]), .A(n285), .Y(n286) );
  OAI21X1 U457 ( .B(n223), .C(n224), .A(n170), .Y(N749) );
  NOR21XL U458 ( .B(n225), .A(n226), .Y(n224) );
  AOI211X1 U459 ( .C(n442), .D(fsmsta[1]), .A(n227), .B(n9), .Y(n223) );
  OAI211X1 U460 ( .C(fsmsta[4]), .D(n228), .A(n229), .B(n71), .Y(n227) );
  OAI21X1 U461 ( .B(n108), .C(n82), .A(n109), .Y(n507) );
  NOR3XL U462 ( .A(sdai_ff_reg0[0]), .B(sdai_ff_reg0[2]), .C(sdai_ff_reg0[1]), 
        .Y(n108) );
  AOI31X1 U463 ( .A(sdai_ff_reg0[1]), .B(sdai_ff_reg0[0]), .C(sdai_ff_reg0[2]), 
        .D(n22), .Y(n109) );
  OAI21X1 U464 ( .B(n284), .C(n35), .A(n187), .Y(N494) );
  XNOR2XL U465 ( .A(n94), .B(framesync[2]), .Y(n284) );
  AOI32X1 U466 ( .A(n93), .B(n294), .C(n334), .D(starto_en), .E(n76), .Y(n346)
         );
  NOR2X1 U467 ( .A(n240), .B(n233), .Y(N747) );
  AOI221XL U468 ( .A(n238), .B(n33), .C(fsmsync[1]), .D(n241), .E(n242), .Y(
        n240) );
  OAI211X1 U469 ( .C(n47), .D(n68), .A(n247), .B(n67), .Y(n241) );
  AOI211X1 U470 ( .C(n68), .D(n243), .A(fsmsync[2]), .B(fsmsync[1]), .Y(n242)
         );
  AOI211X1 U471 ( .C(n45), .D(n221), .A(n222), .B(n107), .Y(n490) );
  INVX1 U472 ( .A(starto_en), .Y(n45) );
  NAND21X1 U473 ( .B(n178), .A(busfree), .Y(n222) );
  INVX1 U474 ( .A(clkint), .Y(n64) );
  GEN2XL U475 ( .D(n62), .E(n53), .C(N469), .B(indelay[2]), .A(n295), .Y(N471)
         );
  NOR4XL U476 ( .A(indelay[2]), .B(n53), .C(n296), .D(n54), .Y(n295) );
  INVX1 U477 ( .A(indelay[1]), .Y(n53) );
  OAI21X1 U478 ( .B(n177), .C(n178), .A(n179), .Y(n498) );
  NAND41X1 U479 ( .D(n180), .A(n177), .B(nedetect), .C(n27), .Y(n179) );
  NOR3XL U480 ( .A(n250), .B(sdaint), .C(n221), .Y(n338) );
  AOI22X1 U481 ( .A(n184), .B(n185), .C(i2ccon_o[4]), .D(n77), .Y(n496) );
  NAND2X1 U482 ( .A(n188), .B(n24), .Y(n184) );
  OAI211X1 U483 ( .C(n72), .D(n7), .A(n187), .B(adrcompen), .Y(n185) );
  AOI21X1 U484 ( .B(n248), .C(n249), .A(n233), .Y(N746) );
  AOI211X1 U485 ( .C(n226), .D(n251), .A(n252), .B(n253), .Y(n249) );
  AOI22X1 U486 ( .A(n238), .B(n254), .C(n234), .D(n32), .Y(n248) );
  AOI211X1 U487 ( .C(sdaint), .D(n68), .A(n67), .B(n63), .Y(n253) );
  AOI21X1 U488 ( .B(n231), .C(n232), .A(n233), .Y(N748) );
  AOI22X1 U489 ( .A(n238), .B(n239), .C(fsmsync[2]), .D(fsmsync[1]), .Y(n231)
         );
  AOI22X1 U490 ( .A(n234), .B(n235), .C(n236), .D(n71), .Y(n232) );
  ENOX1 U491 ( .A(fsmsync[0]), .B(n67), .C(n226), .D(n47), .Y(n236) );
  AOI21X1 U492 ( .B(n339), .C(n340), .A(n332), .Y(N1125) );
  AOI22X1 U493 ( .A(n334), .B(n32), .C(n341), .D(nedetect), .Y(n339) );
  OAI2B11X1 U494 ( .D(test_so2), .C(sclint), .A(n37), .B(n24), .Y(N332) );
  OAI211X1 U495 ( .C(n244), .D(n245), .A(sclint), .B(n246), .Y(n243) );
  AOI22X1 U496 ( .A(fsmmod[2]), .B(n80), .C(fsmmod[1]), .D(fsmmod[0]), .Y(n245) );
  OAI211X1 U497 ( .C(n302), .D(n303), .A(n298), .B(n304), .Y(N409) );
  AOI32X1 U498 ( .A(fsmsta[3]), .B(n444), .C(n98), .D(n302), .E(n441), .Y(n304) );
  NOR2X1 U499 ( .A(n230), .B(n438), .Y(n302) );
  INVX1 U500 ( .A(clk_count1[3]), .Y(n74) );
  AOI31X1 U501 ( .A(n329), .B(n330), .C(n331), .D(n332), .Y(N1126) );
  OAI21X1 U502 ( .B(n221), .C(n71), .A(n130), .Y(n330) );
  AOI32X1 U503 ( .A(sclint), .B(n336), .C(n143), .D(n337), .E(n338), .Y(n329)
         );
  AOI222XL U504 ( .A(n244), .B(n72), .C(n107), .D(n333), .E(n334), .F(n335), 
        .Y(n331) );
  AOI31X1 U505 ( .A(n342), .B(n343), .C(n344), .D(n332), .Y(N1124) );
  AOI22X1 U506 ( .A(n107), .B(n333), .C(n341), .D(n72), .Y(n344) );
  OAI21BBX1 U507 ( .A(n336), .B(sclint), .C(n143), .Y(n342) );
  NAND42X1 U508 ( .C(n346), .D(n239), .A(n56), .B(i2ccon_o[5]), .Y(n343) );
  INVX1 U509 ( .A(scli_ff_reg0[0]), .Y(n50) );
  NAND2X1 U510 ( .A(i2ccon_o[4]), .B(n33), .Y(n254) );
  INVX1 U511 ( .A(scli_ff_reg0[1]), .Y(n49) );
  NAND2X1 U512 ( .A(framesync[2]), .B(n94), .Y(n281) );
  NOR2X1 U513 ( .A(setup_counter_r[1]), .B(setup_counter_r[0]), .Y(n314) );
  INVX1 U514 ( .A(indelay[0]), .Y(n54) );
  NOR2X1 U515 ( .A(n296), .B(indelay[0]), .Y(N469) );
  NAND2X1 U516 ( .A(n25), .B(n183), .Y(n176) );
  NAND4X1 U517 ( .A(scli_ff_reg0[2]), .B(scli_ff_reg0[1]), .C(scli_ff_reg0[0]), 
        .D(n177), .Y(n183) );
  INVX1 U518 ( .A(scli_ff_reg0[2]), .Y(n44) );
  INVX1 U519 ( .A(i2cadr_o[0]), .Y(n448) );
  INVX1 U520 ( .A(bsd7_tmp), .Y(n52) );
  NOR32XL U521 ( .B(starto_en), .C(i2ccon_o[5]), .A(n239), .Y(n337) );
  NOR2X1 U522 ( .A(n347), .B(n178), .Y(N1065) );
  AOI221XL U523 ( .A(fsmdet[1]), .B(sdaint), .C(fsmdet[2]), .D(n95), .E(n188), 
        .Y(n347) );
  NOR3XL U524 ( .A(n68), .B(fsmsync[1]), .C(n67), .Y(n238) );
  NOR4XL U525 ( .A(n57), .B(n63), .C(fsmsync[0]), .D(fsmsync[2]), .Y(n234) );
  INVX1 U526 ( .A(fsmsync[2]), .Y(n67) );
  NOR3XL U527 ( .A(n225), .B(sclint), .C(fsmsync[2]), .Y(n252) );
  NOR3XL U528 ( .A(n279), .B(n22), .C(n120), .Y(N511) );
  XNOR2XL U529 ( .A(bclkcnt[1]), .B(bclkcnt[0]), .Y(n279) );
  NOR3XL U530 ( .A(n120), .B(n22), .C(bclkcnt[0]), .Y(N510) );
  NAND3X1 U531 ( .A(n27), .B(n71), .C(test_so2), .Y(n313) );
  AOI21BX1 U532 ( .C(n352), .B(n353), .A(n178), .Y(N1063) );
  NAND2X1 U533 ( .A(n350), .B(n82), .Y(n353) );
  OAI32X1 U534 ( .A(n350), .B(fsmdet[0]), .C(n82), .D(n351), .E(fsmdet[2]), 
        .Y(n352) );
  INVX1 U535 ( .A(i2ccon_o[4]), .Y(n447) );
  INVX1 U536 ( .A(nedetect), .Y(n72) );
  NAND2X1 U540 ( .A(sclscl), .B(pedetect), .Y(n333) );
  INVX1 U541 ( .A(clk_count2[1]), .Y(n48) );
  INVX1 U542 ( .A(clk_count2[0]), .Y(n51) );
  NOR2X1 U543 ( .A(n348), .B(n178), .Y(N1064) );
  AOI221XL U544 ( .A(fsmdet[2]), .B(fsmdet[0]), .C(n349), .D(n82), .E(n350), 
        .Y(n348) );
  OAI21X1 U545 ( .B(fsmdet[2]), .C(fsmdet[0]), .A(n351), .Y(n349) );
  NOR2X1 U546 ( .A(n297), .B(n296), .Y(N470) );
  XNOR2XL U547 ( .A(indelay[1]), .B(indelay[0]), .Y(n297) );
  OR2X1 U548 ( .A(scli_ff), .B(n23), .Y(N412) );
  OR2X1 U549 ( .A(sdai_ff_reg0[0]), .B(n23), .Y(N432) );
  OR2X1 U550 ( .A(sdai_ff), .B(n23), .Y(N431) );
  OR2X1 U551 ( .A(sdai_ff_reg0[1]), .B(n23), .Y(N433) );
  INVX1 U552 ( .A(n106), .Y(n46) );
  OAI211X1 U553 ( .C(sclscl), .D(pedetect), .A(n107), .B(n24), .Y(n106) );
  INVX1 U554 ( .A(bsd7), .Y(n41) );
  INVX1 U555 ( .A(setup_counter_r[2]), .Y(n38) );
  INVX1 U556 ( .A(clk_count1_ov), .Y(n40) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module extint_a0 ( clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, 
        int2ff, iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, 
        int6ff, iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, 
        ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7, 
        iex8, iex9, iex10, iex11, iex12, sfraddr, sfrdatai, sfrwe, test_si, 
        test_se );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, int2ff,
         iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, int6ff,
         iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, sfrwe,
         test_si, test_se;
  output ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12;
  wire   int0_ff1, int0_fall, int0_clr, N23, int1_ff1, int1_fall, int1_clr,
         N51, int2_ff1, iex2_set, N71, int3_ff1, iex3_set, N90, iex4_set,
         int4_ff1, iex5_set, int5_ff1, iex6_set, int6_ff1, iex7_set, int7_ff1,
         iex8_set, int8_ff1, iex9_set, int9_ff1, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n85, n86, n87, n88, n89, n90, n91, n92, n93;

  SDFFQX1 int4_ff1_reg ( .D(n23), .SIN(int3_ff1), .SMC(test_se), .C(clkper), 
        .Q(int4_ff1) );
  SDFFQX1 int5_ff1_reg ( .D(n16), .SIN(int4_ff1), .SMC(test_se), .C(clkper), 
        .Q(int5_ff1) );
  SDFFQX1 int6_ff1_reg ( .D(n13), .SIN(int5_ff1), .SMC(test_se), .C(clkper), 
        .Q(int6_ff1) );
  SDFFQX1 int7_ff1_reg ( .D(n15), .SIN(int6_ff1), .SMC(test_se), .C(clkper), 
        .Q(int7_ff1) );
  SDFFQX1 int8_ff1_reg ( .D(n93), .SIN(int7_ff1), .SMC(test_se), .C(clkper), 
        .Q(int8_ff1) );
  SDFFQX1 int9_ff1_reg ( .D(n14), .SIN(int8_ff1), .SMC(test_se), .C(clkper), 
        .Q(int9_ff1) );
  SDFFQX1 iex6_set_reg ( .D(n101), .SIN(iex6), .SMC(test_se), .C(clkper), .Q(
        iex6_set) );
  SDFFQX1 iex7_set_reg ( .D(n99), .SIN(iex7), .SMC(test_se), .C(clkper), .Q(
        iex7_set) );
  SDFFQX1 iex8_set_reg ( .D(n97), .SIN(iex8), .SMC(test_se), .C(clkper), .Q(
        iex8_set) );
  SDFFQX1 iex9_set_reg ( .D(n95), .SIN(iex9), .SMC(test_se), .C(clkper), .Q(
        iex9_set) );
  SDFFQX1 iex4_set_reg ( .D(n105), .SIN(iex4), .SMC(test_se), .C(clkper), .Q(
        iex4_set) );
  SDFFQX1 iex5_set_reg ( .D(n103), .SIN(iex5), .SMC(test_se), .C(clkper), .Q(
        iex5_set) );
  SDFFQX1 int0_ff1_reg ( .D(N23), .SIN(int0_fall), .SMC(test_se), .C(clkper), 
        .Q(int0_ff1) );
  SDFFQX1 int1_ff1_reg ( .D(N51), .SIN(int1_fall), .SMC(test_se), .C(clkper), 
        .Q(int1_ff1) );
  SDFFQX1 iex2_set_reg ( .D(n110), .SIN(iex2), .SMC(test_se), .C(clkper), .Q(
        iex2_set) );
  SDFFQX1 iex3_set_reg ( .D(n107), .SIN(iex3), .SMC(test_se), .C(clkper), .Q(
        iex3_set) );
  SDFFQX1 int0_clr_reg ( .D(n118), .SIN(iex9_set), .SMC(test_se), .C(clkper), 
        .Q(int0_clr) );
  SDFFQX1 int1_clr_reg ( .D(n114), .SIN(int0_ff1), .SMC(test_se), .C(clkper), 
        .Q(int1_clr) );
  SDFFQX1 int2_ff1_reg ( .D(N71), .SIN(int1_ff1), .SMC(test_se), .C(clkper), 
        .Q(int2_ff1) );
  SDFFQX1 int3_ff1_reg ( .D(N90), .SIN(int2_ff1), .SMC(test_se), .C(clkper), 
        .Q(int3_ff1) );
  SDFFQX1 int0_fall_reg ( .D(n116), .SIN(int0_clr), .SMC(test_se), .C(clkper), 
        .Q(int0_fall) );
  SDFFQX1 int1_fall_reg ( .D(n112), .SIN(int1_clr), .SMC(test_se), .C(clkper), 
        .Q(int1_fall) );
  SDFFQX1 i3fr_s_reg ( .D(n108), .SIN(i2fr), .SMC(test_se), .C(clkper), .Q(
        i3fr) );
  SDFFQX1 i2fr_s_reg ( .D(n17), .SIN(test_si), .SMC(test_se), .C(clkper), .Q(
        i2fr) );
  SDFFQX1 iex6_s_reg ( .D(n100), .SIN(iex5_set), .SMC(test_se), .C(clkper), 
        .Q(iex6) );
  SDFFQX1 iex9_s_reg ( .D(n94), .SIN(iex8_set), .SMC(test_se), .C(clkper), .Q(
        iex9) );
  SDFFQX1 iex5_s_reg ( .D(n102), .SIN(iex4_set), .SMC(test_se), .C(clkper), 
        .Q(iex5) );
  SDFFQX1 iex8_s_reg ( .D(n96), .SIN(iex7_set), .SMC(test_se), .C(clkper), .Q(
        iex8) );
  SDFFQX1 ie1_s_reg ( .D(n111), .SIN(ie0), .SMC(test_se), .C(clkper), .Q(ie1)
         );
  SDFFQX1 iex4_s_reg ( .D(n104), .SIN(iex3_set), .SMC(test_se), .C(clkper), 
        .Q(iex4) );
  SDFFQX1 iex2_s_reg ( .D(n109), .SIN(ie1), .SMC(test_se), .C(clkper), .Q(iex2) );
  SDFFQX1 ie0_s_reg ( .D(n115), .SIN(i3fr), .SMC(test_se), .C(clkper), .Q(ie0)
         );
  SDFFQX1 iex7_s_reg ( .D(n98), .SIN(iex6_set), .SMC(test_se), .C(clkper), .Q(
        iex7) );
  SDFFQX1 iex3_s_reg ( .D(n106), .SIN(iex2_set), .SMC(test_se), .C(clkper), 
        .Q(iex3) );
  SDFFQX1 it1_s_reg ( .D(n113), .SIN(it0), .SMC(test_se), .C(clkper), .Q(it1)
         );
  SDFFQX1 it0_s_reg ( .D(n117), .SIN(int9_ff1), .SMC(test_se), .C(clkper), .Q(
        it0) );
  INVX1 U3 ( .A(1'b1), .Y(iex12) );
  INVX1 U5 ( .A(1'b1), .Y(iex11) );
  INVX1 U7 ( .A(1'b1), .Y(iex10) );
  INVX1 U9 ( .A(n46), .Y(n18) );
  INVX1 U10 ( .A(n11), .Y(n9) );
  NOR2X1 U11 ( .A(n82), .B(n10), .Y(n46) );
  AND2X1 U12 ( .A(n82), .B(n9), .Y(n48) );
  INVX1 U13 ( .A(n59), .Y(n20) );
  INVX1 U14 ( .A(n57), .Y(n19) );
  INVX1 U15 ( .A(n51), .Y(n21) );
  INVX1 U16 ( .A(n12), .Y(n10) );
  INVX1 U17 ( .A(n12), .Y(n11) );
  NOR43XL U18 ( .B(sfrwe), .C(n75), .D(sfraddr[3]), .A(sfraddr[0]), .Y(n70) );
  NOR4XL U19 ( .A(sfraddr[5]), .B(sfraddr[4]), .C(sfraddr[2]), .D(sfraddr[1]), 
        .Y(n75) );
  NAND21X1 U20 ( .B(sfraddr[6]), .A(n70), .Y(n59) );
  AOI21X1 U21 ( .B(sfraddr[6]), .C(n70), .A(n11), .Y(n57) );
  NAND2X1 U22 ( .A(n54), .B(n55), .Y(n51) );
  AND4X1 U23 ( .A(sfraddr[2]), .B(sfraddr[3]), .C(sfraddr[4]), .D(sfraddr[5]), 
        .Y(n54) );
  NOR43XL U24 ( .B(sfraddr[1]), .C(sfrwe), .D(sfraddr[0]), .A(sfraddr[6]), .Y(
        n55) );
  NAND4X1 U25 ( .A(sfrwe), .B(sfraddr[6]), .C(n83), .D(n84), .Y(n82) );
  NOR2X1 U26 ( .A(sfraddr[1]), .B(sfraddr[0]), .Y(n83) );
  NOR4XL U27 ( .A(sfraddr[5]), .B(sfraddr[4]), .C(sfraddr[3]), .D(sfraddr[2]), 
        .Y(n84) );
  INVX1 U28 ( .A(n60), .Y(n22) );
  INVX1 U29 ( .A(sfrdatai[1]), .Y(n7) );
  INVX1 U30 ( .A(sfrdatai[3]), .Y(n8) );
  INVX1 U31 ( .A(n45), .Y(n15) );
  INVX1 U32 ( .A(rst), .Y(n12) );
  INVX1 U33 ( .A(iex8ack), .Y(n89) );
  INVX1 U34 ( .A(iex9ack), .Y(n90) );
  INVX1 U35 ( .A(n44), .Y(n93) );
  INVX1 U36 ( .A(n43), .Y(n16) );
  INVX1 U37 ( .A(n41), .Y(n23) );
  INVX1 U38 ( .A(n42), .Y(n14) );
  NOR2X1 U39 ( .A(n10), .B(newinstr), .Y(n60) );
  OAI22X1 U40 ( .A(n11), .B(n37), .C(n22), .D(n33), .Y(n114) );
  OAI22X1 U41 ( .A(n11), .B(n36), .C(n22), .D(n32), .Y(n118) );
  NAND2X1 U42 ( .A(int7ff), .B(n9), .Y(n45) );
  NAND21X1 U43 ( .B(int2ff), .A(n9), .Y(N71) );
  NAND21X1 U44 ( .B(int3ff), .A(n9), .Y(N90) );
  INVX1 U45 ( .A(int0ack), .Y(n36) );
  INVX1 U46 ( .A(int1ack), .Y(n37) );
  INVX1 U47 ( .A(iex3ack), .Y(n85) );
  INVX1 U48 ( .A(iex2ack), .Y(n39) );
  INVX1 U49 ( .A(n40), .Y(n13) );
  NAND2X1 U50 ( .A(int8ff), .B(n9), .Y(n44) );
  NOR2X1 U51 ( .A(n10), .B(n92), .Y(N23) );
  NOR2X1 U52 ( .A(n11), .B(n91), .Y(N51) );
  NAND2X1 U53 ( .A(int5ff), .B(n9), .Y(n43) );
  OAI32X1 U54 ( .A(n31), .B(iex5ack), .C(n22), .D(int5_ff1), .E(n43), .Y(n103)
         );
  INVX1 U55 ( .A(iex5_set), .Y(n31) );
  NAND2X1 U56 ( .A(int9ff), .B(n9), .Y(n42) );
  NAND2X1 U57 ( .A(int4ff), .B(n9), .Y(n41) );
  OAI32X1 U58 ( .A(n30), .B(iex4ack), .C(n22), .D(int4_ff1), .E(n41), .Y(n105)
         );
  INVX1 U59 ( .A(iex4_set), .Y(n30) );
  OAI32X1 U60 ( .A(n27), .B(iex9ack), .C(n22), .D(int9_ff1), .E(n42), .Y(n95)
         );
  INVX1 U61 ( .A(iex9_set), .Y(n27) );
  NOR2X1 U62 ( .A(n10), .B(n58), .Y(n117) );
  AOI22X1 U63 ( .A(n20), .B(sfrdatai[0]), .C(it0), .D(n59), .Y(n58) );
  NOR2X1 U64 ( .A(n10), .B(n65), .Y(n113) );
  AOI22X1 U65 ( .A(sfrdatai[2]), .B(n20), .C(it1), .D(n59), .Y(n65) );
  NOR21XL U66 ( .B(n61), .A(n10), .Y(n115) );
  OAI22X1 U67 ( .A(n7), .B(n59), .C(n20), .D(n62), .Y(n61) );
  AOI32X1 U68 ( .A(n32), .B(n36), .C(n63), .D(n92), .E(n35), .Y(n62) );
  ENOX1 U69 ( .A(n64), .B(n35), .C(n92), .D(int0_ff1), .Y(n63) );
  NOR21XL U70 ( .B(n66), .A(n10), .Y(n111) );
  OAI22X1 U71 ( .A(n59), .B(n8), .C(n20), .D(n67), .Y(n66) );
  AOI32X1 U72 ( .A(n33), .B(n37), .C(n68), .D(n91), .E(n34), .Y(n67) );
  ENOX1 U73 ( .A(n69), .B(n34), .C(n91), .D(int1_ff1), .Y(n68) );
  OAI21X1 U74 ( .B(n18), .C(n7), .A(n73), .Y(n109) );
  OAI211X1 U75 ( .C(iex2), .D(iex2_set), .A(n39), .B(n48), .Y(n73) );
  OAI21X1 U76 ( .B(n18), .C(n8), .A(n79), .Y(n104) );
  OAI211X1 U77 ( .C(iex4), .D(iex4_set), .A(n86), .B(n48), .Y(n79) );
  INVX1 U78 ( .A(iex4ack), .Y(n86) );
  AOI21X1 U79 ( .B(n52), .C(n53), .A(n11), .Y(n94) );
  NAND2X1 U80 ( .A(sfrdatai[1]), .B(n21), .Y(n52) );
  OAI211X1 U81 ( .C(iex9), .D(iex9_set), .A(n51), .B(n90), .Y(n53) );
  AOI21X1 U82 ( .B(n49), .C(n50), .A(n10), .Y(n96) );
  NAND2X1 U83 ( .A(n21), .B(sfrdatai[0]), .Y(n49) );
  OAI211X1 U84 ( .C(iex8), .D(iex8_set), .A(n51), .B(n89), .Y(n50) );
  OAI21BBX1 U85 ( .A(n46), .B(sfrdatai[5]), .C(n81), .Y(n100) );
  OAI211X1 U86 ( .C(iex6), .D(iex6_set), .A(n88), .B(n48), .Y(n81) );
  INVX1 U87 ( .A(iex6ack), .Y(n88) );
  OAI21BBX1 U88 ( .A(sfrdatai[4]), .B(n46), .C(n80), .Y(n102) );
  OAI211X1 U89 ( .C(iex5), .D(iex5_set), .A(n87), .B(n48), .Y(n80) );
  INVX1 U90 ( .A(iex5ack), .Y(n87) );
  OAI21BBX1 U91 ( .A(n46), .B(sfrdatai[2]), .C(n78), .Y(n106) );
  OAI211X1 U92 ( .C(iex3), .D(iex3_set), .A(n85), .B(n48), .Y(n78) );
  OAI21BBX1 U93 ( .A(n46), .B(sfrdatai[0]), .C(n47), .Y(n98) );
  OAI211X1 U94 ( .C(iex7), .D(iex7_set), .A(n38), .B(n48), .Y(n47) );
  INVX1 U95 ( .A(iex7ack), .Y(n38) );
  OAI21BBX1 U96 ( .A(n57), .B(i3fr), .C(n74), .Y(n108) );
  NAND3X1 U97 ( .A(n19), .B(n12), .C(sfrdatai[6]), .Y(n74) );
  INVX1 U98 ( .A(n56), .Y(n17) );
  AOI32X1 U99 ( .A(sfrdatai[5]), .B(n9), .C(n19), .D(n57), .E(i2fr), .Y(n56)
         );
  AO33X1 U100 ( .A(int1_ff1), .B(n12), .C(n91), .D(int1_fall), .E(n37), .F(n60), .Y(n112) );
  AO33X1 U101 ( .A(int0_ff1), .B(n12), .C(n92), .D(int0_fall), .E(n36), .F(n60), .Y(n116) );
  OAI32X1 U102 ( .A(n25), .B(iex7ack), .C(n22), .D(int7_ff1), .E(n45), .Y(n99)
         );
  INVX1 U103 ( .A(iex7_set), .Y(n25) );
  OAI32X1 U104 ( .A(n26), .B(iex8ack), .C(n22), .D(int8_ff1), .E(n44), .Y(n97)
         );
  INVX1 U105 ( .A(iex8_set), .Y(n26) );
  OAI32X1 U106 ( .A(n24), .B(iex6ack), .C(n22), .D(int6_ff1), .E(n40), .Y(n101) );
  INVX1 U107 ( .A(iex6_set), .Y(n24) );
  OAI31XL U108 ( .A(n29), .B(i3fr), .C(N90), .D(n76), .Y(n107) );
  INVX1 U109 ( .A(int3_ff1), .Y(n29) );
  AOI33X1 U110 ( .A(int3ff), .B(i3fr), .C(n77), .D(n60), .E(n85), .F(iex3_set), 
        .Y(n76) );
  NOR2X1 U111 ( .A(n10), .B(int3_ff1), .Y(n77) );
  OAI31XL U112 ( .A(n28), .B(i2fr), .C(N71), .D(n71), .Y(n110) );
  INVX1 U113 ( .A(int2_ff1), .Y(n28) );
  AOI33X1 U114 ( .A(int2ff), .B(i2fr), .C(n72), .D(n60), .E(n39), .F(iex2_set), 
        .Y(n71) );
  NOR2X1 U115 ( .A(n10), .B(int2_ff1), .Y(n72) );
  NAND2X1 U119 ( .A(int6ff), .B(n9), .Y(n40) );
  INVX1 U120 ( .A(int1ff), .Y(n91) );
  INVX1 U121 ( .A(int0ff), .Y(n92) );
  NOR2X1 U122 ( .A(ie0), .B(int0_fall), .Y(n64) );
  NOR2X1 U123 ( .A(ie1), .B(int1_fall), .Y(n69) );
  INVX1 U124 ( .A(it0), .Y(n35) );
  INVX1 U125 ( .A(it1), .Y(n34) );
  INVX1 U126 ( .A(int0_clr), .Y(n32) );
  INVX1 U127 ( .A(int1_clr), .Y(n33) );
endmodule


module isr_a0 ( clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, 
        t0ff, int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff, 
        int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b, 
        int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, int_vect_ab, irq, intvect, int_ack_03, int_ack_0b, 
        int_ack_13, int_ack_1b, int_ack_43, int_ack_4b, int_ack_53, int_ack_5b, 
        int_ack_63, int_ack_6b, int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, 
        int_ack_ab, is_reg, ip0, ip1, ien0, ien1, ien2, isr_tm, sfraddr, 
        sfrdatai, sfrwe, test_si, test_se );
  output [4:0] intvect;
  output [3:0] is_reg;
  output [5:0] ip0;
  output [5:0] ip1;
  output [7:0] ien0;
  output [5:0] ien1;
  output [5:0] ien2;
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, t0ff,
         int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff,
         int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b,
         int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b,
         int_vect_a3, int_vect_ab, sfrwe, test_si, test_se;
  output irq, int_ack_03, int_ack_0b, int_ack_13, int_ack_1b, int_ack_43,
         int_ack_4b, int_ack_53, int_ack_5b, int_ack_63, int_ack_6b,
         int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, int_ack_ab, isr_tm;
  wire   N38, N39, N40, N41, N42, N43, N44, N45, N49, N50, N51, N52, N53, N54,
         N55, N58, N59, N60, N61, N62, N63, N64, N67, N68, N69, N70, N71, N72,
         N73, N76, N77, N78, N79, N80, N81, N82, irq_r, N200, N207, N209, N210,
         N211, N212, net12078, net12084, net12089, net12094, net12099,
         net12104, n196, n197, n198, n199, n200, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n201, n202, n203, n204, n205, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n206, n207;

  SNPS_CLOCK_GATE_HIGH_isr_a0_0 clk_gate_ien0_reg_reg ( .CLK(clkper), .EN(N38), 
        .ENCLK(net12078), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_5 clk_gate_ien1_reg_reg ( .CLK(clkper), .EN(N49), 
        .ENCLK(net12084), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_4 clk_gate_ien2_reg_reg ( .CLK(clkper), .EN(N58), 
        .ENCLK(net12089), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_3 clk_gate_ip0_reg_reg ( .CLK(clkper), .EN(N67), 
        .ENCLK(net12094), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_2 clk_gate_ip1_reg_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12099), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_1 clk_gate_intvect_reg_reg ( .CLK(clkper), .EN(
        N207), .ENCLK(net12104), .TE(test_se) );
  SDFFQX1 intvect_reg_reg_1_ ( .D(N209), .SIN(intvect[0]), .SMC(test_se), .C(
        net12104), .Q(intvect[1]) );
  SDFFQX1 intvect_reg_reg_3_ ( .D(N211), .SIN(intvect[2]), .SMC(test_se), .C(
        net12104), .Q(intvect[3]) );
  SDFFQX1 intvect_reg_reg_0_ ( .D(n16), .SIN(ien2[5]), .SMC(test_se), .C(
        net12104), .Q(intvect[0]) );
  SDFFQX1 intvect_reg_reg_4_ ( .D(N212), .SIN(intvect[3]), .SMC(test_se), .C(
        net12104), .Q(intvect[4]) );
  SDFFQX1 intvect_reg_reg_2_ ( .D(N210), .SIN(intvect[1]), .SMC(test_se), .C(
        net12104), .Q(intvect[2]) );
  SDFFQX1 is_reg_s_reg_0_ ( .D(n199), .SIN(irq_r), .SMC(test_se), .C(clkper), 
        .Q(is_reg[0]) );
  SDFFQX1 is_reg_s_reg_1_ ( .D(n196), .SIN(is_reg[0]), .SMC(test_se), .C(
        clkper), .Q(is_reg[1]) );
  SDFFQX1 ien2_reg_reg_5_ ( .D(N64), .SIN(ien2[4]), .SMC(test_se), .C(net12089), .Q(ien2[5]) );
  SDFFQX1 ien2_reg_reg_4_ ( .D(N63), .SIN(ien2[3]), .SMC(test_se), .C(net12089), .Q(ien2[4]) );
  SDFFQX1 ip1_reg_reg_5_ ( .D(N82), .SIN(ip1[4]), .SMC(test_se), .C(net12099), 
        .Q(ip1[5]) );
  SDFFQX1 ip0_reg_reg_5_ ( .D(N73), .SIN(ip0[4]), .SMC(test_se), .C(net12094), 
        .Q(ip0[5]) );
  SDFFQX1 is_reg_s_reg_2_ ( .D(n197), .SIN(is_reg[1]), .SMC(test_se), .C(
        clkper), .Q(is_reg[2]) );
  SDFFQX1 ien0_reg_reg_5_ ( .D(N44), .SIN(ien0[4]), .SMC(test_se), .C(net12078), .Q(ien0[5]) );
  SDFFQX1 ien1_reg_reg_5_ ( .D(N55), .SIN(ien1[4]), .SMC(test_se), .C(net12084), .Q(ien1[5]) );
  SDFFQX1 ip1_reg_reg_4_ ( .D(N81), .SIN(ip1[3]), .SMC(test_se), .C(net12099), 
        .Q(ip1[4]) );
  SDFFQX1 ip0_reg_reg_4_ ( .D(N72), .SIN(ip0[3]), .SMC(test_se), .C(net12094), 
        .Q(ip0[4]) );
  SDFFQX1 is_reg_s_reg_3_ ( .D(n198), .SIN(is_reg[2]), .SMC(test_se), .C(
        clkper), .Q(is_reg[3]) );
  SDFFQX1 ien0_reg_reg_4_ ( .D(N43), .SIN(ien0[3]), .SMC(test_se), .C(net12078), .Q(ien0[4]) );
  SDFFQX1 ien1_reg_reg_4_ ( .D(N54), .SIN(ien1[3]), .SMC(test_se), .C(net12084), .Q(ien1[4]) );
  SDFFQX1 ien0_reg_reg_3_ ( .D(N42), .SIN(ien0[2]), .SMC(test_se), .C(net12078), .Q(ien0[3]) );
  SDFFQX1 isr_tm_reg_reg ( .D(n200), .SIN(is_reg[3]), .SMC(test_se), .C(clkper), .Q(isr_tm) );
  SDFFQX1 ip0_reg_reg_3_ ( .D(N71), .SIN(ip0[2]), .SMC(test_se), .C(net12094), 
        .Q(ip0[3]) );
  SDFFQX1 ien1_reg_reg_3_ ( .D(N53), .SIN(ien1[2]), .SMC(test_se), .C(net12084), .Q(ien1[3]) );
  SDFFQX1 ien2_reg_reg_3_ ( .D(N62), .SIN(ien2[2]), .SMC(test_se), .C(net12089), .Q(ien2[3]) );
  SDFFQX1 ip1_reg_reg_3_ ( .D(N80), .SIN(ip1[2]), .SMC(test_se), .C(net12099), 
        .Q(ip1[3]) );
  SDFFQX1 irq_r_reg ( .D(N200), .SIN(ip1[5]), .SMC(test_se), .C(clkper), .Q(
        irq_r) );
  SDFFQX1 ien0_reg_reg_6_ ( .D(N45), .SIN(ien0[5]), .SMC(test_se), .C(net12078), .Q(ien0[7]) );
  SDFFQX1 ien0_reg_reg_1_ ( .D(N40), .SIN(ien0[0]), .SMC(test_se), .C(net12078), .Q(ien0[1]) );
  SDFFQX1 ien1_reg_reg_1_ ( .D(N51), .SIN(ien1[0]), .SMC(test_se), .C(net12084), .Q(ien1[1]) );
  SDFFQX1 ien2_reg_reg_1_ ( .D(N60), .SIN(ien2[0]), .SMC(test_se), .C(net12089), .Q(ien2[1]) );
  SDFFQX1 ip1_reg_reg_1_ ( .D(N78), .SIN(ip1[0]), .SMC(test_se), .C(net12099), 
        .Q(ip1[1]) );
  SDFFQX1 ip0_reg_reg_0_ ( .D(N68), .SIN(intvect[4]), .SMC(test_se), .C(
        net12094), .Q(ip0[0]) );
  SDFFQX1 ip0_reg_reg_1_ ( .D(N69), .SIN(ip0[0]), .SMC(test_se), .C(net12094), 
        .Q(ip0[1]) );
  SDFFQX1 ien1_reg_reg_0_ ( .D(N50), .SIN(ien0[7]), .SMC(test_se), .C(net12084), .Q(ien1[0]) );
  SDFFQX1 ien2_reg_reg_2_ ( .D(N61), .SIN(ien2[1]), .SMC(test_se), .C(net12089), .Q(ien2[2]) );
  SDFFQX1 ien1_reg_reg_2_ ( .D(N52), .SIN(ien1[1]), .SMC(test_se), .C(net12084), .Q(ien1[2]) );
  SDFFQX1 ien0_reg_reg_2_ ( .D(N41), .SIN(ien0[1]), .SMC(test_se), .C(net12078), .Q(ien0[2]) );
  SDFFQX1 ip1_reg_reg_2_ ( .D(N79), .SIN(ip1[1]), .SMC(test_se), .C(net12099), 
        .Q(ip1[2]) );
  SDFFQX1 ip1_reg_reg_0_ ( .D(N77), .SIN(ip0[5]), .SMC(test_se), .C(net12099), 
        .Q(ip1[0]) );
  SDFFQX1 ip0_reg_reg_2_ ( .D(N70), .SIN(ip0[1]), .SMC(test_se), .C(net12094), 
        .Q(ip0[2]) );
  SDFFQX1 ien2_reg_reg_0_ ( .D(N59), .SIN(ien1[5]), .SMC(test_se), .C(net12089), .Q(ien2[0]) );
  SDFFQX1 ien0_reg_reg_0_ ( .D(N39), .SIN(test_si), .SMC(test_se), .C(net12078), .Q(ien0[0]) );
  INVX1 U3 ( .A(1'b1), .Y(ien0[6]) );
  AND2XL U5 ( .A(sfrwe), .B(sfraddr[3]), .Y(n101) );
  INVXL U6 ( .A(sfraddr[5]), .Y(n5) );
  AOI221XL U7 ( .A(ien0[2]), .B(int_vect_13), .C(ien1[2]), .D(int_vect_53), 
        .E(n39), .Y(n179) );
  AOI221XL U8 ( .A(n33), .B(ip1[4]), .C(n183), .D(ip1[3]), .E(n31), .Y(n159)
         );
  AOI221XL U9 ( .A(n32), .B(ip1[4]), .C(ip0[4]), .D(n182), .E(n165), .Y(n153)
         );
  AOI221XL U10 ( .A(n167), .B(ip1[1]), .C(ip0[1]), .D(n22), .E(n168), .Y(n124)
         );
  NAND3X1 U11 ( .A(n3), .B(n4), .C(n94), .Y(n100) );
  NAND3X1 U12 ( .A(n94), .B(n3), .C(sfraddr[4]), .Y(n99) );
  NAND4X1 U13 ( .A(n3), .B(n5), .C(sfraddr[1]), .D(n97), .Y(n96) );
  NOR2X1 U14 ( .A(n98), .B(n4), .Y(n97) );
  NOR3XL U15 ( .A(n98), .B(sfraddr[1]), .C(n5), .Y(n94) );
  NOR2X1 U16 ( .A(n93), .B(n7), .Y(N78) );
  NOR2X1 U17 ( .A(n93), .B(n6), .Y(N77) );
  NOR2X1 U18 ( .A(n93), .B(n8), .Y(N79) );
  NOR2X1 U19 ( .A(n93), .B(n9), .Y(N80) );
  NOR2X1 U20 ( .A(n93), .B(n10), .Y(N81) );
  NOR2X1 U21 ( .A(n7), .B(n96), .Y(N60) );
  NOR2X1 U22 ( .A(n8), .B(n96), .Y(N61) );
  NOR2X1 U23 ( .A(n6), .B(n96), .Y(N59) );
  NOR2X1 U24 ( .A(n9), .B(n96), .Y(N62) );
  NOR2X1 U25 ( .A(n10), .B(n96), .Y(N63) );
  NOR2X1 U26 ( .A(n11), .B(n96), .Y(N64) );
  NOR2X1 U27 ( .A(n11), .B(n93), .Y(N82) );
  NOR2X1 U28 ( .A(n7), .B(n99), .Y(N51) );
  NOR2X1 U29 ( .A(n8), .B(n99), .Y(N52) );
  NOR2X1 U30 ( .A(n6), .B(n99), .Y(N50) );
  NOR2X1 U31 ( .A(n9), .B(n99), .Y(N53) );
  NOR2X1 U32 ( .A(n10), .B(n99), .Y(N54) );
  NOR2X1 U33 ( .A(n11), .B(n99), .Y(N55) );
  NOR2X1 U34 ( .A(n8), .B(n95), .Y(N70) );
  NOR2X1 U35 ( .A(n7), .B(n95), .Y(N69) );
  NOR2X1 U36 ( .A(n6), .B(n95), .Y(N68) );
  NOR2X1 U37 ( .A(n9), .B(n95), .Y(N71) );
  NOR2X1 U38 ( .A(n10), .B(n95), .Y(N72) );
  NOR2X1 U39 ( .A(n11), .B(n95), .Y(N73) );
  NOR2X1 U40 ( .A(n6), .B(n100), .Y(N39) );
  NOR2X1 U41 ( .A(n8), .B(n100), .Y(N41) );
  NOR2X1 U42 ( .A(n7), .B(n100), .Y(N40) );
  NOR2X1 U43 ( .A(n9), .B(n100), .Y(N42) );
  NOR2X1 U44 ( .A(n11), .B(n100), .Y(N44) );
  NOR2X1 U45 ( .A(n10), .B(n100), .Y(N43) );
  NAND2X1 U46 ( .A(n12), .B(n96), .Y(N58) );
  NAND2X1 U47 ( .A(n12), .B(n93), .Y(N76) );
  NAND2X1 U48 ( .A(n12), .B(n95), .Y(N67) );
  NAND2X1 U49 ( .A(n12), .B(n99), .Y(N49) );
  NAND2X1 U50 ( .A(n12), .B(n100), .Y(N38) );
  INVX1 U51 ( .A(n111), .Y(n17) );
  INVX1 U52 ( .A(sfraddr[4]), .Y(n4) );
  NAND2X1 U53 ( .A(n207), .B(n12), .Y(n67) );
  NAND42XL U54 ( .C(sfraddr[2]), .D(sfraddr[6]), .A(n12), .B(n101), .Y(n98) );
  AND4XL U55 ( .A(sfrwe), .B(sfraddr[1]), .C(sfraddr[2]), .D(sfraddr[0]), .Y(
        n61) );
  NOR21XL U56 ( .B(sfrdatai[7]), .A(n100), .Y(N45) );
  NAND3X1 U57 ( .A(sfraddr[0]), .B(n4), .C(n94), .Y(n95) );
  NAND3X1 U58 ( .A(n94), .B(sfraddr[0]), .C(sfraddr[4]), .Y(n93) );
  NAND21X1 U59 ( .B(n136), .A(n117), .Y(n111) );
  INVX1 U60 ( .A(n132), .Y(n19) );
  NOR2X1 U61 ( .A(rst), .B(n102), .Y(N212) );
  NAND3X1 U62 ( .A(n102), .B(n15), .C(n131), .Y(N207) );
  NOR3XL U63 ( .A(n132), .B(rst), .C(n126), .Y(n131) );
  INVX1 U64 ( .A(n168), .Y(n27) );
  NAND31X1 U65 ( .C(n126), .A(n127), .B(n128), .Y(n108) );
  INVX1 U66 ( .A(n134), .Y(n15) );
  OAI211X1 U67 ( .C(n24), .D(n111), .A(n128), .B(n135), .Y(n134) );
  AOI22X1 U68 ( .A(n117), .B(n136), .C(n137), .D(n19), .Y(n135) );
  NOR2X1 U69 ( .A(rst), .B(n15), .Y(N211) );
  INVX1 U70 ( .A(n143), .Y(n24) );
  INVX1 U71 ( .A(n119), .Y(n16) );
  OAI31XL U72 ( .A(n118), .B(n108), .C(n18), .D(n12), .Y(n119) );
  INVX1 U73 ( .A(n120), .Y(n18) );
  AOI211X1 U74 ( .C(n121), .D(n117), .A(n122), .B(n20), .Y(n120) );
  INVX1 U75 ( .A(sfrdatai[4]), .Y(n10) );
  INVX1 U76 ( .A(sfrdatai[5]), .Y(n11) );
  INVX1 U77 ( .A(sfraddr[0]), .Y(n3) );
  INVX1 U78 ( .A(sfrdatai[1]), .Y(n7) );
  INVX1 U79 ( .A(sfrdatai[2]), .Y(n8) );
  INVX1 U80 ( .A(sfrdatai[0]), .Y(n6) );
  INVX1 U81 ( .A(sfrdatai[3]), .Y(n9) );
  INVX1 U82 ( .A(n189), .Y(n29) );
  NAND32X1 U83 ( .B(retiinstr), .C(rst), .A(n62), .Y(n68) );
  INVX1 U84 ( .A(n71), .Y(n42) );
  INVX1 U85 ( .A(intcall), .Y(n207) );
  INVX1 U86 ( .A(rst), .Y(n12) );
  NAND2X1 U87 ( .A(intcall), .B(n12), .Y(n62) );
  OAI32X1 U88 ( .A(n56), .B(rst), .C(n59), .D(n13), .E(n11), .Y(n200) );
  INVX1 U89 ( .A(n59), .Y(n13) );
  NOR43XL U90 ( .B(n60), .C(n61), .D(n12), .A(sfraddr[3]), .Y(n59) );
  NOR3XL U91 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n60) );
  NOR32XL U92 ( .B(n133), .C(n19), .A(n137), .Y(n117) );
  NAND32X1 U93 ( .B(n109), .C(n107), .A(n106), .Y(n132) );
  NOR4XL U94 ( .A(n183), .B(n38), .C(n171), .D(n27), .Y(n165) );
  NOR2X1 U95 ( .A(n184), .B(n158), .Y(n168) );
  NOR42XL U96 ( .C(n127), .D(n104), .A(n122), .B(n139), .Y(n102) );
  OAI21X1 U97 ( .B(n130), .C(n129), .A(n113), .Y(n139) );
  OAI211X1 U98 ( .C(n185), .D(n53), .A(n49), .B(n166), .Y(n158) );
  AOI211X1 U99 ( .C(n21), .D(n34), .A(n138), .B(n149), .Y(n141) );
  INVX1 U100 ( .A(n142), .Y(n34) );
  NAND2X1 U101 ( .A(n24), .B(n17), .Y(n149) );
  NAND3X1 U102 ( .A(n39), .B(n140), .C(n141), .Y(n113) );
  INVX1 U103 ( .A(n159), .Y(n30) );
  INVX1 U104 ( .A(n169), .Y(n40) );
  INVX1 U105 ( .A(n188), .Y(n31) );
  INVX1 U106 ( .A(n174), .Y(n37) );
  OAI222XL U107 ( .A(n111), .B(n112), .C(n129), .D(n130), .E(n109), .F(n106), 
        .Y(n118) );
  OAI21BBX1 U108 ( .A(n140), .B(n39), .C(n141), .Y(n129) );
  NAND2X1 U109 ( .A(n110), .B(n112), .Y(n143) );
  OAI21X1 U110 ( .B(n124), .C(n125), .A(n116), .Y(n136) );
  AOI211X1 U111 ( .C(n26), .D(n54), .A(n23), .B(n129), .Y(n145) );
  INVX1 U112 ( .A(n130), .Y(n23) );
  NOR4XL U113 ( .A(n142), .B(n111), .C(n143), .D(n124), .Y(n122) );
  INVX1 U114 ( .A(n153), .Y(n26) );
  NAND3X1 U115 ( .A(n17), .B(n24), .C(n138), .Y(n128) );
  AOI21X1 U116 ( .B(n145), .C(n148), .A(n67), .Y(N200) );
  NAND2X1 U117 ( .A(n147), .B(n146), .Y(n148) );
  INVX1 U118 ( .A(n124), .Y(n21) );
  INVX1 U119 ( .A(n179), .Y(n38) );
  AOI31X1 U120 ( .A(n113), .B(n114), .C(n115), .D(rst), .Y(N209) );
  AOI21BX1 U121 ( .C(n116), .B(n117), .A(n118), .Y(n115) );
  AOI31X1 U122 ( .A(n103), .B(n104), .C(n105), .D(rst), .Y(N210) );
  NAND32X1 U123 ( .B(n110), .C(n111), .A(n112), .Y(n103) );
  AOI31X1 U124 ( .A(n14), .B(n106), .C(n107), .D(n108), .Y(n105) );
  INVX1 U125 ( .A(n109), .Y(n14) );
  INVX1 U126 ( .A(n162), .Y(n39) );
  NOR2X1 U127 ( .A(n52), .B(n185), .Y(n189) );
  NOR2X1 U128 ( .A(n133), .B(n132), .Y(n126) );
  NOR21XL U129 ( .B(n150), .A(n151), .Y(n137) );
  INVX1 U130 ( .A(n176), .Y(n22) );
  NOR2X1 U131 ( .A(n124), .B(n125), .Y(n121) );
  INVX1 U132 ( .A(n123), .Y(n20) );
  INVX1 U133 ( .A(n181), .Y(n36) );
  NOR21XL U134 ( .B(n64), .A(n62), .Y(n71) );
  NOR2X1 U135 ( .A(n82), .B(n89), .Y(int_ack_43) );
  NOR2X1 U136 ( .A(n91), .B(n86), .Y(int_ack_1b) );
  OAI32X1 U137 ( .A(n62), .B(n41), .C(n64), .D(n72), .E(n50), .Y(n196) );
  AOI21BBXL U138 ( .B(n67), .C(n66), .A(n71), .Y(n72) );
  INVX1 U139 ( .A(n63), .Y(n41) );
  NAND2X1 U140 ( .A(n90), .B(n48), .Y(n91) );
  OAI211X1 U141 ( .C(n82), .D(n83), .A(n44), .B(n45), .Y(n75) );
  INVX1 U142 ( .A(int_ack_43), .Y(n45) );
  INVX1 U143 ( .A(int_ack_03), .Y(n44) );
  OAI22X1 U144 ( .A(n63), .B(n42), .C(n69), .D(n51), .Y(n197) );
  AOI21BX1 U145 ( .C(n67), .B(n70), .A(n71), .Y(n69) );
  OAI22X1 U146 ( .A(n68), .B(n55), .C(n41), .D(n42), .Y(n198) );
  OAI31XL U147 ( .A(n62), .B(n63), .C(n64), .D(n65), .Y(n199) );
  GEN2XL U148 ( .D(n66), .E(n50), .C(n67), .B(n62), .A(n49), .Y(n65) );
  NAND2X1 U149 ( .A(n55), .B(n68), .Y(n70) );
  NOR21XL U150 ( .B(n84), .A(n82), .Y(n74) );
  NOR2X1 U151 ( .A(n78), .B(n83), .Y(int_ack_8b) );
  NOR2X1 U152 ( .A(n78), .B(n91), .Y(int_ack_0b) );
  NAND2X1 U153 ( .A(n47), .B(n46), .Y(n82) );
  NOR2X1 U154 ( .A(n91), .B(n87), .Y(int_ack_13) );
  NOR2X1 U155 ( .A(n89), .B(n87), .Y(int_ack_53) );
  NOR2X1 U156 ( .A(n78), .B(n89), .Y(int_ack_4b) );
  NOR21XL U157 ( .B(n84), .A(n78), .Y(n73) );
  NOR2X1 U158 ( .A(n89), .B(n86), .Y(int_ack_5b) );
  NOR2X1 U159 ( .A(n83), .B(n87), .Y(int_ack_93) );
  NOR2X1 U160 ( .A(n78), .B(n88), .Y(int_ack_6b) );
  NOR2X1 U161 ( .A(n82), .B(n88), .Y(int_ack_63) );
  NAND42X1 U162 ( .C(n129), .D(n144), .A(n26), .B(n130), .Y(n104) );
  NAND3X1 U163 ( .A(n145), .B(n146), .C(n147), .Y(n127) );
  NOR3XL U164 ( .A(n85), .B(n82), .C(n43), .Y(int_ack_a3) );
  NOR3XL U165 ( .A(n85), .B(n78), .C(n43), .Y(int_ack_ab) );
  NOR2X1 U166 ( .A(n83), .B(n86), .Y(int_ack_9b) );
  INVX1 U167 ( .A(n144), .Y(n54) );
  AND2X1 U168 ( .A(irq_r), .B(ien0[7]), .Y(irq) );
  NOR21XL U169 ( .B(n194), .A(n181), .Y(n161) );
  AOI33X1 U170 ( .A(ip1[4]), .B(n33), .C(ip0[4]), .D(ip1[3]), .E(n183), .F(
        ip0[3]), .Y(n194) );
  INVX1 U171 ( .A(n190), .Y(n32) );
  AOI31X1 U172 ( .A(ip0[4]), .B(n57), .C(n36), .D(n191), .Y(n190) );
  AOI21X1 U173 ( .B(ip1[3]), .C(n183), .A(n192), .Y(n191) );
  AOI211X1 U174 ( .C(n38), .D(ip1[2]), .A(n37), .B(n170), .Y(n188) );
  NAND3X1 U175 ( .A(n125), .B(n142), .C(n205), .Y(n171) );
  NAND3X1 U176 ( .A(ien0[1]), .B(n56), .C(int_vect_0b), .Y(n205) );
  OAI21BBX1 U177 ( .A(ien0[0]), .B(int_vect_03), .C(n151), .Y(n184) );
  OAI221X1 U178 ( .A(isr_tm), .B(int_vect_43), .C(sdaiff), .D(n56), .E(ien1[0]), .Y(n151) );
  NAND2X1 U179 ( .A(int_vect_8b), .B(ien2[1]), .Y(n142) );
  NAND2X1 U180 ( .A(n203), .B(n40), .Y(n181) );
  AOI32X1 U181 ( .A(ip1[2]), .B(n38), .C(ip0[2]), .D(n37), .E(ip0[1]), .Y(n203) );
  NAND3X1 U182 ( .A(n29), .B(n50), .C(n187), .Y(n176) );
  AOI21X1 U183 ( .B(ip0[0]), .C(n184), .A(n30), .Y(n187) );
  INVX1 U184 ( .A(isr_tm), .Y(n56) );
  NAND3X1 U185 ( .A(n204), .B(n55), .C(ien0[7]), .Y(n169) );
  NAND3X1 U186 ( .A(ip1[0]), .B(n184), .C(ip0[0]), .Y(n204) );
  NAND2X1 U187 ( .A(ip1[1]), .B(n171), .Y(n174) );
  AOI211X1 U188 ( .C(n56), .D(n206), .A(n153), .B(n154), .Y(n107) );
  OAI21X1 U189 ( .B(n56), .C(rxd0ff), .A(ien0[4]), .Y(n154) );
  AOI21X1 U190 ( .B(n183), .C(ip0[3]), .A(n28), .Y(n182) );
  AOI21AX1 U191 ( .B(n33), .C(ip0[4]), .A(n182), .Y(n166) );
  NAND4X1 U192 ( .A(int_vect_4b), .B(ien1[1]), .C(n142), .D(n56), .Y(n125) );
  NAND4X1 U193 ( .A(n161), .B(n193), .C(n160), .D(n51), .Y(n170) );
  NAND2X1 U194 ( .A(ip1[0]), .B(n184), .Y(n193) );
  INVX1 U195 ( .A(n195), .Y(n33) );
  AOI221XL U196 ( .A(n201), .B(ien0[4]), .C(ien1[4]), .D(int_vect_63), .E(n54), 
        .Y(n195) );
  ENOX1 U197 ( .A(n206), .B(isr_tm), .C(rxd0ff), .D(isr_tm), .Y(n201) );
  INVX1 U198 ( .A(n186), .Y(n28) );
  AOI221XL U199 ( .A(n171), .B(ip0[1]), .C(n38), .D(ip0[2]), .E(n176), .Y(n186) );
  INVX1 U200 ( .A(int_vect_23), .Y(n206) );
  NOR43XL U201 ( .B(int_vect_6b), .C(ien1[5]), .D(n146), .A(n147), .Y(n138) );
  OAI21X1 U202 ( .B(n169), .C(n58), .A(n170), .Y(n167) );
  OAI21X1 U203 ( .B(n27), .C(n171), .A(n172), .Y(n140) );
  AOI32X1 U204 ( .A(n173), .B(n174), .C(ip1[2]), .D(ip0[2]), .E(n175), .Y(n172) );
  OAI21BBX1 U205 ( .A(ip0[2]), .B(n40), .C(n170), .Y(n173) );
  OAI22X1 U206 ( .A(n176), .B(n171), .C(ip0[1]), .D(n177), .Y(n175) );
  OAI21BBX1 U207 ( .A(ien2[3]), .B(int_vect_9b), .C(n202), .Y(n183) );
  AOI32X1 U208 ( .A(ien0[3]), .B(n56), .C(int_vect_1b), .D(int_vect_5b), .E(
        ien1[3]), .Y(n202) );
  OAI21X1 U209 ( .B(n57), .C(n28), .A(n178), .Y(n152) );
  AOI32X1 U210 ( .A(n35), .B(n168), .C(n179), .D(ip1[3]), .E(n180), .Y(n178)
         );
  INVX1 U211 ( .A(n171), .Y(n35) );
  OAI21X1 U212 ( .B(n57), .C(n181), .A(n31), .Y(n180) );
  NAND3X1 U213 ( .A(n114), .B(n123), .C(n155), .Y(n109) );
  NAND3X1 U214 ( .A(ien0[0]), .B(n150), .C(int_vect_03), .Y(n155) );
  NAND4X1 U215 ( .A(int_vect_0b), .B(ien0[1]), .C(n21), .D(n56), .Y(n123) );
  NAND2X1 U216 ( .A(int_vect_93), .B(ien2[2]), .Y(n162) );
  NAND3X1 U217 ( .A(int_vect_5b), .B(ien1[3]), .C(n163), .Y(n112) );
  AOI21AX1 U218 ( .B(int_vect_9b), .C(ien2[3]), .A(n152), .Y(n163) );
  OAI2B11X1 U219 ( .D(ip1[0]), .C(n156), .A(n157), .B(n158), .Y(n150) );
  AOI33X1 U220 ( .A(n160), .B(n51), .C(n161), .D(ip0[0]), .E(n55), .F(ien0[7]), 
        .Y(n156) );
  NAND4X1 U221 ( .A(n159), .B(ip0[0]), .C(n29), .D(n50), .Y(n157) );
  NAND4X1 U222 ( .A(int_vect_1b), .B(ien0[3]), .C(n152), .D(n56), .Y(n106) );
  NAND4X1 U223 ( .A(int_vect_63), .B(ien1[4]), .C(n26), .D(n144), .Y(n110) );
  NAND3X1 U224 ( .A(i2c_int), .B(n146), .C(ien0[5]), .Y(n133) );
  NAND4X1 U225 ( .A(int_vect_53), .B(ien1[2]), .C(n140), .D(n162), .Y(n116) );
  NAND3X1 U226 ( .A(ien0[2]), .B(n140), .C(int_vect_13), .Y(n114) );
  OAI222XL U227 ( .A(n164), .B(n53), .C(n52), .D(n30), .E(n25), .F(n33), .Y(
        n146) );
  AOI21X1 U228 ( .B(n161), .C(ip1[5]), .A(n166), .Y(n164) );
  INVX1 U229 ( .A(n165), .Y(n25) );
  AOI221XL U230 ( .A(i2c_int), .B(ien0[5]), .C(ien1[5]), .D(int_vect_6b), .E(
        n147), .Y(n185) );
  NAND2X1 U231 ( .A(n189), .B(ip0[5]), .Y(n160) );
  INVX1 U232 ( .A(is_reg[3]), .Y(n55) );
  INVX1 U233 ( .A(is_reg[2]), .Y(n51) );
  AOI21X1 U234 ( .B(n40), .C(ip1[2]), .A(n22), .Y(n177) );
  INVX1 U235 ( .A(ip1[5]), .Y(n52) );
  AOI21X1 U236 ( .B(n36), .C(ip0[4]), .A(n188), .Y(n192) );
  INVX1 U237 ( .A(is_reg[1]), .Y(n50) );
  INVX1 U238 ( .A(ip0[5]), .Y(n53) );
  INVX1 U239 ( .A(ip0[1]), .Y(n58) );
  INVX1 U240 ( .A(is_reg[0]), .Y(n49) );
  INVX1 U241 ( .A(ip0[3]), .Y(n57) );
  OAI22X1 U242 ( .A(n82), .B(n91), .C(n92), .D(n207), .Y(int_ack_03) );
  AOI22X1 U243 ( .A(intvect[2]), .B(intvect[1]), .C(intvect[4]), .D(intvect[3]), .Y(n92) );
  AO2222XL U244 ( .A(ip0[5]), .B(n73), .C(ip0[4]), .D(n74), .E(ip0[0]), .F(n75), .G(n76), .H(n80), .Y(n63) );
  OAI22X1 U245 ( .A(n78), .B(n58), .C(n81), .D(n46), .Y(n80) );
  AOI22X1 U246 ( .A(ip0[2]), .B(n47), .C(ip0[3]), .D(intvect[0]), .Y(n81) );
  AO2222XL U247 ( .A(ip1[5]), .B(n73), .C(ip1[4]), .D(n74), .E(ip1[0]), .F(n75), .G(n76), .H(n77), .Y(n64) );
  OAI22AX1 U248 ( .D(ip1[1]), .C(n78), .A(n79), .B(n46), .Y(n77) );
  AOI22X1 U249 ( .A(ip1[2]), .B(n47), .C(ip1[3]), .D(intvect[0]), .Y(n79) );
  NOR3XL U250 ( .A(intvect[2]), .B(intvect[4]), .C(n207), .Y(n90) );
  NAND2X1 U251 ( .A(n90), .B(intvect[3]), .Y(n89) );
  OR2X1 U252 ( .A(n85), .B(intvect[2]), .Y(n83) );
  NAND3X1 U253 ( .A(intcall), .B(n48), .C(intvect[4]), .Y(n85) );
  NOR2X1 U254 ( .A(n70), .B(is_reg[2]), .Y(n66) );
  NAND2X1 U255 ( .A(intvect[0]), .B(n46), .Y(n78) );
  AOI21X1 U256 ( .B(intvect[3]), .C(intvect[4]), .A(n43), .Y(n84) );
  NAND2X1 U257 ( .A(intvect[1]), .B(intvect[0]), .Y(n86) );
  INVX1 U258 ( .A(intvect[0]), .Y(n47) );
  INVX1 U259 ( .A(intvect[1]), .Y(n46) );
  INVX1 U260 ( .A(intvect[3]), .Y(n48) );
  INVX1 U261 ( .A(intvect[2]), .Y(n43) );
  NAND41X1 U262 ( .D(intvect[4]), .A(intvect[2]), .B(intvect[3]), .C(intcall), 
        .Y(n88) );
  AOI21X1 U263 ( .B(intvect[3]), .C(intvect[4]), .A(intvect[2]), .Y(n76) );
  NAND2X1 U264 ( .A(intvect[1]), .B(n47), .Y(n87) );
  AND2X1 U265 ( .A(int_vect_ab), .B(ien2[5]), .Y(n147) );
  NAND3X1 U267 ( .A(ien2[3]), .B(n152), .C(int_vect_9b), .Y(n130) );
  NAND2X1 U268 ( .A(int_vect_a3), .B(ien2[4]), .Y(n144) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module watchdog_a0 ( wdt_slow, clkwdt, clkper, resetff, newinstr, wdts_s, wdts, 
        ip0wdts, wdt_tm, sfrdatai, sfraddr, sfrwe, wdtrel, test_si, test_se );
  output [1:0] wdts_s;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] wdtrel;
  input wdt_slow, clkwdt, clkper, resetff, newinstr, sfrwe, test_si, test_se;
  output wdts, ip0wdts, wdt_tm;
  wire   wdt_tm_sync, wdt_act_sync, wdt_act, wdtrefresh_sync, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N67, N68, N69, N70, N71, pres_2, N112,
         N113, N114, N115, N116, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, wdt_normal, wdt_normal_ff, N212, net12127, net12133,
         net12138, net12143, net12148, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n125, n135, n136, n137;
  wire   [1:0] pres_8;
  wire   [3:0] cycles_reg;
  wire   [3:0] pres_16;
  wire   [6:0] wdth;
  wire   [7:0] wdtl;

  SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 clk_gate_wdtrel_s_reg ( .CLK(clkper), 
        .EN(N26), .ENCLK(net12127), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 clk_gate_cycles_reg_reg ( .CLK(clkwdt), 
        .EN(N67), .ENCLK(net12133), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 clk_gate_pres_16_reg ( .CLK(clkwdt), .EN(
        N112), .ENCLK(net12138), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 clk_gate_wdth_reg ( .CLK(clkwdt), .EN(
        N165), .ENCLK(net12143), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 clk_gate_wdtl_reg ( .CLK(clkwdt), .EN(
        n124), .ENCLK(net12148), .TE(test_se) );
  watchdog_a0_DW01_inc_0 add_278 ( .A(wdtl), .SUM({N144, N143, N142, N141, 
        N140, N139, N138, N137}) );
  watchdog_a0_DW01_inc_1 add_272 ( .A(wdth), .SUM({N136, N135, N134, N133, 
        N132, N131, N130}) );
  SDFFQX1 wdt_act_reg ( .D(n130), .SIN(pres_16[3]), .SMC(test_se), .C(clkper), 
        .Q(wdt_act) );
  SDFFQX1 wdts_reg ( .D(wdts_s[0]), .SIN(wdtrel[7]), .SMC(test_se), .C(clkper), 
        .Q(wdts) );
  SDFFQX1 wdts_s_reg_1_ ( .D(n126), .SIN(wdts_s[0]), .SMC(test_se), .C(
        net12148), .Q(wdts_s[1]) );
  SDFFQX1 wdts_s_reg_0_ ( .D(n132), .SIN(wdts), .SMC(test_se), .C(net12148), 
        .Q(wdts_s[0]) );
  SDFFQX1 wdt_normal_ff_reg ( .D(n123), .SIN(wdt_act_sync), .SMC(test_se), .C(
        clkper), .Q(wdt_normal_ff) );
  SDFFQX1 wdt_normal_reg ( .D(n133), .SIN(wdt_normal_ff), .SMC(test_se), .C(
        clkper), .Q(wdt_normal) );
  SDFFQX1 wdt_act_sync_reg ( .D(wdt_act), .SIN(wdt_act), .SMC(test_se), .C(
        clkwdt), .Q(wdt_act_sync) );
  SDFFQX1 pres_16_reg_3_ ( .D(N116), .SIN(pres_16[2]), .SMC(test_se), .C(
        net12138), .Q(pres_16[3]) );
  SDFFQX1 wdth_reg_6_ ( .D(N172), .SIN(wdth[5]), .SMC(test_se), .C(net12143), 
        .Q(wdth[6]) );
  SDFFQX1 pres_16_reg_2_ ( .D(N115), .SIN(pres_16[1]), .SMC(test_se), .C(
        net12138), .Q(pres_16[2]) );
  SDFFQX1 pres_8_reg_1_ ( .D(n128), .SIN(pres_8[0]), .SMC(test_se), .C(
        net12133), .Q(pres_8[1]) );
  SDFFQX1 pres_2_reg ( .D(n127), .SIN(ip0wdts), .SMC(test_se), .C(net12133), 
        .Q(pres_2) );
  SDFFQX1 pres_8_reg_0_ ( .D(n129), .SIN(pres_2), .SMC(test_se), .C(net12133), 
        .Q(pres_8[0]) );
  SDFFQX1 wdt_tm_sync_reg ( .D(wdt_tm), .SIN(wdt_tm), .SMC(test_se), .C(clkwdt), .Q(wdt_tm_sync) );
  SDFFQX1 pres_16_reg_1_ ( .D(N114), .SIN(pres_16[0]), .SMC(test_se), .C(
        net12138), .Q(pres_16[1]) );
  SDFFQX1 cycles_reg_reg_2_ ( .D(N70), .SIN(cycles_reg[1]), .SMC(test_se), .C(
        net12133), .Q(cycles_reg[2]) );
  SDFFQX1 pres_16_reg_0_ ( .D(N113), .SIN(pres_8[1]), .SMC(test_se), .C(
        net12138), .Q(pres_16[0]) );
  SDFFQX1 wdth_reg_3_ ( .D(N169), .SIN(wdth[2]), .SMC(test_se), .C(net12143), 
        .Q(wdth[3]) );
  SDFFQX1 wdth_reg_1_ ( .D(N167), .SIN(wdth[0]), .SMC(test_se), .C(net12143), 
        .Q(wdth[1]) );
  SDFFQX1 wdtl_reg_2_ ( .D(N175), .SIN(wdtl[1]), .SMC(test_se), .C(net12148), 
        .Q(wdtl[2]) );
  SDFFQX1 wdth_reg_4_ ( .D(N170), .SIN(wdth[3]), .SMC(test_se), .C(net12143), 
        .Q(wdth[4]) );
  SDFFQX1 cycles_reg_reg_3_ ( .D(N71), .SIN(cycles_reg[2]), .SMC(test_se), .C(
        net12133), .Q(cycles_reg[3]) );
  SDFFQX1 wdtl_reg_4_ ( .D(N177), .SIN(wdtl[3]), .SMC(test_se), .C(net12148), 
        .Q(wdtl[4]) );
  SDFFQX1 wdtrefresh_reg ( .D(N212), .SIN(wdtl[7]), .SMC(test_se), .C(clkper), 
        .Q(wdtrefresh_sync) );
  SDFFQX1 wdth_reg_0_ ( .D(N166), .SIN(wdt_tm_sync), .SMC(test_se), .C(
        net12143), .Q(wdth[0]) );
  SDFFQX1 cycles_reg_reg_1_ ( .D(N69), .SIN(cycles_reg[0]), .SMC(test_se), .C(
        net12133), .Q(cycles_reg[1]) );
  SDFFQX1 cycles_reg_reg_0_ ( .D(N68), .SIN(test_si), .SMC(test_se), .C(
        net12133), .Q(cycles_reg[0]) );
  SDFFQX1 wdth_reg_2_ ( .D(N168), .SIN(wdth[1]), .SMC(test_se), .C(net12143), 
        .Q(wdth[2]) );
  SDFFQX1 wdtl_reg_6_ ( .D(N179), .SIN(wdtl[5]), .SMC(test_se), .C(net12148), 
        .Q(wdtl[6]) );
  SDFFQX1 wdth_reg_5_ ( .D(N171), .SIN(wdth[4]), .SMC(test_se), .C(net12143), 
        .Q(wdth[5]) );
  SDFFQX1 wdtl_reg_1_ ( .D(N174), .SIN(wdtl[0]), .SMC(test_se), .C(net12148), 
        .Q(wdtl[1]) );
  SDFFQX1 wdtl_reg_7_ ( .D(N180), .SIN(wdtl[6]), .SMC(test_se), .C(net12148), 
        .Q(wdtl[7]) );
  SDFFQX1 wdtl_reg_3_ ( .D(N176), .SIN(wdtl[2]), .SMC(test_se), .C(net12148), 
        .Q(wdtl[3]) );
  SDFFQX1 wdtl_reg_5_ ( .D(N178), .SIN(wdtl[4]), .SMC(test_se), .C(net12148), 
        .Q(wdtl[5]) );
  SDFFQX1 wdtl_reg_0_ ( .D(N173), .SIN(wdth[6]), .SMC(test_se), .C(net12148), 
        .Q(wdtl[0]) );
  SDFFQX1 wdtrel_s_reg_7_ ( .D(N34), .SIN(wdtrel[6]), .SMC(test_se), .C(
        net12127), .Q(wdtrel[7]) );
  SDFFQX1 ip0wdts_reg ( .D(n131), .SIN(cycles_reg[3]), .SMC(test_se), .C(
        clkper), .Q(ip0wdts) );
  SDFFQX1 wdt_tm_s_reg ( .D(n134), .SIN(wdt_normal), .SMC(test_se), .C(clkper), 
        .Q(wdt_tm) );
  SDFFQX1 wdtrel_s_reg_6_ ( .D(N33), .SIN(wdtrel[5]), .SMC(test_se), .C(
        net12127), .Q(wdtrel[6]) );
  SDFFQX1 wdtrel_s_reg_4_ ( .D(N31), .SIN(wdtrel[3]), .SMC(test_se), .C(
        net12127), .Q(wdtrel[4]) );
  SDFFQX1 wdtrel_s_reg_5_ ( .D(N32), .SIN(wdtrel[4]), .SMC(test_se), .C(
        net12127), .Q(wdtrel[5]) );
  SDFFQX1 wdtrel_s_reg_3_ ( .D(N30), .SIN(wdtrel[2]), .SMC(test_se), .C(
        net12127), .Q(wdtrel[3]) );
  SDFFQX1 wdtrel_s_reg_1_ ( .D(N28), .SIN(wdtrel[0]), .SMC(test_se), .C(
        net12127), .Q(wdtrel[1]) );
  SDFFQX1 wdtrel_s_reg_2_ ( .D(N29), .SIN(wdtrel[1]), .SMC(test_se), .C(
        net12127), .Q(wdtrel[2]) );
  SDFFQX1 wdtrel_s_reg_0_ ( .D(N27), .SIN(wdtrefresh_sync), .SMC(test_se), .C(
        net12127), .Q(wdtrel[0]) );
  BUFX3 U3 ( .A(n136), .Y(n1) );
  NOR2X1 U4 ( .A(n65), .B(wdtrefresh_sync), .Y(n2) );
  NAND4XL U5 ( .A(sfraddr[1]), .B(n39), .C(sfraddr[2]), .D(n106), .Y(n105) );
  NAND2X1 U6 ( .A(n41), .B(n4), .Y(n40) );
  INVX1 U7 ( .A(sfraddr[4]), .Y(n7) );
  INVX1 U8 ( .A(n6), .Y(n5) );
  INVX1 U9 ( .A(sfraddr[5]), .Y(n8) );
  INVX1 U10 ( .A(n118), .Y(n13) );
  AND4X1 U11 ( .A(sfraddr[5]), .B(n39), .C(n56), .D(n5), .Y(n41) );
  NOR2X1 U12 ( .A(sfraddr[2]), .B(sfraddr[1]), .Y(n56) );
  INVX1 U13 ( .A(n32), .Y(n10) );
  NAND4XL U14 ( .A(sfrwe), .B(n4), .C(n107), .D(n108), .Y(n57) );
  NOR3XL U15 ( .A(sfraddr[1]), .B(sfraddr[6]), .C(sfraddr[2]), .Y(n107) );
  NOR4XL U16 ( .A(n6), .B(n8), .C(n9), .D(n7), .Y(n108) );
  INVX1 U17 ( .A(n4), .Y(n3) );
  INVX1 U18 ( .A(sfraddr[0]), .Y(n4) );
  INVX1 U19 ( .A(sfrdatai[6]), .Y(n9) );
  INVX1 U20 ( .A(sfraddr[3]), .Y(n6) );
  NAND2X1 U21 ( .A(n68), .B(n14), .Y(n118) );
  NOR32XL U22 ( .B(n136), .C(n40), .A(newinstr), .Y(n32) );
  NOR21XL U23 ( .B(sfrdatai[1]), .A(n105), .Y(N28) );
  NOR21XL U24 ( .B(sfrdatai[0]), .A(n105), .Y(N27) );
  NOR21XL U25 ( .B(sfrdatai[2]), .A(n105), .Y(N29) );
  NOR21XL U26 ( .B(sfrdatai[3]), .A(n105), .Y(N30) );
  NOR21XL U27 ( .B(sfrdatai[5]), .A(n105), .Y(N32) );
  NOR21XL U28 ( .B(sfrdatai[4]), .A(n105), .Y(N31) );
  NOR21XL U29 ( .B(sfrdatai[7]), .A(n105), .Y(N34) );
  NOR2X1 U30 ( .A(n9), .B(n105), .Y(N33) );
  NAND2X1 U31 ( .A(n1), .B(n105), .Y(N26) );
  NAND2X1 U32 ( .A(n92), .B(n125), .Y(n94) );
  INVX1 U33 ( .A(n84), .Y(n30) );
  NOR32XL U34 ( .B(n47), .C(n19), .A(n68), .Y(n67) );
  XNOR2XL U35 ( .A(n27), .B(n137), .Y(n52) );
  NOR3XL U36 ( .A(n18), .B(n17), .C(n21), .Y(n68) );
  INVX1 U37 ( .A(n64), .Y(n21) );
  INVX1 U38 ( .A(n110), .Y(n22) );
  NAND2X1 U39 ( .A(n33), .B(n46), .Y(n43) );
  NOR21XL U40 ( .B(N143), .A(n43), .Y(N179) );
  NOR21XL U41 ( .B(N142), .A(n43), .Y(N178) );
  NOR21XL U42 ( .B(N141), .A(n43), .Y(N177) );
  NOR21XL U43 ( .B(N140), .A(n43), .Y(N176) );
  NOR21XL U44 ( .B(N138), .A(n43), .Y(N174) );
  NOR21XL U45 ( .B(N139), .A(n43), .Y(N175) );
  OAI21X1 U46 ( .B(n120), .C(n118), .A(n60), .Y(N115) );
  XNOR2XL U47 ( .A(n119), .B(n15), .Y(n120) );
  ENOX1 U48 ( .A(n31), .B(n35), .C(N135), .D(n2), .Y(N171) );
  NAND2X1 U49 ( .A(n33), .B(n22), .Y(n101) );
  NOR2X1 U50 ( .A(n15), .B(n119), .Y(n113) );
  OAI211X1 U51 ( .C(n46), .D(n109), .A(n35), .B(n136), .Y(N165) );
  NAND21X1 U52 ( .B(n34), .A(n33), .Y(n109) );
  INVX1 U53 ( .A(n65), .Y(n14) );
  OAI2B11X1 U54 ( .D(n2), .C(n34), .A(n35), .B(n136), .Y(n124) );
  ENOX1 U55 ( .A(n125), .B(n35), .C(N132), .D(n33), .Y(N168) );
  INVX1 U56 ( .A(n102), .Y(n23) );
  NAND2X1 U57 ( .A(n1), .B(n65), .Y(N67) );
  OAI32X1 U58 ( .A(n40), .B(resetff), .C(n9), .D(n12), .E(n10), .Y(n133) );
  OAI32X1 U59 ( .A(n12), .B(resetff), .C(n32), .D(n10), .E(n11), .Y(n123) );
  OAI21X1 U60 ( .B(n36), .C(n9), .A(n37), .Y(n134) );
  NAND3X1 U61 ( .A(n36), .B(n136), .C(wdt_tm), .Y(n37) );
  NAND4XL U62 ( .A(sfraddr[1]), .B(n3), .C(sfraddr[2]), .D(n38), .Y(n36) );
  AND4X1 U63 ( .A(n8), .B(n6), .C(n39), .D(n136), .Y(n38) );
  AOI21X1 U64 ( .B(n53), .C(n54), .A(resetff), .Y(n131) );
  OAI21X1 U65 ( .B(ip0wdts), .C(wdts_s[0]), .A(n55), .Y(n54) );
  NAND21X1 U66 ( .B(n55), .A(sfrdatai[6]), .Y(n53) );
  NAND2X1 U67 ( .A(n3), .B(n41), .Y(n55) );
  NOR4XL U68 ( .A(sfraddr[5]), .B(n5), .C(n3), .D(resetff), .Y(n106) );
  OAI31XL U69 ( .A(n57), .B(wdts_s[0]), .C(resetff), .D(n58), .Y(n130) );
  OAI21X1 U70 ( .B(wdts_s[0]), .C(n136), .A(wdt_act), .Y(n58) );
  NOR3XL U71 ( .A(n57), .B(resetff), .C(n11), .Y(N212) );
  NOR3XL U72 ( .A(wdtrel[3]), .B(wdtrel[4]), .C(n94), .Y(n84) );
  AOI211X1 U73 ( .C(n77), .D(wdtrel[5]), .A(n78), .B(n79), .Y(n76) );
  XNOR2XL U74 ( .A(n84), .B(wdth[4]), .Y(n77) );
  AOI21AX1 U75 ( .B(wdth[4]), .C(n80), .A(n81), .Y(n79) );
  OAI211X1 U76 ( .C(n81), .D(n82), .A(n83), .B(n24), .Y(n78) );
  OAI22X1 U77 ( .A(n69), .B(n70), .C(n43), .D(n71), .Y(n126) );
  NAND2X1 U78 ( .A(wdts_s[1]), .B(n47), .Y(n70) );
  OAI2B11X1 U79 ( .D(wdtl[2]), .C(n72), .A(n71), .B(n46), .Y(n69) );
  OR2X1 U80 ( .A(n49), .B(n51), .Y(n72) );
  NOR2X1 U81 ( .A(wdtrel[1]), .B(wdtrel[0]), .Y(n92) );
  NAND4X1 U82 ( .A(n73), .B(n74), .C(n75), .D(n76), .Y(n71) );
  AOI221XL U83 ( .A(n85), .B(n137), .C(wdt_slow), .D(n86), .E(n87), .Y(n75) );
  NOR3XL U84 ( .A(n88), .B(n89), .C(n90), .Y(n74) );
  NOR42XL U85 ( .C(wdtl[2]), .D(wdtl[0]), .A(n95), .B(n96), .Y(n73) );
  NOR2X1 U86 ( .A(n30), .B(wdtrel[5]), .Y(n81) );
  NAND3X1 U87 ( .A(n30), .B(n31), .C(wdth[4]), .Y(n83) );
  NAND4X1 U88 ( .A(n114), .B(n115), .C(wdtl[0]), .D(n116), .Y(n51) );
  NOR2X1 U89 ( .A(n24), .B(n25), .Y(n116) );
  XNOR2XL U90 ( .A(n137), .B(wdtl[6]), .Y(n115) );
  XNOR2XL U91 ( .A(n137), .B(wdtl[5]), .Y(n114) );
  XNOR2XL U92 ( .A(wdth[0]), .B(n91), .Y(n90) );
  AOI21X1 U93 ( .B(wdtrel[1]), .C(wdtrel[0]), .A(n92), .Y(n91) );
  XNOR2XL U94 ( .A(n29), .B(wdth[5]), .Y(n80) );
  XNOR2XL U95 ( .A(wdtrel[6]), .B(wdth[5]), .Y(n82) );
  XOR2X1 U96 ( .A(n98), .B(wdth[3]), .Y(n95) );
  NAND2X1 U97 ( .A(n99), .B(n30), .Y(n98) );
  OAI21X1 U98 ( .B(wdtrel[3]), .C(n94), .A(wdtrel[4]), .Y(n99) );
  XOR2X1 U99 ( .A(n94), .B(n97), .Y(n96) );
  XNOR2XL U100 ( .A(wdtrel[3]), .B(wdth[2]), .Y(n97) );
  NOR3XL U101 ( .A(n102), .B(cycles_reg[2]), .C(n26), .Y(n110) );
  OAI22BX1 U102 ( .B(n42), .A(n43), .D(wdts_s[0]), .C(n42), .Y(n132) );
  OAI211X1 U103 ( .C(n44), .D(n45), .A(n46), .B(n47), .Y(n42) );
  NAND4X1 U104 ( .A(wdth[6]), .B(wdth[5]), .C(n48), .D(wdth[4]), .Y(n45) );
  NAND4X1 U105 ( .A(n49), .B(wdth[0]), .C(wdth[1]), .D(n50), .Y(n44) );
  NOR2X1 U106 ( .A(n22), .B(wdtrefresh_sync), .Y(n64) );
  NAND2X1 U107 ( .A(cycles_reg[1]), .B(cycles_reg[0]), .Y(n102) );
  OAI32X1 U108 ( .A(n66), .B(resetff), .C(n67), .D(n20), .E(n16), .Y(n127) );
  INVX1 U109 ( .A(pres_2), .Y(n20) );
  AOI21BBXL U110 ( .B(pres_2), .C(wdtrefresh_sync), .A(wdt_tm_sync), .Y(n66)
         );
  INVX1 U111 ( .A(n67), .Y(n16) );
  XOR2X1 U112 ( .A(n93), .B(wdth[1]), .Y(n89) );
  OAI21X1 U113 ( .B(n92), .C(n125), .A(n94), .Y(n93) );
  NOR3XL U114 ( .A(n51), .B(wdtl[2]), .C(n52), .Y(n50) );
  INVX1 U115 ( .A(wdtrel[2]), .Y(n125) );
  INVX1 U116 ( .A(wdtl[7]), .Y(n27) );
  INVX1 U117 ( .A(wdtl[3]), .Y(n25) );
  INVX1 U118 ( .A(wdtl[1]), .Y(n24) );
  INVX1 U119 ( .A(wdtrel[6]), .Y(n29) );
  INVX1 U120 ( .A(wdtrel[5]), .Y(n31) );
  NAND2X1 U121 ( .A(n60), .B(n121), .Y(N114) );
  OAI211X1 U122 ( .C(pres_16[1]), .D(pres_16[0]), .A(n119), .B(n13), .Y(n121)
         );
  NAND3X1 U123 ( .A(n60), .B(n136), .C(n122), .Y(N112) );
  AOI22X1 U124 ( .A(n13), .B(pres_2), .C(n14), .D(wdtrefresh_sync), .Y(n122)
         );
  NAND42X1 U125 ( .C(n52), .D(n51), .A(wdtl[4]), .B(wdtl[2]), .Y(n46) );
  NAND31X1 U126 ( .C(n59), .A(n60), .B(n61), .Y(n129) );
  NAND4X1 U127 ( .A(n47), .B(pres_8[0]), .C(n21), .D(n19), .Y(n61) );
  NOR21XL U128 ( .B(N137), .A(n43), .Y(N173) );
  NOR21XL U129 ( .B(N144), .A(n43), .Y(N180) );
  NOR2X1 U130 ( .A(n65), .B(wdtrefresh_sync), .Y(n33) );
  XNOR2XL U131 ( .A(wdtl[4]), .B(wdt_slow), .Y(n49) );
  INVX1 U132 ( .A(resetff), .Y(n136) );
  AO22AXL U133 ( .A(N134), .B(n2), .C(wdtrel[4]), .D(n35), .Y(N170) );
  NAND2X1 U134 ( .A(wdt_act_sync), .B(n136), .Y(n65) );
  AND2X1 U135 ( .A(wdth[2]), .B(wdth[3]), .Y(n48) );
  OAI22X1 U136 ( .A(wdtrel[0]), .B(wdtl[4]), .C(n28), .D(n25), .Y(n87) );
  NOR3XL U137 ( .A(n65), .B(pres_8[0]), .C(n21), .Y(n59) );
  OAI21X1 U138 ( .B(pres_16[0]), .C(n118), .A(n60), .Y(N113) );
  OAI21X1 U139 ( .B(n117), .C(n118), .A(n60), .Y(N116) );
  XNOR2XL U140 ( .A(pres_16[3]), .B(n113), .Y(n117) );
  OAI21X1 U141 ( .B(n100), .C(n101), .A(n60), .Y(N71) );
  AOI32X1 U142 ( .A(n23), .B(n26), .C(cycles_reg[2]), .D(cycles_reg[3]), .E(
        n102), .Y(n100) );
  OAI21X1 U143 ( .B(cycles_reg[0]), .C(n101), .A(n60), .Y(N68) );
  NAND2X1 U144 ( .A(pres_16[1]), .B(pres_16[0]), .Y(n119) );
  ENOX1 U145 ( .A(n27), .B(n135), .C(n28), .D(wdtl[6]), .Y(n88) );
  ENOX1 U146 ( .A(n29), .B(n35), .C(N136), .D(n2), .Y(N172) );
  OAI211X1 U147 ( .C(wdtrel[0]), .D(wdtl[7]), .A(wdtl[6]), .B(wdtl[4]), .Y(n85) );
  OAI211X1 U148 ( .C(n62), .D(n18), .A(n63), .B(n60), .Y(n128) );
  NAND4X1 U149 ( .A(n64), .B(n14), .C(pres_8[0]), .D(n18), .Y(n63) );
  AOI31X1 U150 ( .A(n21), .B(n19), .C(n47), .D(n59), .Y(n62) );
  NAND4X1 U151 ( .A(n110), .B(n111), .C(pres_2), .D(n112), .Y(n34) );
  NOR2X1 U152 ( .A(n17), .B(n18), .Y(n112) );
  OAI21BBX1 U153 ( .A(n113), .B(pres_16[3]), .C(wdtrel[7]), .Y(n111) );
  INVX1 U154 ( .A(wdtrel[0]), .Y(n135) );
  INVX1 U155 ( .A(wdtl[5]), .Y(n28) );
  INVX1 U156 ( .A(cycles_reg[3]), .Y(n26) );
  AO22AXL U157 ( .A(N133), .B(n33), .C(wdtrel[3]), .D(n35), .Y(N169) );
  AO22AXL U158 ( .A(N131), .B(n2), .C(wdtrel[1]), .D(n35), .Y(N167) );
  NAND2X1 U159 ( .A(wdt_tm_sync), .B(n14), .Y(n60) );
  NOR2X1 U160 ( .A(wdtrefresh_sync), .B(resetff), .Y(n47) );
  NAND2X1 U161 ( .A(wdtrefresh_sync), .B(n136), .Y(n35) );
  OAI21X1 U162 ( .B(n101), .C(n104), .A(n60), .Y(N69) );
  OAI21X1 U163 ( .B(cycles_reg[1]), .C(cycles_reg[0]), .A(n102), .Y(n104) );
  INVX1 U164 ( .A(wdt_tm_sync), .Y(n19) );
  NOR3XL U165 ( .A(n101), .B(wdt_tm_sync), .C(n103), .Y(N70) );
  XNOR2XL U166 ( .A(n23), .B(cycles_reg[2]), .Y(n103) );
  INVX1 U167 ( .A(pres_8[1]), .Y(n18) );
  ENOX1 U168 ( .A(n135), .B(n35), .C(N130), .D(n33), .Y(N166) );
  INVX1 U169 ( .A(pres_8[0]), .Y(n17) );
  INVX1 U170 ( .A(pres_16[2]), .Y(n15) );
  INVX1 U171 ( .A(wdt_normal), .Y(n12) );
  INVX1 U172 ( .A(wdt_normal_ff), .Y(n11) );
  OAI2B11X1 U173 ( .D(wdtl[4]), .C(n135), .A(n27), .B(wdtl[3]), .Y(n86) );
  INVX1 U174 ( .A(wdt_slow), .Y(n137) );
  NOR32XL U175 ( .B(n7), .C(sfrwe), .A(sfraddr[6]), .Y(n39) );
endmodule


module watchdog_a0_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module watchdog_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer1_a0 ( clkper, rst, newinstr, t1ff, t1ack, int1ff, t1_tf1, t1ov, 
        sfrdatai, sfraddr, sfrwe, t1_tmod, t1_tr1, tl1, th1, test_si, test_se
 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t1_tmod;
  output [7:0] tl1;
  output [7:0] th1;
  input clkper, rst, newinstr, t1ff, t1ack, int1ff, sfrwe, test_si, test_se;
  output t1_tf1, t1ov, t1_tr1;
  wire   t1clr, th1_ov_ff, tl1_ov_ff, N31, N32, N33, N34, N35, N36, N37, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N95, N97, N98, clk_ov12, N100, net12165,
         net12171, net12176, n54, n55, n56, n57, n58, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n59, n60, n61, n62, n63, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n64;
  wire   [1:0] t0_mode;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer1_a0_0 clk_gate_t1_mode_reg ( .CLK(clkper), .EN(
        N31), .ENCLK(net12165), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_2 clk_gate_tl1_s_reg ( .CLK(clkper), .EN(N50), 
        .ENCLK(net12171), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_1 clk_gate_th1_s_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12176), .TE(test_se) );
  timer1_a0_DW01_inc_0 add_278 ( .A(th1), .SUM({N75, N74, N73, N72, N71, N70, 
        N69, N68}) );
  timer1_a0_DW01_inc_1 add_244 ( .A(tl1), .SUM({N49, N48, N47, N46, N45, N44, 
        N43, N42}) );
  SDFFQX1 clk_count_reg_3_ ( .D(N98), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 clk_count_reg_2_ ( .D(N97), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 tl1_ov_ff_reg ( .D(n56), .SIN(th1[7]), .SMC(test_se), .C(clkper), 
        .Q(tl1_ov_ff) );
  SDFFQX1 clk_count_reg_1_ ( .D(n12), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 t1clr_reg ( .D(n57), .SIN(t1_tr1), .SMC(test_se), .C(clkper), .Q(
        t1clr) );
  SDFFQX1 clk_count_reg_0_ ( .D(N95), .SIN(test_si), .SMC(test_se), .C(clkper), 
        .Q(clk_count[0]) );
  SDFFQX1 th1_ov_ff_reg ( .D(n55), .SIN(t1clr), .SMC(test_se), .C(clkper), .Q(
        th1_ov_ff) );
  SDFFQX1 clk_ov12_reg ( .D(N100), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 t0_mode_reg_0_ ( .D(N36), .SIN(clk_ov12), .SMC(test_se), .C(net12165), .Q(t0_mode[0]) );
  SDFFQX1 t0_mode_reg_1_ ( .D(N37), .SIN(t0_mode[0]), .SMC(test_se), .C(
        net12165), .Q(t0_mode[1]) );
  SDFFQX1 th1_s_reg_7_ ( .D(N84), .SIN(th1[6]), .SMC(test_se), .C(net12176), 
        .Q(th1[7]) );
  SDFFQX1 t1_gate_reg ( .D(N32), .SIN(t1_tmod[2]), .SMC(test_se), .C(net12165), 
        .Q(t1_tmod[3]) );
  SDFFQX1 t1_ct_reg ( .D(N33), .SIN(t0_mode[1]), .SMC(test_se), .C(net12165), 
        .Q(t1_tmod[2]) );
  SDFFQX1 tl1_s_reg_7_ ( .D(N58), .SIN(tl1[6]), .SMC(test_se), .C(net12171), 
        .Q(tl1[7]) );
  SDFFQX1 tl1_s_reg_6_ ( .D(N57), .SIN(tl1[5]), .SMC(test_se), .C(net12171), 
        .Q(tl1[6]) );
  SDFFQX1 th1_s_reg_6_ ( .D(N83), .SIN(th1[5]), .SMC(test_se), .C(net12176), 
        .Q(th1[6]) );
  SDFFQX1 tl1_s_reg_5_ ( .D(N56), .SIN(tl1[4]), .SMC(test_se), .C(net12171), 
        .Q(tl1[5]) );
  SDFFQX1 th1_s_reg_5_ ( .D(N82), .SIN(th1[4]), .SMC(test_se), .C(net12176), 
        .Q(th1[5]) );
  SDFFQX1 th1_s_reg_4_ ( .D(N81), .SIN(th1[3]), .SMC(test_se), .C(net12176), 
        .Q(th1[4]) );
  SDFFQX1 tl1_s_reg_4_ ( .D(N55), .SIN(tl1[3]), .SMC(test_se), .C(net12171), 
        .Q(tl1[4]) );
  SDFFQX1 t1_mode_reg_1_ ( .D(N35), .SIN(t1_tmod[0]), .SMC(test_se), .C(
        net12165), .Q(t1_tmod[1]) );
  SDFFQX1 t1_mode_reg_0_ ( .D(N34), .SIN(t1_tmod[3]), .SMC(test_se), .C(
        net12165), .Q(t1_tmod[0]) );
  SDFFQX1 tl1_s_reg_3_ ( .D(N54), .SIN(tl1[2]), .SMC(test_se), .C(net12171), 
        .Q(tl1[3]) );
  SDFFQX1 th1_s_reg_3_ ( .D(N80), .SIN(th1[2]), .SMC(test_se), .C(net12176), 
        .Q(th1[3]) );
  SDFFQX1 t1_tr1_s_reg ( .D(n58), .SIN(t1_tf1), .SMC(test_se), .C(clkper), .Q(
        t1_tr1) );
  SDFFQX1 t1_tf1_s_reg ( .D(n54), .SIN(t1_tmod[1]), .SMC(test_se), .C(clkper), 
        .Q(t1_tf1) );
  SDFFQX1 tl1_s_reg_1_ ( .D(N52), .SIN(tl1[0]), .SMC(test_se), .C(net12171), 
        .Q(tl1[1]) );
  SDFFQX1 th1_s_reg_1_ ( .D(N78), .SIN(th1[0]), .SMC(test_se), .C(net12176), 
        .Q(th1[1]) );
  SDFFQX1 tl1_s_reg_2_ ( .D(N53), .SIN(tl1[1]), .SMC(test_se), .C(net12171), 
        .Q(tl1[2]) );
  SDFFQX1 th1_s_reg_2_ ( .D(N79), .SIN(th1[1]), .SMC(test_se), .C(net12176), 
        .Q(th1[2]) );
  SDFFQX1 tl1_s_reg_0_ ( .D(N51), .SIN(tl1_ov_ff), .SMC(test_se), .C(net12171), 
        .Q(tl1[0]) );
  SDFFQX1 th1_s_reg_0_ ( .D(N77), .SIN(th1_ov_ff), .SMC(test_se), .C(net12176), 
        .Q(th1[0]) );
  INVX1 U3 ( .A(n22), .Y(n10) );
  AND2X1 U4 ( .A(sfraddr[1]), .B(n50), .Y(n48) );
  NAND21X1 U5 ( .B(n44), .A(n8), .Y(n42) );
  NAND21X1 U6 ( .B(sfraddr[1]), .A(n50), .Y(n62) );
  NOR2X1 U7 ( .A(n4), .B(n62), .Y(N35) );
  NOR2X1 U8 ( .A(n3), .B(n62), .Y(N34) );
  NOR2X1 U9 ( .A(n5), .B(n62), .Y(N33) );
  NOR2X1 U10 ( .A(n6), .B(n62), .Y(N32) );
  NOR2X1 U11 ( .A(n1), .B(n62), .Y(N36) );
  NOR2X1 U12 ( .A(n2), .B(n62), .Y(N37) );
  NAND2X1 U13 ( .A(n8), .B(n62), .Y(N31) );
  INVX1 U14 ( .A(n8), .Y(n7) );
  NOR43XL U15 ( .B(sfrwe), .C(n63), .D(sfraddr[3]), .A(sfraddr[2]), .Y(n32) );
  NOR3XL U16 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n63) );
  NAND32X1 U17 ( .B(sfraddr[0]), .C(sfraddr[1]), .A(n32), .Y(n22) );
  NOR32XL U18 ( .B(n32), .C(sfraddr[0]), .A(n7), .Y(n50) );
  NAND4X1 U19 ( .A(sfraddr[2]), .B(sfraddr[0]), .C(n45), .D(n46), .Y(n44) );
  NOR4XL U20 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[4]), .D(sfraddr[1]), 
        .Y(n46) );
  AND2X1 U21 ( .A(sfraddr[3]), .B(sfrwe), .Y(n45) );
  INVX1 U22 ( .A(n52), .Y(n9) );
  AOI31X1 U23 ( .A(sfraddr[1]), .B(n32), .C(sfraddr[0]), .D(n7), .Y(n52) );
  NAND3X1 U24 ( .A(n42), .B(n8), .C(n43), .Y(N76) );
  INVX1 U25 ( .A(n43), .Y(n11) );
  INVX1 U26 ( .A(sfrdatai[4]), .Y(n3) );
  INVX1 U27 ( .A(sfrdatai[6]), .Y(n5) );
  INVX1 U28 ( .A(sfrdatai[7]), .Y(n6) );
  INVX1 U29 ( .A(sfrdatai[5]), .Y(n4) );
  INVX1 U30 ( .A(sfrdatai[0]), .Y(n1) );
  INVX1 U31 ( .A(sfrdatai[1]), .Y(n2) );
  INVX1 U32 ( .A(rst), .Y(n8) );
  INVX1 U33 ( .A(n38), .Y(n13) );
  OAI22BX1 U34 ( .B(N70), .A(n43), .D(sfrdatai[2]), .C(n42), .Y(N79) );
  OAI22BX1 U35 ( .B(N71), .A(n43), .D(sfrdatai[3]), .C(n42), .Y(N80) );
  NOR3XL U36 ( .A(n24), .B(n20), .C(n9), .Y(n47) );
  OR4X1 U37 ( .A(n49), .B(n47), .C(n48), .D(n7), .Y(N50) );
  NAND4X1 U38 ( .A(n18), .B(n44), .C(n8), .D(n20), .Y(n43) );
  ENOX1 U39 ( .A(n42), .B(n2), .C(N69), .D(n11), .Y(N78) );
  ENOX1 U40 ( .A(n42), .B(n3), .C(N72), .D(n11), .Y(N81) );
  ENOX1 U41 ( .A(n42), .B(n4), .C(N73), .D(n11), .Y(N82) );
  ENOX1 U42 ( .A(n5), .B(n42), .C(N74), .D(n11), .Y(N83) );
  OAI22X1 U43 ( .A(n7), .B(n25), .C(n23), .D(n15), .Y(n55) );
  OR2X1 U44 ( .A(newinstr), .B(n7), .Y(n23) );
  OAI21X1 U45 ( .B(n20), .C(n24), .A(n25), .Y(t1ov) );
  INVX1 U46 ( .A(n24), .Y(n18) );
  NAND2X1 U47 ( .A(n8), .B(n41), .Y(n38) );
  NAND2X1 U48 ( .A(n13), .B(n39), .Y(n36) );
  INVX1 U49 ( .A(n39), .Y(n14) );
  NOR2X1 U50 ( .A(n7), .B(n41), .Y(N100) );
  GEN3XL U51 ( .F(tl1_ov_ff), .G(n19), .E(n20), .D(n30), .C(t1ov), .B(n28), 
        .A(n10), .Y(n29) );
  NAND2X1 U52 ( .A(n20), .B(n15), .Y(n30) );
  AOI211X1 U53 ( .C(t0_mode[0]), .D(t0_mode[1]), .A(n10), .B(n31), .Y(n28) );
  NAND32X1 U54 ( .B(t1ack), .C(t1clr), .A(n8), .Y(n31) );
  ENOX1 U55 ( .A(n26), .B(n27), .C(t1_tf1), .D(n26), .Y(n54) );
  AOI31X1 U56 ( .A(n10), .B(n8), .C(sfrdatai[7]), .D(n28), .Y(n27) );
  NOR4XL U57 ( .A(n29), .B(t1clr), .C(n7), .D(t1ack), .Y(n26) );
  AO222X1 U58 ( .A(n47), .B(th1[0]), .C(n48), .D(sfrdatai[0]), .E(N42), .F(n49), .Y(N51) );
  AO222X1 U59 ( .A(n47), .B(th1[1]), .C(n48), .D(sfrdatai[1]), .E(N43), .F(n49), .Y(N52) );
  AO222X1 U60 ( .A(n47), .B(th1[2]), .C(n48), .D(sfrdatai[2]), .E(N44), .F(n49), .Y(N53) );
  AO222X1 U61 ( .A(n47), .B(th1[3]), .C(n48), .D(sfrdatai[3]), .E(N45), .F(n49), .Y(N54) );
  AO222X1 U62 ( .A(n47), .B(th1[4]), .C(n48), .D(sfrdatai[4]), .E(N46), .F(n49), .Y(N55) );
  AO222X1 U63 ( .A(n47), .B(th1[5]), .C(n48), .D(sfrdatai[5]), .E(N47), .F(n49), .Y(N56) );
  AO222X1 U64 ( .A(n47), .B(th1[6]), .C(n48), .D(sfrdatai[6]), .E(N48), .F(n49), .Y(N57) );
  AO222X1 U65 ( .A(n47), .B(th1[7]), .C(n48), .D(sfrdatai[7]), .E(N49), .F(n49), .Y(N58) );
  AOI211X1 U66 ( .C(t1_tmod[1]), .D(n18), .A(n51), .B(n9), .Y(n49) );
  NOR2X1 U67 ( .A(n7), .B(n21), .Y(n58) );
  AOI22X1 U68 ( .A(sfrdatai[6]), .B(n10), .C(t1_tr1), .D(n22), .Y(n21) );
  ENOX1 U69 ( .A(n42), .B(n1), .C(N68), .D(n11), .Y(N77) );
  ENOX1 U70 ( .A(n6), .B(n42), .C(N75), .D(n11), .Y(N84) );
  OAI22BX1 U71 ( .B(t1ack), .A(n7), .D(t1clr), .C(n23), .Y(n57) );
  OAI22AX1 U72 ( .D(tl1_ov_ff), .C(n23), .A(n7), .B(n24), .Y(n56) );
  NAND4X1 U73 ( .A(th1[2]), .B(th1[1]), .C(n33), .D(n34), .Y(n25) );
  NOR32XL U74 ( .B(th1[7]), .C(th1[6]), .A(n35), .Y(n34) );
  NOR32XL U75 ( .B(th1[0]), .C(n20), .A(n24), .Y(n33) );
  NAND3X1 U76 ( .A(th1[4]), .B(th1[3]), .C(th1[5]), .Y(n35) );
  NAND4X1 U77 ( .A(tl1[3]), .B(tl1[2]), .C(tl1[4]), .D(n53), .Y(n24) );
  NOR42XL U78 ( .C(tl1[1]), .D(tl1[0]), .A(n51), .B(n59), .Y(n53) );
  AOI32X1 U79 ( .A(tl1[6]), .B(tl1[5]), .C(tl1[7]), .D(n20), .E(n19), .Y(n59)
         );
  OAI211X1 U80 ( .C(n19), .D(n20), .A(clk_ov12), .B(n60), .Y(n51) );
  AOI211X1 U81 ( .C(t1_tmod[3]), .D(n64), .A(t1_tmod[2]), .B(n61), .Y(n60) );
  INVX1 U82 ( .A(int1ff), .Y(n64) );
  AOI21X1 U83 ( .B(t0_mode[1]), .C(t0_mode[0]), .A(t1_tr1), .Y(n61) );
  INVX1 U84 ( .A(t1_tmod[1]), .Y(n20) );
  INVX1 U85 ( .A(t1_tmod[0]), .Y(n19) );
  NAND2X1 U86 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n39) );
  OAI32X1 U87 ( .A(n38), .B(clk_count[2]), .C(n39), .D(n16), .E(n36), .Y(N97)
         );
  NAND3X1 U88 ( .A(n14), .B(n16), .C(clk_count[3]), .Y(n41) );
  OAI21X1 U89 ( .B(n17), .C(n36), .A(n37), .Y(N98) );
  NAND4X1 U90 ( .A(clk_count[2]), .B(n13), .C(n14), .D(n17), .Y(n37) );
  INVX1 U91 ( .A(clk_count[3]), .Y(n17) );
  INVX1 U92 ( .A(th1_ov_ff), .Y(n15) );
  INVX1 U93 ( .A(clk_count[2]), .Y(n16) );
  NOR2X1 U94 ( .A(clk_count[0]), .B(n38), .Y(N95) );
  INVX1 U95 ( .A(n40), .Y(n12) );
  OAI211X1 U96 ( .C(clk_count[0]), .D(clk_count[1]), .A(n13), .B(n39), .Y(n40)
         );
endmodule


module timer1_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module timer1_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer0_a0 ( clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, t0_tf0, 
        t0_tf1, sfrdatai, sfraddr, sfrwe, t0_tmod, t0_tr0, t0_tr1, tl0, th0, 
        test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t0_tmod;
  output [7:0] tl0;
  output [7:0] th0;
  input clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, sfrwe, test_si,
         test_se;
  output t0_tf0, t0_tf1, t0_tr0, t0_tr1;
  wire   t0clr, th0_ov_ff, tl0_ov_ff, t1clr, N39, N40, N41, N42, N43, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N101, N103, N104, clk_ov12, N106, net12193,
         net12199, net12204, n60, n61, n62, n63, n64, n65, n66, n67, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n68, n69, n70, n71, n72, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n73, n74, n75, n76, n77;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer0_a0_0 clk_gate_t0_ct_reg ( .CLK(clkper), .EN(N39), 
        .ENCLK(net12193), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_2 clk_gate_th0_s_reg ( .CLK(clkper), .EN(N55), 
        .ENCLK(net12199), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_1 clk_gate_tl0_s_reg ( .CLK(clkper), .EN(N79), 
        .ENCLK(net12204), .TE(test_se) );
  timer0_a0_DW01_inc_0 add_347 ( .A(tl0), .SUM({N78, N77, N76, N75, N74, N73, 
        N72, N71}) );
  timer0_a0_DW01_inc_1 add_309 ( .A(th0), .SUM({N54, N53, N52, N51, N50, N49, 
        N48, N47}) );
  SDFFQX1 tl0_ov_ff_reg ( .D(n64), .SIN(th0[7]), .SMC(test_se), .C(clkper), 
        .Q(tl0_ov_ff) );
  SDFFQX1 t1clr_reg ( .D(n63), .SIN(t0clr), .SMC(test_se), .C(clkper), .Q(
        t1clr) );
  SDFFQX1 t0clr_reg ( .D(n65), .SIN(t0_tr1), .SMC(test_se), .C(clkper), .Q(
        t0clr) );
  SDFFQX1 th0_ov_ff_reg ( .D(n61), .SIN(t1clr), .SMC(test_se), .C(clkper), .Q(
        th0_ov_ff) );
  SDFFQX1 clk_count_reg_3_ ( .D(N104), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 clk_count_reg_2_ ( .D(N103), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 clk_count_reg_1_ ( .D(n20), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 clk_count_reg_0_ ( .D(N101), .SIN(test_si), .SMC(test_se), .C(clkper), .Q(clk_count[0]) );
  SDFFQX1 clk_ov12_reg ( .D(N106), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 tl0_s_reg_7_ ( .D(N87), .SIN(tl0[6]), .SMC(test_se), .C(net12204), 
        .Q(tl0[7]) );
  SDFFQX1 th0_s_reg_7_ ( .D(N63), .SIN(th0[6]), .SMC(test_se), .C(net12199), 
        .Q(th0[7]) );
  SDFFQX1 tl0_s_reg_6_ ( .D(N86), .SIN(tl0[5]), .SMC(test_se), .C(net12204), 
        .Q(tl0[6]) );
  SDFFQX1 th0_s_reg_6_ ( .D(N62), .SIN(th0[5]), .SMC(test_se), .C(net12199), 
        .Q(th0[6]) );
  SDFFQX1 tl0_s_reg_5_ ( .D(N85), .SIN(tl0[4]), .SMC(test_se), .C(net12204), 
        .Q(tl0[5]) );
  SDFFQX1 th0_s_reg_5_ ( .D(N61), .SIN(th0[4]), .SMC(test_se), .C(net12199), 
        .Q(th0[5]) );
  SDFFQX1 th0_s_reg_4_ ( .D(N60), .SIN(th0[3]), .SMC(test_se), .C(net12199), 
        .Q(th0[4]) );
  SDFFQX1 tl0_s_reg_4_ ( .D(N84), .SIN(tl0[3]), .SMC(test_se), .C(net12204), 
        .Q(tl0[4]) );
  SDFFQX1 t0_gate_reg ( .D(N40), .SIN(t0_tmod[2]), .SMC(test_se), .C(net12193), 
        .Q(t0_tmod[3]) );
  SDFFQX1 tl0_s_reg_3_ ( .D(N83), .SIN(tl0[2]), .SMC(test_se), .C(net12204), 
        .Q(tl0[3]) );
  SDFFQX1 th0_s_reg_3_ ( .D(N59), .SIN(th0[2]), .SMC(test_se), .C(net12199), 
        .Q(th0[3]) );
  SDFFQX1 t0_tr1_s_reg ( .D(n66), .SIN(t0_tr0), .SMC(test_se), .C(clkper), .Q(
        t0_tr1) );
  SDFFQX1 t0_tr0_s_reg ( .D(n67), .SIN(t0_tf1), .SMC(test_se), .C(clkper), .Q(
        t0_tr0) );
  SDFFQX1 t0_tf0_s_reg ( .D(n60), .SIN(t0_tmod[1]), .SMC(test_se), .C(clkper), 
        .Q(t0_tf0) );
  SDFFQX1 t0_tf1_s_reg ( .D(n62), .SIN(t0_tf0), .SMC(test_se), .C(clkper), .Q(
        t0_tf1) );
  SDFFQX1 t0_ct_reg ( .D(N41), .SIN(clk_ov12), .SMC(test_se), .C(net12193), 
        .Q(t0_tmod[2]) );
  SDFFQX1 th0_s_reg_1_ ( .D(N57), .SIN(th0[0]), .SMC(test_se), .C(net12199), 
        .Q(th0[1]) );
  SDFFQX1 tl0_s_reg_2_ ( .D(N82), .SIN(tl0[1]), .SMC(test_se), .C(net12204), 
        .Q(tl0[2]) );
  SDFFQX1 tl0_s_reg_1_ ( .D(N81), .SIN(tl0[0]), .SMC(test_se), .C(net12204), 
        .Q(tl0[1]) );
  SDFFQX1 t0_mode_reg_1_ ( .D(N43), .SIN(t0_tmod[0]), .SMC(test_se), .C(
        net12193), .Q(t0_tmod[1]) );
  SDFFQX1 th0_s_reg_2_ ( .D(N58), .SIN(th0[1]), .SMC(test_se), .C(net12199), 
        .Q(th0[2]) );
  SDFFQX1 t0_mode_reg_0_ ( .D(N42), .SIN(t0_tmod[3]), .SMC(test_se), .C(
        net12193), .Q(t0_tmod[0]) );
  SDFFQX1 tl0_s_reg_0_ ( .D(N80), .SIN(tl0_ov_ff), .SMC(test_se), .C(net12204), 
        .Q(tl0[0]) );
  SDFFQX1 th0_s_reg_0_ ( .D(N56), .SIN(th0_ov_ff), .SMC(test_se), .C(net12199), 
        .Q(th0[0]) );
  NAND4XL U3 ( .A(sfraddr[2]), .B(sfrwe), .C(n55), .D(n56), .Y(n50) );
  INVX1 U4 ( .A(n25), .Y(n16) );
  NAND2X1 U5 ( .A(n17), .B(n10), .Y(n25) );
  INVX1 U6 ( .A(n31), .Y(n17) );
  NAND3X1 U7 ( .A(n2), .B(n1), .C(n41), .Y(n31) );
  NOR2X1 U8 ( .A(n11), .B(n16), .Y(n26) );
  AND4X1 U9 ( .A(sfraddr[1]), .B(n41), .C(n10), .D(n2), .Y(n44) );
  OR2X1 U10 ( .A(n50), .B(n15), .Y(n49) );
  AOI31X1 U11 ( .A(sfraddr[1]), .B(n2), .C(n41), .D(n12), .Y(n46) );
  NOR2X1 U12 ( .A(n4), .B(n57), .Y(N43) );
  NOR2X1 U13 ( .A(n3), .B(n57), .Y(N42) );
  NOR2X1 U14 ( .A(n5), .B(n57), .Y(N41) );
  NOR2X1 U15 ( .A(n6), .B(n57), .Y(N40) );
  NAND2X1 U16 ( .A(n10), .B(n57), .Y(N39) );
  INVX1 U17 ( .A(sfraddr[1]), .Y(n1) );
  INVX1 U18 ( .A(n11), .Y(n10) );
  NOR43XL U19 ( .B(sfrwe), .C(n58), .D(sfraddr[3]), .A(sfraddr[2]), .Y(n41) );
  NOR3XL U20 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n58) );
  OR4X1 U21 ( .A(n43), .B(n44), .C(n42), .D(n13), .Y(N79) );
  NAND4X1 U22 ( .A(sfraddr[0]), .B(n41), .C(n10), .D(n1), .Y(n57) );
  NOR4XL U23 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[4]), .D(sfraddr[1]), 
        .Y(n56) );
  AND2X1 U24 ( .A(sfraddr[3]), .B(n2), .Y(n55) );
  INVX1 U25 ( .A(n48), .Y(n18) );
  NAND3X1 U26 ( .A(n48), .B(n10), .C(n49), .Y(N55) );
  INVX1 U27 ( .A(sfraddr[0]), .Y(n2) );
  INVX1 U28 ( .A(sfrdatai[4]), .Y(n7) );
  INVX1 U29 ( .A(sfrdatai[6]), .Y(n9) );
  INVX1 U30 ( .A(sfrdatai[0]), .Y(n3) );
  INVX1 U31 ( .A(sfrdatai[1]), .Y(n4) );
  INVX1 U32 ( .A(sfrdatai[2]), .Y(n5) );
  INVX1 U33 ( .A(sfrdatai[3]), .Y(n6) );
  INVX1 U34 ( .A(sfrdatai[5]), .Y(n8) );
  BUFX3 U35 ( .A(rst), .Y(n11) );
  INVX1 U36 ( .A(t0ack), .Y(n19) );
  BUFX3 U37 ( .A(rst), .Y(n12) );
  BUFX3 U38 ( .A(rst), .Y(n15) );
  INVX1 U39 ( .A(n70), .Y(n21) );
  BUFX3 U40 ( .A(rst), .Y(n14) );
  BUFX3 U41 ( .A(rst), .Y(n13) );
  AOI31X1 U42 ( .A(n33), .B(n73), .C(n77), .D(n17), .Y(n37) );
  NOR32XL U43 ( .B(n47), .C(n46), .A(n45), .Y(n43) );
  AND2X1 U44 ( .A(n45), .B(n46), .Y(n42) );
  NAND3X1 U45 ( .A(n50), .B(n10), .C(n40), .Y(n48) );
  ENOX1 U46 ( .A(n4), .B(n49), .C(N48), .D(n18), .Y(N57) );
  ENOX1 U47 ( .A(n5), .B(n49), .C(N49), .D(n18), .Y(N58) );
  ENOX1 U48 ( .A(n6), .B(n49), .C(N50), .D(n18), .Y(N59) );
  ENOX1 U49 ( .A(n7), .B(n49), .C(N51), .D(n18), .Y(N60) );
  ENOX1 U50 ( .A(n9), .B(n49), .C(N53), .D(n18), .Y(N62) );
  ENOX1 U51 ( .A(n8), .B(n49), .C(N52), .D(n18), .Y(N61) );
  OAI22X1 U52 ( .A(n14), .B(n19), .C(n27), .D(n24), .Y(n65) );
  OAI22X1 U53 ( .A(n14), .B(n33), .C(n27), .D(n73), .Y(n61) );
  OR2X1 U54 ( .A(newinstr), .B(n15), .Y(n27) );
  INVX1 U55 ( .A(n28), .Y(n75) );
  NAND2X1 U56 ( .A(n10), .B(n59), .Y(n70) );
  NAND2X1 U57 ( .A(n21), .B(n71), .Y(n68) );
  INVX1 U58 ( .A(n71), .Y(n22) );
  NOR2X1 U59 ( .A(n12), .B(n59), .Y(N106) );
  OAI22BX1 U60 ( .B(n29), .A(n30), .D(t0_tf1), .C(n29), .Y(n62) );
  AOI32X1 U61 ( .A(n31), .B(n10), .C(n32), .D(sfrdatai[7]), .E(n16), .Y(n30)
         );
  OAI211X1 U62 ( .C(n77), .D(n33), .A(n26), .B(n32), .Y(n29) );
  NOR2X1 U63 ( .A(t1clr), .B(t1ack), .Y(n32) );
  ENOX1 U64 ( .A(n25), .B(n9), .C(n26), .D(t0_tr1), .Y(n66) );
  ENOX1 U65 ( .A(n25), .B(n7), .C(n26), .D(t0_tr0), .Y(n67) );
  OAI211X1 U66 ( .C(n25), .D(n8), .A(n34), .B(n35), .Y(n60) );
  NAND4X1 U67 ( .A(t0_tf0), .B(n26), .C(n19), .D(n24), .Y(n34) );
  NAND42X1 U68 ( .C(n36), .D(t0ack), .A(n24), .B(n10), .Y(n35) );
  OAI31XL U69 ( .A(n75), .B(tl0_ov_ff), .C(n77), .D(n37), .Y(n36) );
  AO222X1 U70 ( .A(n42), .B(th0[0]), .C(N71), .D(n43), .E(sfrdatai[0]), .F(n44), .Y(N80) );
  AO222X1 U71 ( .A(n42), .B(th0[1]), .C(N72), .D(n43), .E(sfrdatai[1]), .F(n44), .Y(N81) );
  AO222X1 U72 ( .A(n42), .B(th0[2]), .C(N73), .D(n43), .E(sfrdatai[2]), .F(n44), .Y(N82) );
  AO222X1 U73 ( .A(n42), .B(th0[3]), .C(N74), .D(n43), .E(sfrdatai[3]), .F(n44), .Y(N83) );
  AO222X1 U74 ( .A(n42), .B(th0[4]), .C(N75), .D(n43), .E(n44), .F(sfrdatai[4]), .Y(N84) );
  AO222X1 U75 ( .A(n42), .B(th0[5]), .C(N76), .D(n43), .E(n44), .F(sfrdatai[5]), .Y(N85) );
  AO222X1 U76 ( .A(n42), .B(th0[6]), .C(N77), .D(n43), .E(n44), .F(sfrdatai[6]), .Y(N86) );
  AO222X1 U77 ( .A(n42), .B(th0[7]), .C(N78), .D(n43), .E(n44), .F(sfrdatai[7]), .Y(N87) );
  OAI22BX1 U78 ( .B(N54), .A(n48), .D(sfrdatai[7]), .C(n49), .Y(N63) );
  ENOX1 U79 ( .A(n3), .B(n49), .C(N47), .D(n18), .Y(N56) );
  OAI22BX1 U80 ( .B(t1ack), .A(n13), .D(t1clr), .C(n27), .Y(n63) );
  OAI22AX1 U81 ( .D(tl0_ov_ff), .C(n27), .A(n14), .B(n28), .Y(n64) );
  NOR43XL U82 ( .B(t0_tr0), .C(n54), .D(clk_ov12), .A(t0_tmod[2]), .Y(n47) );
  NAND21X1 U83 ( .B(int0ff), .A(t0_tmod[3]), .Y(n54) );
  NAND4X1 U84 ( .A(tl0[3]), .B(tl0[2]), .C(tl0[4]), .D(n52), .Y(n28) );
  NOR43XL U85 ( .B(tl0[1]), .C(tl0[0]), .D(n47), .A(n53), .Y(n52) );
  AOI32X1 U86 ( .A(tl0[6]), .B(tl0[5]), .C(tl0[7]), .D(n77), .E(n76), .Y(n53)
         );
  INVX1 U87 ( .A(t0_tmod[0]), .Y(n76) );
  AOI21X1 U88 ( .B(n77), .C(n28), .A(n51), .Y(n40) );
  AOI31X1 U89 ( .A(t0_tmod[0]), .B(t0_tr1), .C(clk_ov12), .D(n77), .Y(n51) );
  NAND4X1 U90 ( .A(th0[3]), .B(th0[2]), .C(n38), .D(n39), .Y(n33) );
  AND4X1 U91 ( .A(th0[4]), .B(th0[5]), .C(th0[6]), .D(th0[7]), .Y(n39) );
  AND3X1 U92 ( .A(th0[1]), .B(n40), .C(th0[0]), .Y(n38) );
  NOR3XL U93 ( .A(n28), .B(t0_tmod[0]), .C(n77), .Y(n45) );
  INVX1 U94 ( .A(t0_tmod[1]), .Y(n77) );
  NAND2X1 U95 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n71) );
  OAI32X1 U96 ( .A(n70), .B(clk_count[2]), .C(n71), .D(n23), .E(n68), .Y(N103)
         );
  NAND3X1 U97 ( .A(n22), .B(n23), .C(clk_count[3]), .Y(n59) );
  OAI21X1 U98 ( .B(n74), .C(n68), .A(n69), .Y(N104) );
  NAND4X1 U99 ( .A(clk_count[2]), .B(n21), .C(n22), .D(n74), .Y(n69) );
  INVX1 U100 ( .A(clk_count[3]), .Y(n74) );
  INVX1 U101 ( .A(n72), .Y(n20) );
  OAI211X1 U102 ( .C(clk_count[0]), .D(clk_count[1]), .A(n21), .B(n71), .Y(n72) );
  INVX1 U103 ( .A(t0clr), .Y(n24) );
  INVX1 U104 ( .A(clk_count[2]), .Y(n23) );
  NOR2X1 U105 ( .A(clk_count[0]), .B(n70), .Y(N101) );
  INVX1 U106 ( .A(th0_ov_ff), .Y(n73) );
endmodule


module timer0_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module timer0_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module serial0_a0 ( t_shift_clk, r_shift_clk, clkper, rst, newinstr, rxd0ff, 
        t1ov, rxd0o, rxd0oe, txd0, sfrdatai, sfraddr, sfrwe, s0con, s0buf, 
        s0rell, s0relh, smod, bd, test_si, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] s0con;
  output [7:0] s0buf;
  output [7:0] s0rell;
  output [7:0] s0relh;
  input clkper, rst, newinstr, rxd0ff, t1ov, sfrwe, test_si, test_se;
  output t_shift_clk, r_shift_clk, rxd0o, rxd0oe, txd0, smod, bd;
  wire   r_clk_ov2, t1ov_ff, N59, ri_tmp, rxd0_val, s0con2_val, s0con2_tmp,
         ti_tmp, N109, N110, N111, N112, N113, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, baud_rate_ov, N142, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N166, N169, N170, N185, N186, N187, N188,
         N190, clk_ov12, N191, r_start, baud_r_count, baud_r2_clk, N207,
         t_baud_ov, t_start, N223, N224, N225, N227, N230, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N281, N282,
         N283, N284, N303, rxd0_fall, rxd0_ff, rxd0_fall_fl, receive_11_bits,
         N306, N307, N324, N325, N326, N327, N333, ri0_fall, ri0_ff, N360,
         N361, N362, N363, N364, N375, N376, N377, N378, N379, N380, N381,
         N382, N424, N425, N426, N427, N428, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, net12232, net12238, net12243, net12248,
         net12253, net12258, net12263, net12268, net12273, net12278, net12283,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n29, n67, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n246, n247, n248;
  wire   [3:0] r_baud_count;
  wire   [3:0] r_shift_count;
  wire   [3:0] t_shift_count;
  wire   [9:0] tim_baud;
  wire   [3:0] clk_count;
  wire   [3:0] t_baud_count;
  wire   [10:0] t_shift_reg;
  wire   [1:0] fluctuation_conter;
  wire   [2:0] rxd0_vec;
  wire   [7:0] r_shift_reg;

  MAJ3X1 U331 ( .A(rxd0_vec[1]), .B(rxd0_vec[0]), .C(rxd0_vec[2]), .Y(n172) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_0 clk_gate_s0con_s_reg ( .CLK(clkper), .EN(
        n67), .ENCLK(net12232), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_10 clk_gate_s0rell_s_reg ( .CLK(clkper), 
        .EN(N117), .ENCLK(net12238), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_9 clk_gate_s0relh_s_reg ( .CLK(clkper), .EN(
        N128), .ENCLK(net12243), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_8 clk_gate_tim_baud_reg ( .CLK(clkper), .EN(
        N166), .ENCLK(net12248), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_7 clk_gate_t_baud_count_reg ( .CLK(clkper), 
        .EN(N223), .ENCLK(net12253), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_6 clk_gate_t_shift_reg_reg ( .CLK(clkper), 
        .EN(N257), .ENCLK(net12258), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_5 clk_gate_rxd0_vec_reg ( .CLK(clkper), .EN(
        N324), .ENCLK(net12263), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_4 clk_gate_r_baud_count_reg ( .CLK(clkper), 
        .EN(N360), .ENCLK(net12268), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_3 clk_gate_r_shift_reg_reg ( .CLK(clkper), 
        .EN(n29), .ENCLK(net12273), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_2 clk_gate_r_shift_count_reg ( .CLK(clkper), 
        .EN(N428), .ENCLK(net12278), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_1 clk_gate_s0buf_r_reg ( .CLK(clkper), .EN(
        N471), .ENCLK(net12283), .TE(test_se) );
  serial0_a0_DW01_inc_0 add_584 ( .A(tim_baud), .SUM({N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145}) );
  SDFFQX1 r_shift_reg_reg_0_ ( .D(N375), .SIN(r_shift_count[3]), .SMC(test_se), 
        .C(net12273), .Q(r_shift_reg[0]) );
  SDFFQX1 t_shift_reg_reg_10_ ( .D(N268), .SIN(t_shift_reg[9]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[10]) );
  SDFFQX1 t_shift_reg_reg_1_ ( .D(N259), .SIN(t_shift_reg[0]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[1]) );
  SDFFQX1 ti_tmp_reg ( .D(n242), .SIN(t_start), .SMC(test_se), .C(clkper), .Q(
        ti_tmp) );
  SDFFQX1 t_shift_reg_reg_2_ ( .D(N260), .SIN(t_shift_reg[1]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[2]) );
  SDFFQX1 receive_11_bits_reg ( .D(n229), .SIN(r_start), .SMC(test_se), .C(
        clkper), .Q(receive_11_bits) );
  SDFFQX1 ri_tmp_reg ( .D(n238), .SIN(ri0_ff), .SMC(test_se), .C(clkper), .Q(
        ri_tmp) );
  SDFFQX1 baud_r_count_reg ( .D(n245), .SIN(baud_r2_clk), .SMC(test_se), .C(
        clkper), .Q(baud_r_count) );
  SDFFQX1 t_shift_reg_reg_0_ ( .D(N258), .SIN(t_shift_count[3]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[0]) );
  SDFFQX1 r_shift_reg_reg_7_ ( .D(N382), .SIN(r_shift_reg[6]), .SMC(test_se), 
        .C(net12273), .Q(r_shift_reg[7]) );
  SDFFQX1 r_shift_reg_reg_6_ ( .D(N381), .SIN(r_shift_reg[5]), .SMC(test_se), 
        .C(net12273), .Q(r_shift_reg[6]) );
  SDFFQX1 r_shift_reg_reg_5_ ( .D(N380), .SIN(r_shift_reg[4]), .SMC(test_se), 
        .C(net12273), .Q(r_shift_reg[5]) );
  SDFFQX1 r_shift_reg_reg_4_ ( .D(N379), .SIN(r_shift_reg[3]), .SMC(test_se), 
        .C(net12273), .Q(r_shift_reg[4]) );
  SDFFQX1 r_shift_reg_reg_3_ ( .D(N378), .SIN(r_shift_reg[2]), .SMC(test_se), 
        .C(net12273), .Q(r_shift_reg[3]) );
  SDFFQX1 r_shift_reg_reg_2_ ( .D(N377), .SIN(r_shift_reg[1]), .SMC(test_se), 
        .C(net12273), .Q(r_shift_reg[2]) );
  SDFFQX1 r_shift_reg_reg_1_ ( .D(N376), .SIN(r_shift_reg[0]), .SMC(test_se), 
        .C(net12273), .Q(r_shift_reg[1]) );
  SDFFQX1 fluctuation_conter_reg_1_ ( .D(n233), .SIN(fluctuation_conter[0]), 
        .SMC(test_se), .C(clkper), .Q(fluctuation_conter[1]) );
  SDFFQX1 t_shift_reg_reg_9_ ( .D(N267), .SIN(t_shift_reg[8]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[9]) );
  SDFFQX1 t_shift_reg_reg_8_ ( .D(N266), .SIN(t_shift_reg[7]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[8]) );
  SDFFQX1 t_shift_reg_reg_7_ ( .D(N265), .SIN(t_shift_reg[6]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[7]) );
  SDFFQX1 t_shift_reg_reg_6_ ( .D(N264), .SIN(t_shift_reg[5]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[6]) );
  SDFFQX1 t_shift_reg_reg_5_ ( .D(N263), .SIN(t_shift_reg[4]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[5]) );
  SDFFQX1 t_shift_reg_reg_4_ ( .D(N262), .SIN(t_shift_reg[3]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[4]) );
  SDFFQX1 t_shift_reg_reg_3_ ( .D(N261), .SIN(t_shift_reg[2]), .SMC(test_se), 
        .C(net12258), .Q(t_shift_reg[3]) );
  SDFFQX1 rxd0_vec_reg_2_ ( .D(N327), .SIN(rxd0_vec[1]), .SMC(test_se), .C(
        net12263), .Q(rxd0_vec[2]) );
  SDFFQX1 rxd0_vec_reg_1_ ( .D(N326), .SIN(rxd0_vec[0]), .SMC(test_se), .C(
        net12263), .Q(rxd0_vec[1]) );
  SDFFQX1 rxd0_ff_reg ( .D(N307), .SIN(rxd0_fall), .SMC(test_se), .C(clkper), 
        .Q(rxd0_ff) );
  SDFFQX1 rxd0_vec_reg_0_ ( .D(N325), .SIN(rxd0_val), .SMC(test_se), .C(
        net12263), .Q(rxd0_vec[0]) );
  SDFFQX1 ri0_ff_reg ( .D(n218), .SIN(ri0_fall), .SMC(test_se), .C(clkper), 
        .Q(ri0_ff) );
  SDFFQX1 rxd0_fall_fl_reg ( .D(n235), .SIN(ri_tmp), .SMC(test_se), .C(clkper), 
        .Q(rxd0_fall_fl) );
  SDFFQX1 ri0_fall_reg ( .D(n236), .SIN(receive_11_bits), .SMC(test_se), .C(
        clkper), .Q(ri0_fall) );
  SDFFQX1 t_shift_count_reg_3_ ( .D(N284), .SIN(t_shift_count[2]), .SMC(
        test_se), .C(net12258), .Q(t_shift_count[3]) );
  SDFFQX1 fluctuation_conter_reg_0_ ( .D(n234), .SIN(clk_ov12), .SMC(test_se), 
        .C(clkper), .Q(fluctuation_conter[0]) );
  SDFFQX1 s0con2_val_reg ( .D(n231), .SIN(s0con2_tmp), .SMC(test_se), .C(
        net12263), .Q(s0con2_val) );
  SDFFQX1 s0con2_tmp_reg ( .D(n232), .SIN(s0buf[7]), .SMC(test_se), .C(clkper), 
        .Q(s0con2_tmp) );
  SDFFQX1 clk_count_reg_2_ ( .D(N187), .SIN(clk_count[1]), .SMC(test_se), .C(
        clkper), .Q(clk_count[2]) );
  SDFFQX1 clk_count_reg_3_ ( .D(N188), .SIN(clk_count[2]), .SMC(test_se), .C(
        clkper), .Q(clk_count[3]) );
  SDFFQX1 clk_ov12_reg ( .D(N191), .SIN(clk_count[3]), .SMC(test_se), .C(
        clkper), .Q(clk_ov12) );
  SDFFQX1 t_baud_ov_reg ( .D(N230), .SIN(t_baud_count[3]), .SMC(test_se), .C(
        clkper), .Q(t_baud_ov) );
  SDFFQX1 tim_baud_reg_9_ ( .D(n64), .SIN(tim_baud[8]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[9]) );
  SDFFQX1 tim_baud_reg_8_ ( .D(n65), .SIN(tim_baud[7]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[8]) );
  SDFFQX1 t_shift_count_reg_1_ ( .D(N282), .SIN(t_shift_count[0]), .SMC(
        test_se), .C(net12258), .Q(t_shift_count[1]) );
  SDFFQX1 r_shift_count_reg_3_ ( .D(N427), .SIN(r_shift_count[2]), .SMC(
        test_se), .C(net12278), .Q(r_shift_count[3]) );
  SDFFQX1 t_shift_count_reg_0_ ( .D(N281), .SIN(t_baud_ov), .SMC(test_se), .C(
        net12258), .Q(t_shift_count[0]) );
  SDFFQX1 r_shift_count_reg_1_ ( .D(N425), .SIN(r_shift_count[0]), .SMC(
        test_se), .C(net12278), .Q(r_shift_count[1]) );
  SDFFQX1 t_shift_count_reg_2_ ( .D(N283), .SIN(t_shift_count[1]), .SMC(
        test_se), .C(net12258), .Q(t_shift_count[2]) );
  SDFFQX1 r_shift_count_reg_2_ ( .D(N426), .SIN(r_shift_count[1]), .SMC(
        test_se), .C(net12278), .Q(r_shift_count[2]) );
  SDFFQX1 t_baud_count_reg_3_ ( .D(N227), .SIN(t_baud_count[2]), .SMC(test_se), 
        .C(net12253), .Q(t_baud_count[3]) );
  SDFFQX1 t_baud_count_reg_1_ ( .D(N225), .SIN(t_baud_count[0]), .SMC(test_se), 
        .C(net12253), .Q(t_baud_count[1]) );
  SDFFQX1 clk_count_reg_1_ ( .D(N186), .SIN(clk_count[0]), .SMC(test_se), .C(
        clkper), .Q(clk_count[1]) );
  SDFFQX1 rxd0_val_reg ( .D(N333), .SIN(rxd0_ff), .SMC(test_se), .C(clkper), 
        .Q(rxd0_val) );
  SDFFQX1 t_baud_count_reg_0_ ( .D(N224), .SIN(t1ov_ff), .SMC(test_se), .C(
        net12253), .Q(t_baud_count[0]) );
  SDFFQX1 t_baud_count_reg_2_ ( .D(n61), .SIN(t_baud_count[1]), .SMC(test_se), 
        .C(net12253), .Q(t_baud_count[2]) );
  SDFFQX1 clk_count_reg_0_ ( .D(N185), .SIN(bd), .SMC(test_se), .C(clkper), 
        .Q(clk_count[0]) );
  SDFFQX1 rxd0_fall_reg ( .D(N306), .SIN(rxd0_fall_fl), .SMC(test_se), .C(
        clkper), .Q(rxd0_fall) );
  SDFFQX1 r_start_reg ( .D(n240), .SIN(r_shift_reg[7]), .SMC(test_se), .C(
        clkper), .Q(r_start) );
  SDFFQX1 baud_r2_clk_reg ( .D(N207), .SIN(test_si), .SMC(test_se), .C(clkper), 
        .Q(baud_r2_clk) );
  SDFFQX1 tim_baud_reg_2_ ( .D(N169), .SIN(tim_baud[1]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[2]) );
  SDFFQX1 tim_baud_reg_7_ ( .D(n66), .SIN(tim_baud[6]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[7]) );
  SDFFQX1 tim_baud_reg_5_ ( .D(n69), .SIN(tim_baud[4]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[5]) );
  SDFFQX1 tim_baud_reg_1_ ( .D(n71), .SIN(tim_baud[0]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[1]) );
  SDFFQX1 tim_baud_reg_6_ ( .D(n68), .SIN(tim_baud[5]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[6]) );
  SDFFQX1 tim_baud_reg_3_ ( .D(N170), .SIN(tim_baud[2]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[3]) );
  SDFFQX1 tim_baud_reg_4_ ( .D(n70), .SIN(tim_baud[3]), .SMC(test_se), .C(
        net12248), .Q(tim_baud[4]) );
  SDFFQX1 r_baud_count_reg_1_ ( .D(N362), .SIN(r_baud_count[0]), .SMC(test_se), 
        .C(net12268), .Q(r_baud_count[1]) );
  SDFFQX1 r_shift_count_reg_0_ ( .D(N424), .SIN(r_clk_ov2), .SMC(test_se), .C(
        net12278), .Q(r_shift_count[0]) );
  SDFFQX1 r_baud_count_reg_3_ ( .D(N364), .SIN(r_baud_count[2]), .SMC(test_se), 
        .C(net12268), .Q(r_baud_count[3]) );
  SDFFQX1 tim_baud_reg_0_ ( .D(n72), .SIN(ti_tmp), .SMC(test_se), .C(net12248), 
        .Q(tim_baud[0]) );
  SDFFQX1 r_baud_count_reg_0_ ( .D(N361), .SIN(fluctuation_conter[1]), .SMC(
        test_se), .C(net12268), .Q(r_baud_count[0]) );
  SDFFQX1 r_baud_count_reg_2_ ( .D(N363), .SIN(r_baud_count[1]), .SMC(test_se), 
        .C(net12268), .Q(r_baud_count[2]) );
  SDFFQX1 t1ov_ff_reg ( .D(N59), .SIN(smod), .SMC(test_se), .C(clkper), .Q(
        t1ov_ff) );
  SDFFQX1 baud_rate_ov_reg ( .D(N142), .SIN(baud_r_count), .SMC(test_se), .C(
        clkper), .Q(baud_rate_ov) );
  SDFFQX1 r_clk_ov2_reg ( .D(N190), .SIN(r_baud_count[3]), .SMC(test_se), .C(
        clkper), .Q(r_clk_ov2) );
  SDFFQX1 s0buf_r_reg_6_ ( .D(N478), .SIN(s0buf[5]), .SMC(test_se), .C(
        net12283), .Q(s0buf[6]) );
  SDFFQX1 s0buf_r_reg_7_ ( .D(N479), .SIN(s0buf[6]), .SMC(test_se), .C(
        net12283), .Q(s0buf[7]) );
  SDFFQX1 s0rell_s_reg_7_ ( .D(N125), .SIN(s0rell[6]), .SMC(test_se), .C(
        net12238), .Q(s0rell[7]) );
  SDFFQX1 s0rell_s_reg_6_ ( .D(N124), .SIN(s0rell[5]), .SMC(test_se), .C(
        net12238), .Q(s0rell[6]) );
  SDFFQX1 bd_s_reg ( .D(n25), .SIN(baud_rate_ov), .SMC(test_se), .C(clkper), 
        .Q(bd) );
  SDFFQX1 smod_s_reg ( .D(n244), .SIN(s0rell[7]), .SMC(test_se), .C(clkper), 
        .Q(smod) );
  SDFFQX1 s0relh_s_reg_7_ ( .D(N136), .SIN(s0relh[6]), .SMC(test_se), .C(
        net12243), .Q(s0relh[7]) );
  SDFFQX1 s0relh_s_reg_5_ ( .D(N134), .SIN(s0relh[4]), .SMC(test_se), .C(
        net12243), .Q(s0relh[5]) );
  SDFFQX1 s0buf_r_reg_5_ ( .D(N477), .SIN(s0buf[4]), .SMC(test_se), .C(
        net12283), .Q(s0buf[5]) );
  SDFFQX1 s0buf_r_reg_4_ ( .D(N476), .SIN(s0buf[3]), .SMC(test_se), .C(
        net12283), .Q(s0buf[4]) );
  SDFFQX1 s0relh_s_reg_6_ ( .D(N135), .SIN(s0relh[5]), .SMC(test_se), .C(
        net12243), .Q(s0relh[6]) );
  SDFFQX1 s0relh_s_reg_4_ ( .D(N133), .SIN(s0relh[3]), .SMC(test_se), .C(
        net12243), .Q(s0relh[4]) );
  SDFFQX1 s0rell_s_reg_5_ ( .D(N123), .SIN(s0rell[4]), .SMC(test_se), .C(
        net12238), .Q(s0rell[5]) );
  SDFFQX1 s0rell_s_reg_4_ ( .D(N122), .SIN(s0rell[3]), .SMC(test_se), .C(
        net12238), .Q(s0rell[4]) );
  SDFFQX1 s0con_s_reg_5_ ( .D(N111), .SIN(s0con[4]), .SMC(test_se), .C(
        net12232), .Q(s0con[5]) );
  SDFFQX1 s0con_s_reg_4_ ( .D(N110), .SIN(s0con[3]), .SMC(test_se), .C(
        net12232), .Q(s0con[4]) );
  SDFFQX1 s0relh_s_reg_3_ ( .D(N132), .SIN(s0relh[2]), .SMC(test_se), .C(
        net12243), .Q(s0relh[3]) );
  SDFFQX1 s0buf_r_reg_3_ ( .D(N475), .SIN(s0buf[2]), .SMC(test_se), .C(
        net12283), .Q(s0buf[3]) );
  SDFFQX1 s0rell_s_reg_3_ ( .D(N121), .SIN(s0rell[2]), .SMC(test_se), .C(
        net12238), .Q(s0rell[3]) );
  SDFFQX1 s0con_s_reg_3_ ( .D(N109), .SIN(s0con[2]), .SMC(test_se), .C(
        net12232), .Q(s0con[3]) );
  SDFFQX1 rxd0o_reg ( .D(N303), .SIN(rxd0_vec[2]), .SMC(test_se), .C(clkper), 
        .Q(rxd0o) );
  SDFFQX1 txd0_reg ( .D(n239), .SIN(tim_baud[9]), .SMC(test_se), .C(clkper), 
        .Q(txd0) );
  SDFFQX1 t_start_reg ( .D(n243), .SIN(t_shift_reg[10]), .SMC(test_se), .C(
        clkper), .Q(t_start) );
  SDFFQX1 s0con_s_reg_7_ ( .D(N113), .SIN(s0con[6]), .SMC(test_se), .C(
        net12232), .Q(s0con[7]) );
  SDFFQX1 s0con_s_reg_6_ ( .D(N112), .SIN(s0con[5]), .SMC(test_se), .C(
        net12232), .Q(s0con[6]) );
  SDFFQX1 s0rell_s_reg_2_ ( .D(N120), .SIN(s0rell[1]), .SMC(test_se), .C(
        net12238), .Q(s0rell[2]) );
  SDFFQX1 s0rell_s_reg_0_ ( .D(N118), .SIN(s0relh[7]), .SMC(test_se), .C(
        net12238), .Q(s0rell[0]) );
  SDFFQX1 s0con_s_reg_1_ ( .D(n241), .SIN(s0con[0]), .SMC(test_se), .C(clkper), 
        .Q(s0con[1]) );
  SDFFQX1 s0buf_r_reg_1_ ( .D(N473), .SIN(s0buf[0]), .SMC(test_se), .C(
        net12283), .Q(s0buf[1]) );
  SDFFQX1 s0rell_s_reg_1_ ( .D(N119), .SIN(s0rell[0]), .SMC(test_se), .C(
        net12238), .Q(s0rell[1]) );
  SDFFQX1 s0relh_s_reg_1_ ( .D(N130), .SIN(s0relh[0]), .SMC(test_se), .C(
        net12243), .Q(s0relh[1]) );
  SDFFQX1 s0relh_s_reg_2_ ( .D(N131), .SIN(s0relh[1]), .SMC(test_se), .C(
        net12243), .Q(s0relh[2]) );
  SDFFQX1 s0buf_r_reg_2_ ( .D(N474), .SIN(s0buf[1]), .SMC(test_se), .C(
        net12283), .Q(s0buf[2]) );
  SDFFQX1 s0buf_r_reg_0_ ( .D(N472), .SIN(rxd0o), .SMC(test_se), .C(net12283), 
        .Q(s0buf[0]) );
  SDFFQX1 s0relh_s_reg_0_ ( .D(N129), .SIN(s0con[7]), .SMC(test_se), .C(
        net12243), .Q(s0relh[0]) );
  SDFFQX1 s0con_s_reg_2_ ( .D(n230), .SIN(s0con[1]), .SMC(test_se), .C(clkper), 
        .Q(s0con[2]) );
  SDFFQX1 s0con_s_reg_0_ ( .D(n237), .SIN(s0con2_val), .SMC(test_se), .C(
        clkper), .Q(s0con[0]) );
  NAND2XL U3 ( .A(n214), .B(sfraddr[4]), .Y(n213) );
  NAND21XL U4 ( .B(sfraddr[4]), .A(n214), .Y(n215) );
  BUFX3 U5 ( .A(n83), .Y(n1) );
  BUFX3 U6 ( .A(n82), .Y(n2) );
  BUFX3 U7 ( .A(n227), .Y(n3) );
  AOI22AXL U8 ( .A(baud_r2_clk), .B(n223), .D(n95), .C(smod), .Y(n153) );
  AOI221XL U9 ( .A(n227), .B(r_shift_clk), .C(r_start), .D(n112), .E(n22), .Y(
        n149) );
  NOR41XL U10 ( .D(r_shift_count[0]), .A(r_shift_count[3]), .B(
        r_shift_count[1]), .C(r_shift_count[2]), .Y(n111) );
  INVX1 U11 ( .A(n126), .Y(n32) );
  INVX1 U12 ( .A(n103), .Y(n31) );
  INVX1 U13 ( .A(n104), .Y(n67) );
  NOR2X1 U14 ( .A(n143), .B(n20), .Y(n103) );
  NOR2X1 U15 ( .A(n21), .B(n103), .Y(n104) );
  NAND2X1 U16 ( .A(n143), .B(n15), .Y(n126) );
  INVX1 U17 ( .A(n180), .Y(n28) );
  NAND2X1 U18 ( .A(n16), .B(n215), .Y(N117) );
  NAND2X1 U19 ( .A(n15), .B(n213), .Y(N128) );
  INVX1 U20 ( .A(n20), .Y(n15) );
  INVX1 U21 ( .A(n21), .Y(n16) );
  INVX1 U22 ( .A(n20), .Y(n17) );
  INVX1 U23 ( .A(n20), .Y(n18) );
  NOR2X1 U24 ( .A(n192), .B(n19), .Y(n180) );
  INVX1 U25 ( .A(n175), .Y(n30) );
  NAND3X1 U26 ( .A(n4), .B(n6), .C(n93), .Y(n143) );
  OAI21X1 U27 ( .B(n31), .C(n13), .A(n24), .Y(N112) );
  NOR2X1 U28 ( .A(n31), .B(n10), .Y(N109) );
  NOR2X1 U29 ( .A(n31), .B(n11), .Y(N110) );
  NOR2X1 U30 ( .A(n31), .B(n12), .Y(N111) );
  NOR2X1 U31 ( .A(n14), .B(n31), .Y(N113) );
  NAND3X1 U32 ( .A(n28), .B(n17), .C(n175), .Y(N257) );
  INVX1 U33 ( .A(n184), .Y(n27) );
  OAI21X1 U34 ( .B(n8), .C(n213), .A(n24), .Y(N130) );
  OAI21X1 U35 ( .B(n7), .C(n213), .A(n24), .Y(N129) );
  OAI21X1 U36 ( .B(n7), .C(n215), .A(n18), .Y(N118) );
  OAI21X1 U37 ( .B(n10), .C(n215), .A(n24), .Y(N121) );
  OAI21X1 U38 ( .B(n11), .C(n215), .A(n24), .Y(N122) );
  OAI21X1 U39 ( .B(n13), .C(n215), .A(n24), .Y(N124) );
  OAI21X1 U40 ( .B(n14), .C(n215), .A(n24), .Y(N125) );
  NOR2X1 U41 ( .A(n9), .B(n215), .Y(N120) );
  NOR2X1 U42 ( .A(n8), .B(n215), .Y(N119) );
  NOR2X1 U43 ( .A(n12), .B(n215), .Y(N123) );
  NOR2X1 U44 ( .A(n9), .B(n213), .Y(N131) );
  NOR2X1 U45 ( .A(n10), .B(n213), .Y(N132) );
  NOR2X1 U46 ( .A(n11), .B(n213), .Y(N133) );
  NOR2X1 U47 ( .A(n14), .B(n213), .Y(N136) );
  NOR2X1 U48 ( .A(n12), .B(n213), .Y(N134) );
  NOR2X1 U49 ( .A(n13), .B(n213), .Y(N135) );
  INVX1 U50 ( .A(n6), .Y(n5) );
  INVX1 U51 ( .A(n150), .Y(n63) );
  INVX1 U52 ( .A(n24), .Y(n20) );
  INVX1 U53 ( .A(n18), .Y(n19) );
  INVX1 U54 ( .A(n23), .Y(n21) );
  INVX1 U55 ( .A(n23), .Y(n22) );
  NOR32XL U56 ( .B(sfraddr[3]), .C(sfrwe), .A(sfraddr[2]), .Y(n216) );
  NOR2X1 U57 ( .A(n28), .B(n227), .Y(n184) );
  NAND3X1 U58 ( .A(n192), .B(n17), .C(t_shift_clk), .Y(n175) );
  NAND3X1 U59 ( .A(n93), .B(n6), .C(sfraddr[0]), .Y(n192) );
  INVX1 U60 ( .A(n178), .Y(n26) );
  NOR3XL U61 ( .A(n22), .B(n5), .C(sfraddr[0]), .Y(n217) );
  INVX1 U62 ( .A(sfraddr[0]), .Y(n4) );
  INVX1 U63 ( .A(sfraddr[6]), .Y(n6) );
  INVX1 U64 ( .A(sfrdatai[4]), .Y(n11) );
  INVX1 U65 ( .A(sfrdatai[7]), .Y(n14) );
  INVX1 U66 ( .A(sfrdatai[6]), .Y(n13) );
  INVX1 U67 ( .A(sfrdatai[5]), .Y(n12) );
  INVX1 U68 ( .A(sfrdatai[3]), .Y(n10) );
  INVX1 U69 ( .A(sfrdatai[2]), .Y(n9) );
  INVX1 U70 ( .A(sfrdatai[0]), .Y(n7) );
  INVX1 U71 ( .A(sfrdatai[1]), .Y(n8) );
  NAND31X1 U72 ( .C(n138), .A(n227), .B(n15), .Y(n124) );
  NOR3XL U73 ( .A(n138), .B(rst), .C(n112), .Y(n150) );
  OAI211X1 U74 ( .C(n55), .D(n63), .A(n125), .B(n18), .Y(N471) );
  AND2X1 U75 ( .A(t1ov), .B(n16), .Y(N59) );
  INVX1 U76 ( .A(rst), .Y(n24) );
  OR2X1 U77 ( .A(n204), .B(n206), .Y(n205) );
  INVX1 U78 ( .A(n218), .Y(n246) );
  INVX1 U79 ( .A(rst), .Y(n23) );
  INVX1 U80 ( .A(n206), .Y(n52) );
  INVX1 U81 ( .A(n117), .Y(n227) );
  NOR2X1 U82 ( .A(n227), .B(n225), .Y(rxd0oe) );
  NOR2X1 U83 ( .A(n28), .B(n117), .Y(n178) );
  OAI222XL U84 ( .A(n31), .B(n7), .C(n126), .D(n37), .E(n103), .F(n246), .Y(
        n237) );
  OAI32X1 U85 ( .A(n223), .B(n20), .C(n96), .D(n14), .E(n33), .Y(n244) );
  INVX1 U86 ( .A(n96), .Y(n33) );
  NOR43XL U87 ( .B(n97), .C(n98), .D(n17), .A(sfraddr[3]), .Y(n96) );
  NOR3XL U88 ( .A(sfraddr[4]), .B(n5), .C(sfraddr[5]), .Y(n97) );
  INVX1 U89 ( .A(newinstr), .Y(n35) );
  OAI211X1 U90 ( .C(n117), .D(n138), .A(n35), .B(n18), .Y(n123) );
  OAI221X1 U91 ( .A(n123), .B(n37), .C(n55), .D(n124), .E(n125), .Y(n238) );
  OAI22X1 U92 ( .A(n63), .B(n46), .C(n125), .D(n45), .Y(N473) );
  OAI22X1 U93 ( .A(n63), .B(n45), .C(n125), .D(n44), .Y(N474) );
  OAI22X1 U94 ( .A(n63), .B(n44), .C(n125), .D(n43), .Y(N475) );
  OAI22X1 U95 ( .A(n63), .B(n43), .C(n125), .D(n42), .Y(N476) );
  OAI22X1 U96 ( .A(n63), .B(n42), .C(n125), .D(n41), .Y(N477) );
  OAI22X1 U97 ( .A(n63), .B(n41), .C(n125), .D(n40), .Y(N478) );
  OAI22X1 U98 ( .A(n63), .B(n40), .C(n56), .D(n125), .Y(N479) );
  NOR3XL U99 ( .A(n141), .B(n153), .C(n80), .Y(r_shift_clk) );
  NAND3X1 U100 ( .A(n111), .B(n247), .C(r_shift_clk), .Y(n138) );
  INVX1 U101 ( .A(n153), .Y(n60) );
  OAI22X1 U102 ( .A(n194), .B(n195), .C(n196), .D(n73), .Y(N227) );
  AOI21X1 U103 ( .B(n62), .C(n219), .A(n197), .Y(n196) );
  AOI211X1 U104 ( .C(n79), .D(n78), .A(n195), .B(n199), .Y(N225) );
  INVX1 U105 ( .A(n195), .Y(n62) );
  NOR2X1 U106 ( .A(n195), .B(n199), .Y(n197) );
  NOR32XL U107 ( .B(n116), .C(n16), .A(n3), .Y(n164) );
  OAI21X1 U108 ( .B(n57), .C(n52), .A(n23), .Y(n204) );
  NOR2X1 U109 ( .A(n60), .B(n133), .Y(n134) );
  NAND21X1 U110 ( .B(n151), .A(n149), .Y(N428) );
  NOR2X1 U111 ( .A(n247), .B(n19), .Y(n218) );
  OAI21X1 U112 ( .B(n22), .C(n115), .A(N382), .Y(n155) );
  AOI31X1 U113 ( .A(n155), .B(n3), .C(n165), .D(n164), .Y(n160) );
  OAI32X1 U114 ( .A(n58), .B(n52), .C(n204), .D(n57), .E(n205), .Y(N188) );
  NOR2X1 U115 ( .A(n152), .B(n227), .Y(n112) );
  OAI21X1 U116 ( .B(n153), .C(n248), .A(n24), .Y(N325) );
  AOI22AXL U117 ( .A(n111), .B(n112), .D(n113), .C(n108), .Y(n110) );
  NOR4XL U118 ( .A(n193), .B(n79), .C(rst), .D(n153), .Y(N230) );
  NAND3X1 U119 ( .A(n219), .B(n73), .C(n78), .Y(n193) );
  INVX1 U120 ( .A(n111), .Y(n74) );
  NOR2X1 U121 ( .A(n225), .B(n152), .Y(t_shift_clk) );
  OR2X1 U122 ( .A(n165), .B(n117), .Y(n113) );
  NAND2X1 U123 ( .A(n56), .B(n15), .Y(N382) );
  INVX1 U124 ( .A(n149), .Y(n29) );
  NOR2X1 U125 ( .A(n169), .B(n167), .Y(N363) );
  XNOR2XL U126 ( .A(n148), .B(n76), .Y(n169) );
  NAND3X1 U127 ( .A(n17), .B(n59), .C(n167), .Y(N360) );
  INVX1 U128 ( .A(n133), .Y(n50) );
  OAI21X1 U129 ( .B(n3), .C(n116), .A(n113), .Y(n151) );
  NAND32X1 U130 ( .B(n1), .C(n2), .A(n15), .Y(N166) );
  NOR2X1 U131 ( .A(n53), .B(n54), .Y(n206) );
  NAND3X1 U132 ( .A(n112), .B(n17), .C(n111), .Y(n125) );
  AOI21X1 U133 ( .B(n225), .C(n80), .A(n22), .Y(n119) );
  NOR2X1 U134 ( .A(n78), .B(n79), .Y(n199) );
  OAI21X1 U135 ( .B(n153), .C(n225), .A(n24), .Y(N223) );
  AOI211X1 U136 ( .C(n54), .D(n53), .A(n204), .B(n206), .Y(N186) );
  NOR3XL U137 ( .A(n38), .B(n22), .C(n95), .Y(N207) );
  NOR2X1 U138 ( .A(n54), .B(rst), .Y(N190) );
  NOR2X1 U139 ( .A(n20), .B(n94), .Y(n245) );
  XNOR2XL U140 ( .A(n38), .B(n95), .Y(n94) );
  NAND3X1 U141 ( .A(n117), .B(n39), .C(n119), .Y(N303) );
  NAND2X1 U142 ( .A(n153), .B(n15), .Y(N324) );
  INVX1 U143 ( .A(n141), .Y(n75) );
  NOR3XL U144 ( .A(n209), .B(n21), .C(n203), .Y(N142) );
  NAND2X1 U145 ( .A(n16), .B(n45), .Y(N376) );
  NAND2X1 U146 ( .A(n16), .B(n44), .Y(N377) );
  NAND2X1 U147 ( .A(n16), .B(n43), .Y(N378) );
  NAND2X1 U148 ( .A(n16), .B(n42), .Y(N379) );
  NAND2X1 U149 ( .A(n16), .B(n41), .Y(N380) );
  NAND2X1 U150 ( .A(n16), .B(n40), .Y(N381) );
  NAND2X1 U151 ( .A(n16), .B(n46), .Y(N375) );
  NOR2X1 U152 ( .A(n19), .B(n248), .Y(N307) );
  INVX1 U153 ( .A(n137), .Y(n55) );
  NOR2X1 U154 ( .A(s0con[7]), .B(s0con[6]), .Y(n117) );
  INVX1 U155 ( .A(t_start), .Y(n225) );
  AO222X1 U156 ( .A(sfrdatai[1]), .B(n103), .C(n32), .D(ti_tmp), .E(s0con[1]), 
        .F(n104), .Y(n241) );
  OAI21X1 U157 ( .B(n31), .C(n9), .A(n142), .Y(n230) );
  AOI33X1 U158 ( .A(s0con2_tmp), .B(n32), .C(s0con2_val), .D(n104), .E(n36), 
        .F(s0con[2]), .Y(n142) );
  INVX1 U159 ( .A(s0con2_tmp), .Y(n36) );
  OAI211X1 U160 ( .C(n7), .D(n26), .A(n23), .B(n190), .Y(N260) );
  AOI22X1 U161 ( .A(n184), .B(sfrdatai[1]), .C(t_shift_reg[3]), .D(n30), .Y(
        n190) );
  OAI211X1 U162 ( .C(n8), .D(n26), .A(n23), .B(n189), .Y(N261) );
  AOI22X1 U163 ( .A(n184), .B(sfrdatai[2]), .C(t_shift_reg[4]), .D(n30), .Y(
        n189) );
  OAI211X1 U164 ( .C(n26), .D(n12), .A(n23), .B(n185), .Y(N265) );
  AOI22X1 U165 ( .A(n184), .B(sfrdatai[6]), .C(t_shift_reg[8]), .D(n30), .Y(
        n185) );
  OAI211X1 U166 ( .C(n26), .D(n13), .A(n23), .B(n183), .Y(N266) );
  AOI22X1 U167 ( .A(n184), .B(sfrdatai[7]), .C(t_shift_reg[9]), .D(n30), .Y(
        n183) );
  OAI211X1 U168 ( .C(n26), .D(n10), .A(n18), .B(n187), .Y(N263) );
  AOI22X1 U169 ( .A(sfrdatai[4]), .B(n184), .C(t_shift_reg[6]), .D(n30), .Y(
        n187) );
  OAI211X1 U170 ( .C(n26), .D(n11), .A(n23), .B(n186), .Y(N264) );
  AOI22X1 U171 ( .A(sfrdatai[5]), .B(n184), .C(t_shift_reg[7]), .D(n30), .Y(
        n186) );
  OAI211X1 U172 ( .C(n9), .D(n26), .A(n18), .B(n188), .Y(N262) );
  AOI22X1 U173 ( .A(sfrdatai[3]), .B(n184), .C(t_shift_reg[5]), .D(n30), .Y(
        n188) );
  GEN2XL U174 ( .D(t_shift_count[1]), .E(t_shift_count[0]), .C(n177), .B(n30), 
        .A(n178), .Y(N282) );
  INVX1 U175 ( .A(n91), .Y(n25) );
  AOI32X1 U176 ( .A(bd), .B(n17), .C(n92), .D(n34), .E(sfrdatai[7]), .Y(n91)
         );
  INVX1 U177 ( .A(n92), .Y(n34) );
  NAND4X1 U178 ( .A(n5), .B(n93), .C(n15), .D(n4), .Y(n92) );
  OAI21X1 U179 ( .B(t_shift_count[0]), .C(n175), .A(n179), .Y(N281) );
  OAI21X1 U180 ( .B(s0con[7]), .C(n226), .A(n180), .Y(n179) );
  OAI21X1 U181 ( .B(n174), .C(n175), .A(n28), .Y(N284) );
  XOR2X1 U182 ( .A(n100), .B(t_shift_count[3]), .Y(n174) );
  NAND3X1 U183 ( .A(n27), .B(n17), .C(n182), .Y(N267) );
  AOI22X1 U184 ( .A(t_shift_reg[10]), .B(n30), .C(n180), .D(sfrdatai[7]), .Y(
        n182) );
  OAI2B11X1 U185 ( .D(t_shift_reg[1]), .C(n175), .A(n28), .B(n23), .Y(N258) );
  AOI21X1 U186 ( .B(n100), .C(n176), .A(n175), .Y(N283) );
  NAND21X1 U187 ( .B(n177), .A(t_shift_count[2]), .Y(n176) );
  OAI211X1 U188 ( .C(n7), .D(n27), .A(n18), .B(n191), .Y(N259) );
  NAND2X1 U189 ( .A(t_shift_reg[2]), .B(n30), .Y(n191) );
  NAND2X1 U190 ( .A(n28), .B(n99), .Y(n243) );
  OAI211X1 U191 ( .C(t_shift_count[3]), .D(n100), .A(n23), .B(t_start), .Y(n99) );
  NAND3X1 U192 ( .A(n175), .B(n17), .C(n181), .Y(N268) );
  OAI21X1 U193 ( .B(s0con[3]), .C(n228), .A(n180), .Y(n181) );
  NOR2X1 U194 ( .A(n20), .B(n101), .Y(n242) );
  AOI32X1 U195 ( .A(t_shift_count[0]), .B(t_shift_clk), .C(n102), .D(ti_tmp), 
        .E(n35), .Y(n101) );
  NOR3XL U196 ( .A(t_shift_count[1]), .B(t_shift_count[3]), .C(
        t_shift_count[2]), .Y(n102) );
  ENOX1 U197 ( .A(n124), .B(n136), .C(n136), .D(s0con2_tmp), .Y(n232) );
  OAI21X1 U198 ( .B(n124), .C(n137), .A(n123), .Y(n136) );
  OAI22AX1 U199 ( .D(n201), .C(t1ov_ff), .A(n201), .B(n202), .Y(n95) );
  NOR2X1 U200 ( .A(n226), .B(bd), .Y(n201) );
  AOI221XL U201 ( .A(s0con[6]), .B(n221), .C(n203), .D(n226), .E(n117), .Y(
        n202) );
  ENOX1 U202 ( .A(n125), .B(n46), .C(r_shift_reg[0]), .D(n150), .Y(N472) );
  INVX1 U203 ( .A(s0con[6]), .Y(n226) );
  NOR2X1 U204 ( .A(s0relh[7]), .B(r_clk_ov2), .Y(n203) );
  OAI211X1 U205 ( .C(n222), .D(n194), .A(t_start), .B(n200), .Y(n195) );
  NOR2X1 U206 ( .A(rst), .B(n153), .Y(n200) );
  NAND2X1 U207 ( .A(n147), .B(n154), .Y(n141) );
  OAI32X1 U208 ( .A(n77), .B(s0relh[6]), .C(r_baud_count[2]), .D(n76), .E(n222), .Y(n154) );
  OAI32X1 U209 ( .A(n49), .B(n20), .C(n139), .D(n56), .E(n124), .Y(n231) );
  INVX1 U210 ( .A(s0con2_val), .Y(n49) );
  NOR4XL U211 ( .A(n140), .B(n74), .C(n141), .D(n80), .Y(n139) );
  NAND3X1 U212 ( .A(n227), .B(n247), .C(n137), .Y(n140) );
  INVX1 U213 ( .A(s0relh[6]), .Y(n222) );
  OAI21X1 U214 ( .B(n80), .C(n105), .A(n106), .Y(n240) );
  OAI211X1 U215 ( .C(n107), .D(n108), .A(n105), .B(n18), .Y(n106) );
  NAND41X1 U216 ( .D(n107), .A(n17), .B(n109), .C(n110), .Y(n105) );
  NOR3XL U217 ( .A(n227), .B(r_start), .C(n116), .Y(n107) );
  NAND4X1 U218 ( .A(n75), .B(n114), .C(n60), .D(n227), .Y(n109) );
  OAI21BBX1 U219 ( .A(n115), .B(rxd0_val), .C(n74), .Y(n114) );
  NOR2X1 U220 ( .A(t_baud_count[0]), .B(n195), .Y(N224) );
  INVX1 U221 ( .A(baud_rate_ov), .Y(n221) );
  INVX1 U222 ( .A(n198), .Y(n61) );
  AOI32X1 U223 ( .A(n62), .B(n219), .C(n199), .D(t_baud_count[2]), .E(n197), 
        .Y(n198) );
  NAND31X1 U224 ( .C(n152), .A(ri0_fall), .B(s0con[4]), .Y(n116) );
  OAI22X1 U225 ( .A(s0relh[7]), .B(n221), .C(n209), .D(n224), .Y(n82) );
  AOI21X1 U226 ( .B(n224), .C(r_clk_ov2), .A(n82), .Y(n83) );
  GEN2XL U227 ( .D(n50), .E(n47), .C(n134), .B(fluctuation_conter[1]), .A(n135), .Y(n233) );
  NOR4XL U228 ( .A(fluctuation_conter[1]), .B(n134), .C(n133), .D(n47), .Y(
        n135) );
  INVX1 U229 ( .A(n84), .Y(n65) );
  AOI221XL U230 ( .A(s0relh[0]), .B(n82), .C(N153), .D(n83), .E(n22), .Y(n84)
         );
  OAI22X1 U231 ( .A(t_baud_ov), .B(n117), .C(clk_ov12), .D(n227), .Y(n152) );
  NAND2X1 U232 ( .A(rxd0_fall_fl), .B(n15), .Y(n133) );
  NAND4X1 U233 ( .A(r_start), .B(n60), .C(n15), .D(n59), .Y(n167) );
  OAI32X1 U234 ( .A(n204), .B(clk_count[2]), .C(n52), .D(n58), .E(n205), .Y(
        N187) );
  OAI32X1 U235 ( .A(n133), .B(fluctuation_conter[0]), .C(n134), .D(n51), .E(
        n47), .Y(n234) );
  INVX1 U236 ( .A(n134), .Y(n51) );
  OAI32X1 U237 ( .A(n47), .B(n59), .C(n133), .D(r_baud_count[0]), .E(n167), 
        .Y(N361) );
  OAI32X1 U238 ( .A(n48), .B(n59), .C(n133), .D(n170), .E(n167), .Y(N362) );
  INVX1 U239 ( .A(fluctuation_conter[1]), .Y(n48) );
  AOI21X1 U240 ( .B(r_baud_count[1]), .C(n220), .A(n147), .Y(n170) );
  NOR2X1 U241 ( .A(n220), .B(r_baud_count[1]), .Y(n147) );
  NOR4XL U242 ( .A(rxd0_fall), .B(receive_11_bits), .C(r_start), .D(n173), .Y(
        N306) );
  AOI31X1 U243 ( .A(n17), .B(n248), .C(rxd0_ff), .D(n50), .Y(n173) );
  INVX1 U244 ( .A(r_baud_count[2]), .Y(n76) );
  OAI22AX1 U245 ( .D(n155), .C(n156), .A(n21), .B(n157), .Y(N427) );
  AOI21BBXL U246 ( .B(n3), .C(n156), .A(n151), .Y(n157) );
  AOI21X1 U247 ( .B(n158), .C(r_shift_count[3]), .A(n108), .Y(n156) );
  OAI22X1 U248 ( .A(n20), .B(n113), .C(n162), .D(n163), .Y(N425) );
  AOI21X1 U249 ( .B(r_shift_count[0]), .C(r_shift_count[1]), .A(n161), .Y(n162) );
  AOI21X1 U250 ( .B(n155), .C(n3), .A(n164), .Y(n163) );
  OAI21BX1 U251 ( .C(ri0_fall), .B(n127), .A(n128), .Y(n236) );
  NAND4X1 U252 ( .A(ri0_ff), .B(n127), .C(n15), .D(n247), .Y(n128) );
  GEN2XL U253 ( .D(ri0_ff), .E(n117), .C(n19), .B(n246), .A(n112), .Y(n127) );
  AOI21X1 U254 ( .B(n158), .C(n159), .A(n160), .Y(N426) );
  NAND21X1 U255 ( .B(n161), .A(r_shift_count[2]), .Y(n159) );
  NAND41X1 U256 ( .D(n210), .A(tim_baud[8]), .B(tim_baud[9]), .C(n211), .Y(
        n209) );
  NAND3X1 U257 ( .A(tim_baud[6]), .B(tim_baud[5]), .C(tim_baud[7]), .Y(n210)
         );
  NOR32XL U258 ( .B(tim_baud[4]), .C(tim_baud[3]), .A(n212), .Y(n211) );
  NAND3X1 U259 ( .A(tim_baud[1]), .B(tim_baud[0]), .C(tim_baud[2]), .Y(n212)
         );
  OAI21BBX1 U260 ( .A(n60), .B(rxd0_vec[0]), .C(n18), .Y(N326) );
  OAI21BBX1 U261 ( .A(n60), .B(rxd0_vec[1]), .C(n18), .Y(N327) );
  INVX1 U262 ( .A(r_baud_count[3]), .Y(n77) );
  INVX1 U263 ( .A(r_baud_count[0]), .Y(n220) );
  NOR2X1 U264 ( .A(n166), .B(n167), .Y(N364) );
  XNOR2XL U265 ( .A(r_baud_count[3]), .B(n168), .Y(n166) );
  NOR2X1 U266 ( .A(n76), .B(n148), .Y(n168) );
  NOR2X1 U267 ( .A(rst), .B(n208), .Y(N169) );
  AOI22X1 U268 ( .A(N147), .B(n83), .C(s0rell[2]), .D(n2), .Y(n208) );
  NOR2X1 U269 ( .A(n19), .B(n207), .Y(N170) );
  AOI22X1 U270 ( .A(N148), .B(n1), .C(s0rell[3]), .D(n2), .Y(n207) );
  NOR2X1 U271 ( .A(r_shift_count[0]), .B(n160), .Y(N424) );
  INVX1 U272 ( .A(smod), .Y(n223) );
  INVX1 U273 ( .A(n81), .Y(n64) );
  AOI221XL U274 ( .A(s0relh[1]), .B(n82), .C(N154), .D(n83), .E(n22), .Y(n81)
         );
  INVX1 U275 ( .A(n89), .Y(n68) );
  AOI221XL U276 ( .A(s0rell[6]), .B(n82), .C(N151), .D(n83), .E(n21), .Y(n89)
         );
  INVX1 U277 ( .A(n86), .Y(n71) );
  AOI221XL U278 ( .A(s0rell[1]), .B(n82), .C(N146), .D(n83), .E(n21), .Y(n86)
         );
  INVX1 U279 ( .A(n88), .Y(n69) );
  AOI221XL U280 ( .A(s0rell[5]), .B(n82), .C(N150), .D(n83), .E(n21), .Y(n88)
         );
  INVX1 U281 ( .A(n90), .Y(n66) );
  AOI221XL U282 ( .A(s0rell[7]), .B(n82), .C(N152), .D(n83), .E(n22), .Y(n90)
         );
  INVX1 U283 ( .A(n87), .Y(n70) );
  AOI221XL U284 ( .A(s0rell[4]), .B(n82), .C(N149), .D(n83), .E(n21), .Y(n87)
         );
  INVX1 U285 ( .A(n85), .Y(n72) );
  AOI221XL U286 ( .A(s0rell[0]), .B(n82), .C(N145), .D(n83), .E(n21), .Y(n85)
         );
  NAND21X1 U287 ( .B(r_shift_count[2]), .A(n161), .Y(n158) );
  AND4X1 U288 ( .A(n58), .B(n53), .C(N190), .D(clk_count[3]), .Y(N191) );
  NAND2X1 U289 ( .A(s0con[5]), .B(n56), .Y(n137) );
  AND2X1 U290 ( .A(rxd0_ff), .B(n111), .Y(n132) );
  NOR42XL U291 ( .C(r_shift_count[3]), .D(r_shift_count[1]), .A(
        r_shift_count[0]), .B(r_shift_count[2]), .Y(n115) );
  NOR2X1 U292 ( .A(r_shift_count[0]), .B(r_shift_count[1]), .Y(n161) );
  NOR31X1 U293 ( .C(t_shift_count[0]), .A(t_shift_count[2]), .B(
        t_shift_count[1]), .Y(n122) );
  OAI21X1 U294 ( .B(n3), .C(n248), .A(n171), .Y(N333) );
  AOI21X1 U295 ( .B(n172), .C(n3), .A(n22), .Y(n171) );
  AOI211X1 U296 ( .C(n129), .D(n130), .A(n131), .B(n21), .Y(n235) );
  AOI22X1 U297 ( .A(s0relh[6]), .B(r_baud_count[2]), .C(r_baud_count[3]), .D(
        n222), .Y(n131) );
  OAI21BBX1 U298 ( .A(rxd0_fall), .B(n108), .C(rxd0_fall_fl), .Y(n129) );
  NAND4X1 U299 ( .A(n248), .B(n228), .C(s0con[6]), .D(n132), .Y(n130) );
  NOR2X1 U300 ( .A(n158), .B(r_shift_count[3]), .Y(n108) );
  INVX1 U301 ( .A(s0con[0]), .Y(n247) );
  INVX1 U302 ( .A(rxd0_val), .Y(n56) );
  NOR3XL U303 ( .A(n228), .B(n22), .C(n144), .Y(n229) );
  AOI32X1 U304 ( .A(n145), .B(n146), .C(receive_11_bits), .D(n111), .E(n75), 
        .Y(n144) );
  NAND31X1 U305 ( .C(n148), .A(s0relh[6]), .B(n76), .Y(n145) );
  NAND4X1 U306 ( .A(n147), .B(r_baud_count[2]), .C(n77), .D(n222), .Y(n146) );
  INVX1 U307 ( .A(r_start), .Y(n80) );
  OAI211X1 U308 ( .C(n117), .D(n39), .A(n118), .B(n119), .Y(n239) );
  OAI21BBX1 U309 ( .A(n120), .B(n121), .C(n117), .Y(n118) );
  OAI31XL U310 ( .A(clk_count[0]), .B(clk_count[2]), .C(clk_count[1]), .D(
        clk_count[3]), .Y(n121) );
  AOI33X1 U311 ( .A(txd0), .B(t_shift_count[3]), .C(n122), .D(n58), .E(n57), 
        .F(n52), .Y(n120) );
  INVX1 U312 ( .A(clk_count[0]), .Y(n54) );
  INVX1 U313 ( .A(t_baud_count[0]), .Y(n79) );
  NAND2X1 U314 ( .A(rxd0_fall), .B(s0con[4]), .Y(n165) );
  NAND3X1 U315 ( .A(n199), .B(n73), .C(t_baud_count[2]), .Y(n194) );
  INVX1 U316 ( .A(clk_count[1]), .Y(n53) );
  INVX1 U317 ( .A(t_baud_count[1]), .Y(n78) );
  INVX1 U318 ( .A(t_baud_count[3]), .Y(n73) );
  INVX1 U319 ( .A(s0relh[7]), .Y(n224) );
  NOR2X1 U320 ( .A(clk_count[0]), .B(n204), .Y(N185) );
  NAND21X1 U321 ( .B(t_shift_count[2]), .A(n177), .Y(n100) );
  NOR2X1 U322 ( .A(t_shift_count[1]), .B(t_shift_count[0]), .Y(n177) );
  INVX1 U323 ( .A(rxd0ff), .Y(n248) );
  NAND2X1 U324 ( .A(r_baud_count[1]), .B(r_baud_count[0]), .Y(n148) );
  INVX1 U325 ( .A(rxd0_fall), .Y(n59) );
  INVX1 U326 ( .A(s0con[7]), .Y(n228) );
  INVX1 U327 ( .A(fluctuation_conter[0]), .Y(n47) );
  INVX1 U328 ( .A(clk_count[2]), .Y(n58) );
  INVX1 U329 ( .A(t_baud_count[2]), .Y(n219) );
  INVX1 U330 ( .A(clk_count[3]), .Y(n57) );
  INVX1 U332 ( .A(r_shift_reg[1]), .Y(n46) );
  INVX1 U333 ( .A(r_shift_reg[2]), .Y(n45) );
  INVX1 U334 ( .A(r_shift_reg[3]), .Y(n44) );
  INVX1 U335 ( .A(r_shift_reg[4]), .Y(n43) );
  INVX1 U336 ( .A(r_shift_reg[5]), .Y(n42) );
  INVX1 U337 ( .A(r_shift_reg[6]), .Y(n41) );
  INVX1 U338 ( .A(r_shift_reg[7]), .Y(n40) );
  INVX1 U339 ( .A(baud_r_count), .Y(n38) );
  INVX1 U340 ( .A(t_shift_reg[0]), .Y(n39) );
  INVX1 U341 ( .A(ri_tmp), .Y(n37) );
  AND4XL U342 ( .A(sfraddr[1]), .B(n216), .C(sfraddr[5]), .D(n217), .Y(n214)
         );
  AND4XL U343 ( .A(sfrwe), .B(sfraddr[2]), .C(sfraddr[1]), .D(sfraddr[0]), .Y(
        n98) );
  NOR42XL U344 ( .C(sfraddr[4]), .D(n216), .A(sfraddr[1]), .B(sfraddr[5]), .Y(
        n93) );
endmodule


module serial0_a0_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ports_a0 ( clkper, rst, port0, sfrdatai, sfraddr, sfrwe, test_si, 
        test_se );
  output [7:0] port0;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkper, rst, sfrwe, test_si, test_se;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, net12300, n2, n3, n4, n1;

  SNPS_CLOCK_GATE_HIGH_ports_a0 clk_gate_p0_reg ( .CLK(clkper), .EN(N2), 
        .ENCLK(net12300), .TE(test_se) );
  SDFFQX1 p0_reg_7_ ( .D(N10), .SIN(port0[6]), .SMC(test_se), .C(net12300), 
        .Q(port0[7]) );
  SDFFQX1 p0_reg_6_ ( .D(N9), .SIN(port0[5]), .SMC(test_se), .C(net12300), .Q(
        port0[6]) );
  SDFFQX1 p0_reg_4_ ( .D(N7), .SIN(port0[3]), .SMC(test_se), .C(net12300), .Q(
        port0[4]) );
  SDFFQX1 p0_reg_5_ ( .D(N8), .SIN(port0[4]), .SMC(test_se), .C(net12300), .Q(
        port0[5]) );
  SDFFQX1 p0_reg_3_ ( .D(N6), .SIN(port0[2]), .SMC(test_se), .C(net12300), .Q(
        port0[3]) );
  SDFFQX1 p0_reg_2_ ( .D(N5), .SIN(port0[1]), .SMC(test_se), .C(net12300), .Q(
        port0[2]) );
  SDFFQX1 p0_reg_1_ ( .D(N4), .SIN(port0[0]), .SMC(test_se), .C(net12300), .Q(
        port0[1]) );
  SDFFQX1 p0_reg_0_ ( .D(N3), .SIN(test_si), .SMC(test_se), .C(net12300), .Q(
        port0[0]) );
  NOR21XL U2 ( .B(sfrdatai[1]), .A(n2), .Y(N4) );
  NOR21XL U3 ( .B(sfrdatai[2]), .A(n2), .Y(N5) );
  NOR21XL U4 ( .B(sfrdatai[0]), .A(n2), .Y(N3) );
  NOR21XL U5 ( .B(sfrdatai[3]), .A(n2), .Y(N6) );
  NOR21XL U6 ( .B(sfrdatai[5]), .A(n2), .Y(N8) );
  NOR21XL U7 ( .B(sfrdatai[4]), .A(n2), .Y(N7) );
  NOR21XL U8 ( .B(sfrdatai[6]), .A(n2), .Y(N9) );
  NOR21XL U9 ( .B(sfrdatai[7]), .A(n2), .Y(N10) );
  NAND2X1 U10 ( .A(n1), .B(n2), .Y(N2) );
  INVX1 U11 ( .A(rst), .Y(n1) );
  NAND42X1 U12 ( .C(sfraddr[3]), .D(sfraddr[2]), .A(n3), .B(n4), .Y(n2) );
  NOR3XL U13 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n3) );
  NOR42XL U14 ( .C(sfrwe), .D(n1), .A(sfraddr[1]), .B(sfraddr[0]), .Y(n4) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ports_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mdu_a0 ( clkper, rst, mdubsy, sfrdatai, sfraddr, sfrwe, sfroe, arcon, 
        md0, md1, md2, md3, md4, md5, test_si, test_so, test_se );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] arcon;
  output [7:0] md0;
  output [7:0] md1;
  output [7:0] md2;
  output [7:0] md3;
  output [7:0] md4;
  output [7:0] md5;
  input clkper, rst, sfrwe, sfroe, test_si, test_se;
  output mdubsy, test_so;
  wire   N104, N105, N106, N107, N108, N109, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N332, N333, N334, N335, N336, N337, N338, N339, N340,
         N405, N406, N407, N408, N409, N410, N411, N412, N413, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N566, N567, N568, N569, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N610,
         N674, N675, N676, N677, N678, set_div16, set_div32, N802, N892, N893,
         N894, N895, net12318, net12324, net12329, net12334, net12339,
         net12344, net12349, n408, n410, n411, n412, n413, n414, n119, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n409, n1, n2, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2;
  wire   [3:0] oper_reg;
  wire   [4:1] counter_st;
  wire   [17:1] sum1;
  wire   [17:1] sum;
  wire   [15:0] norm_reg;
  wire   [1:0] mdu_op;
  wire   [17:1] arg_a;
  wire   [16:1] arg_b;
  wire   [17:0] arg_c;
  wire   [16:1] arg_d;

  SNPS_CLOCK_GATE_HIGH_mdu_a0_0 clk_gate_arcon_s_reg ( .CLK(clkper), .EN(N104), 
        .ENCLK(net12318), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_6 clk_gate_md0_s_reg ( .CLK(clkper), .EN(N190), 
        .ENCLK(net12324), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_5 clk_gate_md1_s_reg ( .CLK(clkper), .EN(N258), 
        .ENCLK(net12329), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_4 clk_gate_md2_s_reg ( .CLK(clkper), .EN(N332), 
        .ENCLK(net12334), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_3 clk_gate_md3_s_reg ( .CLK(clkper), .EN(N405), 
        .ENCLK(net12339), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_2 clk_gate_md4_s_reg ( .CLK(clkper), .EN(N453), 
        .ENCLK(net12344), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_1 clk_gate_md5_s_reg ( .CLK(clkper), .EN(N483), 
        .ENCLK(net12349), .TE(test_se) );
  mdu_a0_DW01_add_0 add_1040 ( .A(arg_c), .B({1'b0, arg_d, n409}), .CI(1'b0), 
        .SUM({sum, SYNOPSYS_UNCONNECTED_1}), .CO() );
  mdu_a0_DW01_add_1 add_961 ( .A({arg_a, n119}), .B({1'b0, arg_b, n409}), .CI(
        1'b0), .SUM({sum1, SYNOPSYS_UNCONNECTED_2}), .CO() );
  SDFFQX1 set_div16_reg ( .D(n414), .SIN(oper_reg[3]), .SMC(test_se), .C(
        clkper), .Q(set_div16) );
  SDFFQX1 setmdef_reg ( .D(N802), .SIN(set_div32), .SMC(test_se), .C(clkper), 
        .Q(test_so) );
  SDFFQX1 set_div32_reg ( .D(n413), .SIN(set_div16), .SMC(test_se), .C(clkper), 
        .Q(set_div32) );
  SDFFQX1 counter_st_reg_0_ ( .D(N674), .SIN(arcon[7]), .SMC(test_se), .C(
        clkper), .Q(N610) );
  SDFFQX1 counter_st_reg_4_ ( .D(N678), .SIN(counter_st[3]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[4]) );
  SDFFQX1 counter_st_reg_1_ ( .D(N675), .SIN(N610), .SMC(test_se), .C(clkper), 
        .Q(counter_st[1]) );
  SDFFQX1 counter_st_reg_3_ ( .D(N677), .SIN(counter_st[2]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[3]) );
  SDFFQX1 counter_st_reg_2_ ( .D(N676), .SIN(counter_st[1]), .SMC(test_se), 
        .C(clkper), .Q(counter_st[2]) );
  SDFFQX1 oper_reg_reg_0_ ( .D(N892), .SIN(norm_reg[15]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[0]) );
  SDFFQX1 oper_reg_reg_3_ ( .D(N895), .SIN(oper_reg[2]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[3]) );
  SDFFQX1 oper_reg_reg_2_ ( .D(N894), .SIN(oper_reg[1]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[2]) );
  SDFFQX1 oper_reg_reg_1_ ( .D(N893), .SIN(oper_reg[0]), .SMC(test_se), .C(
        clkper), .Q(oper_reg[1]) );
  SDFFQX1 arcon_s_reg_7_ ( .D(n410), .SIN(arcon[6]), .SMC(test_se), .C(clkper), 
        .Q(arcon[7]) );
  SDFFQX1 md0_s_reg_7_ ( .D(N198), .SIN(md0[6]), .SMC(test_se), .C(net12324), 
        .Q(md0[7]) );
  SDFFQX1 arcon_s_reg_6_ ( .D(n408), .SIN(arcon[5]), .SMC(test_se), .C(clkper), 
        .Q(arcon[6]) );
  SDFFQX1 arcon_s_reg_5_ ( .D(n50), .SIN(arcon[4]), .SMC(test_se), .C(net12318), .Q(arcon[5]) );
  SDFFQX1 md1_s_reg_5_ ( .D(N264), .SIN(md1[4]), .SMC(test_se), .C(net12329), 
        .Q(md1[5]) );
  SDFFQX1 md0_s_reg_6_ ( .D(N197), .SIN(md0[5]), .SMC(test_se), .C(net12324), 
        .Q(md0[6]) );
  SDFFQX1 md1_s_reg_4_ ( .D(N263), .SIN(md1[3]), .SMC(test_se), .C(net12329), 
        .Q(md1[4]) );
  SDFFQX1 arcon_s_reg_4_ ( .D(N109), .SIN(arcon[3]), .SMC(test_se), .C(
        net12318), .Q(arcon[4]) );
  SDFFQX1 md0_s_reg_5_ ( .D(N196), .SIN(md0[4]), .SMC(test_se), .C(net12324), 
        .Q(md0[5]) );
  SDFFQX1 md0_s_reg_4_ ( .D(N195), .SIN(md0[3]), .SMC(test_se), .C(net12324), 
        .Q(md0[4]) );
  SDFFQX1 md1_s_reg_6_ ( .D(N265), .SIN(md1[5]), .SMC(test_se), .C(net12329), 
        .Q(md1[6]) );
  SDFFQX1 norm_reg_reg_15_ ( .D(N581), .SIN(norm_reg[14]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[15]) );
  SDFFQX1 arcon_s_reg_3_ ( .D(N108), .SIN(arcon[2]), .SMC(test_se), .C(
        net12318), .Q(arcon[3]) );
  SDFFQX1 md0_s_reg_3_ ( .D(N194), .SIN(md0[2]), .SMC(test_se), .C(net12324), 
        .Q(md0[3]) );
  SDFFQX1 norm_reg_reg_14_ ( .D(N580), .SIN(norm_reg[13]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[14]) );
  SDFFQX1 norm_reg_reg_13_ ( .D(N579), .SIN(norm_reg[12]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[13]) );
  SDFFQX1 md1_s_reg_3_ ( .D(N262), .SIN(md1[2]), .SMC(test_se), .C(net12329), 
        .Q(md1[3]) );
  SDFFQX1 md5_s_reg_6_ ( .D(N490), .SIN(md5[5]), .SMC(test_se), .C(net12349), 
        .Q(md5[6]) );
  SDFFQX1 md5_s_reg_7_ ( .D(N491), .SIN(md5[6]), .SMC(test_se), .C(net12349), 
        .Q(md5[7]) );
  SDFFQX1 md3_s_reg_6_ ( .D(N412), .SIN(md3[5]), .SMC(test_se), .C(net12339), 
        .Q(md3[6]) );
  SDFFQX1 md3_s_reg_5_ ( .D(N411), .SIN(md3[4]), .SMC(test_se), .C(net12339), 
        .Q(md3[5]) );
  SDFFQX1 norm_reg_reg_12_ ( .D(N578), .SIN(norm_reg[11]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[12]) );
  SDFFQX1 md5_s_reg_5_ ( .D(N489), .SIN(md5[4]), .SMC(test_se), .C(net12349), 
        .Q(md5[5]) );
  SDFFQX1 norm_reg_reg_10_ ( .D(N576), .SIN(norm_reg[9]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[10]) );
  SDFFQX1 norm_reg_reg_11_ ( .D(N577), .SIN(norm_reg[10]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[11]) );
  SDFFQX1 md3_s_reg_3_ ( .D(N409), .SIN(md3[2]), .SMC(test_se), .C(net12339), 
        .Q(md3[3]) );
  SDFFQX1 md3_s_reg_4_ ( .D(N410), .SIN(md3[3]), .SMC(test_se), .C(net12339), 
        .Q(md3[4]) );
  SDFFQX1 md5_s_reg_3_ ( .D(N487), .SIN(md5[2]), .SMC(test_se), .C(net12349), 
        .Q(md5[3]) );
  SDFFQX1 md5_s_reg_4_ ( .D(N488), .SIN(md5[3]), .SMC(test_se), .C(net12349), 
        .Q(md5[4]) );
  SDFFQX1 norm_reg_reg_9_ ( .D(N575), .SIN(norm_reg[8]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[9]) );
  SDFFQX1 norm_reg_reg_8_ ( .D(N574), .SIN(norm_reg[7]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[8]) );
  SDFFQX1 norm_reg_reg_7_ ( .D(N573), .SIN(norm_reg[6]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[7]) );
  SDFFQX1 norm_reg_reg_6_ ( .D(N572), .SIN(norm_reg[5]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[6]) );
  SDFFQX1 md2_s_reg_7_ ( .D(N340), .SIN(md2[6]), .SMC(test_se), .C(net12334), 
        .Q(md2[7]) );
  SDFFQX1 md4_s_reg_7_ ( .D(N461), .SIN(md4[6]), .SMC(test_se), .C(net12344), 
        .Q(md4[7]) );
  SDFFQX1 norm_reg_reg_4_ ( .D(N570), .SIN(norm_reg[3]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[4]) );
  SDFFQX1 norm_reg_reg_5_ ( .D(N571), .SIN(norm_reg[4]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[5]) );
  SDFFQX1 md2_s_reg_6_ ( .D(N339), .SIN(md2[5]), .SMC(test_se), .C(net12334), 
        .Q(md2[6]) );
  SDFFQX1 md2_s_reg_5_ ( .D(N338), .SIN(md2[4]), .SMC(test_se), .C(net12334), 
        .Q(md2[5]) );
  SDFFQX1 md4_s_reg_6_ ( .D(N460), .SIN(md4[5]), .SMC(test_se), .C(net12344), 
        .Q(md4[6]) );
  SDFFQX1 md4_s_reg_5_ ( .D(N459), .SIN(md4[4]), .SMC(test_se), .C(net12344), 
        .Q(md4[5]) );
  SDFFQX1 norm_reg_reg_3_ ( .D(N569), .SIN(norm_reg[2]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[3]) );
  SDFFQX1 md2_s_reg_4_ ( .D(N337), .SIN(md2[3]), .SMC(test_se), .C(net12334), 
        .Q(md2[4]) );
  SDFFQX1 md4_s_reg_4_ ( .D(N458), .SIN(md4[3]), .SMC(test_se), .C(net12344), 
        .Q(md4[4]) );
  SDFFQX1 norm_reg_reg_2_ ( .D(N568), .SIN(norm_reg[1]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[2]) );
  SDFFQX1 norm_reg_reg_1_ ( .D(N567), .SIN(norm_reg[0]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[1]) );
  SDFFQX1 md4_s_reg_3_ ( .D(N457), .SIN(md4[2]), .SMC(test_se), .C(net12344), 
        .Q(md4[3]) );
  SDFFQX1 md2_s_reg_3_ ( .D(N336), .SIN(md2[2]), .SMC(test_se), .C(net12334), 
        .Q(md2[3]) );
  SDFFQX1 norm_reg_reg_0_ ( .D(N566), .SIN(mdu_op[1]), .SMC(test_se), .C(
        clkper), .Q(norm_reg[0]) );
  SDFFQX1 md1_s_reg_7_ ( .D(N266), .SIN(md1[6]), .SMC(test_se), .C(net12329), 
        .Q(md1[7]) );
  SDFFQX1 md3_s_reg_7_ ( .D(N413), .SIN(md3[6]), .SMC(test_se), .C(net12339), 
        .Q(md3[7]) );
  SDFFQX1 mdu_op_reg_0_ ( .D(n411), .SIN(md5[7]), .SMC(test_se), .C(clkper), 
        .Q(mdu_op[0]) );
  SDFFQX1 mdu_op_reg_1_ ( .D(n412), .SIN(mdu_op[0]), .SMC(test_se), .C(clkper), 
        .Q(mdu_op[1]) );
  SDFFQX1 md0_s_reg_1_ ( .D(N192), .SIN(md0[0]), .SMC(test_se), .C(net12324), 
        .Q(md0[1]) );
  SDFFQX1 md1_s_reg_2_ ( .D(N261), .SIN(md1[1]), .SMC(test_se), .C(net12329), 
        .Q(md1[2]) );
  SDFFQX1 md5_s_reg_1_ ( .D(N485), .SIN(md5[0]), .SMC(test_se), .C(net12349), 
        .Q(md5[1]) );
  SDFFQX1 arcon_s_reg_1_ ( .D(N106), .SIN(arcon[0]), .SMC(test_se), .C(
        net12318), .Q(arcon[1]) );
  SDFFQX1 md2_s_reg_2_ ( .D(N335), .SIN(md2[1]), .SMC(test_se), .C(net12334), 
        .Q(md2[2]) );
  SDFFQX1 md4_s_reg_1_ ( .D(N455), .SIN(md4[0]), .SMC(test_se), .C(net12344), 
        .Q(md4[1]) );
  SDFFQX1 md2_s_reg_1_ ( .D(N334), .SIN(md2[0]), .SMC(test_se), .C(net12334), 
        .Q(md2[1]) );
  SDFFQX1 md3_s_reg_1_ ( .D(N407), .SIN(md3[0]), .SMC(test_se), .C(net12339), 
        .Q(md3[1]) );
  SDFFQX1 md1_s_reg_1_ ( .D(N260), .SIN(md1[0]), .SMC(test_se), .C(net12329), 
        .Q(md1[1]) );
  SDFFQX1 md0_s_reg_2_ ( .D(N193), .SIN(md0[1]), .SMC(test_se), .C(net12324), 
        .Q(md0[2]) );
  SDFFQX1 md0_s_reg_0_ ( .D(N191), .SIN(counter_st[4]), .SMC(test_se), .C(
        net12324), .Q(md0[0]) );
  SDFFQX1 arcon_s_reg_0_ ( .D(N105), .SIN(test_si), .SMC(test_se), .C(net12318), .Q(arcon[0]) );
  SDFFQX1 arcon_s_reg_2_ ( .D(N107), .SIN(arcon[1]), .SMC(test_se), .C(
        net12318), .Q(arcon[2]) );
  SDFFQX1 md1_s_reg_0_ ( .D(N259), .SIN(md0[7]), .SMC(test_se), .C(net12329), 
        .Q(md1[0]) );
  SDFFQX1 md2_s_reg_0_ ( .D(N333), .SIN(md1[7]), .SMC(test_se), .C(net12334), 
        .Q(md2[0]) );
  SDFFQX1 md3_s_reg_2_ ( .D(N408), .SIN(md3[1]), .SMC(test_se), .C(net12339), 
        .Q(md3[2]) );
  SDFFQX1 md5_s_reg_2_ ( .D(N486), .SIN(md5[1]), .SMC(test_se), .C(net12349), 
        .Q(md5[2]) );
  SDFFQX1 md5_s_reg_0_ ( .D(N484), .SIN(md4[7]), .SMC(test_se), .C(net12349), 
        .Q(md5[0]) );
  SDFFQX1 md4_s_reg_2_ ( .D(N456), .SIN(md4[1]), .SMC(test_se), .C(net12344), 
        .Q(md4[2]) );
  SDFFQX1 md4_s_reg_0_ ( .D(N454), .SIN(md3[7]), .SMC(test_se), .C(net12344), 
        .Q(md4[0]) );
  SDFFQX1 md3_s_reg_0_ ( .D(N406), .SIN(md2[7]), .SMC(test_se), .C(net12339), 
        .Q(md3[0]) );
  NAND2X1 U5 ( .A(n275), .B(n54), .Y(n1) );
  NAND2X1 U6 ( .A(n244), .B(n275), .Y(n2) );
  INVX1 U7 ( .A(n298), .Y(n5) );
  INVX1 U8 ( .A(n55), .Y(n6) );
  BUFX3 U9 ( .A(n300), .Y(n7) );
  NAND2X1 U10 ( .A(n20), .B(n259), .Y(n8) );
  NAND2X1 U11 ( .A(n112), .B(arg_c[0]), .Y(n9) );
  INVX1 U12 ( .A(n340), .Y(n10) );
  BUFX3 U13 ( .A(n257), .Y(n11) );
  BUFX3 U14 ( .A(n189), .Y(n12) );
  BUFX3 U15 ( .A(n295), .Y(n13) );
  INVX1 U16 ( .A(n97), .Y(n14) );
  INVX1 U17 ( .A(n23), .Y(n15) );
  BUFX3 U18 ( .A(n256), .Y(n16) );
  NAND2X1 U19 ( .A(sum1[17]), .B(arg_c[0]), .Y(n17) );
  BUFX3 U20 ( .A(n195), .Y(n18) );
  INVX1 U21 ( .A(n67), .Y(n19) );
  INVX1 U22 ( .A(n96), .Y(n20) );
  INVX1 U23 ( .A(n51), .Y(n21) );
  INVX1 U24 ( .A(n371), .Y(n22) );
  BUFX3 U25 ( .A(n304), .Y(n23) );
  INVX1 U26 ( .A(n119), .Y(n24) );
  INVX1 U27 ( .A(sum[17]), .Y(n25) );
  INVX1 U28 ( .A(n25), .Y(n26) );
  INVX1 U29 ( .A(n25), .Y(n27) );
  INVX1 U30 ( .A(n168), .Y(n51) );
  NAND2X1 U31 ( .A(n315), .B(n161), .Y(N405) );
  NAND2X1 U32 ( .A(n315), .B(n162), .Y(N332) );
  INVX1 U33 ( .A(n332), .Y(n54) );
  INVX1 U34 ( .A(n371), .Y(n66) );
  INVX1 U35 ( .A(n33), .Y(n31) );
  INVX1 U36 ( .A(n409), .Y(n36) );
  INVX1 U37 ( .A(n33), .Y(n32) );
  INVX1 U38 ( .A(n409), .Y(n35) );
  NAND2X1 U39 ( .A(n56), .B(n275), .Y(n166) );
  NAND2X1 U40 ( .A(n52), .B(n275), .Y(n168) );
  NAND2X1 U41 ( .A(n244), .B(n275), .Y(n161) );
  NAND2X1 U42 ( .A(n275), .B(n54), .Y(n162) );
  NAND2X1 U43 ( .A(n275), .B(n53), .Y(n239) );
  NAND2X1 U44 ( .A(n165), .B(n275), .Y(n357) );
  OR2X1 U45 ( .A(n242), .B(n48), .Y(n159) );
  NAND2X1 U46 ( .A(n47), .B(n242), .Y(n278) );
  NAND3X1 U47 ( .A(n274), .B(n47), .C(n159), .Y(N453) );
  NAND3X1 U48 ( .A(n274), .B(n47), .C(n6), .Y(N483) );
  NAND3X1 U49 ( .A(n276), .B(n28), .C(n37), .Y(n332) );
  INVX1 U50 ( .A(n229), .Y(n52) );
  INVX1 U51 ( .A(n354), .Y(n53) );
  INVX1 U52 ( .A(n246), .Y(n56) );
  OR2X1 U53 ( .A(n334), .B(n335), .Y(n292) );
  NAND2X1 U54 ( .A(n67), .B(n336), .Y(n371) );
  INVX1 U55 ( .A(n302), .Y(n67) );
  NOR32XL U56 ( .B(n336), .C(n337), .A(n334), .Y(n315) );
  INVX1 U57 ( .A(rst), .Y(n47) );
  NAND2X1 U58 ( .A(n20), .B(n259), .Y(n255) );
  INVX1 U59 ( .A(n409), .Y(n34) );
  INVX1 U60 ( .A(n427), .Y(n33) );
  INVX1 U61 ( .A(n262), .Y(n96) );
  NAND42X1 U62 ( .C(n245), .D(sfraddr[1]), .A(n37), .B(n289), .Y(n242) );
  NOR2X1 U63 ( .A(n28), .B(n57), .Y(n289) );
  OAI21X1 U64 ( .B(n164), .C(n354), .A(n47), .Y(n158) );
  OAI21X1 U65 ( .B(n164), .C(n246), .A(n47), .Y(n230) );
  OAI21BX1 U66 ( .C(n244), .B(n164), .A(n49), .Y(n291) );
  OAI21BX1 U67 ( .C(n165), .B(n164), .A(n49), .Y(n359) );
  OAI21X1 U68 ( .B(n164), .C(n332), .A(n47), .Y(n317) );
  NOR2X1 U69 ( .A(n57), .B(n48), .Y(n275) );
  OAI21AX1 U70 ( .B(n164), .C(n229), .A(n230), .Y(n198) );
  NAND2X1 U71 ( .A(n407), .B(n82), .Y(n380) );
  NAND4X1 U72 ( .A(n379), .B(n380), .C(n168), .D(n47), .Y(N104) );
  NAND2X1 U73 ( .A(n356), .B(n357), .Y(N190) );
  NAND2X1 U74 ( .A(n356), .B(n239), .Y(N258) );
  NOR21XL U75 ( .B(sfraddr[1]), .A(n245), .Y(n276) );
  NAND3X1 U76 ( .A(n276), .B(n38), .C(sfraddr[2]), .Y(n246) );
  NOR4XL U77 ( .A(n28), .B(n245), .C(n37), .D(sfraddr[1]), .Y(n244) );
  NAND3X1 U78 ( .A(n37), .B(n276), .C(sfraddr[2]), .Y(n229) );
  NAND3X1 U79 ( .A(n38), .B(n28), .C(n276), .Y(n354) );
  OAI31XL U80 ( .A(n38), .B(sfraddr[1]), .C(n245), .D(n246), .Y(n243) );
  INVX1 U81 ( .A(n38), .Y(n37) );
  NOR4XL U82 ( .A(n38), .B(n245), .C(sfraddr[1]), .D(sfraddr[2]), .Y(n165) );
  INVX1 U83 ( .A(sfraddr[2]), .Y(n28) );
  OAI31XL U84 ( .A(n265), .B(n78), .C(n261), .D(n274), .Y(n334) );
  NAND3X1 U85 ( .A(n78), .B(n261), .C(n75), .Y(n274) );
  NOR2X1 U86 ( .A(n378), .B(n68), .Y(n302) );
  NAND3X1 U87 ( .A(n261), .B(n265), .C(n78), .Y(n296) );
  NAND3X1 U88 ( .A(n77), .B(n265), .C(n78), .Y(n378) );
  INVX1 U89 ( .A(n261), .Y(n77) );
  NOR2X1 U90 ( .A(n377), .B(n68), .Y(n335) );
  INVX1 U91 ( .A(n374), .Y(n74) );
  INVX1 U92 ( .A(n265), .Y(n75) );
  NAND3X1 U93 ( .A(n78), .B(n77), .C(n75), .Y(n336) );
  INVX1 U94 ( .A(n298), .Y(n69) );
  NOR43XL U95 ( .B(n296), .C(n377), .D(n378), .A(n48), .Y(n337) );
  NOR3XL U96 ( .A(n78), .B(rst), .C(n265), .Y(n259) );
  INVX1 U97 ( .A(n49), .Y(n48) );
  NOR2X1 U98 ( .A(n112), .B(n26), .Y(n262) );
  NAND2X1 U99 ( .A(n26), .B(n259), .Y(n257) );
  NAND2X1 U100 ( .A(n112), .B(arg_c[0]), .Y(n191) );
  NAND2X1 U101 ( .A(n259), .B(n260), .Y(n256) );
  INVX1 U102 ( .A(n196), .Y(n427) );
  INVX1 U103 ( .A(n260), .Y(n97) );
  INVX1 U104 ( .A(n409), .Y(n428) );
  INVX1 U105 ( .A(n196), .Y(n119) );
  INVX1 U106 ( .A(sfrwe), .Y(n57) );
  NAND21X1 U107 ( .B(n406), .A(n407), .Y(n379) );
  AOI21X1 U108 ( .B(sfrwe), .C(n52), .A(n48), .Y(n407) );
  NOR2X1 U109 ( .A(n48), .B(sfrwe), .Y(n164) );
  OAI31XL U110 ( .A(n56), .B(n52), .C(n165), .D(sfrwe), .Y(n241) );
  AOI31X1 U111 ( .A(n2), .B(n1), .C(n236), .D(n237), .Y(N802) );
  AOI21AX1 U112 ( .B(n238), .C(n49), .A(n239), .Y(n236) );
  OAI2B11X1 U113 ( .D(sfroe), .C(n240), .A(n241), .B(n242), .Y(n238) );
  NOR4XL U114 ( .A(n243), .B(n244), .C(n53), .D(n54), .Y(n240) );
  NAND41X1 U115 ( .D(sfraddr[4]), .A(sfraddr[5]), .B(sfraddr[3]), .C(
        sfraddr[6]), .Y(n245) );
  INVX1 U116 ( .A(sfraddr[0]), .Y(n38) );
  INVX1 U117 ( .A(sfrdatai[4]), .Y(n43) );
  INVX1 U118 ( .A(sfrdatai[7]), .Y(n46) );
  INVX1 U119 ( .A(sfrdatai[6]), .Y(n45) );
  INVX1 U120 ( .A(sfrdatai[0]), .Y(n39) );
  INVX1 U121 ( .A(sfrdatai[1]), .Y(n40) );
  INVX1 U122 ( .A(sfrdatai[2]), .Y(n41) );
  INVX1 U123 ( .A(sfrdatai[3]), .Y(n42) );
  INVX1 U124 ( .A(sfrdatai[5]), .Y(n44) );
  NOR32XL U125 ( .B(n202), .C(n399), .A(n79), .Y(n401) );
  NAND3X1 U126 ( .A(n210), .B(n181), .C(n401), .Y(n261) );
  NOR42XL U127 ( .C(n405), .D(n406), .A(n85), .B(n237), .Y(n399) );
  NOR2X1 U128 ( .A(n178), .B(n84), .Y(n405) );
  INVX1 U129 ( .A(n183), .Y(n84) );
  OAI21X1 U130 ( .B(n261), .C(n376), .A(n75), .Y(n374) );
  NAND2X1 U131 ( .A(n404), .B(n401), .Y(n265) );
  INVX1 U132 ( .A(n376), .Y(n78) );
  NOR2X1 U133 ( .A(n396), .B(n378), .Y(n29) );
  NOR2X1 U134 ( .A(n396), .B(n377), .Y(n293) );
  NAND3X1 U135 ( .A(n265), .B(n376), .C(n77), .Y(n377) );
  INVX1 U136 ( .A(n23), .Y(n70) );
  NOR2X1 U137 ( .A(n396), .B(n378), .Y(n30) );
  NOR2X1 U138 ( .A(n396), .B(n378), .Y(n298) );
  INVX1 U139 ( .A(n340), .Y(n65) );
  NAND2X1 U140 ( .A(n208), .B(n210), .Y(n254) );
  INVX1 U141 ( .A(n182), .Y(n79) );
  NOR32XL U142 ( .B(n337), .C(n13), .A(n74), .Y(n356) );
  INVX1 U143 ( .A(n396), .Y(n68) );
  INVX1 U144 ( .A(n404), .Y(n82) );
  INVX1 U145 ( .A(rst), .Y(n49) );
  INVX1 U146 ( .A(n207), .Y(n64) );
  INVX1 U147 ( .A(n215), .Y(n83) );
  INVX1 U148 ( .A(n210), .Y(n80) );
  OAI21X1 U149 ( .B(n431), .C(n430), .A(n409), .Y(n196) );
  OAI22X1 U150 ( .A(n17), .B(n116), .C(n191), .D(n117), .Y(arg_c[17]) );
  NOR2X1 U151 ( .A(sum[17]), .B(sum1[17]), .Y(n260) );
  INVX1 U152 ( .A(sum[15]), .Y(n99) );
  INVX1 U153 ( .A(sum[16]), .Y(n98) );
  NAND2X1 U154 ( .A(sum1[17]), .B(arg_c[0]), .Y(n190) );
  INVX1 U155 ( .A(sum1[17]), .Y(n112) );
  NAND2X1 U156 ( .A(n430), .B(n431), .Y(n409) );
  OAI222XL U157 ( .A(n422), .B(n255), .C(n423), .D(n256), .E(n257), .F(n111), 
        .Y(N568) );
  OAI222XL U158 ( .A(n419), .B(n8), .C(n420), .D(n256), .E(n257), .F(n110), 
        .Y(N569) );
  OAI222XL U159 ( .A(n155), .B(n255), .C(n157), .D(n256), .E(n257), .F(n108), 
        .Y(N571) );
  OAI222XL U160 ( .A(n416), .B(n8), .C(n418), .D(n256), .E(n257), .F(n109), 
        .Y(N570) );
  OAI222XL U161 ( .A(n149), .B(n255), .C(n150), .D(n256), .E(n257), .F(n107), 
        .Y(N572) );
  OAI222XL U162 ( .A(n147), .B(n8), .C(n151), .D(n256), .E(n257), .F(n106), 
        .Y(N573) );
  OAI222XL U163 ( .A(n143), .B(n255), .C(n145), .D(n256), .E(n257), .F(n105), 
        .Y(N574) );
  OAI222XL U164 ( .A(n141), .B(n8), .C(n142), .D(n256), .E(n257), .F(n104), 
        .Y(N575) );
  OAI222XL U165 ( .A(n137), .B(n255), .C(n138), .D(n256), .E(n257), .F(n102), 
        .Y(N577) );
  OAI222XL U166 ( .A(n139), .B(n8), .C(n140), .D(n16), .E(n11), .F(n103), .Y(
        N576) );
  OAI222XL U167 ( .A(n130), .B(n255), .C(n133), .D(n16), .E(n11), .F(n101), 
        .Y(N578) );
  OAI222XL U168 ( .A(n129), .B(n8), .C(n134), .D(n16), .E(n11), .F(n100), .Y(
        N579) );
  OAI222XL U169 ( .A(n126), .B(n255), .C(n127), .D(n16), .E(n11), .F(n99), .Y(
        N580) );
  OAI222XL U170 ( .A(n120), .B(n8), .C(n122), .D(n16), .E(n11), .F(n98), .Y(
        N581) );
  OAI22X1 U171 ( .A(n40), .B(n159), .C(n284), .D(n278), .Y(N455) );
  AOI222XL U172 ( .A(sum[2]), .B(n26), .C(n14), .D(n285), .E(n262), .F(sum1[1]), .Y(n284) );
  OAI22X1 U173 ( .A(n193), .B(n426), .C(n429), .D(n424), .Y(n285) );
  OAI22X1 U174 ( .A(n39), .B(n159), .C(n286), .D(n278), .Y(N454) );
  AOI22X1 U175 ( .A(n287), .B(n288), .C(sum[1]), .D(n26), .Y(n286) );
  OAI22X1 U176 ( .A(n193), .B(n125), .C(n429), .D(n115), .Y(n288) );
  NAND2X1 U177 ( .A(n96), .B(n97), .Y(n287) );
  INVX1 U178 ( .A(n193), .Y(n429) );
  INVX1 U179 ( .A(sum[14]), .Y(n100) );
  INVX1 U180 ( .A(sum[12]), .Y(n102) );
  INVX1 U181 ( .A(sum[13]), .Y(n101) );
  INVX1 U182 ( .A(sum[11]), .Y(n103) );
  INVX1 U183 ( .A(sum[10]), .Y(n104) );
  INVX1 U184 ( .A(sum[9]), .Y(n105) );
  INVX1 U185 ( .A(sum[8]), .Y(n106) );
  INVX1 U186 ( .A(sum[6]), .Y(n108) );
  INVX1 U187 ( .A(sum[7]), .Y(n107) );
  INVX1 U188 ( .A(sum[5]), .Y(n109) );
  INVX1 U189 ( .A(sum[3]), .Y(n111) );
  INVX1 U190 ( .A(sum[4]), .Y(n110) );
  INVX1 U191 ( .A(sum1[2]), .Y(n422) );
  INVX1 U192 ( .A(sum1[3]), .Y(n419) );
  INVX1 U193 ( .A(sum1[4]), .Y(n416) );
  INVX1 U194 ( .A(sum1[5]), .Y(n155) );
  INVX1 U195 ( .A(sum1[6]), .Y(n149) );
  INVX1 U196 ( .A(sum1[7]), .Y(n147) );
  INVX1 U197 ( .A(sum1[8]), .Y(n143) );
  INVX1 U198 ( .A(sum1[9]), .Y(n141) );
  INVX1 U199 ( .A(sum1[10]), .Y(n139) );
  INVX1 U200 ( .A(sum1[11]), .Y(n137) );
  INVX1 U201 ( .A(sum1[12]), .Y(n130) );
  INVX1 U202 ( .A(sum1[13]), .Y(n129) );
  INVX1 U203 ( .A(sum1[14]), .Y(n126) );
  INVX1 U204 ( .A(sum1[15]), .Y(n120) );
  INVX1 U205 ( .A(sum[2]), .Y(n113) );
  INVX1 U206 ( .A(sum1[16]), .Y(n116) );
  OAI222XL U207 ( .A(n379), .B(n391), .C(n250), .D(n380), .E(n168), .F(n41), 
        .Y(N107) );
  OAI222XL U208 ( .A(n168), .B(n39), .C(n252), .D(n380), .E(n62), .F(n379), 
        .Y(N105) );
  OAI222XL U209 ( .A(n379), .B(n63), .C(n251), .D(n380), .E(n168), .F(n40), 
        .Y(N106) );
  INVX1 U210 ( .A(n394), .Y(n63) );
  OAI222XL U211 ( .A(n379), .B(n389), .C(n249), .D(n380), .E(n21), .F(n42), 
        .Y(N108) );
  OAI222XL U212 ( .A(n379), .B(n61), .C(n247), .D(n380), .E(n168), .F(n43), 
        .Y(N109) );
  INVX1 U213 ( .A(n381), .Y(n61) );
  OAI211X1 U214 ( .C(n197), .D(n198), .A(n166), .B(n168), .Y(N895) );
  AOI211X1 U215 ( .C(n79), .D(n199), .A(n200), .B(n201), .Y(n197) );
  OAI32X1 U216 ( .A(n202), .B(n426), .C(n203), .D(n409), .E(n204), .Y(n201) );
  OAI222XL U217 ( .A(n205), .B(n206), .C(n207), .D(n208), .E(n209), .F(n210), 
        .Y(n200) );
  OAI211X1 U218 ( .C(n160), .D(n58), .A(n161), .B(n162), .Y(n413) );
  NOR2X1 U219 ( .A(n163), .B(n164), .Y(n160) );
  NOR4XL U220 ( .A(rst), .B(n52), .C(n165), .D(n56), .Y(n163) );
  AOI31X1 U221 ( .A(n218), .B(n219), .C(n220), .D(n198), .Y(N893) );
  AOI22BXL U222 ( .B(n206), .A(n205), .D(n208), .C(n64), .Y(n219) );
  NOR32XL U223 ( .B(n221), .C(n210), .A(n222), .Y(n220) );
  AOI21X1 U224 ( .B(n224), .C(n214), .A(n225), .Y(n218) );
  INVX1 U225 ( .A(sum1[1]), .Y(n425) );
  NAND2X1 U226 ( .A(n193), .B(n194), .Y(arg_c[0]) );
  INVX1 U227 ( .A(sum[1]), .Y(n114) );
  NAND2X1 U228 ( .A(n234), .B(n402), .Y(n183) );
  AOI21BBXL U229 ( .B(n125), .C(n296), .A(n293), .Y(n304) );
  NAND42X1 U230 ( .C(n254), .D(n224), .A(n399), .B(n202), .Y(n376) );
  AOI211X1 U231 ( .C(n125), .D(n76), .A(n74), .B(n335), .Y(n340) );
  INVX1 U232 ( .A(n296), .Y(n76) );
  OAI31XL U233 ( .A(n397), .B(n29), .C(n293), .D(n385), .Y(n382) );
  NOR3XL U234 ( .A(n125), .B(n75), .C(n77), .Y(n397) );
  AND2X1 U235 ( .A(n400), .B(n402), .Y(n178) );
  NOR2X1 U236 ( .A(n81), .B(n86), .Y(n403) );
  OAI31XL U237 ( .A(n81), .B(n88), .C(n87), .D(mdubsy), .Y(n237) );
  NAND2X1 U238 ( .A(n398), .B(n400), .Y(mdubsy) );
  NAND2X1 U239 ( .A(n403), .B(n402), .Y(n406) );
  NOR2X1 U240 ( .A(n251), .B(n248), .Y(N675) );
  NOR2X1 U241 ( .A(n249), .B(n248), .Y(N677) );
  NOR2X1 U242 ( .A(n250), .B(n248), .Y(N676) );
  NOR2X1 U243 ( .A(n247), .B(n248), .Y(N678) );
  NOR2X1 U244 ( .A(n252), .B(n248), .Y(N674) );
  INVX1 U245 ( .A(n204), .Y(n85) );
  NAND21X1 U246 ( .B(n336), .A(n221), .Y(n295) );
  AOI21X1 U247 ( .B(n234), .C(n233), .A(n224), .Y(n404) );
  NAND2X1 U248 ( .A(n233), .B(n403), .Y(n182) );
  NAND2X1 U249 ( .A(n398), .B(n403), .Y(n210) );
  NAND2X1 U250 ( .A(n398), .B(n234), .Y(n202) );
  NAND2X1 U251 ( .A(n402), .B(n86), .Y(n181) );
  NAND2X1 U252 ( .A(n233), .B(n400), .Y(n208) );
  NAND42X1 U253 ( .C(n254), .D(n82), .A(n206), .B(n182), .Y(n385) );
  NAND2X1 U254 ( .A(n386), .B(n71), .Y(n396) );
  INVX1 U255 ( .A(n393), .Y(n73) );
  NAND21X1 U256 ( .B(n202), .A(n203), .Y(n215) );
  NAND2X1 U257 ( .A(n223), .B(n71), .Y(n207) );
  AOI31X1 U258 ( .A(n217), .B(n72), .C(n62), .D(n68), .Y(n214) );
  NAND2X1 U259 ( .A(n393), .B(n62), .Y(n387) );
  OAI31XL U260 ( .A(n253), .B(n254), .C(n82), .D(n47), .Y(n248) );
  NAND3X1 U261 ( .A(n206), .B(n182), .C(n202), .Y(n253) );
  OAI21X1 U262 ( .B(n231), .C(n72), .A(n387), .Y(n391) );
  NAND4X1 U263 ( .A(n448), .B(n135), .C(n136), .D(n426), .Y(n185) );
  NAND4X1 U264 ( .A(n153), .B(n146), .C(n438), .D(n447), .Y(n186) );
  NOR21XL U265 ( .B(norm_reg[15]), .A(n24), .Y(arg_a[17]) );
  OAI22X1 U266 ( .A(md4[1]), .B(n36), .C(n441), .D(n195), .Y(arg_b[2]) );
  OAI22X1 U267 ( .A(n423), .B(n196), .C(n31), .D(n440), .Y(arg_a[2]) );
  OAI22X1 U268 ( .A(md4[2]), .B(n36), .C(n433), .D(n195), .Y(arg_b[3]) );
  OAI22X1 U269 ( .A(n420), .B(n196), .C(n31), .D(n439), .Y(arg_a[3]) );
  OAI22X1 U270 ( .A(md4[3]), .B(n36), .C(n417), .D(n195), .Y(arg_b[4]) );
  OAI22X1 U271 ( .A(n418), .B(n196), .C(n31), .D(n421), .Y(arg_a[4]) );
  OAI22X1 U272 ( .A(md4[4]), .B(n36), .C(n156), .D(n195), .Y(arg_b[5]) );
  OAI22X1 U273 ( .A(n157), .B(n196), .C(n31), .D(n415), .Y(arg_a[5]) );
  OAI22X1 U274 ( .A(md4[5]), .B(n36), .C(n154), .D(n195), .Y(arg_b[6]) );
  OAI22X1 U275 ( .A(n150), .B(n196), .C(n32), .D(n152), .Y(arg_a[6]) );
  OAI22X1 U276 ( .A(md4[2]), .B(n34), .C(n189), .D(n433), .Y(arg_d[3]) );
  OAI222XL U277 ( .A(n17), .B(n422), .C(n191), .D(n423), .E(n119), .F(n416), 
        .Y(arg_c[3]) );
  OAI22X1 U278 ( .A(md4[6]), .B(n36), .C(n148), .D(n195), .Y(arg_b[7]) );
  OAI22X1 U279 ( .A(n151), .B(n196), .C(n32), .D(n153), .Y(arg_a[7]) );
  OAI22X1 U280 ( .A(md4[3]), .B(n34), .C(n189), .D(n417), .Y(arg_d[4]) );
  OAI222XL U281 ( .A(n190), .B(n419), .C(n9), .D(n420), .E(n119), .F(n155), 
        .Y(arg_c[4]) );
  OAI22X1 U282 ( .A(md4[7]), .B(n36), .C(n144), .D(n195), .Y(arg_b[8]) );
  OAI22X1 U283 ( .A(n145), .B(n196), .C(n427), .D(n146), .Y(arg_a[8]) );
  OAI22X1 U284 ( .A(md4[4]), .B(n34), .C(n189), .D(n156), .Y(arg_d[5]) );
  OAI222XL U285 ( .A(n17), .B(n416), .C(n191), .D(n418), .E(n119), .F(n149), 
        .Y(arg_c[5]) );
  OAI22X1 U286 ( .A(md5[0]), .B(n35), .C(n442), .D(n195), .Y(arg_b[9]) );
  OAI22X1 U287 ( .A(n142), .B(n196), .C(n427), .D(n438), .Y(arg_a[9]) );
  OAI22X1 U288 ( .A(md4[5]), .B(n34), .C(n189), .D(n154), .Y(arg_d[6]) );
  OAI222XL U289 ( .A(n190), .B(n155), .C(n9), .D(n157), .E(n119), .F(n147), 
        .Y(arg_c[6]) );
  OAI22X1 U290 ( .A(md5[1]), .B(n34), .C(n449), .D(n18), .Y(arg_b[10]) );
  OAI22X1 U291 ( .A(n140), .B(n24), .C(n31), .D(n447), .Y(arg_a[10]) );
  OAI22X1 U292 ( .A(md4[6]), .B(n35), .C(n189), .D(n148), .Y(arg_d[7]) );
  OAI222XL U293 ( .A(n17), .B(n149), .C(n191), .D(n150), .E(n119), .F(n143), 
        .Y(arg_c[7]) );
  OAI22X1 U294 ( .A(md5[2]), .B(n428), .C(n444), .D(n18), .Y(arg_b[11]) );
  OAI22X1 U295 ( .A(n138), .B(n24), .C(n31), .D(n448), .Y(arg_a[11]) );
  OAI22X1 U296 ( .A(md4[7]), .B(n34), .C(n189), .D(n144), .Y(arg_d[8]) );
  OAI222XL U297 ( .A(n190), .B(n147), .C(n9), .D(n151), .E(n119), .F(n141), 
        .Y(arg_c[8]) );
  OAI22X1 U298 ( .A(md5[3]), .B(n428), .C(n131), .D(n18), .Y(arg_b[12]) );
  OAI22X1 U299 ( .A(n133), .B(n24), .C(n31), .D(n135), .Y(arg_a[12]) );
  OAI22X1 U300 ( .A(md5[0]), .B(n35), .C(n189), .D(n442), .Y(arg_d[9]) );
  OAI222XL U301 ( .A(n17), .B(n143), .C(n191), .D(n145), .E(n427), .F(n139), 
        .Y(arg_c[9]) );
  OAI22X1 U302 ( .A(md5[4]), .B(n428), .C(n132), .D(n18), .Y(arg_b[13]) );
  OAI22X1 U303 ( .A(n134), .B(n24), .C(n31), .D(n136), .Y(arg_a[13]) );
  OAI22X1 U304 ( .A(md5[1]), .B(n35), .C(n12), .D(n449), .Y(arg_d[10]) );
  OAI222XL U305 ( .A(n190), .B(n141), .C(n9), .D(n142), .E(n427), .F(n137), 
        .Y(arg_c[10]) );
  ENOX1 U306 ( .A(n127), .B(n24), .C(n24), .D(md3[5]), .Y(arg_a[14]) );
  OAI22X1 U307 ( .A(md5[5]), .B(n428), .C(n128), .D(n18), .Y(arg_b[14]) );
  OAI22X1 U308 ( .A(md5[2]), .B(n35), .C(n12), .D(n444), .Y(arg_d[11]) );
  OAI222XL U309 ( .A(n17), .B(n139), .C(n191), .D(n140), .E(n427), .F(n130), 
        .Y(arg_c[11]) );
  OAI22X1 U310 ( .A(md5[6]), .B(n36), .C(n121), .D(n18), .Y(arg_b[15]) );
  OAI22X1 U311 ( .A(n122), .B(n24), .C(n31), .D(n125), .Y(arg_a[15]) );
  OAI22X1 U312 ( .A(md5[3]), .B(n35), .C(n12), .D(n131), .Y(arg_d[12]) );
  OAI222XL U313 ( .A(n190), .B(n137), .C(n9), .D(n138), .E(n427), .F(n129), 
        .Y(arg_c[12]) );
  OAI22X1 U314 ( .A(md5[4]), .B(n35), .C(n12), .D(n132), .Y(arg_d[13]) );
  OAI222XL U315 ( .A(n17), .B(n130), .C(n191), .D(n133), .E(n427), .F(n126), 
        .Y(arg_c[13]) );
  OAI22X1 U316 ( .A(md5[5]), .B(n35), .C(n12), .D(n128), .Y(arg_d[14]) );
  OAI222XL U317 ( .A(n190), .B(n129), .C(n9), .D(n134), .E(n427), .F(n120), 
        .Y(arg_c[14]) );
  OAI22X1 U318 ( .A(md5[6]), .B(n35), .C(n12), .D(n121), .Y(arg_d[15]) );
  OAI222XL U319 ( .A(n17), .B(n126), .C(n191), .D(n127), .E(n32), .F(n116), 
        .Y(arg_c[15]) );
  OAI22X1 U320 ( .A(md4[0]), .B(n36), .C(n432), .D(n195), .Y(arg_b[1]) );
  OAI21X1 U321 ( .B(n32), .C(n443), .A(n192), .Y(arg_a[1]) );
  OAI22X1 U322 ( .A(md5[7]), .B(n36), .C(n124), .D(n18), .Y(arg_b[16]) );
  OAI22X1 U323 ( .A(n117), .B(n24), .C(n31), .D(n426), .Y(arg_a[16]) );
  OAI22X1 U324 ( .A(md5[7]), .B(n35), .C(n12), .D(n124), .Y(arg_d[16]) );
  OAI222XL U325 ( .A(n190), .B(n120), .C(n9), .D(n122), .E(n32), .F(n112), .Y(
        arg_c[16]) );
  NAND2X1 U326 ( .A(md0[0]), .B(n34), .Y(n195) );
  NAND2X1 U327 ( .A(mdu_op[1]), .B(n430), .Y(n193) );
  OAI22X1 U328 ( .A(md4[1]), .B(n34), .C(n189), .D(n441), .Y(arg_d[2]) );
  OAI222XL U329 ( .A(n190), .B(n425), .C(sum1[17]), .D(n192), .E(n119), .F(
        n419), .Y(arg_c[2]) );
  OAI22X1 U330 ( .A(n44), .B(n161), .C(n301), .D(n291), .Y(N411) );
  AOI221XL U331 ( .A(n302), .B(md3[7]), .C(n30), .D(md3[6]), .E(n303), .Y(n301) );
  OAI222XL U332 ( .A(n300), .B(n135), .C(n99), .D(n295), .E(n304), .F(n136), 
        .Y(n303) );
  OAI222XL U333 ( .A(n425), .B(n255), .C(n258), .D(n16), .E(n11), .F(n113), 
        .Y(N567) );
  AOI22X1 U334 ( .A(n77), .B(md3[7]), .C(md1[7]), .D(n261), .Y(n258) );
  AOI22AXL U335 ( .A(n429), .B(md3[7]), .D(n194), .C(md1[7]), .Y(n192) );
  OAI22X1 U336 ( .A(n39), .B(n357), .C(n375), .D(n359), .Y(N191) );
  AOI222XL U337 ( .A(n30), .B(md0[1]), .C(md0[2]), .D(n371), .E(n74), .F(n27), 
        .Y(n375) );
  OAI22X1 U338 ( .A(n166), .B(n40), .C(n272), .D(n230), .Y(N485) );
  AOI222XL U339 ( .A(sum[10]), .B(n26), .C(n260), .D(norm_reg[7]), .E(n262), 
        .F(sum1[9]), .Y(n272) );
  OAI22X1 U340 ( .A(n166), .B(n41), .C(n271), .D(n230), .Y(N486) );
  AOI222XL U341 ( .A(sum[11]), .B(n27), .C(n260), .D(norm_reg[8]), .E(n262), 
        .F(sum1[10]), .Y(n271) );
  OAI22X1 U342 ( .A(n166), .B(n39), .C(n273), .D(n230), .Y(N484) );
  AOI222XL U343 ( .A(sum[9]), .B(n26), .C(n260), .D(norm_reg[6]), .E(n262), 
        .F(sum1[8]), .Y(n273) );
  OAI22X1 U344 ( .A(n41), .B(n159), .C(n283), .D(n278), .Y(N456) );
  AOI222XL U345 ( .A(sum[3]), .B(n27), .C(n14), .D(norm_reg[0]), .E(n20), .F(
        sum1[2]), .Y(n283) );
  OAI22X1 U346 ( .A(n42), .B(n159), .C(n282), .D(n278), .Y(N457) );
  AOI222XL U347 ( .A(sum[4]), .B(n26), .C(n14), .D(norm_reg[1]), .E(n20), .F(
        sum1[3]), .Y(n282) );
  OAI22X1 U348 ( .A(n43), .B(n159), .C(n281), .D(n278), .Y(N458) );
  AOI222XL U349 ( .A(sum[5]), .B(n27), .C(n14), .D(norm_reg[2]), .E(n20), .F(
        sum1[4]), .Y(n281) );
  OAI22X1 U350 ( .A(n44), .B(n159), .C(n280), .D(n278), .Y(N459) );
  AOI222XL U351 ( .A(sum[6]), .B(n26), .C(n14), .D(norm_reg[3]), .E(n20), .F(
        sum1[5]), .Y(n280) );
  OAI22X1 U352 ( .A(n45), .B(n159), .C(n279), .D(n278), .Y(N460) );
  AOI222XL U353 ( .A(sum[7]), .B(n27), .C(n14), .D(norm_reg[4]), .E(n20), .F(
        sum1[6]), .Y(n279) );
  OAI22X1 U354 ( .A(n46), .B(n159), .C(n277), .D(n278), .Y(N461) );
  AOI222XL U355 ( .A(sum[8]), .B(n27), .C(n14), .D(norm_reg[5]), .E(n20), .F(
        sum1[7]), .Y(n277) );
  OAI22X1 U356 ( .A(n166), .B(n43), .C(n269), .D(n230), .Y(N488) );
  AOI222XL U357 ( .A(sum[13]), .B(n27), .C(n260), .D(norm_reg[10]), .E(n262), 
        .F(sum1[12]), .Y(n269) );
  OAI22X1 U358 ( .A(n166), .B(n42), .C(n270), .D(n230), .Y(N487) );
  AOI222XL U359 ( .A(sum[12]), .B(n26), .C(n260), .D(norm_reg[9]), .E(n262), 
        .F(sum1[11]), .Y(n270) );
  OAI22X1 U360 ( .A(n6), .B(n44), .C(n268), .D(n230), .Y(N489) );
  AOI222XL U361 ( .A(sum[14]), .B(n27), .C(n260), .D(norm_reg[11]), .E(n262), 
        .F(sum1[13]), .Y(n268) );
  OAI22X1 U362 ( .A(n6), .B(n46), .C(n266), .D(n230), .Y(N491) );
  AOI222XL U363 ( .A(sum[16]), .B(n26), .C(n260), .D(norm_reg[13]), .E(n262), 
        .F(sum1[15]), .Y(n266) );
  OAI22X1 U364 ( .A(n6), .B(n45), .C(n267), .D(n230), .Y(N490) );
  AOI222XL U365 ( .A(sum[15]), .B(n27), .C(n260), .D(norm_reg[12]), .E(n262), 
        .F(sum1[14]), .Y(n267) );
  OAI22X1 U366 ( .A(n45), .B(n2), .C(n297), .D(n291), .Y(N412) );
  AOI221XL U367 ( .A(md3[5]), .B(n15), .C(n298), .D(md3[7]), .E(n299), .Y(n297) );
  OAI22X1 U368 ( .A(n7), .B(n136), .C(n98), .D(n13), .Y(n299) );
  OAI22X1 U369 ( .A(n46), .B(n161), .C(n290), .D(n291), .Y(N413) );
  AOI221XL U370 ( .A(md3[5]), .B(n292), .C(n293), .D(md3[6]), .E(n294), .Y(
        n290) );
  OAI22AX1 U371 ( .D(n27), .C(n13), .A(n187), .B(n296), .Y(n294) );
  INVX1 U372 ( .A(mdu_op[0]), .Y(n430) );
  NAND2X1 U373 ( .A(mdu_op[0]), .B(n431), .Y(n194) );
  OAI21X1 U374 ( .B(n11), .C(n114), .A(n263), .Y(N566) );
  OAI211X1 U375 ( .C(md1[6]), .D(n77), .A(n259), .B(n264), .Y(n263) );
  AOI22X1 U376 ( .A(n97), .B(n96), .C(n77), .D(n125), .Y(n264) );
  INVX1 U377 ( .A(mdu_op[1]), .Y(n431) );
  OAI22X1 U378 ( .A(n43), .B(n2), .C(n305), .D(n291), .Y(N410) );
  AOI221XL U379 ( .A(n302), .B(md3[6]), .C(n29), .D(md3[5]), .E(n306), .Y(n305) );
  OAI222XL U380 ( .A(n300), .B(n448), .C(n100), .D(n295), .E(n304), .F(n135), 
        .Y(n306) );
  INVX1 U381 ( .A(md2[0]), .Y(n443) );
  INVX1 U382 ( .A(md4[0]), .Y(n432) );
  OAI22X1 U383 ( .A(n41), .B(n161), .C(n309), .D(n291), .Y(N408) );
  AOI221XL U384 ( .A(n302), .B(md3[4]), .C(n29), .D(md3[3]), .E(n310), .Y(n309) );
  OAI222XL U385 ( .A(n300), .B(n438), .C(n102), .D(n295), .E(n304), .F(n447), 
        .Y(n310) );
  OAI22X1 U386 ( .A(n42), .B(n2), .C(n307), .D(n291), .Y(N409) );
  AOI221XL U387 ( .A(n302), .B(md3[5]), .C(n30), .D(md3[4]), .E(n308), .Y(n307) );
  OAI222XL U388 ( .A(n300), .B(n447), .C(n101), .D(n295), .E(n304), .F(n448), 
        .Y(n308) );
  INVX1 U389 ( .A(md2[1]), .Y(n440) );
  INVX1 U390 ( .A(md4[1]), .Y(n441) );
  INVX1 U391 ( .A(norm_reg[0]), .Y(n423) );
  OAI22X1 U392 ( .A(n40), .B(n161), .C(n311), .D(n291), .Y(N407) );
  AOI221XL U393 ( .A(n302), .B(md3[3]), .C(n30), .D(md3[2]), .E(n312), .Y(n311) );
  OAI222XL U394 ( .A(n300), .B(n146), .C(n103), .D(n295), .E(n304), .F(n438), 
        .Y(n312) );
  INVX1 U395 ( .A(md2[3]), .Y(n421) );
  INVX1 U396 ( .A(md2[2]), .Y(n439) );
  INVX1 U397 ( .A(md4[3]), .Y(n417) );
  INVX1 U398 ( .A(md4[2]), .Y(n433) );
  INVX1 U399 ( .A(norm_reg[1]), .Y(n420) );
  INVX1 U400 ( .A(norm_reg[2]), .Y(n418) );
  OAI22X1 U401 ( .A(n39), .B(n2), .C(n313), .D(n291), .Y(N406) );
  AOI221XL U402 ( .A(n302), .B(md3[2]), .C(n29), .D(md3[1]), .E(n314), .Y(n313) );
  OAI222XL U403 ( .A(n300), .B(n153), .C(n104), .D(n295), .E(n304), .F(n146), 
        .Y(n314) );
  OAI22X1 U404 ( .A(n46), .B(n162), .C(n316), .D(n317), .Y(N340) );
  AOI221XL U405 ( .A(n302), .B(md3[1]), .C(n30), .D(md3[0]), .E(n318), .Y(n316) );
  OAI222XL U406 ( .A(n300), .B(n152), .C(n105), .D(n295), .E(n304), .F(n153), 
        .Y(n318) );
  INVX1 U407 ( .A(md2[4]), .Y(n415) );
  INVX1 U408 ( .A(md4[4]), .Y(n156) );
  INVX1 U409 ( .A(norm_reg[3]), .Y(n157) );
  OAI22X1 U410 ( .A(n45), .B(n1), .C(n319), .D(n317), .Y(N339) );
  AOI221XL U411 ( .A(n19), .B(md3[0]), .C(n29), .D(md2[7]), .E(n320), .Y(n319)
         );
  OAI222XL U412 ( .A(n300), .B(n415), .C(n106), .D(n295), .E(n304), .F(n152), 
        .Y(n320) );
  INVX1 U413 ( .A(md2[6]), .Y(n153) );
  INVX1 U414 ( .A(md2[5]), .Y(n152) );
  INVX1 U415 ( .A(md4[5]), .Y(n154) );
  INVX1 U416 ( .A(md4[6]), .Y(n148) );
  INVX1 U417 ( .A(norm_reg[4]), .Y(n150) );
  INVX1 U418 ( .A(norm_reg[5]), .Y(n151) );
  OAI22X1 U419 ( .A(n43), .B(n162), .C(n323), .D(n317), .Y(N337) );
  AOI221XL U420 ( .A(n19), .B(md2[6]), .C(n29), .D(md2[5]), .E(n324), .Y(n323)
         );
  OAI222XL U421 ( .A(n300), .B(n439), .C(n108), .D(n295), .E(n304), .F(n421), 
        .Y(n324) );
  OAI22X1 U422 ( .A(n44), .B(n1), .C(n321), .D(n317), .Y(N338) );
  AOI221XL U423 ( .A(n19), .B(md2[7]), .C(n30), .D(md2[6]), .E(n322), .Y(n321)
         );
  OAI222XL U424 ( .A(n7), .B(n421), .C(n107), .D(n13), .E(n23), .F(n415), .Y(
        n322) );
  INVX1 U425 ( .A(md2[7]), .Y(n146) );
  INVX1 U426 ( .A(md4[7]), .Y(n144) );
  INVX1 U427 ( .A(norm_reg[6]), .Y(n145) );
  OAI22X1 U428 ( .A(n42), .B(n162), .C(n325), .D(n317), .Y(N336) );
  AOI221XL U429 ( .A(n19), .B(md2[5]), .C(n30), .D(md2[4]), .E(n326), .Y(n325)
         );
  OAI222XL U430 ( .A(n7), .B(n440), .C(n109), .D(n13), .E(n23), .F(n439), .Y(
        n326) );
  INVX1 U431 ( .A(md3[1]), .Y(n447) );
  INVX1 U432 ( .A(md3[0]), .Y(n438) );
  INVX1 U433 ( .A(md5[1]), .Y(n449) );
  INVX1 U434 ( .A(md5[0]), .Y(n442) );
  INVX1 U435 ( .A(norm_reg[7]), .Y(n142) );
  INVX1 U436 ( .A(norm_reg[8]), .Y(n140) );
  OAI22X1 U437 ( .A(n40), .B(n1), .C(n329), .D(n317), .Y(N334) );
  AOI221XL U438 ( .A(n19), .B(md2[3]), .C(n30), .D(md2[2]), .E(n330), .Y(n329)
         );
  OAI222XL U439 ( .A(n7), .B(n424), .C(n111), .D(n13), .E(n23), .F(n443), .Y(
        n330) );
  OAI22X1 U440 ( .A(n41), .B(n162), .C(n327), .D(n317), .Y(N335) );
  AOI221XL U441 ( .A(n19), .B(md2[4]), .C(n29), .D(md2[3]), .E(n328), .Y(n327)
         );
  OAI222XL U442 ( .A(n7), .B(n443), .C(n110), .D(n13), .E(n23), .F(n440), .Y(
        n328) );
  INVX1 U443 ( .A(md3[2]), .Y(n448) );
  INVX1 U444 ( .A(md5[2]), .Y(n444) );
  INVX1 U445 ( .A(norm_reg[9]), .Y(n138) );
  OAI22X1 U446 ( .A(md4[0]), .B(n34), .C(n189), .D(n432), .Y(arg_d[1]) );
  OAI222XL U447 ( .A(n193), .B(n125), .C(n194), .D(n115), .E(n119), .F(n422), 
        .Y(arg_c[1]) );
  OAI22X1 U448 ( .A(n39), .B(n1), .C(n331), .D(n317), .Y(N333) );
  AOI221XL U449 ( .A(n19), .B(md2[2]), .C(n29), .D(md2[1]), .E(n333), .Y(n331)
         );
  OAI222XL U450 ( .A(n7), .B(n115), .C(n113), .D(n13), .E(n23), .F(n424), .Y(
        n333) );
  OAI22X1 U451 ( .A(n40), .B(n357), .C(n372), .D(n359), .Y(N192) );
  AOI221XL U452 ( .A(md0[0]), .B(n15), .C(md0[3]), .D(n371), .E(n373), .Y(n372) );
  ENOX1 U453 ( .A(n112), .B(n374), .C(n29), .D(md0[2]), .Y(n373) );
  OAI22X1 U454 ( .A(n41), .B(n357), .C(n369), .D(n359), .Y(N193) );
  AOI221XL U455 ( .A(md0[0]), .B(n65), .C(md0[1]), .D(n70), .E(n370), .Y(n369)
         );
  ENOX1 U456 ( .A(n22), .B(n95), .C(n30), .D(md0[3]), .Y(n370) );
  OAI22X1 U457 ( .A(n42), .B(n357), .C(n367), .D(n359), .Y(N194) );
  AOI221XL U458 ( .A(md0[1]), .B(n65), .C(md0[2]), .D(n70), .E(n368), .Y(n367)
         );
  OAI22X1 U459 ( .A(n69), .B(n95), .C(n66), .D(n92), .Y(n368) );
  OAI22X1 U460 ( .A(n43), .B(n357), .C(n365), .D(n359), .Y(N195) );
  AOI221XL U461 ( .A(md0[2]), .B(n65), .C(md0[3]), .D(n70), .E(n366), .Y(n365)
         );
  OAI22X1 U462 ( .A(n69), .B(n92), .C(n66), .D(n89), .Y(n366) );
  OAI22X1 U463 ( .A(n44), .B(n357), .C(n363), .D(n359), .Y(N196) );
  AOI221XL U464 ( .A(md0[3]), .B(n65), .C(md0[4]), .D(n70), .E(n364), .Y(n363)
         );
  OAI22X1 U465 ( .A(n69), .B(n89), .C(n66), .D(n90), .Y(n364) );
  OAI22X1 U466 ( .A(n46), .B(n357), .C(n358), .D(n359), .Y(N198) );
  AOI221XL U467 ( .A(md0[5]), .B(n10), .C(md0[6]), .D(n15), .E(n360), .Y(n358)
         );
  OAI22X1 U468 ( .A(n69), .B(n434), .C(n66), .D(n446), .Y(n360) );
  OAI22X1 U469 ( .A(n45), .B(n357), .C(n361), .D(n359), .Y(N197) );
  AOI221XL U470 ( .A(md0[4]), .B(n10), .C(md0[5]), .D(n15), .E(n362), .Y(n361)
         );
  OAI22X1 U471 ( .A(n69), .B(n90), .C(n22), .D(n434), .Y(n362) );
  OAI22X1 U472 ( .A(n40), .B(n239), .C(n351), .D(n158), .Y(N260) );
  AOI221XL U473 ( .A(md0[7]), .B(n65), .C(md1[0]), .D(n70), .E(n352), .Y(n351)
         );
  OAI22X1 U474 ( .A(n69), .B(n445), .C(n66), .D(n123), .Y(n352) );
  OAI22X1 U475 ( .A(n41), .B(n239), .C(n349), .D(n158), .Y(N261) );
  AOI221XL U476 ( .A(md1[0]), .B(n65), .C(md1[1]), .D(n70), .E(n350), .Y(n349)
         );
  OAI22X1 U477 ( .A(n69), .B(n123), .C(n66), .D(n93), .Y(n350) );
  OAI22X1 U478 ( .A(n39), .B(n239), .C(n353), .D(n158), .Y(N259) );
  AOI221XL U479 ( .A(md0[6]), .B(n65), .C(md0[7]), .D(n70), .E(n355), .Y(n353)
         );
  OAI22X1 U480 ( .A(n69), .B(n446), .C(n66), .D(n445), .Y(n355) );
  OAI22X1 U481 ( .A(n46), .B(n239), .C(n338), .D(n158), .Y(N266) );
  AOI221XL U482 ( .A(n302), .B(md2[1]), .C(n30), .D(md2[0]), .E(n339), .Y(n338) );
  OAI222XL U483 ( .A(n23), .B(n115), .C(n340), .D(n91), .E(n114), .F(n336), 
        .Y(n339) );
  OAI22X1 U484 ( .A(n42), .B(n239), .C(n347), .D(n158), .Y(N262) );
  AOI221XL U485 ( .A(md1[1]), .B(n65), .C(md1[2]), .D(n70), .E(n348), .Y(n347)
         );
  OAI22X1 U486 ( .A(n69), .B(n93), .C(n66), .D(n91), .Y(n348) );
  OAI22X1 U487 ( .A(n45), .B(n239), .C(n341), .D(n158), .Y(N265) );
  AOI221XL U488 ( .A(n302), .B(md2[0]), .C(n29), .D(md1[7]), .E(n342), .Y(n341) );
  OAI222XL U489 ( .A(n23), .B(n91), .C(n340), .D(n93), .E(n425), .F(n336), .Y(
        n342) );
  OAI22X1 U490 ( .A(n43), .B(n239), .C(n345), .D(n158), .Y(N263) );
  AOI221XL U491 ( .A(md1[2]), .B(n65), .C(md1[3]), .D(n70), .E(n346), .Y(n345)
         );
  OAI22X1 U492 ( .A(n69), .B(n91), .C(n66), .D(n115), .Y(n346) );
  OAI22X1 U493 ( .A(n44), .B(n239), .C(n343), .D(n158), .Y(N264) );
  AOI221XL U494 ( .A(md1[3]), .B(n65), .C(md1[4]), .D(n70), .E(n344), .Y(n343)
         );
  OAI22X1 U495 ( .A(n115), .B(n5), .C(n66), .D(n424), .Y(n344) );
  OAI21BX1 U496 ( .C(set_div16), .B(n158), .A(n159), .Y(n414) );
  OAI31XL U497 ( .A(n430), .B(n48), .C(n55), .D(n169), .Y(n411) );
  AOI31X1 U498 ( .A(set_div16), .B(n58), .C(n55), .D(n51), .Y(n169) );
  INVX1 U499 ( .A(n166), .Y(n55) );
  OAI211X1 U500 ( .C(n58), .D(n166), .A(n167), .B(n168), .Y(n412) );
  NAND3X1 U501 ( .A(n166), .B(n47), .C(mdu_op[1]), .Y(n167) );
  OAI211X1 U502 ( .C(n211), .D(n198), .A(n166), .B(n168), .Y(N894) );
  AOI211X1 U503 ( .C(n85), .D(n430), .A(n212), .B(n213), .Y(n211) );
  OAI221X1 U504 ( .A(n182), .B(n199), .C(n64), .D(n208), .E(n215), .Y(n212) );
  ENOX1 U505 ( .A(md3[7]), .B(n202), .C(n82), .D(n214), .Y(n213) );
  INVX1 U506 ( .A(md3[4]), .Y(n136) );
  INVX1 U507 ( .A(md3[3]), .Y(n135) );
  AOI31X1 U508 ( .A(n226), .B(n227), .C(n228), .D(n198), .Y(N892) );
  OR2X1 U509 ( .A(n205), .B(n206), .Y(n227) );
  AOI32X1 U510 ( .A(n233), .B(n234), .C(n214), .D(n83), .E(arcon[5]), .Y(n226)
         );
  AOI221XL U511 ( .A(n80), .B(n209), .C(n85), .D(n193), .E(n225), .Y(n228) );
  INVX1 U512 ( .A(md5[4]), .Y(n132) );
  INVX1 U513 ( .A(md5[3]), .Y(n131) );
  INVX1 U514 ( .A(norm_reg[10]), .Y(n133) );
  INVX1 U515 ( .A(norm_reg[11]), .Y(n134) );
  INVX1 U516 ( .A(n171), .Y(n50) );
  AOI32X1 U517 ( .A(arcon[5]), .B(n47), .C(n168), .D(n51), .E(sfrdatai[5]), 
        .Y(n171) );
  INVX1 U518 ( .A(md5[5]), .Y(n128) );
  INVX1 U519 ( .A(norm_reg[12]), .Y(n127) );
  INVX1 U520 ( .A(md3[6]), .Y(n125) );
  INVX1 U521 ( .A(md3[7]), .Y(n426) );
  INVX1 U522 ( .A(md5[6]), .Y(n121) );
  INVX1 U523 ( .A(md5[7]), .Y(n124) );
  INVX1 U524 ( .A(norm_reg[13]), .Y(n122) );
  INVX1 U525 ( .A(norm_reg[14]), .Y(n117) );
  NAND2X1 U526 ( .A(md0[1]), .B(n34), .Y(n189) );
  AOI211X1 U527 ( .C(sfroe), .D(n52), .A(n170), .B(n48), .Y(n410) );
  NOR2X1 U528 ( .A(arcon[7]), .B(test_so), .Y(n170) );
  INVX1 U529 ( .A(md1[6]), .Y(n115) );
  AOI21BBXL U530 ( .B(md3[6]), .C(n296), .A(n292), .Y(n300) );
  NOR2X1 U531 ( .A(n88), .B(oper_reg[2]), .Y(n402) );
  NOR2X1 U532 ( .A(n86), .B(oper_reg[1]), .Y(n234) );
  OA222X1 U533 ( .A(counter_st[1]), .B(n384), .C(n394), .D(n382), .E(n385), 
        .F(n435), .Y(n251) );
  OA222X1 U534 ( .A(n60), .B(n382), .C(n390), .D(n384), .E(n385), .F(n118), 
        .Y(n249) );
  INVX1 U535 ( .A(arcon[3]), .Y(n118) );
  AOI21X1 U536 ( .B(counter_st[3]), .C(n73), .A(n386), .Y(n390) );
  INVX1 U537 ( .A(n389), .Y(n60) );
  OA222X1 U538 ( .A(n59), .B(n382), .C(n392), .D(n384), .E(n385), .F(n437), 
        .Y(n250) );
  AOI21X1 U539 ( .B(counter_st[2]), .C(counter_st[1]), .A(n393), .Y(n392) );
  INVX1 U540 ( .A(n391), .Y(n59) );
  OA222X1 U541 ( .A(n381), .B(n382), .C(n383), .D(n384), .E(n385), .F(n94), 
        .Y(n247) );
  INVX1 U542 ( .A(arcon[4]), .Y(n94) );
  AOI21BBXL U543 ( .B(n71), .C(n386), .A(n68), .Y(n383) );
  OA222X1 U544 ( .A(N610), .B(n382), .C(n384), .D(n62), .E(n385), .F(n436), 
        .Y(n252) );
  OAI31XL U545 ( .A(n395), .B(n335), .C(n75), .D(n385), .Y(n384) );
  OAI21X1 U546 ( .B(md3[6]), .C(n77), .A(n67), .Y(n395) );
  NAND3X1 U547 ( .A(n400), .B(oper_reg[3]), .C(oper_reg[2]), .Y(n204) );
  NOR2X1 U548 ( .A(oper_reg[3]), .B(oper_reg[2]), .Y(n398) );
  NOR2X1 U549 ( .A(oper_reg[1]), .B(oper_reg[0]), .Y(n400) );
  INVX1 U550 ( .A(oper_reg[0]), .Y(n86) );
  INVX1 U551 ( .A(oper_reg[1]), .Y(n81) );
  INVX1 U552 ( .A(oper_reg[3]), .Y(n88) );
  INVX1 U553 ( .A(oper_reg[2]), .Y(n87) );
  NOR32XL U554 ( .B(oper_reg[1]), .C(n233), .A(oper_reg[0]), .Y(n224) );
  NOR2X1 U555 ( .A(n87), .B(oper_reg[3]), .Y(n233) );
  NOR2X1 U556 ( .A(counter_st[2]), .B(counter_st[1]), .Y(n393) );
  NOR2X1 U557 ( .A(n73), .B(counter_st[3]), .Y(n386) );
  NOR32XL U558 ( .B(n231), .C(counter_st[2]), .A(counter_st[3]), .Y(n223) );
  XNOR2XL U559 ( .A(n387), .B(counter_st[3]), .Y(n389) );
  AOI22BXL U560 ( .B(n387), .A(n217), .D(n388), .C(counter_st[4]), .Y(n381) );
  NOR2X1 U561 ( .A(counter_st[3]), .B(n387), .Y(n388) );
  INVX1 U562 ( .A(N610), .Y(n62) );
  NAND3X1 U563 ( .A(oper_reg[1]), .B(n86), .C(n398), .Y(n206) );
  NOR2X1 U564 ( .A(counter_st[3]), .B(counter_st[4]), .Y(n217) );
  NAND3X1 U565 ( .A(n234), .B(oper_reg[3]), .C(oper_reg[2]), .Y(n221) );
  INVX1 U566 ( .A(counter_st[4]), .Y(n71) );
  NOR2X1 U567 ( .A(counter_st[1]), .B(N610), .Y(n231) );
  NAND2X1 U568 ( .A(n187), .B(n216), .Y(n199) );
  NAND4X1 U569 ( .A(counter_st[1]), .B(n217), .C(n62), .D(n72), .Y(n216) );
  NAND2X1 U570 ( .A(counter_st[4]), .B(n223), .Y(n209) );
  AOI21X1 U571 ( .B(counter_st[1]), .C(N610), .A(n231), .Y(n394) );
  OAI22X1 U572 ( .A(n194), .B(n204), .C(arcon[5]), .D(n215), .Y(n222) );
  OAI31XL U573 ( .A(n202), .B(md3[7]), .C(n203), .D(n182), .Y(n225) );
  NOR2X1 U574 ( .A(md3[6]), .B(md3[5]), .Y(n187) );
  NAND4X1 U575 ( .A(n436), .B(n435), .C(n235), .D(n437), .Y(n203) );
  NOR2X1 U576 ( .A(arcon[4]), .B(arcon[3]), .Y(n235) );
  NOR4XL U577 ( .A(md4[2]), .B(md4[1]), .C(md4[0]), .D(n181), .Y(n175) );
  NOR4XL U578 ( .A(n179), .B(n180), .C(md5[4]), .D(md5[3]), .Y(n177) );
  NAND4X1 U579 ( .A(n144), .B(n442), .C(n449), .D(n444), .Y(n179) );
  NAND3X1 U580 ( .A(n121), .B(n124), .C(n128), .Y(n180) );
  NAND4X1 U581 ( .A(counter_st[4]), .B(counter_st[1]), .C(n232), .D(n62), .Y(
        n205) );
  NOR2X1 U582 ( .A(counter_st[3]), .B(counter_st[2]), .Y(n232) );
  INVX1 U583 ( .A(counter_st[2]), .Y(n72) );
  AOI31X1 U584 ( .A(n172), .B(n173), .C(n174), .D(n48), .Y(n408) );
  NAND4X1 U585 ( .A(arcon[6]), .B(n182), .C(n183), .D(n181), .Y(n173) );
  OAI31XL U586 ( .A(n184), .B(n185), .C(n186), .D(n84), .Y(n172) );
  AOI31X1 U587 ( .A(n175), .B(n176), .C(n177), .D(n178), .Y(n174) );
  INVX1 U588 ( .A(md1[7]), .Y(n424) );
  NAND4X1 U589 ( .A(n443), .B(n440), .C(n187), .D(n188), .Y(n184) );
  NOR4XL U590 ( .A(md2[5]), .B(md2[4]), .C(md2[3]), .D(md2[2]), .Y(n188) );
  INVX1 U591 ( .A(arcon[1]), .Y(n435) );
  INVX1 U592 ( .A(md1[5]), .Y(n91) );
  INVX1 U593 ( .A(arcon[2]), .Y(n437) );
  INVX1 U594 ( .A(md1[4]), .Y(n93) );
  INVX1 U595 ( .A(arcon[0]), .Y(n436) );
  NOR4XL U596 ( .A(md4[6]), .B(md4[5]), .C(md4[4]), .D(md4[3]), .Y(n176) );
  INVX1 U597 ( .A(md1[1]), .Y(n446) );
  INVX1 U598 ( .A(set_div32), .Y(n58) );
  INVX1 U599 ( .A(md0[4]), .Y(n95) );
  INVX1 U600 ( .A(md1[3]), .Y(n123) );
  INVX1 U601 ( .A(md0[6]), .Y(n89) );
  INVX1 U602 ( .A(md0[7]), .Y(n90) );
  INVX1 U603 ( .A(md0[5]), .Y(n92) );
  INVX1 U604 ( .A(md1[2]), .Y(n445) );
  INVX1 U605 ( .A(md1[0]), .Y(n434) );
endmodule


module mdu_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module mdu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module wakeupctrl_a0 ( irq, int0ff, int1ff, it0, it1, isreg, intprior0, 
        intprior1, eal, eint0, eint1, pmuintreq );
  input [3:0] isreg;
  input [1:0] intprior0;
  input [1:0] intprior1;
  input irq, int0ff, int1ff, it0, it1, eal, eint0, eint1;
  output pmuintreq;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n1;

  NAND42X1 U1 ( .C(it0), .D(int0ff), .A(eint0), .B(n9), .Y(n3) );
  OAI2B11X1 U2 ( .D(intprior0[0]), .C(n6), .A(n10), .B(n8), .Y(n9) );
  OAI21X1 U3 ( .B(intprior0[0]), .C(n1), .A(intprior1[0]), .Y(n10) );
  AO21X1 U4 ( .B(n2), .C(eal), .A(irq), .Y(pmuintreq) );
  AOI21X1 U5 ( .B(n3), .C(n4), .A(isreg[3]), .Y(n2) );
  NAND42X1 U6 ( .C(it1), .D(int1ff), .A(eint1), .B(n5), .Y(n4) );
  OAI2B11X1 U7 ( .D(intprior0[1]), .C(n6), .A(n7), .B(n8), .Y(n5) );
  OAI21X1 U8 ( .B(intprior0[1]), .C(n1), .A(intprior1[1]), .Y(n7) );
  OR2X1 U9 ( .A(isreg[1]), .B(isreg[2]), .Y(n6) );
  OR2X1 U10 ( .A(isreg[0]), .B(n6), .Y(n8) );
  INVX1 U11 ( .A(isreg[2]), .Y(n1) );
endmodule


module pmurstctrl_a0 ( resetff, wdts, srst, pmuintreq, stop, idle, clkcpu_en, 
        clkper_en, cpu_resume, rsttowdt, rsttosrst, rst );
  input resetff, wdts, srst, pmuintreq, stop, idle;
  output clkcpu_en, clkper_en, cpu_resume, rsttowdt, rsttosrst, rst;
  wire   n2;

  OAI21X1 U1 ( .B(stop), .C(idle), .A(n2), .Y(clkcpu_en) );
  NAND2X1 U2 ( .A(stop), .B(n2), .Y(clkper_en) );
  BUFX3 U3 ( .A(pmuintreq), .Y(cpu_resume) );
  INVX1 U4 ( .A(pmuintreq), .Y(n2) );
  OR2X1 U5 ( .A(srst), .B(resetff), .Y(rsttowdt) );
  OR2X1 U6 ( .A(wdts), .B(rsttowdt), .Y(rst) );
  OR2X1 U7 ( .A(resetff), .B(wdts), .Y(rsttosrst) );
endmodule


module sfrmux_a0 ( isfrwait, sfraddr, c, ac, f0, rs, ov, f1, p, acc, b, dpl, 
        dph, dps, dpc, p2, sp, smod, pmw, p2sel, gf0, stop, idle, ckcon, port0, 
        port0ff, rmwinstr, arcon, md0, md1, md2, md3, md4, md5, t0_tmod, 
        t0_tf0, t0_tf1, t0_tr0, t0_tr1, tl0, th0, t1_tmod, t1_tf1, t1_tr1, tl1, 
        th1, wdtrel, ip0wdts, wdt_tm, t2con, s0con, s0buf, s0rell, s0relh, bd, 
        ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9, 
        iex10, iex11, iex12, ien0, ien1, ien2, ip0, ip1, isr_tm, i2c_int, 
        i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o, sfrdatai, tf1_gate, riti0_gate, 
        iex7_gate, iex2_gate, srstflag, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, ext_sfr_sel, sfrdatao );
  input [6:0] sfraddr;
  input [1:0] rs;
  input [7:0] acc;
  input [7:0] b;
  input [7:0] dpl;
  input [7:0] dph;
  input [3:0] dps;
  input [5:0] dpc;
  input [7:0] p2;
  input [7:0] sp;
  input [7:0] ckcon;
  input [7:0] port0;
  input [7:0] port0ff;
  input [7:0] arcon;
  input [7:0] md0;
  input [7:0] md1;
  input [7:0] md2;
  input [7:0] md3;
  input [7:0] md4;
  input [7:0] md5;
  input [3:0] t0_tmod;
  input [7:0] tl0;
  input [7:0] th0;
  input [3:0] t1_tmod;
  input [7:0] tl1;
  input [7:0] th1;
  input [7:0] wdtrel;
  input [7:0] t2con;
  input [7:0] s0con;
  input [7:0] s0buf;
  input [7:0] s0rell;
  input [7:0] s0relh;
  input [7:0] ien0;
  input [5:0] ien1;
  input [5:0] ien2;
  input [5:0] ip0;
  input [5:0] ip1;
  input [7:0] i2cdat_o;
  input [7:0] i2cadr_o;
  input [7:0] i2ccon_o;
  input [7:0] i2csta_o;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  input isfrwait, c, ac, f0, ov, f1, p, smod, pmw, p2sel, gf0, stop, idle,
         rmwinstr, t0_tf0, t0_tf1, t0_tr0, t0_tr1, t1_tf1, t1_tr1, ip0wdts,
         wdt_tm, bd, ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12, isr_tm, i2c_int, srstflag;
  output tf1_gate, riti0_gate, iex7_gate, iex2_gate, int_vect_8b, int_vect_93,
         int_vect_9b, int_vect_a3, ext_sfr_sel;
  wire   n34, n35, n36, n37, n72, n73, n74, n75, n94, n95, n96, n97, n116,
         n117, n118, n119, n136, n137, n138, n139, net83096, net83100,
         net83124, net83162, net83163, net83249, net83252, net83253, net83264,
         net83318, net83319, net83320, net83322, net83333, net83334, net83339,
         net83346, net83348, net83357, net83359, net83362, net83365, net83372,
         net83389, net83393, net83394, net87439, net87461, net87609, net88957,
         net89060, net95004, net96039, net97663, net97744, net97764, net97776,
         net97837, net97856, net97864, net98352, net98374, net98635, net99166,
         net99226, net99404, net99568, net99800, net100030, net100109,
         net100143, net100193, net101202, net101395, net101453, net101493,
         net101591, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356;

  NOR6X1 U2 ( .A(net83357), .B(net97776), .C(net99568), .D(net87439), .E(
        net87609), .F(net101202), .Y(net97837) );
  NOR21X1 U3 ( .B(net97864), .A(net83362), .Y(net101453) );
  NOR2X1 U4 ( .A(net96039), .B(n132), .Y(net97864) );
  AND4X2 U5 ( .A(n9), .B(net83320), .C(net83322), .D(net83319), .Y(net83318)
         );
  NAND31X1 U6 ( .C(sfraddr[0]), .A(sfraddr[1]), .B(net89060), .Y(net83359) );
  INVX1 U7 ( .A(n164), .Y(n341) );
  AOI221X1 U8 ( .A(s0rell[2]), .B(n319), .C(dph[2]), .D(n322), .E(n249), .Y(
        n256) );
  NAND42X1 U9 ( .C(net98635), .D(sfraddr[5]), .A(net101202), .B(n6), .Y(n8) );
  NAND21X2 U10 ( .B(net100030), .A(n46), .Y(n160) );
  INVX2 U11 ( .A(sfraddr[2]), .Y(net89060) );
  INVXL U12 ( .A(n127), .Y(n126) );
  INVX1 U13 ( .A(md2[0]), .Y(n71) );
  INVX1 U14 ( .A(md3[0]), .Y(n76) );
  INVX1 U15 ( .A(th0[0]), .Y(n77) );
  INVXL U16 ( .A(net83359), .Y(net98352) );
  NOR2X2 U17 ( .A(net99166), .B(sfraddr[1]), .Y(net95004) );
  INVX2 U18 ( .A(sfraddr[1]), .Y(net97856) );
  BUFX3 U19 ( .A(net97776), .Y(net97663) );
  NAND32X1 U20 ( .B(net97856), .C(n14), .A(net89060), .Y(net100030) );
  NAND21X1 U21 ( .B(net89060), .A(net99226), .Y(n40) );
  INVXL U22 ( .A(n61), .Y(n21) );
  INVX1 U23 ( .A(sp[2]), .Y(n78) );
  INVX1 U24 ( .A(port0ff[2]), .Y(n80) );
  INVX1 U25 ( .A(dpl[2]), .Y(n79) );
  INVX1 U26 ( .A(n163), .Y(n343) );
  INVX1 U27 ( .A(n201), .Y(n295) );
  INVX1 U28 ( .A(n207), .Y(n317) );
  OA222X1 U29 ( .A(n16), .B(n220), .C(n17), .D(n219), .E(n18), .F(net83264), 
        .Y(net83319) );
  INVX1 U30 ( .A(n243), .Y(n38) );
  INVX1 U31 ( .A(net99226), .Y(net100193) );
  NAND32X1 U32 ( .B(net87609), .C(n25), .A(n122), .Y(n162) );
  NAND31X1 U33 ( .C(net89060), .A(n24), .B(net100143), .Y(n164) );
  INVX1 U34 ( .A(net97837), .Y(net83348) );
  EORX1 U35 ( .A(dpl[1]), .B(n323), .C(n33), .D(n261), .Y(n89) );
  INVX1 U36 ( .A(port0ff[1]), .Y(n33) );
  NAND32X1 U37 ( .B(sfraddr[5]), .C(n134), .A(net99568), .Y(net83252) );
  INVX1 U38 ( .A(i2ccon_o[0]), .Y(n17) );
  INVX1 U39 ( .A(s0relh[0]), .Y(n18) );
  INVX1 U40 ( .A(i2cdat_o[0]), .Y(n16) );
  NOR2X1 U41 ( .A(n83), .B(n261), .Y(n64) );
  INVX1 U42 ( .A(net83264), .Y(net83096) );
  NOR3X1 U43 ( .A(n11), .B(n12), .C(net97776), .Y(net97764) );
  INVX1 U44 ( .A(n15), .Y(net83100) );
  INVX1 U45 ( .A(net101453), .Y(net83334) );
  INVX1 U46 ( .A(n29), .Y(n154) );
  INVX1 U47 ( .A(ov), .Y(n22) );
  INVX1 U48 ( .A(port0[2]), .Y(n20) );
  AOI221X1 U49 ( .A(tl0[2]), .B(n346), .C(t0_tmod[2]), .D(n66), .E(n244), .Y(
        n259) );
  INVX1 U50 ( .A(md2[2]), .Y(n57) );
  INVX1 U51 ( .A(md1[2]), .Y(n58) );
  NAND31X1 U52 ( .C(n215), .A(n214), .B(n213), .Y(n216) );
  AND3X1 U53 ( .A(n205), .B(n204), .C(n203), .Y(n214) );
  NOR43XL U54 ( .B(n194), .C(n193), .D(n192), .A(n191), .Y(n217) );
  NOR43XL U55 ( .B(n229), .C(n228), .D(n227), .A(n226), .Y(n240) );
  NAND32X1 U56 ( .B(net101395), .C(n156), .A(rmwinstr), .Y(n184) );
  INVX1 U57 ( .A(n125), .Y(n158) );
  NAND2X2 U58 ( .A(n67), .B(n68), .Y(sfrdatao[0]) );
  NAND2X1 U59 ( .A(n184), .B(n158), .Y(n261) );
  INVXL U60 ( .A(sfraddr[6]), .Y(net96039) );
  NOR2X1 U61 ( .A(n30), .B(n222), .Y(n1) );
  NOR2X1 U62 ( .A(n31), .B(n221), .Y(n2) );
  NOR2X1 U63 ( .A(n32), .B(n159), .Y(n3) );
  NOR3XL U64 ( .A(n1), .B(n2), .C(n3), .Y(net83320) );
  INVX1 U65 ( .A(s0buf[0]), .Y(n30) );
  INVX1 U66 ( .A(acc[0]), .Y(n31) );
  NAND32XL U67 ( .B(net87439), .C(n134), .A(net99568), .Y(n221) );
  INVX1 U68 ( .A(i2csta_o[0]), .Y(n32) );
  AND2X1 U69 ( .A(ip1[0]), .B(net83163), .Y(n4) );
  AND2X1 U70 ( .A(iex7), .B(net83162), .Y(n5) );
  NOR3X1 U71 ( .A(n4), .B(n5), .C(n10), .Y(n9) );
  INVX3 U72 ( .A(n160), .Y(n345) );
  INVX1 U73 ( .A(sfraddr[3]), .Y(net101591) );
  INVXL U74 ( .A(n157), .Y(n323) );
  NAND21XL U75 ( .B(net83359), .A(n143), .Y(n157) );
  NAND21X1 U76 ( .B(net83359), .A(net97864), .Y(n233) );
  INVX1 U77 ( .A(n69), .Y(n122) );
  INVX1 U78 ( .A(n182), .Y(n320) );
  INVX1 U79 ( .A(n234), .Y(n351) );
  INVX1 U80 ( .A(n183), .Y(n321) );
  OR3X2 U81 ( .A(net97776), .B(net89060), .C(sfraddr[1]), .Y(n69) );
  BUFX1 U82 ( .A(sfraddr[2]), .Y(n7) );
  AO222X1 U83 ( .A(md0[0]), .B(net101453), .C(i2cadr_o[0]), .D(net97764), .E(
        t2con[0]), .F(net83100), .Y(n10) );
  BUFXL U84 ( .A(n8), .Y(n15) );
  NAND21XL U85 ( .B(n15), .A(t2con[1]), .Y(net83249) );
  INVX1 U86 ( .A(net83252), .Y(net83162) );
  INVXL U87 ( .A(net83253), .Y(net83163) );
  BUFX3 U88 ( .A(iex7), .Y(iex7_gate) );
  INVX3 U89 ( .A(sfraddr[6]), .Y(net97776) );
  OR3X4 U90 ( .A(net97856), .B(n14), .C(n7), .Y(n12) );
  INVX2 U91 ( .A(sfraddr[0]), .Y(n14) );
  INVX1 U92 ( .A(n14), .Y(net99800) );
  OR3X2 U93 ( .A(n14), .B(sfraddr[1]), .C(sfraddr[2]), .Y(net83362) );
  NAND32X1 U94 ( .B(n13), .C(net87461), .A(net87439), .Y(n11) );
  INVX3 U95 ( .A(sfraddr[5]), .Y(net87439) );
  INVX3 U96 ( .A(sfraddr[4]), .Y(net87461) );
  INVX1 U97 ( .A(sfraddr[3]), .Y(n13) );
  AND4X1 U98 ( .A(net83348), .B(net83264), .C(net83346), .D(n8), .Y(net83372)
         );
  BUFX2 U99 ( .A(net97744), .Y(n6) );
  INVXL U100 ( .A(n6), .Y(net83389) );
  NAND21X4 U101 ( .B(sfraddr[2]), .A(net95004), .Y(net83339) );
  BUFX8 U102 ( .A(sfraddr[0]), .Y(net99166) );
  INVXL U103 ( .A(sfraddr[0]), .Y(net87609) );
  BUFX3 U104 ( .A(sfraddr[4]), .Y(net98635) );
  BUFX2 U105 ( .A(sfraddr[4]), .Y(net99404) );
  INVX1 U106 ( .A(net83362), .Y(net83394) );
  NAND42X1 U107 ( .C(net99404), .D(sfraddr[6]), .A(net87439), .B(net101202), 
        .Y(n133) );
  BUFXL U108 ( .A(net83339), .Y(net101395) );
  NOR31XL U109 ( .C(net99166), .A(n156), .B(n27), .Y(n44) );
  NOR3X1 U110 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[3]), .Y(n87) );
  NAND2X2 U111 ( .A(n49), .B(n50), .Y(sfrdatao[2]) );
  INVX1 U112 ( .A(n220), .Y(n353) );
  NAND32XL U113 ( .B(net96039), .C(net83359), .A(n325), .Y(n220) );
  INVX1 U114 ( .A(n219), .Y(n352) );
  INVX1 U115 ( .A(n19), .Y(n255) );
  INVXL U116 ( .A(net101202), .Y(net101493) );
  BUFX3 U117 ( .A(sfraddr[3]), .Y(net101202) );
  OAI221X1 U118 ( .A(n20), .B(n21), .C(n22), .D(n183), .E(n23), .Y(n19) );
  OA222X1 U119 ( .A(n78), .B(n182), .C(n79), .D(n157), .E(n80), .F(n261), .Y(
        n23) );
  INVX1 U120 ( .A(n54), .Y(n24) );
  NAND42X1 U121 ( .C(net98635), .D(sfraddr[6]), .A(net87439), .B(net101202), 
        .Y(n54) );
  INVX3 U122 ( .A(n133), .Y(n128) );
  INVXL U123 ( .A(n221), .Y(n349) );
  NAND32X1 U124 ( .B(net101591), .C(net87461), .A(net87439), .Y(n47) );
  NAND2X1 U125 ( .A(sfrdatai[1]), .B(n92), .Y(n39) );
  NAND3X1 U126 ( .A(sfraddr[3]), .B(sfraddr[5]), .C(net87461), .Y(n25) );
  NAND3XL U127 ( .A(sfraddr[3]), .B(sfraddr[5]), .C(net87461), .Y(n132) );
  INVXL U128 ( .A(n45), .Y(n26) );
  NAND21X1 U129 ( .B(net89060), .A(net99226), .Y(n27) );
  NAND21X1 U130 ( .B(net89060), .A(net99226), .Y(net83357) );
  OR2XL U131 ( .A(n127), .B(n134), .Y(n196) );
  NOR43XL U132 ( .B(n160), .C(n163), .D(n176), .A(n346), .Y(n129) );
  NOR3XL U133 ( .A(net87609), .B(n156), .C(net83357), .Y(n28) );
  NOR3X2 U134 ( .A(n55), .B(net83359), .C(net88957), .Y(n29) );
  INVX3 U135 ( .A(n151), .Y(n331) );
  INVXL U136 ( .A(n28), .Y(n161) );
  BUFX1 U137 ( .A(sfraddr[1]), .Y(net99226) );
  INVX3 U138 ( .A(n176), .Y(n45) );
  INVX1 U139 ( .A(n222), .Y(n324) );
  NAND21X1 U140 ( .B(net83362), .A(n128), .Y(n163) );
  NAND21X2 U141 ( .B(net83339), .A(n128), .Y(n176) );
  NAND21XL U142 ( .B(n177), .A(tl0[1]), .Y(n178) );
  NOR21X1 U143 ( .B(n93), .A(n262), .Y(n92) );
  NAND4X2 U144 ( .A(n39), .B(n38), .C(n242), .D(n241), .Y(sfrdatao[1]) );
  INVXL U145 ( .A(net83357), .Y(net83365) );
  NAND21XL U146 ( .B(net101395), .A(n143), .Y(n125) );
  INVXL U147 ( .A(net83339), .Y(net83393) );
  NAND21X1 U148 ( .B(n131), .A(net83393), .Y(n188) );
  INVXL U149 ( .A(n184), .Y(n333) );
  BUFXL U150 ( .A(net95004), .Y(net100143) );
  NAND32XL U151 ( .B(n55), .C(net83362), .A(net97663), .Y(n222) );
  INVXL U152 ( .A(net83394), .Y(net100109) );
  NAND21X1 U153 ( .B(net87461), .A(sfraddr[5]), .Y(n127) );
  NAND31XL U154 ( .C(n25), .A(net83394), .B(net97663), .Y(n206) );
  NAND32X1 U155 ( .B(net99568), .C(n134), .A(net87439), .Y(n183) );
  BUFX1 U156 ( .A(n262), .Y(n41) );
  NOR21XL U157 ( .B(n93), .A(n41), .Y(n48) );
  NOR21X2 U158 ( .B(n93), .A(n262), .Y(n42) );
  NOR21XL U159 ( .B(n93), .A(n41), .Y(n43) );
  OR3X4 U160 ( .A(n40), .B(n156), .C(net99800), .Y(n208) );
  NAND32X2 U161 ( .B(n55), .C(net83339), .A(net97663), .Y(net83346) );
  INVX3 U162 ( .A(net83346), .Y(net83124) );
  AO222X1 U163 ( .A(ien1[2]), .B(n290), .C(ien0[2]), .D(n318), .E(ien2[2]), 
        .F(n29), .Y(n249) );
  NAND32X2 U164 ( .B(net83339), .C(n25), .A(net97663), .Y(n153) );
  INVX2 U165 ( .A(net98635), .Y(net99568) );
  INVXL U166 ( .A(n26), .Y(n347) );
  AND4X1 U167 ( .A(net83372), .B(n140), .C(n135), .D(net83252), .Y(n141) );
  NAND32X1 U168 ( .B(net88957), .C(net101591), .A(n126), .Y(n131) );
  INVX2 U169 ( .A(net97776), .Y(net88957) );
  NAND42X4 U170 ( .C(n148), .D(n149), .A(n147), .B(n146), .Y(n262) );
  NAND32X1 U171 ( .B(n27), .C(n54), .A(net87609), .Y(n195) );
  INVXL U172 ( .A(n54), .Y(n46) );
  NAND6X1 U173 ( .A(n255), .B(n258), .C(n257), .D(n256), .E(n259), .F(n254), 
        .Y(n260) );
  INVX2 U174 ( .A(n177), .Y(n346) );
  NAND2X1 U175 ( .A(tl0[0]), .B(n346), .Y(n52) );
  INVXL U176 ( .A(net97764), .Y(net83333) );
  NOR21X2 U177 ( .B(sfraddr[6]), .A(net83339), .Y(net97744) );
  NAND21X1 U178 ( .B(net83359), .A(n128), .Y(n177) );
  OR3X2 U179 ( .A(n47), .B(n69), .C(net99166), .Y(n219) );
  NAND32X2 U180 ( .B(net99568), .C(net83359), .A(n124), .Y(n200) );
  AND4X1 U181 ( .A(n195), .B(n162), .C(n164), .D(n151), .Y(n135) );
  INVX2 U182 ( .A(n196), .Y(n330) );
  NAND2X1 U183 ( .A(sfrdatai[2]), .B(n48), .Y(n49) );
  INVX1 U184 ( .A(n56), .Y(n258) );
  INVX3 U185 ( .A(n153), .Y(n318) );
  INVX1 U186 ( .A(n189), .Y(n322) );
  INVX1 U187 ( .A(n260), .Y(n50) );
  AO222X1 U188 ( .A(gf0), .B(n28), .C(it1), .D(n347), .E(tl1[2]), .F(n345), 
        .Y(n244) );
  NAND2XL U189 ( .A(md4[0]), .B(n344), .Y(n51) );
  NAND2XL U190 ( .A(t0_tmod[0]), .B(n343), .Y(n53) );
  AND3X1 U191 ( .A(n51), .B(n52), .C(n53), .Y(n167) );
  INVXL U192 ( .A(net89060), .Y(net98374) );
  NAND32X2 U193 ( .B(net101591), .C(net87461), .A(net87439), .Y(n55) );
  OAI221X1 U194 ( .A(n57), .B(n234), .C(n58), .D(n233), .E(n59), .Y(n56) );
  AOI222XL U195 ( .A(md3[2]), .B(n70), .C(md4[2]), .D(n344), .E(th0[2]), .F(
        n341), .Y(n59) );
  INVX1 U196 ( .A(n174), .Y(n68) );
  AND4XL U197 ( .A(n154), .B(n222), .C(n233), .D(n150), .Y(n146) );
  INVX1 U198 ( .A(n47), .Y(n325) );
  NAND4X2 U199 ( .A(n128), .B(net100193), .C(net98374), .D(net99166), .Y(n151)
         );
  BUFXL U200 ( .A(n28), .Y(n60) );
  NAND21X2 U201 ( .B(n131), .A(net98352), .Y(net83264) );
  BUFXL U202 ( .A(n333), .Y(n61) );
  NAND6X1 U203 ( .A(n171), .B(n173), .C(n169), .D(n172), .E(net83318), .F(n170), .Y(n174) );
  NOR2X1 U204 ( .A(n81), .B(n182), .Y(n62) );
  NOR2X1 U205 ( .A(n82), .B(n157), .Y(n63) );
  NOR3X1 U206 ( .A(n62), .B(n63), .C(n64), .Y(n84) );
  INVX1 U207 ( .A(sp[0]), .Y(n81) );
  INVX1 U208 ( .A(dpl[0]), .Y(n82) );
  INVX1 U209 ( .A(port0ff[0]), .Y(n83) );
  AND3X1 U210 ( .A(n84), .B(n86), .C(n85), .Y(n169) );
  INVXL U211 ( .A(n26), .Y(n65) );
  INVXL U212 ( .A(n261), .Y(n332) );
  BUFXL U213 ( .A(n343), .Y(n66) );
  INVX3 U214 ( .A(n188), .Y(n290) );
  NAND2X2 U215 ( .A(sfrdatai[0]), .B(n42), .Y(n67) );
  INVX2 U216 ( .A(n195), .Y(n335) );
  INVX3 U217 ( .A(n162), .Y(n344) );
  NOR3XL U218 ( .A(n69), .B(net99800), .C(n25), .Y(n70) );
  OA21X1 U219 ( .B(net83389), .C(n55), .A(n219), .Y(n130) );
  OR3X2 U220 ( .A(n69), .B(n25), .C(net99800), .Y(n232) );
  NAND21X1 U221 ( .B(n219), .A(i2ccon_o[1]), .Y(n229) );
  OA222X1 U222 ( .A(n71), .B(n234), .C(n76), .D(n232), .E(n164), .F(n77), .Y(
        n166) );
  NAND21X1 U223 ( .B(net100030), .A(net97864), .Y(n234) );
  NAND21X1 U224 ( .B(net100109), .A(n143), .Y(n182) );
  NAND32X1 U225 ( .B(net83359), .C(n25), .A(net97663), .Y(n190) );
  NAND21X2 U226 ( .B(net99404), .A(n87), .Y(n156) );
  NAND2XL U227 ( .A(port0[0]), .B(n333), .Y(n85) );
  NAND2XL U228 ( .A(p), .B(n321), .Y(n86) );
  NOR32X2 U229 ( .B(n218), .C(n217), .A(n216), .Y(n242) );
  INVX1 U230 ( .A(n198), .Y(n88) );
  INVXL U231 ( .A(n158), .Y(n93) );
  INVX3 U232 ( .A(n208), .Y(n334) );
  INVXL U233 ( .A(n156), .Y(n143) );
  INVX2 U234 ( .A(n202), .Y(n336) );
  INVX2 U235 ( .A(n150), .Y(n337) );
  INVXL U236 ( .A(n159), .Y(n350) );
  INVXL U237 ( .A(n123), .Y(n124) );
  AND3X2 U238 ( .A(n240), .B(n239), .C(n238), .Y(n241) );
  NAND32X1 U239 ( .B(n199), .C(n88), .A(n197), .Y(n215) );
  AND4XL U240 ( .A(n187), .B(n186), .C(n185), .D(n89), .Y(n218) );
  AND4X1 U241 ( .A(n237), .B(n236), .C(n235), .D(n90), .Y(n238) );
  AOI22XL U242 ( .A(md4[1]), .B(n344), .C(th0[1]), .D(n341), .Y(n90) );
  AND4X1 U243 ( .A(n231), .B(n230), .C(net83249), .D(n91), .Y(n239) );
  AOI22XL U244 ( .A(i2cadr_o[1]), .B(net97764), .C(md0[1]), .D(net101453), .Y(
        n91) );
  AOI21BXL U245 ( .C(n26), .B(ie0), .A(n175), .Y(n179) );
  AND4X1 U246 ( .A(n157), .B(n182), .C(n202), .D(n144), .Y(n147) );
  NAND6XL U247 ( .A(n188), .B(net83253), .C(n220), .D(n207), .E(n234), .F(
        net83334), .Y(n149) );
  NAND32XL U248 ( .B(net99568), .C(net100030), .A(n124), .Y(n201) );
  AND4X1 U249 ( .A(n190), .B(n206), .C(n232), .D(n153), .Y(n140) );
  INVX1 U250 ( .A(n233), .Y(n342) );
  INVX1 U251 ( .A(n200), .Y(n267) );
  NAND21XL U252 ( .B(n131), .A(net83394), .Y(net83253) );
  NAND21XL U253 ( .B(net100030), .A(n143), .Y(n189) );
  AND4XL U254 ( .A(n200), .B(net83333), .C(n189), .D(n161), .Y(n144) );
  INVX1 U255 ( .A(n190), .Y(n319) );
  INVX1 U256 ( .A(n206), .Y(n305) );
  NAND32XL U257 ( .B(n47), .C(net87609), .A(n122), .Y(n159) );
  OR2X1 U258 ( .A(net97776), .B(n25), .Y(n145) );
  NAND32XL U259 ( .B(net87609), .C(n145), .A(net83365), .Y(n202) );
  NAND32XL U260 ( .B(n145), .C(n27), .A(net87609), .Y(n150) );
  NAND5XL U261 ( .A(net83393), .B(sfraddr[5]), .C(net97663), .D(net101493), 
        .E(net99568), .Y(n207) );
  AND4X1 U262 ( .A(n129), .B(n201), .C(n130), .D(n159), .Y(n142) );
  NAND21XL U263 ( .B(n201), .A(dpc[1]), .Y(n204) );
  NAND42X1 U264 ( .C(n181), .D(n180), .A(n179), .B(n178), .Y(n243) );
  AND4X1 U265 ( .A(n253), .B(n252), .C(n251), .D(n250), .Y(n254) );
  NOR43XL U266 ( .B(n212), .C(n211), .D(n210), .A(n209), .Y(n213) );
  OR4X1 U267 ( .A(n136), .B(n137), .C(n138), .D(n139), .Y(sfrdatao[3]) );
  NAND43X1 U268 ( .B(n266), .C(n265), .D(n264), .A(n263), .Y(n136) );
  NAND43X1 U269 ( .B(n271), .C(n270), .D(n269), .A(n268), .Y(n137) );
  NAND43X1 U270 ( .B(n276), .C(n275), .D(n274), .A(n273), .Y(n139) );
  OR4X1 U271 ( .A(n116), .B(n117), .C(n118), .D(n119), .Y(sfrdatao[4]) );
  NAND43X1 U272 ( .B(n280), .C(n279), .D(n278), .A(n277), .Y(n116) );
  NAND43X1 U273 ( .B(n284), .C(n283), .D(n282), .A(n281), .Y(n117) );
  NAND43X1 U274 ( .B(n289), .C(n288), .D(n287), .A(n286), .Y(n119) );
  OR4X1 U275 ( .A(n94), .B(n95), .C(n96), .D(n97), .Y(sfrdatao[5]) );
  NAND43X1 U276 ( .B(n294), .C(n293), .D(n292), .A(n291), .Y(n94) );
  NAND43X1 U277 ( .B(n299), .C(n298), .D(n297), .A(n296), .Y(n95) );
  NAND43X1 U278 ( .B(n304), .C(n303), .D(n302), .A(n301), .Y(n97) );
  OR4X1 U279 ( .A(n72), .B(n73), .C(n74), .D(n75), .Y(sfrdatao[6]) );
  NAND32X1 U280 ( .B(n308), .C(n307), .A(n306), .Y(n72) );
  NAND32X1 U281 ( .B(n311), .C(n310), .A(n309), .Y(n73) );
  NAND32X1 U282 ( .B(n316), .C(n315), .A(n314), .Y(n75) );
  OR4X1 U283 ( .A(n34), .B(n35), .C(n36), .D(n37), .Y(sfrdatao[7]) );
  NAND32X1 U284 ( .B(n340), .C(n339), .A(n338), .Y(n35) );
  NAND43X1 U285 ( .B(n329), .C(n328), .D(n327), .A(n326), .Y(n34) );
  NAND32X1 U286 ( .B(n356), .C(n355), .A(n354), .Y(n37) );
  AO222X1 U287 ( .A(ien1[0]), .B(n290), .C(ien0[0]), .D(n318), .E(ien2[0]), 
        .F(n29), .Y(n155) );
  AOI221X1 U288 ( .A(ip0[0]), .B(n305), .C(p2[0]), .D(n317), .E(n152), .Y(n171) );
  AO222X1 U289 ( .A(s0con[0]), .B(net83124), .C(th1[0]), .D(n331), .E(
        wdtrel[0]), .F(n334), .Y(n152) );
  AOI22X1 U290 ( .A(md1[0]), .B(n342), .C(dps[0]), .D(n267), .Y(n165) );
  AOI222XL U291 ( .A(tl1[0]), .B(n345), .C(it0), .D(n45), .E(n44), .F(idle), 
        .Y(n168) );
  AND4X1 U292 ( .A(n248), .B(n247), .C(n246), .D(n245), .Y(n257) );
  AOI222XL U293 ( .A(i2cdat_o[2]), .B(n353), .C(i2ccon_o[2]), .D(n352), .E(
        s0relh[2]), .F(net83096), .Y(n248) );
  AOI222XL U294 ( .A(t2con[2]), .B(net83100), .C(i2cadr_o[2]), .D(net97764), 
        .E(md0[2]), .F(net101453), .Y(n246) );
  AOI22XL U295 ( .A(ip1[2]), .B(net83163), .C(iex3), .D(net83162), .Y(n245) );
  AOI222XL U296 ( .A(ckcon[0]), .B(n335), .C(dpc[0]), .D(n295), .E(arcon[0]), 
        .F(n336), .Y(n173) );
  AOI222XL U297 ( .A(b[0]), .B(n330), .C(md5[0]), .D(n337), .E(srstflag), .F(
        net97837), .Y(n172) );
  AOI222XL U298 ( .A(wdtrel[2]), .B(n334), .C(th1[2]), .D(n331), .E(s0con[2]), 
        .F(net83124), .Y(n251) );
  AOI222XL U299 ( .A(b[2]), .B(n330), .C(ckcon[2]), .D(n335), .E(md5[2]), .F(
        n337), .Y(n252) );
  AOI222XL U300 ( .A(s0buf[2]), .B(n324), .C(acc[2]), .D(n349), .E(i2csta_o[2]), .F(n350), .Y(n247) );
  AOI22XL U301 ( .A(ip0[2]), .B(n305), .C(p2[2]), .D(n317), .Y(n250) );
  NAND21XL U302 ( .B(n182), .A(sp[1]), .Y(n187) );
  NAND21XL U303 ( .B(n220), .A(i2cdat_o[1]), .Y(n227) );
  NAND21XL U304 ( .B(net83264), .A(s0relh[1]), .Y(n228) );
  NAND21XL U305 ( .B(n189), .A(dph[1]), .Y(n193) );
  NAND21XL U306 ( .B(n190), .A(s0rell[1]), .Y(n192) );
  NAND21XL U307 ( .B(n188), .A(ien1[1]), .Y(n194) );
  NAND21XL U308 ( .B(net83253), .A(ip1[1]), .Y(n231) );
  NAND21XL U309 ( .B(n233), .A(md1[1]), .Y(n236) );
  NAND21XL U310 ( .B(n234), .A(md2[1]), .Y(n235) );
  AND2X1 U311 ( .A(i2csta_o[1]), .B(n350), .Y(n225) );
  NAND21XL U312 ( .B(n222), .A(s0buf[1]), .Y(n223) );
  NAND21XL U313 ( .B(n221), .A(acc[1]), .Y(n224) );
  AND2XL U314 ( .A(tl1[1]), .B(n345), .Y(n175) );
  AO22XL U315 ( .A(ien0[1]), .B(n318), .C(ien2[1]), .D(n29), .Y(n191) );
  AO22XL U316 ( .A(th1[1]), .B(n331), .C(s0con[1]), .D(net83124), .Y(n209) );
  NAND21XL U317 ( .B(n196), .A(b[1]), .Y(n197) );
  NAND21XL U318 ( .B(n195), .A(ckcon[1]), .Y(n198) );
  NAND21XL U319 ( .B(n206), .A(ip0[1]), .Y(n212) );
  NAND21XL U320 ( .B(n232), .A(md3[1]), .Y(n237) );
  NAND21XL U321 ( .B(n183), .A(f1), .Y(n186) );
  NAND21XL U322 ( .B(n208), .A(wdtrel[1]), .Y(n210) );
  NAND21XL U323 ( .B(n207), .A(p2[1]), .Y(n211) );
  NAND21XL U324 ( .B(n202), .A(arcon[1]), .Y(n203) );
  AOI222XL U325 ( .A(arcon[2]), .B(n336), .C(dps[2]), .D(n267), .E(dpc[2]), 
        .F(n295), .Y(n253) );
  AND2XL U326 ( .A(md5[1]), .B(n337), .Y(n199) );
  AND2XL U327 ( .A(t0_tmod[1]), .B(n343), .Y(n180) );
  NAND21XL U328 ( .B(n200), .A(dps[1]), .Y(n205) );
  AND2XL U329 ( .A(stop), .B(n28), .Y(n181) );
  AOI222XL U330 ( .A(p2sel), .B(n60), .C(sfrdatai[3]), .D(n43), .E(ie1), .F(
        n65), .Y(n272) );
  NAND4X1 U331 ( .A(n98), .B(n99), .C(n100), .D(n272), .Y(n138) );
  AOI22XL U332 ( .A(md1[3]), .B(n342), .C(md2[3]), .D(n351), .Y(n98) );
  AOI222XL U333 ( .A(md3[3]), .B(n70), .C(md4[3]), .D(n344), .E(th0[3]), .F(
        n341), .Y(n99) );
  AOI222XL U334 ( .A(tl0[3]), .B(n346), .C(tl1[3]), .D(n345), .E(t0_tmod[3]), 
        .F(n66), .Y(n100) );
  AO222XL U335 ( .A(th1[3]), .B(n331), .C(b[3]), .D(n330), .E(s0con[3]), .F(
        net83124), .Y(n270) );
  AO222XL U336 ( .A(md0[3]), .B(net101453), .C(i2cadr_o[3]), .D(net97764), .E(
        t2con[3]), .F(net83100), .Y(n275) );
  AO222XL U337 ( .A(dpl[3]), .B(n323), .C(dph[3]), .D(n322), .E(sp[3]), .F(
        n320), .Y(n265) );
  AO222XL U338 ( .A(i2csta_o[3]), .B(n350), .C(acc[3]), .D(n349), .E(s0buf[3]), 
        .F(n324), .Y(n274) );
  AO222XL U339 ( .A(ien2[3]), .B(n29), .C(ien1[3]), .D(n290), .E(s0rell[3]), 
        .F(n319), .Y(n264) );
  AO22XL U340 ( .A(iex4), .B(net83162), .C(ip1[3]), .D(net83163), .Y(n276) );
  AO22XL U341 ( .A(rs[0]), .B(n321), .C(port0ff[3]), .D(n332), .Y(n266) );
  AO22XL U342 ( .A(md5[3]), .B(n337), .C(ckcon[3]), .D(n335), .Y(n269) );
  AOI222XL U343 ( .A(ien0[3]), .B(n318), .C(ip0[3]), .D(n305), .E(p2[3]), .F(
        n317), .Y(n263) );
  AOI222XL U344 ( .A(arcon[3]), .B(n336), .C(dps[3]), .D(n267), .E(dpc[3]), 
        .F(n295), .Y(n268) );
  AOI222XL U345 ( .A(i2cdat_o[3]), .B(n353), .C(i2ccon_o[3]), .D(n352), .E(
        s0relh[3]), .F(net83096), .Y(n273) );
  AOI222XL U346 ( .A(pmw), .B(n60), .C(sfrdatai[4]), .D(n43), .E(t0_tr0), .F(
        n65), .Y(n285) );
  NAND4X1 U347 ( .A(n101), .B(n102), .C(n103), .D(n285), .Y(n118) );
  AOI22XL U348 ( .A(md1[4]), .B(n342), .C(md2[4]), .D(n351), .Y(n101) );
  AOI222XL U349 ( .A(md3[4]), .B(n70), .C(md4[4]), .D(n344), .E(th0[4]), .F(
        n341), .Y(n102) );
  AOI222XL U350 ( .A(tl0[4]), .B(n346), .C(tl1[4]), .D(n345), .E(t1_tmod[0]), 
        .F(n66), .Y(n103) );
  AOI222XL U351 ( .A(isr_tm), .B(n60), .C(sfrdatai[5]), .D(n43), .E(t0_tf0), 
        .F(n65), .Y(n300) );
  NAND4X1 U352 ( .A(n104), .B(n105), .C(n106), .D(n300), .Y(n96) );
  AOI22XL U353 ( .A(md1[5]), .B(n342), .C(md2[5]), .D(n351), .Y(n104) );
  AOI222XL U354 ( .A(md3[5]), .B(n70), .C(md4[5]), .D(n344), .E(th0[5]), .F(
        n341), .Y(n105) );
  AOI222XL U355 ( .A(tl0[5]), .B(n346), .C(tl1[5]), .D(n345), .E(t1_tmod[1]), 
        .F(n66), .Y(n106) );
  NAND4X1 U356 ( .A(n107), .B(n108), .C(n109), .D(n313), .Y(n74) );
  AOI22XL U357 ( .A(md1[6]), .B(n342), .C(th0[6]), .D(n341), .Y(n107) );
  AOI222XL U358 ( .A(md4[6]), .B(n344), .C(t1_tmod[2]), .D(n66), .E(md3[6]), 
        .F(n70), .Y(n108) );
  AOI22XL U359 ( .A(tl0[6]), .B(n346), .C(tl1[6]), .D(n345), .Y(n109) );
  AOI221XL U360 ( .A(wdt_tm), .B(n60), .C(sfrdatai[6]), .D(n43), .E(n312), .Y(
        n313) );
  OA21XL U361 ( .B(t1_tr1), .C(t0_tr1), .A(n65), .Y(n312) );
  AOI222XL U362 ( .A(smod), .B(n60), .C(sfrdatai[7]), .D(n48), .E(tf1_gate), 
        .F(n65), .Y(n348) );
  AO222XL U363 ( .A(md0[5]), .B(net101453), .C(i2cadr_o[5]), .D(net97764), .E(
        t2con[5]), .F(net83100), .Y(n303) );
  AO222XL U364 ( .A(md0[4]), .B(net101453), .C(i2cadr_o[4]), .D(net97764), .E(
        t2con[4]), .F(net83100), .Y(n288) );
  AO222XL U365 ( .A(s0con[4]), .B(net83124), .C(th1[4]), .D(n331), .E(
        wdtrel[4]), .F(n334), .Y(n283) );
  AO222XL U366 ( .A(dph[4]), .B(n322), .C(s0rell[4]), .D(n319), .E(dpl[4]), 
        .F(n323), .Y(n279) );
  AO222XL U367 ( .A(ien1[4]), .B(n290), .C(ien0[4]), .D(n318), .E(ien2[4]), 
        .F(n29), .Y(n278) );
  NAND4X1 U368 ( .A(n110), .B(n111), .C(n112), .D(n348), .Y(n36) );
  AOI22XL U369 ( .A(md1[7]), .B(n342), .C(th0[7]), .D(n341), .Y(n110) );
  AOI222XL U370 ( .A(md4[7]), .B(n344), .C(t1_tmod[3]), .D(n66), .E(md3[7]), 
        .F(n70), .Y(n111) );
  AOI22XL U371 ( .A(tl0[7]), .B(n346), .C(tl1[7]), .D(n345), .Y(n112) );
  AO22XL U372 ( .A(iex6), .B(net83162), .C(ip1[5]), .D(net83163), .Y(n304) );
  AO22XL U373 ( .A(iex5), .B(net83162), .C(ip1[4]), .D(net83163), .Y(n289) );
  AO22XL U374 ( .A(rs[1]), .B(n321), .C(sp[4]), .D(n320), .Y(n280) );
  AO22XL U375 ( .A(b[5]), .B(n330), .C(md5[5]), .D(n337), .Y(n297) );
  AO22XL U376 ( .A(b[4]), .B(n330), .C(md5[4]), .D(n337), .Y(n282) );
  AO22XL U377 ( .A(i2csta_o[5]), .B(n350), .C(acc[5]), .D(n349), .Y(n302) );
  AO22XL U378 ( .A(i2csta_o[4]), .B(n350), .C(acc[4]), .D(n349), .Y(n287) );
  AOI222XL U379 ( .A(i2cdat_o[4]), .B(n353), .C(i2ccon_o[4]), .D(n352), .E(
        s0relh[4]), .F(net83096), .Y(n286) );
  AOI222XL U380 ( .A(ckcon[4]), .B(n335), .C(dpc[4]), .D(n295), .E(arcon[4]), 
        .F(n336), .Y(n281) );
  AO222XL U381 ( .A(s0con[5]), .B(net83124), .C(th1[5]), .D(n331), .E(
        wdtrel[5]), .F(n334), .Y(n298) );
  AO222XL U382 ( .A(dph[5]), .B(n322), .C(s0rell[5]), .D(n319), .E(dpl[5]), 
        .F(n323), .Y(n293) );
  AO222XL U383 ( .A(ien1[5]), .B(n290), .C(ien0[5]), .D(n318), .E(ien2[5]), 
        .F(n29), .Y(n292) );
  AO2222XL U384 ( .A(md0[6]), .B(net101453), .C(i2cadr_o[6]), .D(net97764), 
        .E(md2[6]), .F(n351), .G(t2con[6]), .H(net83100), .Y(n315) );
  AO2222XL U385 ( .A(dpl[6]), .B(n323), .C(dph[6]), .D(n322), .E(ac), .F(n321), 
        .G(sp[6]), .H(n320), .Y(n307) );
  AO22XL U386 ( .A(f0), .B(n321), .C(sp[5]), .D(n320), .Y(n294) );
  AO22XL U387 ( .A(th1[6]), .B(n331), .C(b[6]), .D(n330), .Y(n311) );
  AO22XL U388 ( .A(i2csta_o[6]), .B(n350), .C(acc[6]), .D(n349), .Y(n316) );
  AOI222XL U389 ( .A(p2[5]), .B(n317), .C(s0buf[5]), .D(n324), .E(ip0[5]), .F(
        n305), .Y(n291) );
  AOI222XL U390 ( .A(p2[4]), .B(n317), .C(s0buf[4]), .D(n324), .E(ip0[4]), .F(
        n305), .Y(n277) );
  AOI222XL U391 ( .A(i2cdat_o[5]), .B(n353), .C(i2ccon_o[5]), .D(n352), .E(
        s0relh[5]), .F(net83096), .Y(n301) );
  AOI222XL U392 ( .A(ckcon[5]), .B(n335), .C(dpc[5]), .D(n295), .E(arcon[5]), 
        .F(n336), .Y(n296) );
  AOI222XL U393 ( .A(i2cdat_o[6]), .B(n353), .C(i2ccon_o[6]), .D(n352), .E(
        s0relh[6]), .F(net83096), .Y(n314) );
  AO2222XL U394 ( .A(dpl[7]), .B(n323), .C(dph[7]), .D(n322), .E(c), .F(n321), 
        .G(sp[7]), .H(n320), .Y(n327) );
  AO2222XL U395 ( .A(md0[7]), .B(net101453), .C(i2cadr_o[7]), .D(net97764), 
        .E(md2[7]), .F(n351), .G(t2con[7]), .H(net83100), .Y(n355) );
  AO22XL U396 ( .A(s0rell[7]), .B(n319), .C(ien0[7]), .D(n318), .Y(n328) );
  AO22XL U397 ( .A(th1[7]), .B(n331), .C(b[7]), .D(n330), .Y(n340) );
  AO22XL U398 ( .A(i2csta_o[7]), .B(n350), .C(acc[7]), .D(n349), .Y(n356) );
  AO22XL U399 ( .A(s0rell[6]), .B(n319), .C(ien0[6]), .D(n318), .Y(n308) );
  AOI222XL U400 ( .A(p2[6]), .B(n317), .C(s0buf[6]), .D(n324), .E(ip0wdts), 
        .F(n305), .Y(n306) );
  AOI222XL U401 ( .A(i2cdat_o[7]), .B(n353), .C(i2ccon_o[7]), .D(n352), .E(
        s0relh[7]), .F(net83096), .Y(n354) );
  AOI222XL U402 ( .A(md5[6]), .B(n337), .C(arcon[6]), .D(n336), .E(ckcon[6]), 
        .F(n335), .Y(n309) );
  AOI222XL U403 ( .A(md5[7]), .B(n337), .C(arcon[7]), .D(n336), .E(ckcon[7]), 
        .F(n335), .Y(n338) );
  AND2XL U404 ( .A(p2[7]), .B(n317), .Y(n329) );
  AOI32XL U405 ( .A(bd), .B(n325), .C(n6), .D(s0buf[7]), .E(n324), .Y(n326) );
  BUFX3 U406 ( .A(iex8), .Y(int_vect_8b) );
  BUFX3 U407 ( .A(iex2), .Y(iex2_gate) );
  OR2X1 U408 ( .A(s0con[1]), .B(s0con[0]), .Y(riti0_gate) );
  BUFX3 U409 ( .A(iex9), .Y(int_vect_93) );
  OR2X1 U410 ( .A(t0_tf1), .B(t1_tf1), .Y(tf1_gate) );
  BUFX3 U411 ( .A(iex11), .Y(int_vect_a3) );
  BUFX3 U412 ( .A(iex10), .Y(int_vect_9b) );
  NAND21X2 U413 ( .B(net101202), .A(net97744), .Y(n134) );
  AOI221X1 U414 ( .A(s0rell[0]), .B(n319), .C(dph[0]), .D(n322), .E(n155), .Y(
        n170) );
  INVXL U415 ( .A(n87), .Y(n123) );
  AND4X1 U416 ( .A(n168), .B(n166), .C(n167), .D(n165), .Y(net83322) );
  NAND21XL U417 ( .B(net83252), .A(iex2), .Y(n230) );
  NAND6X1 U418 ( .A(n141), .B(n196), .C(n183), .D(n142), .E(n221), .F(n208), 
        .Y(n148) );
  NAND32XL U419 ( .B(n61), .C(n41), .A(n261), .Y(ext_sfr_sel) );
  AO2222XL U420 ( .A(wdtrel[7]), .B(n334), .C(s0con[7]), .D(net83124), .E(
        port0[7]), .F(n61), .G(port0ff[7]), .H(n332), .Y(n339) );
  AO2222XL U421 ( .A(wdtrel[6]), .B(n334), .C(s0con[6]), .D(net83124), .E(
        port0[6]), .F(n61), .G(port0ff[6]), .H(n332), .Y(n310) );
  AO22XL U422 ( .A(port0[5]), .B(n61), .C(port0ff[5]), .D(n332), .Y(n299) );
  AO22XL U423 ( .A(port0[4]), .B(n61), .C(port0ff[4]), .D(n332), .Y(n284) );
  AO22XL U424 ( .A(port0[3]), .B(n61), .C(wdtrel[3]), .D(n334), .Y(n271) );
  NAND21XL U425 ( .B(n184), .A(port0[1]), .Y(n185) );
  NAND31X4 U426 ( .C(n225), .A(n224), .B(n223), .Y(n226) );
endmodule


module syncneg_a0 ( clk, reset, rsttowdt, rsttosrst, rst, int0, int1, port0i, 
        rxd0i, sdai, int0ff, int1ff, port0ff, t0ff, t1ff, rxd0ff, sdaiff, 
        rsttowdtff, rsttosrstff, rstff, resetff, test_si, test_se );
  input [7:0] port0i;
  output [7:0] port0ff;
  input clk, reset, rsttowdt, rsttosrst, rst, int0, int1, rxd0i, sdai, test_si,
         test_se;
  output int0ff, int1ff, t0ff, t1ff, rxd0ff, sdaiff, rsttowdtff, rsttosrstff,
         rstff, resetff;
  wire   reset_ff1, int0_ff1, int1_ff1, rxd0_ff1, sdai_ff1;
  wire   [7:0] p0_ff1;

  SDFFQX1 reset_ff2_reg ( .D(reset_ff1), .SIN(reset_ff1), .SMC(test_se), .C(
        clk), .Q(resetff) );
  SDFFQX1 rsttosrst_ff1_reg ( .D(rsttosrst), .SIN(rstff), .SMC(test_se), .C(
        clk), .Q(rsttosrstff) );
  SDFFQX1 rsttowdt_ff1_reg ( .D(rsttowdt), .SIN(rsttosrstff), .SMC(test_se), 
        .C(clk), .Q(rsttowdtff) );
  SDFFQX1 int0_ff2_reg ( .D(int0_ff1), .SIN(int0_ff1), .SMC(test_se), .C(clk), 
        .Q(int0ff) );
  SDFFQX1 int1_ff2_reg ( .D(int1_ff1), .SIN(int1_ff1), .SMC(test_se), .C(clk), 
        .Q(int1ff) );
  SDFFQX1 p0_ff2_reg_7_ ( .D(p0_ff1[7]), .SIN(port0ff[6]), .SMC(test_se), .C(
        clk), .Q(port0ff[7]) );
  SDFFQX1 p0_ff2_reg_6_ ( .D(p0_ff1[6]), .SIN(port0ff[5]), .SMC(test_se), .C(
        clk), .Q(port0ff[6]) );
  SDFFQX1 p0_ff2_reg_5_ ( .D(p0_ff1[5]), .SIN(port0ff[4]), .SMC(test_se), .C(
        clk), .Q(port0ff[5]) );
  SDFFQX1 p0_ff2_reg_4_ ( .D(p0_ff1[4]), .SIN(port0ff[3]), .SMC(test_se), .C(
        clk), .Q(port0ff[4]) );
  SDFFQX1 sdai_ff2_reg ( .D(sdai_ff1), .SIN(sdai_ff1), .SMC(test_se), .C(clk), 
        .Q(sdaiff) );
  SDFFQX1 rxd0_ff2_reg ( .D(rxd0_ff1), .SIN(rxd0_ff1), .SMC(test_se), .C(clk), 
        .Q(rxd0ff) );
  SDFFQX1 p0_ff2_reg_3_ ( .D(p0_ff1[3]), .SIN(port0ff[2]), .SMC(test_se), .C(
        clk), .Q(port0ff[3]) );
  SDFFQX1 p0_ff2_reg_1_ ( .D(p0_ff1[1]), .SIN(port0ff[0]), .SMC(test_se), .C(
        clk), .Q(port0ff[1]) );
  SDFFQX1 p0_ff2_reg_0_ ( .D(p0_ff1[0]), .SIN(p0_ff1[7]), .SMC(test_se), .C(
        clk), .Q(port0ff[0]) );
  SDFFQX1 p0_ff2_reg_2_ ( .D(p0_ff1[2]), .SIN(port0ff[1]), .SMC(test_se), .C(
        clk), .Q(port0ff[2]) );
  SDFFQX1 rst_ff1_reg ( .D(rst), .SIN(resetff), .SMC(test_se), .C(clk), .Q(
        rstff) );
  SDFFQX1 int0_ff1_reg ( .D(int0), .SIN(test_si), .SMC(test_se), .C(clk), .Q(
        int0_ff1) );
  SDFFQX1 int1_ff1_reg ( .D(int1), .SIN(int0ff), .SMC(test_se), .C(clk), .Q(
        int1_ff1) );
  SDFFQX1 p0_ff1_reg_6_ ( .D(port0i[6]), .SIN(p0_ff1[5]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[6]) );
  SDFFQX1 p0_ff1_reg_5_ ( .D(port0i[5]), .SIN(p0_ff1[4]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[5]) );
  SDFFQX1 p0_ff1_reg_4_ ( .D(port0i[4]), .SIN(p0_ff1[3]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[4]) );
  SDFFQX1 p0_ff1_reg_3_ ( .D(port0i[3]), .SIN(p0_ff1[2]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[3]) );
  SDFFQX1 p0_ff1_reg_2_ ( .D(port0i[2]), .SIN(p0_ff1[1]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[2]) );
  SDFFQX1 p0_ff1_reg_1_ ( .D(port0i[1]), .SIN(p0_ff1[0]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[1]) );
  SDFFQX1 p0_ff1_reg_0_ ( .D(port0i[0]), .SIN(int1ff), .SMC(test_se), .C(clk), 
        .Q(p0_ff1[0]) );
  SDFFQX1 rxd0_ff1_reg ( .D(rxd0i), .SIN(rsttowdtff), .SMC(test_se), .C(clk), 
        .Q(rxd0_ff1) );
  SDFFQX1 p0_ff1_reg_7_ ( .D(port0i[7]), .SIN(p0_ff1[6]), .SMC(test_se), .C(
        clk), .Q(p0_ff1[7]) );
  SDFFQX1 sdai_ff1_reg ( .D(sdai), .SIN(rxd0ff), .SMC(test_se), .C(clk), .Q(
        sdai_ff1) );
  SDFFQX1 reset_ff1_reg ( .D(reset), .SIN(port0ff[7]), .SMC(test_se), .C(clk), 
        .Q(reset_ff1) );
  INVX1 U5 ( .A(1'b1), .Y(t1ff) );
  INVX1 U7 ( .A(1'b1), .Y(t0ff) );
endmodule


module mcu51_cpu_a0 ( clkcpu, rst, mempsack, memack, memdatai, memaddr, 
        mempsrd, mempswr, memrd, memwr, memaddr_comb, mempsrd_comb, 
        mempswr_comb, memrd_comb, memwr_comb, cpu_hold, cpu_resume, irq, 
        intvect, intcall, retiinstr, newinstr, rmwinstr, waitstaten, ramdatai, 
        sfrdatai, ramsfraddr, ramdatao, ramoe, ramwe, sfroe, sfrwe, sfroe_r, 
        sfrwe_r, sfroe_comb_s, sfrwe_comb_s, pc_o, pc_ini, cs_run, instr, 
        codefetch_s, sfrack, ramsfraddr_comb, ramdatao_comb, ramoe_comb, 
        ramwe_comb, ckcon, pmw, p2sel, gf0, stop, idle, acc, b, rs, c, ac, ov, 
        p, f0, f1, dph, dpl, dps, dpc, p2, sp, test_si, test_so, test_se );
  input [7:0] memdatai;
  output [15:0] memaddr;
  output [15:0] memaddr_comb;
  input [4:0] intvect;
  input [7:0] ramdatai;
  input [7:0] sfrdatai;
  output [7:0] ramsfraddr;
  output [7:0] ramdatao;
  output [15:0] pc_o;
  input [15:0] pc_ini;
  output [7:0] instr;
  output [7:0] ramsfraddr_comb;
  output [7:0] ramdatao_comb;
  output [7:0] ckcon;
  output [7:0] acc;
  output [7:0] b;
  output [1:0] rs;
  output [7:0] dph;
  output [7:0] dpl;
  output [3:0] dps;
  output [5:0] dpc;
  output [7:0] p2;
  output [7:0] sp;
  input clkcpu, rst, mempsack, memack, cpu_hold, cpu_resume, irq, sfrack,
         test_si, test_se;
  output mempsrd, mempswr, memrd, memwr, mempsrd_comb, mempswr_comb,
         memrd_comb, memwr_comb, intcall, retiinstr, newinstr, rmwinstr,
         waitstaten, ramoe, ramwe, sfroe, sfrwe, sfroe_r, sfrwe_r,
         sfroe_comb_s, sfrwe_comb_s, cs_run, codefetch_s, ramoe_comb,
         ramwe_comb, pmw, p2sel, gf0, stop, idle, c, ac, ov, p, f0, f1,
         test_so;
  wire   N343, N344, N345, n2864, finishmul, finishdiv, N370, N371, N372, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491,
         N492, N493, N494, N495, d_hold, idle_r, cpu_resume_fff, stop_r,
         ramsfrwe, N512, N515, N520, pdmode, interrupt, N582, N583, N584, N585,
         N588, N589, N590, phase0_ff, newinstrlock, N670, N671, N672, N673,
         N674, N675, N676, N677, N679, N680, N681, N682, N683, N684, N685,
         N689, N690, accactv, N10562, N10563, N10564, N10565, N10566, N10567,
         N10568, N10569, N10570, N10571, N10572, N10573, N10574, N10575,
         N10576, N10577, N10578, N10581, N10582, N10583, N10584, N10585,
         N10586, N10587, N10588, N10589, N11478, N11479, N11480, N11481,
         N11482, N11483, N11484, N11486, N11487, N11488, N11489, N11491,
         N11498, N11499, N11500, N11501, N11502, N11503, N11504, N11505,
         N12469, N12470, N12472, N12477, N12478, N12479, N12480, N12481,
         N12482, N12483, N12484, N12485, N12486, N12487, N12488, N12489,
         N12490, N12491, N12492, N12493, N12494, N12495, N12496, N12497,
         N12498, N12499, N12500, N12501, N12502, N12503, N12504, N12505,
         N12506, N12507, N12508, N12509, N12510, N12511, N12512, N12513,
         N12514, N12515, N12516, N12517, N12518, N12519, N12520, N12521,
         N12522, N12523, N12524, N12525, N12526, N12527, N12528, N12529,
         N12530, N12531, N12532, N12533, N12534, N12535, N12536, N12537,
         N12538, N12539, N12540, N12541, N12542, N12543, N12544, N12545,
         N12546, N12547, N12548, N12549, N12550, N12551, N12552, N12553,
         N12554, N12555, N12556, N12557, N12558, N12559, N12560, N12561,
         N12562, N12563, N12564, N12566, N12567, N12568, N12569, N12570,
         N12571, N12572, N12573, N12575, N12576, N12577, N12578, N12579,
         N12580, N12581, N12582, N12584, N12585, N12586, N12587, N12588,
         N12589, N12590, N12591, N12593, N12594, N12595, N12596, N12597,
         N12598, N12599, N12600, N12602, N12603, N12604, N12605, N12606,
         N12607, N12608, N12609, N12611, N12612, N12613, N12614, N12615,
         N12616, N12617, N12618, N12620, N12621, N12622, N12623, N12624,
         N12625, N12626, N12627, N12629, N12630, N12631, N12632, N12633,
         N12634, N12635, N12636, N12637, N12644, N12651, N12658, N12665,
         N12672, N12679, N12686, N12690, N12691, N12692, N12693, N12694,
         N12695, N12697, N12698, N12699, N12700, N12701, N12702, N12703,
         N12704, N12705, N12706, N12709, N12710, N12711, N12714, N12715,
         N12716, N12717, N12718, N12719, N12720, N12721, N12722, N12723,
         N12724, N12725, N12726, N12727, N12728, N12729, N12730, N12801,
         N12802, N12803, N12804, N12805, N12806, N12807, N12808, N12824,
         N12825, N12826, N12827, N12828, N12829, N12830, N12831, N12841,
         N12842, N12843, N12844, N12845, N12846, N12847, N12848, N12849,
         N12850, N12851, N12852, N12853, N12854, N12855, N12856, N12905,
         israccess, N12912, waitcnt_1_, waitcnt_0_, N12965, N12966, N12967,
         N12968, N12969, N12970, N12971, N12972, N12974, N12975, N12976,
         N12977, N13014, N13023, N13032, N13041, N13050, N13059, N13068,
         N13077, N13086, N13095, N13104, N13113, N13122, N13131, N13140,
         N13149, N13158, N13167, N13176, N13185, N13194, N13203, N13212,
         N13221, N13230, N13239, N13248, N13257, N13266, N13275, N13284,
         N13293, multemp1_0_, N13324, N13325, N13326, N13327, N13328, N13329,
         N13330, N13331, N13332, N13336, N13337, N13338, N13339, N13340,
         N13341, N13342, N13343, N13345, N13346, N13347, N13348, N13349,
         N13350, N13351, N13352, N13353, N13366, N13367, N13368, N13369,
         N13370, N13371, N13372, N13373, cpu_resume_ff1, N13379, N13380,
         net12372, net12378, net12383, net12388, net12393, net12398, net12403,
         net12408, net12413, net12418, net12423, net12428, net12433, net12438,
         net12443, net12448, net12453, net12458, net12463, net12468, net12473,
         net12478, net12483, net12488, net12493, net12498, net12503, net12508,
         net12513, net12518, net12523, net12528, net12533, net12538, net12543,
         net12548, net12553, net12558, net12563, net12568, net12573, net12578,
         net12583, net12588, net12593, net12598, net12603, net12608, net12613,
         net12618, net12623, net12628, net12633, net12638, net12643, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, N14351, N14350, N14349,
         N14348, N14347, N14346, N14345, N14344, N14343, N14342, N14341,
         N14340, N14339, N14338, N14337, N14336, n2871, n2872, n2870, n2867,
         n2868, n2865, n2869, n2866, n284, n286, n2873, n2446, multemp1_8_,
         multemp1_7_, multemp1_6_, multemp1_5_, multemp1_4_, multemp1_3_,
         multemp1_2_, multemp1_1_, n208, n210, n211, n259, n527, n529, n530,
         n566, n567, n568, n569, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n933, n934,
         n936, n940, n941, n957, n1216, n1225, n1231, n1238, n1239, n1285,
         n1286, n1288, n1293, n1294, n1298, n1299, n1300, n1301, n1302, n1303,
         n1309, n1310, n1311, n1312, n1316, n1317, n1318, n1319, n1320, n1326,
         n1327, n1328, n1329, n1330, n1334, n1335, n1336, n1337, n1350, n1352,
         n1353, n1354, n1355, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1426, n1466, n2069, n2070, n2071, n2072, n2073, n2139, n1, n2,
         n3, n8, n10, n11, n12, n13, n14, n15, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n39, n41, n43, n45, n47, n48, n49, n51, n53, n55, n56, n57, n59, n61,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n122, n123, n124, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n138, n139,
         n140, n141, n142, n143, n145, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n185, n186, n187,
         n188, n189, n191, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n203, n204, n206, n207, n209, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n285, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n418, n419,
         n420, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n528, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n570,
         n571, n572, n573, n574, n575, n576, n577, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n935, n937, n938, n939, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1226, n1227, n1228, n1229, n1230, n1232,
         n1233, n1234, n1235, n1236, n1237, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1287, n1289, n1290, n1291, n1292, n1295, n1296, n1297, n1304, n1305,
         n1306, n1307, n1308, n1313, n1314, n1315, n1321, n1322, n1323, n1324,
         n1325, n1331, n1332, n1333, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1351, n1356, n1357, n1358,
         n1359, n1360, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, SYNOPSYS_UNCONNECTED_1;
  wire   [2:0] state;
  wire   [5:0] phase;
  wire   [15:0] alu_out;
  wire   [15:0] pc_i;
  wire   [7:0] temp;
  wire   [18:0] dec_accop;
  wire   [7:0] dec_cop;
  wire   [9:1] multemp2;
  wire   [7:0] temp2_comb;
  wire   [15:0] dptr_inc;
  wire   [63:0] dpl_reg;
  wire   [63:0] dph_reg;
  wire   [47:0] dpc_tab;
  wire   [255:0] rn_reg;
  wire   [7:0] multempreg;
  wire   [6:0] divtempreg;

  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 clk_gate_finishmul_reg ( .CLK(clkcpu), 
        .EN(N370), .ENCLK(net12372), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 clk_gate_instr_reg ( .CLK(clkcpu), .EN(
        N685), .ENCLK(net12378), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 clk_gate_bitno_reg ( .CLK(clkcpu), .EN(
        N11491), .ENCLK(net12383), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 clk_gate_dph_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N12556), .ENCLK(net12388), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 clk_gate_dph_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N12547), .ENCLK(net12393), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 clk_gate_dph_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N12538), .ENCLK(net12398), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 clk_gate_dph_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N12529), .ENCLK(net12403), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 clk_gate_dph_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N12520), .ENCLK(net12408), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 clk_gate_dph_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N12511), .ENCLK(net12413), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 clk_gate_dph_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N12502), .ENCLK(net12418), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 clk_gate_dph_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N12493), .ENCLK(net12423), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 clk_gate_dpc_tab_reg_7_ ( .CLK(clkcpu), 
        .EN(N12686), .ENCLK(net12428), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 clk_gate_dpc_tab_reg_6_ ( .CLK(clkcpu), 
        .EN(N12679), .ENCLK(net12433), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 clk_gate_dpc_tab_reg_5_ ( .CLK(clkcpu), 
        .EN(N12672), .ENCLK(net12438), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 clk_gate_dpc_tab_reg_4_ ( .CLK(clkcpu), 
        .EN(N12665), .ENCLK(net12443), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 clk_gate_dpc_tab_reg_3_ ( .CLK(clkcpu), 
        .EN(N12658), .ENCLK(net12448), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 clk_gate_dpc_tab_reg_2_ ( .CLK(clkcpu), 
        .EN(N12651), .ENCLK(net12453), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 clk_gate_dpc_tab_reg_1_ ( .CLK(clkcpu), 
        .EN(N12644), .ENCLK(net12458), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 clk_gate_dpc_tab_reg_0_ ( .CLK(clkcpu), 
        .EN(N12637), .ENCLK(net12463), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 clk_gate_temp_reg ( .CLK(clkcpu), .EN(
        N12722), .ENCLK(net12468), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 clk_gate_waitcnt_reg ( .CLK(clkcpu), 
        .EN(N12977), .ENCLK(net12473), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 clk_gate_rn_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N13293), .ENCLK(net12478), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 clk_gate_rn_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N13284), .ENCLK(net12483), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 clk_gate_rn_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N13275), .ENCLK(net12488), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 clk_gate_rn_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N13266), .ENCLK(net12493), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 clk_gate_rn_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N13257), .ENCLK(net12498), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 clk_gate_rn_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N13248), .ENCLK(net12503), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 clk_gate_rn_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N13239), .ENCLK(net12508), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 clk_gate_rn_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N13230), .ENCLK(net12513), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 clk_gate_rn_reg_reg_8_ ( .CLK(clkcpu), 
        .EN(N13221), .ENCLK(net12518), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 clk_gate_rn_reg_reg_9_ ( .CLK(clkcpu), 
        .EN(N13212), .ENCLK(net12523), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 clk_gate_rn_reg_reg_10_ ( .CLK(clkcpu), 
        .EN(N13203), .ENCLK(net12528), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 clk_gate_rn_reg_reg_11_ ( .CLK(clkcpu), 
        .EN(N13194), .ENCLK(net12533), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 clk_gate_rn_reg_reg_12_ ( .CLK(clkcpu), 
        .EN(N13185), .ENCLK(net12538), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 clk_gate_rn_reg_reg_13_ ( .CLK(clkcpu), 
        .EN(N13176), .ENCLK(net12543), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 clk_gate_rn_reg_reg_14_ ( .CLK(clkcpu), 
        .EN(N13167), .ENCLK(net12548), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 clk_gate_rn_reg_reg_15_ ( .CLK(clkcpu), 
        .EN(N13158), .ENCLK(net12553), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 clk_gate_rn_reg_reg_16_ ( .CLK(clkcpu), 
        .EN(N13149), .ENCLK(net12558), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 clk_gate_rn_reg_reg_17_ ( .CLK(clkcpu), 
        .EN(N13140), .ENCLK(net12563), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 clk_gate_rn_reg_reg_18_ ( .CLK(clkcpu), 
        .EN(N13131), .ENCLK(net12568), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 clk_gate_rn_reg_reg_19_ ( .CLK(clkcpu), 
        .EN(N13122), .ENCLK(net12573), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 clk_gate_rn_reg_reg_20_ ( .CLK(clkcpu), 
        .EN(N13113), .ENCLK(net12578), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 clk_gate_rn_reg_reg_21_ ( .CLK(clkcpu), 
        .EN(N13104), .ENCLK(net12583), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 clk_gate_rn_reg_reg_22_ ( .CLK(clkcpu), 
        .EN(N13095), .ENCLK(net12588), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 clk_gate_rn_reg_reg_23_ ( .CLK(clkcpu), 
        .EN(N13086), .ENCLK(net12593), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 clk_gate_rn_reg_reg_24_ ( .CLK(clkcpu), 
        .EN(N13077), .ENCLK(net12598), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 clk_gate_rn_reg_reg_25_ ( .CLK(clkcpu), 
        .EN(N13068), .ENCLK(net12603), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 clk_gate_rn_reg_reg_26_ ( .CLK(clkcpu), 
        .EN(N13059), .ENCLK(net12608), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 clk_gate_rn_reg_reg_27_ ( .CLK(clkcpu), 
        .EN(N13050), .ENCLK(net12613), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 clk_gate_rn_reg_reg_28_ ( .CLK(clkcpu), 
        .EN(N13041), .ENCLK(net12618), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 clk_gate_rn_reg_reg_29_ ( .CLK(clkcpu), 
        .EN(N13032), .ENCLK(net12623), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 clk_gate_rn_reg_reg_30_ ( .CLK(clkcpu), 
        .EN(N13023), .ENCLK(net12628), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 clk_gate_rn_reg_reg_31_ ( .CLK(clkcpu), 
        .EN(N13014), .ENCLK(net12633), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 clk_gate_multempreg_reg ( .CLK(clkcpu), 
        .EN(N13324), .ENCLK(net12638), .TE(test_se) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 clk_gate_divtempreg_reg ( .CLK(clkcpu), 
        .EN(N13366), .ENCLK(net12643), .TE(test_se) );
  mcu51_cpu_a0_DW01_inc_0 add_5525 ( .A({n211, n210, n208, n286, n343, n284, 
        n332, n259}), .SUM({N12808, N12807, N12806, N12805, N12804, N12803, 
        N12802, N12801}) );
  mcu51_cpu_a0_DW01_inc_1 add_5286 ( .A({n2139, n251, n250, n249, n248, n247, 
        n246, n245, n244, n238, n237, n233, n232, n223, n224, n226}), .SUM(
        dptr_inc) );
  mcu51_cpu_a0_DW01_inc_2 r715 ( .A(pc_o), .SUM(pc_i) );
  mcu51_cpu_a0_DW01_add_8 add_5901_aco ( .A({1'b0, multempreg}), .B({1'b0, 
        N14343, N14342, N14341, N14340, N14339, N14338, N14337, N14336}), .CI(
        1'b0), .SUM({multemp1_8_, multemp1_7_, multemp1_6_, multemp1_5_, 
        multemp1_4_, multemp1_3_, multemp1_2_, multemp1_1_, multemp1_0_}), 
        .CO() );
  mcu51_cpu_a0_DW01_add_7 add_5907_aco ( .A({1'b0, multemp1_8_, multemp1_7_, 
        multemp1_6_, multemp1_5_, multemp1_4_, multemp1_3_, multemp1_2_, 
        multemp1_1_}), .B({1'b0, N14351, N14350, N14349, N14348, N14347, 
        N14346, N14345, N14344}), .CI(1'b0), .SUM(multemp2), .CO() );
  mcu51_cpu_a0_DW01_sub_1 sub_5950 ( .A({1'b0, divtempreg, acc[7]}), .B({1'b0, 
        b}), .CI(1'b0), .DIFF({N13343, SYNOPSYS_UNCONNECTED_1, N13342, N13341, 
        N13340, N13339, N13338, N13337, N13336}), .CO() );
  mcu51_cpu_a0_DW01_sub_0 sub_5969 ( .A({1'b0, n335, n322, n323, n314, n316, 
        n315, n312, acc[6]}), .B({1'b0, b}), .CI(1'b0), .DIFF({N13353, N13352, 
        N13351, N13350, N13349, N13348, N13347, N13346, N13345}), .CO() );
  mcu51_cpu_a0_DW01_add_0 add_5586 ( .A({n2826, n2826, n2826, n2826, n2826, 
        n2826, n2826, n2826, N12831, N12830, N12829, N12828, N12827, N12826, 
        N12825, N12824}), .B({N12856, N12855, N12854, N12853, N12852, N12851, 
        N12850, N12849, N12848, N12847, N12846, N12845, N12844, N12843, N12842, 
        N12841}), .CI(1'b0), .SUM(alu_out), .CO() );
  SDFFQX1 pc_reg_5_ ( .D(N485), .SIN(pc_o[4]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[5]) );
  SDFFQX1 pc_reg_6_ ( .D(N486), .SIN(memaddr[5]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[6]) );
  SDFFQX1 pc_reg_7_ ( .D(N487), .SIN(memaddr[6]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[7]) );
  SDFFQX1 pc_reg_8_ ( .D(N488), .SIN(memaddr[7]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[8]) );
  SDFFQX1 pc_reg_9_ ( .D(N489), .SIN(pc_o[8]), .SMC(test_se), .C(net12372), 
        .Q(memaddr[9]) );
  SDFFQX1 pc_reg_10_ ( .D(N490), .SIN(pc_o[9]), .SMC(test_se), .C(net12372), 
        .Q(memaddr[10]) );
  SDFFQX1 pc_reg_11_ ( .D(N491), .SIN(pc_o[10]), .SMC(test_se), .C(net12372), 
        .Q(memaddr[11]) );
  SDFFQX1 pc_reg_12_ ( .D(N492), .SIN(pc_o[11]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[12]) );
  SDFFQX1 pc_reg_13_ ( .D(N493), .SIN(pc_o[12]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[13]) );
  SDFFQX1 pc_reg_14_ ( .D(N494), .SIN(pc_o[13]), .SMC(test_se), .C(net12372), 
        .Q(memaddr[14]) );
  SDFFQX1 pc_reg_15_ ( .D(N495), .SIN(pc_o[14]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[15]) );
  SDFFQX1 cpu_resume_ff1_reg ( .D(N13379), .SIN(ckcon[7]), .SMC(test_se), .C(
        clkcpu), .Q(cpu_resume_ff1) );
  SDFFQX1 newinstrlock_reg ( .D(n1878), .SIN(multempreg[7]), .SMC(test_se), 
        .C(net12372), .Q(newinstrlock) );
  SDFFQX1 phase0_ff_reg ( .D(N689), .SIN(pdmode), .SMC(test_se), .C(net12372), 
        .Q(phase0_ff) );
  SDFFQX1 finishdiv_reg ( .D(N372), .SIN(f1), .SMC(test_se), .C(net12372), .Q(
        finishdiv) );
  SDFFQX1 finishmul_reg ( .D(N371), .SIN(finishdiv), .SMC(test_se), .C(
        net12372), .Q(finishmul) );
  SDFFQX1 multempreg_reg_7_ ( .D(N13332), .SIN(multempreg[6]), .SMC(test_se), 
        .C(net12638), .Q(multempreg[7]) );
  SDFFQX1 multempreg_reg_6_ ( .D(N13331), .SIN(multempreg[5]), .SMC(test_se), 
        .C(net12638), .Q(multempreg[6]) );
  SDFFQX1 multempreg_reg_5_ ( .D(N13330), .SIN(multempreg[4]), .SMC(test_se), 
        .C(net12638), .Q(multempreg[5]) );
  SDFFQX1 multempreg_reg_4_ ( .D(N13329), .SIN(multempreg[3]), .SMC(test_se), 
        .C(net12638), .Q(multempreg[4]) );
  SDFFQX1 multempreg_reg_3_ ( .D(N13328), .SIN(multempreg[2]), .SMC(test_se), 
        .C(net12638), .Q(multempreg[3]) );
  SDFFQX1 multempreg_reg_2_ ( .D(N13327), .SIN(multempreg[1]), .SMC(test_se), 
        .C(net12638), .Q(multempreg[2]) );
  SDFFQX1 pdmode_reg ( .D(n2446), .SIN(pc_o[15]), .SMC(test_se), .C(net12372), 
        .Q(pdmode) );
  SDFFQX1 d_hold_reg ( .D(cpu_hold), .SIN(cpu_resume_fff), .SMC(test_se), .C(
        clkcpu), .Q(d_hold) );
  SDFFQX1 cpu_resume_fff_reg ( .D(N13380), .SIN(cpu_resume_ff1), .SMC(test_se), 
        .C(clkcpu), .Q(cpu_resume_fff) );
  SDFFQX1 p2_reg_reg_6_ ( .D(N12491), .SIN(p2[5]), .SMC(test_se), .C(net12372), 
        .Q(p2[6]) );
  SDFFQX1 p2_reg_reg_7_ ( .D(N12492), .SIN(p2[6]), .SMC(test_se), .C(net12372), 
        .Q(p2[7]) );
  SDFFQX1 f0_reg ( .D(n1882), .SIN(dps[3]), .SMC(test_se), .C(net12372), .Q(f0) );
  SDFFQX1 p2_reg_reg_5_ ( .D(N12490), .SIN(p2[4]), .SMC(test_se), .C(net12372), 
        .Q(p2[5]) );
  SDFFQX1 p2_reg_reg_4_ ( .D(N12489), .SIN(p2[3]), .SMC(test_se), .C(net12372), 
        .Q(p2[4]) );
  SDFFQX1 dpc_tab_reg_5__5_ ( .D(N12692), .SIN(dpc_tab[34]), .SMC(test_se), 
        .C(net12438), .Q(dpc_tab[35]) );
  SDFFQX1 dpc_tab_reg_5__4_ ( .D(n402), .SIN(dpc_tab[33]), .SMC(test_se), .C(
        net12438), .Q(dpc_tab[34]) );
  SDFFQX1 dpc_tab_reg_7__5_ ( .D(N12692), .SIN(dpc_tab[46]), .SMC(test_se), 
        .C(net12428), .Q(dpc_tab[47]) );
  SDFFQX1 dpc_tab_reg_4__5_ ( .D(N12692), .SIN(dpc_tab[28]), .SMC(test_se), 
        .C(net12443), .Q(dpc_tab[29]) );
  SDFFQX1 dpc_tab_reg_4__4_ ( .D(n402), .SIN(dpc_tab[27]), .SMC(test_se), .C(
        net12443), .Q(dpc_tab[28]) );
  SDFFQX1 dpc_tab_reg_6__5_ ( .D(N12692), .SIN(dpc_tab[40]), .SMC(test_se), 
        .C(net12433), .Q(dpc_tab[41]) );
  SDFFQX1 dpc_tab_reg_6__4_ ( .D(N12691), .SIN(dpc_tab[39]), .SMC(test_se), 
        .C(net12433), .Q(dpc_tab[40]) );
  SDFFQX1 dpc_tab_reg_3__5_ ( .D(n2812), .SIN(dpc_tab[22]), .SMC(test_se), .C(
        net12448), .Q(dpc_tab[23]) );
  SDFFQX1 dpc_tab_reg_3__4_ ( .D(N12691), .SIN(dpc_tab[21]), .SMC(test_se), 
        .C(net12448), .Q(dpc_tab[22]) );
  SDFFQX1 dpc_tab_reg_0__5_ ( .D(n2812), .SIN(dpc_tab[4]), .SMC(test_se), .C(
        net12463), .Q(dpc_tab[5]) );
  SDFFQX1 dpc_tab_reg_1__5_ ( .D(n2812), .SIN(dpc_tab[10]), .SMC(test_se), .C(
        net12458), .Q(dpc_tab[11]) );
  SDFFQX1 dpc_tab_reg_1__4_ ( .D(n402), .SIN(dpc_tab[9]), .SMC(test_se), .C(
        net12458), .Q(dpc_tab[10]) );
  SDFFQX1 dpc_tab_reg_2__5_ ( .D(n2812), .SIN(dpc_tab[16]), .SMC(test_se), .C(
        net12453), .Q(dpc_tab[17]) );
  SDFFQX1 dpc_tab_reg_2__4_ ( .D(N12691), .SIN(dpc_tab[15]), .SMC(test_se), 
        .C(net12453), .Q(dpc_tab[16]) );
  SDFFQX1 dpc_tab_reg_7__4_ ( .D(N12691), .SIN(dpc_tab[45]), .SMC(test_se), 
        .C(net12428), .Q(dpc_tab[46]) );
  SDFFQX1 dpc_tab_reg_0__4_ ( .D(n402), .SIN(dpc_tab[3]), .SMC(test_se), .C(
        net12463), .Q(dpc_tab[4]) );
  SDFFQX1 dph_reg_reg_7__7_ ( .D(N12564), .SIN(dph_reg[62]), .SMC(test_se), 
        .C(net12388), .Q(dph_reg[63]) );
  SDFFQX1 dph_reg_reg_4__7_ ( .D(N12537), .SIN(dph_reg[38]), .SMC(test_se), 
        .C(net12403), .Q(dph_reg[39]) );
  SDFFQX1 dph_reg_reg_5__7_ ( .D(N12546), .SIN(dph_reg[46]), .SMC(test_se), 
        .C(net12398), .Q(dph_reg[47]) );
  SDFFQX1 dph_reg_reg_6__7_ ( .D(N12555), .SIN(dph_reg[54]), .SMC(test_se), 
        .C(net12393), .Q(dph_reg[55]) );
  SDFFQX1 dph_reg_reg_3__7_ ( .D(N12528), .SIN(dph_reg[30]), .SMC(test_se), 
        .C(net12408), .Q(dph_reg[31]) );
  SDFFQX1 dph_reg_reg_1__7_ ( .D(N12510), .SIN(dph_reg[14]), .SMC(test_se), 
        .C(net12418), .Q(dph_reg[15]) );
  SDFFQX1 dph_reg_reg_0__7_ ( .D(N12501), .SIN(dph_reg[6]), .SMC(test_se), .C(
        net12423), .Q(dph_reg[7]) );
  SDFFQX1 dph_reg_reg_2__7_ ( .D(N12519), .SIN(dph_reg[22]), .SMC(test_se), 
        .C(net12413), .Q(dph_reg[23]) );
  SDFFQX1 dph_reg_reg_3__6_ ( .D(N12527), .SIN(dph_reg[29]), .SMC(test_se), 
        .C(net12408), .Q(dph_reg[30]) );
  SDFFQX1 dph_reg_reg_7__6_ ( .D(N12563), .SIN(dph_reg[61]), .SMC(test_se), 
        .C(net12388), .Q(dph_reg[62]) );
  SDFFQX1 dph_reg_reg_2__6_ ( .D(N12518), .SIN(dph_reg[21]), .SMC(test_se), 
        .C(net12413), .Q(dph_reg[22]) );
  SDFFQX1 dph_reg_reg_6__6_ ( .D(N12554), .SIN(dph_reg[53]), .SMC(test_se), 
        .C(net12393), .Q(dph_reg[54]) );
  SDFFQX1 dph_reg_reg_3__5_ ( .D(N12526), .SIN(dph_reg[28]), .SMC(test_se), 
        .C(net12408), .Q(dph_reg[29]) );
  SDFFQX1 dph_reg_reg_7__5_ ( .D(N12562), .SIN(dph_reg[60]), .SMC(test_se), 
        .C(net12388), .Q(dph_reg[61]) );
  SDFFQX1 dph_reg_reg_6__5_ ( .D(N12553), .SIN(dph_reg[52]), .SMC(test_se), 
        .C(net12393), .Q(dph_reg[53]) );
  SDFFQX1 dph_reg_reg_5__6_ ( .D(N12545), .SIN(dph_reg[45]), .SMC(test_se), 
        .C(net12398), .Q(dph_reg[46]) );
  SDFFQX1 dph_reg_reg_5__5_ ( .D(N12544), .SIN(dph_reg[44]), .SMC(test_se), 
        .C(net12398), .Q(dph_reg[45]) );
  SDFFQX1 dph_reg_reg_1__6_ ( .D(N12509), .SIN(dph_reg[13]), .SMC(test_se), 
        .C(net12418), .Q(dph_reg[14]) );
  SDFFQX1 dph_reg_reg_1__5_ ( .D(N12508), .SIN(dph_reg[12]), .SMC(test_se), 
        .C(net12418), .Q(dph_reg[13]) );
  SDFFQX1 dph_reg_reg_0__6_ ( .D(N12500), .SIN(dph_reg[5]), .SMC(test_se), .C(
        net12423), .Q(dph_reg[6]) );
  SDFFQX1 dph_reg_reg_0__5_ ( .D(N12499), .SIN(dph_reg[4]), .SMC(test_se), .C(
        net12423), .Q(dph_reg[5]) );
  SDFFQX1 dph_reg_reg_4__6_ ( .D(N12536), .SIN(dph_reg[37]), .SMC(test_se), 
        .C(net12403), .Q(dph_reg[38]) );
  SDFFQX1 dph_reg_reg_4__5_ ( .D(N12535), .SIN(dph_reg[36]), .SMC(test_se), 
        .C(net12403), .Q(dph_reg[37]) );
  SDFFQX1 dph_reg_reg_3__4_ ( .D(N12525), .SIN(dph_reg[27]), .SMC(test_se), 
        .C(net12408), .Q(dph_reg[28]) );
  SDFFQX1 dph_reg_reg_7__4_ ( .D(N12561), .SIN(dph_reg[59]), .SMC(test_se), 
        .C(net12388), .Q(dph_reg[60]) );
  SDFFQX1 dph_reg_reg_2__5_ ( .D(N12517), .SIN(dph_reg[20]), .SMC(test_se), 
        .C(net12413), .Q(dph_reg[21]) );
  SDFFQX1 dph_reg_reg_2__4_ ( .D(N12516), .SIN(dph_reg[19]), .SMC(test_se), 
        .C(net12413), .Q(dph_reg[20]) );
  SDFFQX1 dph_reg_reg_6__4_ ( .D(N12552), .SIN(dph_reg[51]), .SMC(test_se), 
        .C(net12393), .Q(dph_reg[52]) );
  SDFFQX1 dph_reg_reg_5__4_ ( .D(N12543), .SIN(dph_reg[43]), .SMC(test_se), 
        .C(net12398), .Q(dph_reg[44]) );
  SDFFQX1 dph_reg_reg_1__4_ ( .D(N12507), .SIN(dph_reg[11]), .SMC(test_se), 
        .C(net12418), .Q(dph_reg[12]) );
  SDFFQX1 dph_reg_reg_0__4_ ( .D(N12498), .SIN(dph_reg[3]), .SMC(test_se), .C(
        net12423), .Q(dph_reg[4]) );
  SDFFQX1 dph_reg_reg_4__4_ ( .D(N12534), .SIN(dph_reg[35]), .SMC(test_se), 
        .C(net12403), .Q(dph_reg[36]) );
  SDFFQX1 p2sel_s_reg ( .D(N520), .SIN(p2[7]), .SMC(test_se), .C(net12372), 
        .Q(p2sel) );
  SDFFQX1 p2_reg_reg_3_ ( .D(N12488), .SIN(p2[2]), .SMC(test_se), .C(net12372), 
        .Q(p2[3]) );
  SDFFQX1 dpc_tab_reg_5__3_ ( .D(N12690), .SIN(dpc_tab[32]), .SMC(test_se), 
        .C(net12438), .Q(dpc_tab[33]) );
  SDFFQX1 dpc_tab_reg_7__3_ ( .D(N12690), .SIN(dpc_tab[44]), .SMC(test_se), 
        .C(net12428), .Q(dpc_tab[45]) );
  SDFFQX1 dpc_tab_reg_4__3_ ( .D(n390), .SIN(dpc_tab[26]), .SMC(test_se), .C(
        net12443), .Q(dpc_tab[27]) );
  SDFFQX1 dpc_tab_reg_6__3_ ( .D(n390), .SIN(dpc_tab[38]), .SMC(test_se), .C(
        net12433), .Q(dpc_tab[39]) );
  SDFFQX1 dpc_tab_reg_3__3_ ( .D(N12690), .SIN(dpc_tab[20]), .SMC(test_se), 
        .C(net12448), .Q(dpc_tab[21]) );
  SDFFQX1 dpc_tab_reg_0__3_ ( .D(n390), .SIN(dpc_tab[2]), .SMC(test_se), .C(
        net12463), .Q(dpc_tab[3]) );
  SDFFQX1 dpc_tab_reg_1__3_ ( .D(N12690), .SIN(dpc_tab[8]), .SMC(test_se), .C(
        net12458), .Q(dpc_tab[9]) );
  SDFFQX1 dpc_tab_reg_2__3_ ( .D(n390), .SIN(dpc_tab[14]), .SMC(test_se), .C(
        net12453), .Q(dpc_tab[15]) );
  SDFFQX1 dph_reg_reg_3__3_ ( .D(N12524), .SIN(dph_reg[26]), .SMC(test_se), 
        .C(net12408), .Q(dph_reg[27]) );
  SDFFQX1 dph_reg_reg_7__3_ ( .D(N12560), .SIN(dph_reg[58]), .SMC(test_se), 
        .C(net12388), .Q(dph_reg[59]) );
  SDFFQX1 dph_reg_reg_2__3_ ( .D(N12515), .SIN(dph_reg[18]), .SMC(test_se), 
        .C(net12413), .Q(dph_reg[19]) );
  SDFFQX1 dph_reg_reg_6__3_ ( .D(N12551), .SIN(dph_reg[50]), .SMC(test_se), 
        .C(net12393), .Q(dph_reg[51]) );
  SDFFQX1 dph_reg_reg_5__3_ ( .D(N12542), .SIN(dph_reg[42]), .SMC(test_se), 
        .C(net12398), .Q(dph_reg[43]) );
  SDFFQX1 dph_reg_reg_1__3_ ( .D(N12506), .SIN(dph_reg[10]), .SMC(test_se), 
        .C(net12418), .Q(dph_reg[11]) );
  SDFFQX1 dph_reg_reg_0__3_ ( .D(N12497), .SIN(dph_reg[2]), .SMC(test_se), .C(
        net12423), .Q(dph_reg[3]) );
  SDFFQX1 dph_reg_reg_4__3_ ( .D(N12533), .SIN(dph_reg[34]), .SMC(test_se), 
        .C(net12403), .Q(dph_reg[35]) );
  SDFFQX1 dpl_reg_reg_3__7_ ( .D(N12600), .SIN(dpl_reg[30]), .SMC(test_se), 
        .C(net12408), .Q(dpl_reg[31]) );
  SDFFQX1 dpl_reg_reg_7__7_ ( .D(N12636), .SIN(dpl_reg[62]), .SMC(test_se), 
        .C(net12388), .Q(dpl_reg[63]) );
  SDFFQX1 dpl_reg_reg_2__7_ ( .D(N12591), .SIN(dpl_reg[22]), .SMC(test_se), 
        .C(net12413), .Q(dpl_reg[23]) );
  SDFFQX1 dpl_reg_reg_6__7_ ( .D(N12627), .SIN(dpl_reg[54]), .SMC(test_se), 
        .C(net12393), .Q(dpl_reg[55]) );
  SDFFQX1 dpl_reg_reg_5__7_ ( .D(N12618), .SIN(dpl_reg[46]), .SMC(test_se), 
        .C(net12398), .Q(dpl_reg[47]) );
  SDFFQX1 dpl_reg_reg_1__7_ ( .D(N12582), .SIN(dpl_reg[14]), .SMC(test_se), 
        .C(net12418), .Q(dpl_reg[15]) );
  SDFFQX1 dpl_reg_reg_0__7_ ( .D(N12573), .SIN(dpl_reg[6]), .SMC(test_se), .C(
        net12423), .Q(dpl_reg[7]) );
  SDFFQX1 dpl_reg_reg_4__7_ ( .D(N12609), .SIN(dpl_reg[38]), .SMC(test_se), 
        .C(net12403), .Q(dpl_reg[39]) );
  SDFFQX1 ramoe_r_reg ( .D(N11486), .SIN(ramdatao[7]), .SMC(test_se), .C(
        net12372), .Q(ramoe) );
  SDFFQX1 idle_r_reg ( .D(N512), .SIN(gf0), .SMC(test_se), .C(net12372), .Q(
        idle_r) );
  SDFFQX1 stop_r_reg ( .D(N515), .SIN(state[2]), .SMC(test_se), .C(net12372), 
        .Q(stop_r) );
  SDFFQX1 israccess_reg ( .D(N12912), .SIN(interrupt), .SMC(test_se), .C(
        net12372), .Q(israccess) );
  SDFFQX1 phase_reg_5_ ( .D(N684), .SIN(phase[4]), .SMC(test_se), .C(net12372), 
        .Q(phase[5]) );
  SDFFQX1 state_reg_0_ ( .D(N588), .SIN(sp[7]), .SMC(test_se), .C(net12372), 
        .Q(state[0]) );
  SDFFQX1 p_reg ( .D(N12905), .SIN(p2sel), .SMC(test_se), .C(net12372), .Q(p)
         );
  SDFFQX1 state_reg_2_ ( .D(N590), .SIN(state[1]), .SMC(test_se), .C(net12372), 
        .Q(state[2]) );
  SDFFQX1 f1_reg ( .D(n1883), .SIN(f0), .SMC(test_se), .C(net12372), .Q(f1) );
  SDFFQX1 ov_reg_reg ( .D(N12711), .SIN(newinstrlock), .SMC(test_se), .C(
        net12372), .Q(ov) );
  SDFFQX1 state_reg_1_ ( .D(N589), .SIN(state[0]), .SMC(test_se), .C(net12372), 
        .Q(state[1]) );
  SDFFQX1 phase_reg_4_ ( .D(N683), .SIN(phase[3]), .SMC(test_se), .C(net12372), 
        .Q(phase[4]) );
  SDFFQX1 phase_reg_3_ ( .D(N682), .SIN(phase[2]), .SMC(test_se), .C(net12372), 
        .Q(phase[3]) );
  SDFFQX1 p2_reg_reg_1_ ( .D(N12486), .SIN(p2[0]), .SMC(test_se), .C(net12372), 
        .Q(p2[1]) );
  SDFFQX1 stop_s_reg ( .D(n1880), .SIN(stop_r), .SMC(test_se), .C(net12372), 
        .Q(stop) );
  SDFFQX1 gf0_reg ( .D(n1881), .SIN(finishmul), .SMC(test_se), .C(net12372), 
        .Q(gf0) );
  SDFFQX1 dph_reg_reg_3__2_ ( .D(N12523), .SIN(dph_reg[25]), .SMC(test_se), 
        .C(net12408), .Q(dph_reg[26]) );
  SDFFQX1 dph_reg_reg_3__1_ ( .D(N12522), .SIN(dph_reg[24]), .SMC(test_se), 
        .C(net12408), .Q(dph_reg[25]) );
  SDFFQX1 dph_reg_reg_7__2_ ( .D(N12559), .SIN(dph_reg[57]), .SMC(test_se), 
        .C(net12388), .Q(dph_reg[58]) );
  SDFFQX1 dph_reg_reg_7__1_ ( .D(N12558), .SIN(dph_reg[56]), .SMC(test_se), 
        .C(net12388), .Q(dph_reg[57]) );
  SDFFQX1 dph_reg_reg_2__2_ ( .D(N12514), .SIN(dph_reg[17]), .SMC(test_se), 
        .C(net12413), .Q(dph_reg[18]) );
  SDFFQX1 dph_reg_reg_2__1_ ( .D(N12513), .SIN(dph_reg[16]), .SMC(test_se), 
        .C(net12413), .Q(dph_reg[17]) );
  SDFFQX1 dph_reg_reg_6__2_ ( .D(N12550), .SIN(dph_reg[49]), .SMC(test_se), 
        .C(net12393), .Q(dph_reg[50]) );
  SDFFQX1 dph_reg_reg_6__1_ ( .D(N12549), .SIN(dph_reg[48]), .SMC(test_se), 
        .C(net12393), .Q(dph_reg[49]) );
  SDFFQX1 dph_reg_reg_6__0_ ( .D(N12548), .SIN(dph_reg[47]), .SMC(test_se), 
        .C(net12393), .Q(dph_reg[48]) );
  SDFFQX1 dpc_tab_reg_3__1_ ( .D(n401), .SIN(dpc_tab[18]), .SMC(test_se), .C(
        net12448), .Q(dpc_tab[19]) );
  SDFFQX1 dpc_tab_reg_7__1_ ( .D(n2828), .SIN(dpc_tab[42]), .SMC(test_se), .C(
        net12428), .Q(dpc_tab[43]) );
  SDFFQX1 dpc_tab_reg_0__1_ ( .D(n401), .SIN(dpc_tab[0]), .SMC(test_se), .C(
        net12463), .Q(dpc_tab[1]) );
  SDFFQX1 dpc_tab_reg_4__1_ ( .D(n401), .SIN(dpc_tab[24]), .SMC(test_se), .C(
        net12443), .Q(dpc_tab[25]) );
  SDFFQX1 dpc_tab_reg_1__1_ ( .D(n401), .SIN(dpc_tab[6]), .SMC(test_se), .C(
        net12458), .Q(dpc_tab[7]) );
  SDFFQX1 dpc_tab_reg_5__1_ ( .D(n401), .SIN(dpc_tab[30]), .SMC(test_se), .C(
        net12438), .Q(dpc_tab[31]) );
  SDFFQX1 dpc_tab_reg_2__1_ ( .D(n401), .SIN(dpc_tab[12]), .SMC(test_se), .C(
        net12453), .Q(dpc_tab[13]) );
  SDFFQX1 dpc_tab_reg_6__1_ ( .D(n2828), .SIN(dpc_tab[36]), .SMC(test_se), .C(
        net12433), .Q(dpc_tab[37]) );
  SDFFQX1 p2_reg_reg_2_ ( .D(N12487), .SIN(p2[1]), .SMC(test_se), .C(net12372), 
        .Q(p2[2]) );
  SDFFQX1 p2_reg_reg_0_ ( .D(N12485), .SIN(ov), .SMC(test_se), .C(net12372), 
        .Q(p2[0]) );
  SDFFQX1 dpl_reg_reg_5__6_ ( .D(N12617), .SIN(dpl_reg[45]), .SMC(test_se), 
        .C(net12398), .Q(dpl_reg[46]) );
  SDFFQX1 dph_reg_reg_5__2_ ( .D(N12541), .SIN(dph_reg[41]), .SMC(test_se), 
        .C(net12398), .Q(dph_reg[42]) );
  SDFFQX1 dph_reg_reg_5__1_ ( .D(N12540), .SIN(dph_reg[40]), .SMC(test_se), 
        .C(net12398), .Q(dph_reg[41]) );
  SDFFQX1 dph_reg_reg_5__0_ ( .D(N12539), .SIN(dph_reg[39]), .SMC(test_se), 
        .C(net12398), .Q(dph_reg[40]) );
  SDFFQX1 dpl_reg_reg_1__6_ ( .D(N12581), .SIN(dpl_reg[13]), .SMC(test_se), 
        .C(net12418), .Q(dpl_reg[14]) );
  SDFFQX1 dph_reg_reg_1__2_ ( .D(N12505), .SIN(dph_reg[9]), .SMC(test_se), .C(
        net12418), .Q(dph_reg[10]) );
  SDFFQX1 dph_reg_reg_1__1_ ( .D(N12504), .SIN(dph_reg[8]), .SMC(test_se), .C(
        net12418), .Q(dph_reg[9]) );
  SDFFQX1 dpl_reg_reg_0__6_ ( .D(N12572), .SIN(dpl_reg[5]), .SMC(test_se), .C(
        net12423), .Q(dpl_reg[6]) );
  SDFFQX1 dph_reg_reg_0__2_ ( .D(N12496), .SIN(dph_reg[1]), .SMC(test_se), .C(
        net12423), .Q(dph_reg[2]) );
  SDFFQX1 dph_reg_reg_0__1_ ( .D(N12495), .SIN(dph_reg[0]), .SMC(test_se), .C(
        net12423), .Q(dph_reg[1]) );
  SDFFQX1 dpl_reg_reg_4__6_ ( .D(N12608), .SIN(dpl_reg[37]), .SMC(test_se), 
        .C(net12403), .Q(dpl_reg[38]) );
  SDFFQX1 dph_reg_reg_4__2_ ( .D(N12532), .SIN(dph_reg[33]), .SMC(test_se), 
        .C(net12403), .Q(dph_reg[34]) );
  SDFFQX1 dph_reg_reg_4__1_ ( .D(N12531), .SIN(dph_reg[32]), .SMC(test_se), 
        .C(net12403), .Q(dph_reg[33]) );
  SDFFQX1 sfrwe_r_reg ( .D(N11489), .SIN(sfroe_r), .SMC(test_se), .C(net12372), 
        .Q(sfrwe_r) );
  SDFFQX1 sfroe_r_reg ( .D(N11488), .SIN(rs[1]), .SMC(test_se), .C(net12372), 
        .Q(sfroe_r) );
  SDFFQX1 memwr_s_reg ( .D(N585), .SIN(memrd), .SMC(test_se), .C(net12372), 
        .Q(memwr) );
  SDFFQX1 rn_reg_reg_28__6_ ( .D(n415), .SIN(rn_reg[29]), .SMC(test_se), .C(
        net12618), .Q(rn_reg[30]) );
  SDFFQX1 rn_reg_reg_12__6_ ( .D(n414), .SIN(rn_reg[157]), .SMC(test_se), .C(
        net12538), .Q(rn_reg[158]) );
  SDFFQX1 rn_reg_reg_6__6_ ( .D(n414), .SIN(rn_reg[205]), .SMC(test_se), .C(
        net12508), .Q(rn_reg[206]) );
  SDFFQX1 rn_reg_reg_22__6_ ( .D(n413), .SIN(rn_reg[77]), .SMC(test_se), .C(
        net12588), .Q(rn_reg[78]) );
  SDFFQX1 dec_cop_reg_0_ ( .D(N10582), .SIN(dec_accop[18]), .SMC(test_se), .C(
        net12372), .Q(dec_cop[0]) );
  SDFFQX1 rmwinstr_reg ( .D(N690), .SIN(ramwe), .SMC(test_se), .C(net12372), 
        .Q(rmwinstr) );
  SDFFQX1 dpl_reg_reg_3__6_ ( .D(N12599), .SIN(dpl_reg[29]), .SMC(test_se), 
        .C(net12408), .Q(dpl_reg[30]) );
  SDFFQX1 dpl_reg_reg_7__6_ ( .D(N12635), .SIN(dpl_reg[61]), .SMC(test_se), 
        .C(net12388), .Q(dpl_reg[62]) );
  SDFFQX1 dpl_reg_reg_2__6_ ( .D(N12590), .SIN(dpl_reg[21]), .SMC(test_se), 
        .C(net12413), .Q(dpl_reg[22]) );
  SDFFQX1 dpl_reg_reg_6__6_ ( .D(N12626), .SIN(dpl_reg[53]), .SMC(test_se), 
        .C(net12393), .Q(dpl_reg[54]) );
  SDFFQX1 dph_reg_reg_2__0_ ( .D(N12512), .SIN(dph_reg[15]), .SMC(test_se), 
        .C(net12413), .Q(dph_reg[16]) );
  SDFFQX1 dpc_tab_reg_3__2_ ( .D(n394), .SIN(dpc_tab[19]), .SMC(test_se), .C(
        net12448), .Q(dpc_tab[20]) );
  SDFFQX1 dpc_tab_reg_3__0_ ( .D(n409), .SIN(dpc_tab[17]), .SMC(test_se), .C(
        net12448), .Q(dpc_tab[18]) );
  SDFFQX1 dpc_tab_reg_7__0_ ( .D(n409), .SIN(dpc_tab[41]), .SMC(test_se), .C(
        net12428), .Q(dpc_tab[42]) );
  SDFFQX1 dpc_tab_reg_0__2_ ( .D(n394), .SIN(dpc_tab[1]), .SMC(test_se), .C(
        net12463), .Q(dpc_tab[2]) );
  SDFFQX1 dpc_tab_reg_0__0_ ( .D(n409), .SIN(divtempreg[6]), .SMC(test_se), 
        .C(net12463), .Q(dpc_tab[0]) );
  SDFFQX1 dpc_tab_reg_4__0_ ( .D(n409), .SIN(dpc_tab[23]), .SMC(test_se), .C(
        net12443), .Q(dpc_tab[24]) );
  SDFFQX1 dpc_tab_reg_1__2_ ( .D(n395), .SIN(dpc_tab[7]), .SMC(test_se), .C(
        net12458), .Q(dpc_tab[8]) );
  SDFFQX1 dpc_tab_reg_1__0_ ( .D(n409), .SIN(dpc_tab[5]), .SMC(test_se), .C(
        net12458), .Q(dpc_tab[6]) );
  SDFFQX1 dpc_tab_reg_5__0_ ( .D(n409), .SIN(dpc_tab[29]), .SMC(test_se), .C(
        net12438), .Q(dpc_tab[30]) );
  SDFFQX1 dpc_tab_reg_2__2_ ( .D(n394), .SIN(dpc_tab[13]), .SMC(test_se), .C(
        net12453), .Q(dpc_tab[14]) );
  SDFFQX1 dpc_tab_reg_2__0_ ( .D(n409), .SIN(dpc_tab[11]), .SMC(test_se), .C(
        net12453), .Q(dpc_tab[12]) );
  SDFFQX1 dpc_tab_reg_6__0_ ( .D(n409), .SIN(dpc_tab[35]), .SMC(test_se), .C(
        net12433), .Q(dpc_tab[36]) );
  SDFFQX1 dpl_reg_reg_3__5_ ( .D(N12598), .SIN(dpl_reg[28]), .SMC(test_se), 
        .C(net12408), .Q(dpl_reg[29]) );
  SDFFQX1 dpl_reg_reg_7__5_ ( .D(N12634), .SIN(dpl_reg[60]), .SMC(test_se), 
        .C(net12388), .Q(dpl_reg[61]) );
  SDFFQX1 dph_reg_reg_7__0_ ( .D(N12557), .SIN(dph_reg[55]), .SMC(test_se), 
        .C(net12388), .Q(dph_reg[56]) );
  SDFFQX1 dph_reg_reg_3__0_ ( .D(N12521), .SIN(dph_reg[23]), .SMC(test_se), 
        .C(net12408), .Q(dph_reg[24]) );
  SDFFQX1 dpl_reg_reg_2__5_ ( .D(N12589), .SIN(dpl_reg[20]), .SMC(test_se), 
        .C(net12413), .Q(dpl_reg[21]) );
  SDFFQX1 dpl_reg_reg_6__5_ ( .D(N12625), .SIN(dpl_reg[52]), .SMC(test_se), 
        .C(net12393), .Q(dpl_reg[53]) );
  SDFFQX1 rn_reg_reg_7__6_ ( .D(n414), .SIN(rn_reg[197]), .SMC(test_se), .C(
        net12513), .Q(rn_reg[198]) );
  SDFFQX1 rn_reg_reg_3__6_ ( .D(n413), .SIN(rn_reg[229]), .SMC(test_se), .C(
        net12493), .Q(rn_reg[230]) );
  SDFFQX1 rn_reg_reg_19__6_ ( .D(n415), .SIN(rn_reg[101]), .SMC(test_se), .C(
        net12573), .Q(rn_reg[102]) );
  SDFFQX1 rn_reg_reg_23__6_ ( .D(n413), .SIN(rn_reg[69]), .SMC(test_se), .C(
        net12593), .Q(rn_reg[70]) );
  SDFFQX1 dpc_tab_reg_7__2_ ( .D(n394), .SIN(dpc_tab[43]), .SMC(test_se), .C(
        net12428), .Q(dpc_tab[44]) );
  SDFFQX1 rn_reg_reg_27__6_ ( .D(n415), .SIN(rn_reg[37]), .SMC(test_se), .C(
        net12613), .Q(rn_reg[38]) );
  SDFFQX1 rn_reg_reg_31__6_ ( .D(n413), .SIN(rn_reg[5]), .SMC(test_se), .C(
        net12633), .Q(rn_reg[6]) );
  SDFFQX1 rn_reg_reg_11__6_ ( .D(n414), .SIN(rn_reg[165]), .SMC(test_se), .C(
        net12533), .Q(rn_reg[166]) );
  SDFFQX1 rn_reg_reg_15__6_ ( .D(n415), .SIN(rn_reg[133]), .SMC(test_se), .C(
        net12553), .Q(rn_reg[134]) );
  SDFFQX1 rn_reg_reg_0__6_ ( .D(n413), .SIN(rn_reg[253]), .SMC(test_se), .C(
        net12478), .Q(rn_reg[254]) );
  SDFFQX1 rn_reg_reg_4__6_ ( .D(n414), .SIN(rn_reg[221]), .SMC(test_se), .C(
        net12498), .Q(rn_reg[222]) );
  SDFFQX1 rn_reg_reg_16__6_ ( .D(n415), .SIN(rn_reg[125]), .SMC(test_se), .C(
        net12558), .Q(rn_reg[126]) );
  SDFFQX1 rn_reg_reg_20__6_ ( .D(n415), .SIN(rn_reg[93]), .SMC(test_se), .C(
        net12578), .Q(rn_reg[94]) );
  SDFFQX1 dpc_tab_reg_4__2_ ( .D(n394), .SIN(dpc_tab[25]), .SMC(test_se), .C(
        net12443), .Q(dpc_tab[26]) );
  SDFFQX1 rn_reg_reg_24__6_ ( .D(n413), .SIN(rn_reg[61]), .SMC(test_se), .C(
        net12598), .Q(rn_reg[62]) );
  SDFFQX1 rn_reg_reg_8__6_ ( .D(n414), .SIN(rn_reg[189]), .SMC(test_se), .C(
        net12518), .Q(rn_reg[190]) );
  SDFFQX1 rn_reg_reg_5__6_ ( .D(n414), .SIN(rn_reg[213]), .SMC(test_se), .C(
        net12503), .Q(rn_reg[214]) );
  SDFFQX1 rn_reg_reg_1__6_ ( .D(n413), .SIN(rn_reg[245]), .SMC(test_se), .C(
        net12483), .Q(rn_reg[246]) );
  SDFFQX1 rn_reg_reg_17__6_ ( .D(n415), .SIN(rn_reg[117]), .SMC(test_se), .C(
        net12563), .Q(rn_reg[118]) );
  SDFFQX1 rn_reg_reg_21__6_ ( .D(n415), .SIN(rn_reg[85]), .SMC(test_se), .C(
        net12583), .Q(rn_reg[86]) );
  SDFFQX1 dpc_tab_reg_5__2_ ( .D(n394), .SIN(dpc_tab[31]), .SMC(test_se), .C(
        net12438), .Q(dpc_tab[32]) );
  SDFFQX1 rn_reg_reg_25__6_ ( .D(n2833), .SIN(rn_reg[53]), .SMC(test_se), .C(
        net12603), .Q(rn_reg[54]) );
  SDFFQX1 rn_reg_reg_29__6_ ( .D(n2833), .SIN(rn_reg[21]), .SMC(test_se), .C(
        net12623), .Q(rn_reg[22]) );
  SDFFQX1 rn_reg_reg_9__6_ ( .D(n414), .SIN(rn_reg[181]), .SMC(test_se), .C(
        net12523), .Q(rn_reg[182]) );
  SDFFQX1 rn_reg_reg_13__6_ ( .D(n414), .SIN(rn_reg[149]), .SMC(test_se), .C(
        net12543), .Q(rn_reg[150]) );
  SDFFQX1 rn_reg_reg_2__6_ ( .D(n413), .SIN(rn_reg[237]), .SMC(test_se), .C(
        net12488), .Q(rn_reg[238]) );
  SDFFQX1 rn_reg_reg_18__6_ ( .D(n415), .SIN(rn_reg[109]), .SMC(test_se), .C(
        net12568), .Q(rn_reg[110]) );
  SDFFQX1 dpc_tab_reg_6__2_ ( .D(n394), .SIN(dpc_tab[37]), .SMC(test_se), .C(
        net12433), .Q(dpc_tab[38]) );
  SDFFQX1 dpl_reg_reg_3__4_ ( .D(N12597), .SIN(dpl_reg[27]), .SMC(test_se), 
        .C(net12408), .Q(dpl_reg[28]) );
  SDFFQX1 dpl_reg_reg_7__4_ ( .D(N12633), .SIN(dpl_reg[59]), .SMC(test_se), 
        .C(net12388), .Q(dpl_reg[60]) );
  SDFFQX1 dpl_reg_reg_6__4_ ( .D(N12624), .SIN(dpl_reg[51]), .SMC(test_se), 
        .C(net12393), .Q(dpl_reg[52]) );
  SDFFQX1 ckcon_r_reg_6_ ( .D(N12971), .SIN(ckcon[5]), .SMC(test_se), .C(
        net12372), .Q(ckcon[6]) );
  SDFFQX1 dpl_reg_reg_5__5_ ( .D(N12616), .SIN(dpl_reg[44]), .SMC(test_se), 
        .C(net12398), .Q(dpl_reg[45]) );
  SDFFQX1 dpl_reg_reg_5__4_ ( .D(N12615), .SIN(dpl_reg[43]), .SMC(test_se), 
        .C(net12398), .Q(dpl_reg[44]) );
  SDFFQX1 dpl_reg_reg_1__5_ ( .D(N12580), .SIN(dpl_reg[12]), .SMC(test_se), 
        .C(net12418), .Q(dpl_reg[13]) );
  SDFFQX1 dph_reg_reg_1__0_ ( .D(N12503), .SIN(dph_reg[7]), .SMC(test_se), .C(
        net12418), .Q(dph_reg[8]) );
  SDFFQX1 dpl_reg_reg_1__4_ ( .D(N12579), .SIN(dpl_reg[11]), .SMC(test_se), 
        .C(net12418), .Q(dpl_reg[12]) );
  SDFFQX1 dpl_reg_reg_0__5_ ( .D(N12571), .SIN(dpl_reg[4]), .SMC(test_se), .C(
        net12423), .Q(dpl_reg[5]) );
  SDFFQX1 dph_reg_reg_0__0_ ( .D(N12494), .SIN(dpc_tab[47]), .SMC(test_se), 
        .C(net12423), .Q(dph_reg[0]) );
  SDFFQX1 dpl_reg_reg_0__4_ ( .D(N12570), .SIN(dpl_reg[3]), .SMC(test_se), .C(
        net12423), .Q(dpl_reg[4]) );
  SDFFQX1 dpl_reg_reg_4__5_ ( .D(N12607), .SIN(dpl_reg[36]), .SMC(test_se), 
        .C(net12403), .Q(dpl_reg[37]) );
  SDFFQX1 dph_reg_reg_4__0_ ( .D(N12530), .SIN(dph_reg[31]), .SMC(test_se), 
        .C(net12403), .Q(dph_reg[32]) );
  SDFFQX1 dpl_reg_reg_4__4_ ( .D(N12606), .SIN(dpl_reg[35]), .SMC(test_se), 
        .C(net12403), .Q(dpl_reg[36]) );
  SDFFQX1 idle_s_reg ( .D(n1879), .SIN(idle_r), .SMC(test_se), .C(net12372), 
        .Q(idle) );
  SDFFQX1 ckcon_r_reg_0_ ( .D(N12965), .SIN(c), .SMC(test_se), .C(net12372), 
        .Q(ckcon[0]) );
  SDFFQX1 ckcon_r_reg_2_ ( .D(N12967), .SIN(ckcon[1]), .SMC(test_se), .C(
        net12372), .Q(ckcon[2]) );
  SDFFQX1 ckcon_r_reg_1_ ( .D(N12966), .SIN(ckcon[0]), .SMC(test_se), .C(
        net12372), .Q(ckcon[1]) );
  SDFFQX1 waitcnt_reg_2_ ( .D(N12976), .SIN(waitcnt_1_), .SMC(test_se), .C(
        net12473), .Q(test_so) );
  SDFFQX1 mempsrd_r_reg ( .D(N582), .SIN(israccess), .SMC(test_se), .C(
        net12372), .Q(mempsrd) );
  SDFFQX1 mempswr_s_reg ( .D(N583), .SIN(mempsrd), .SMC(test_se), .C(net12372), 
        .Q(n2864) );
  SDFFQX1 rn_reg_reg_28__5_ ( .D(n387), .SIN(rn_reg[28]), .SMC(test_se), .C(
        net12618), .Q(rn_reg[29]) );
  SDFFQX1 rn_reg_reg_28__2_ ( .D(n2813), .SIN(rn_reg[25]), .SMC(test_se), .C(
        net12618), .Q(rn_reg[26]) );
  SDFFQX1 rn_reg_reg_12__5_ ( .D(n388), .SIN(rn_reg[156]), .SMC(test_se), .C(
        net12538), .Q(rn_reg[157]) );
  SDFFQX1 rn_reg_reg_12__2_ ( .D(n396), .SIN(rn_reg[153]), .SMC(test_se), .C(
        net12538), .Q(rn_reg[154]) );
  SDFFQX1 rn_reg_reg_28__7_ ( .D(n2831), .SIN(rn_reg[30]), .SMC(test_se), .C(
        net12618), .Q(rn_reg[31]) );
  SDFFQX1 rn_reg_reg_12__7_ ( .D(n407), .SIN(rn_reg[158]), .SMC(test_se), .C(
        net12538), .Q(rn_reg[159]) );
  SDFFQX1 rn_reg_reg_6__2_ ( .D(n396), .SIN(rn_reg[201]), .SMC(test_se), .C(
        net12508), .Q(rn_reg[202]) );
  SDFFQX1 rn_reg_reg_6__5_ ( .D(n389), .SIN(rn_reg[204]), .SMC(test_se), .C(
        net12508), .Q(rn_reg[205]) );
  SDFFQX1 rn_reg_reg_22__5_ ( .D(n2812), .SIN(rn_reg[76]), .SMC(test_se), .C(
        net12588), .Q(rn_reg[77]) );
  SDFFQX1 rn_reg_reg_22__2_ ( .D(n395), .SIN(rn_reg[73]), .SMC(test_se), .C(
        net12588), .Q(rn_reg[74]) );
  SDFFQX1 rn_reg_reg_6__7_ ( .D(n407), .SIN(rn_reg[206]), .SMC(test_se), .C(
        net12508), .Q(rn_reg[207]) );
  SDFFQX1 rn_reg_reg_22__7_ ( .D(n406), .SIN(rn_reg[78]), .SMC(test_se), .C(
        net12588), .Q(rn_reg[79]) );
  SDFFQX1 multempreg_reg_0_ ( .D(N13325), .SIN(memwr), .SMC(test_se), .C(
        net12638), .Q(multempreg[0]) );
  SDFFQX1 multempreg_reg_1_ ( .D(N13326), .SIN(multempreg[0]), .SMC(test_se), 
        .C(net12638), .Q(multempreg[1]) );
  SDFFQX1 dec_cop_reg_2_ ( .D(N10584), .SIN(dec_cop[1]), .SMC(test_se), .C(
        net12372), .Q(dec_cop[2]) );
  SDFFQX1 rn_reg_reg_26__6_ ( .D(n2833), .SIN(rn_reg[45]), .SMC(test_se), .C(
        net12608), .Q(rn_reg[46]) );
  SDFFQX1 rn_reg_reg_30__6_ ( .D(n413), .SIN(rn_reg[13]), .SMC(test_se), .C(
        net12628), .Q(rn_reg[14]) );
  SDFFQX1 rn_reg_reg_10__6_ ( .D(n414), .SIN(rn_reg[173]), .SMC(test_se), .C(
        net12528), .Q(rn_reg[174]) );
  SDFFQX1 rn_reg_reg_14__6_ ( .D(n415), .SIN(rn_reg[141]), .SMC(test_se), .C(
        net12548), .Q(rn_reg[142]) );
  SDFFQX1 dpl_reg_reg_2__4_ ( .D(N12588), .SIN(dpl_reg[19]), .SMC(test_se), 
        .C(net12413), .Q(dpl_reg[20]) );
  SDFFQX1 rn_reg_reg_3__2_ ( .D(n396), .SIN(rn_reg[225]), .SMC(test_se), .C(
        net12493), .Q(rn_reg[226]) );
  SDFFQX1 rn_reg_reg_7__2_ ( .D(n396), .SIN(rn_reg[193]), .SMC(test_se), .C(
        net12513), .Q(rn_reg[194]) );
  SDFFQX1 rn_reg_reg_3__5_ ( .D(n389), .SIN(rn_reg[228]), .SMC(test_se), .C(
        net12493), .Q(rn_reg[229]) );
  SDFFQX1 rn_reg_reg_19__5_ ( .D(n387), .SIN(rn_reg[100]), .SMC(test_se), .C(
        net12573), .Q(rn_reg[101]) );
  SDFFQX1 rn_reg_reg_19__2_ ( .D(n397), .SIN(rn_reg[97]), .SMC(test_se), .C(
        net12573), .Q(rn_reg[98]) );
  SDFFQX1 rn_reg_reg_23__2_ ( .D(n395), .SIN(rn_reg[65]), .SMC(test_se), .C(
        net12593), .Q(rn_reg[66]) );
  SDFFQX1 rn_reg_reg_27__5_ ( .D(n387), .SIN(rn_reg[36]), .SMC(test_se), .C(
        net12613), .Q(rn_reg[37]) );
  SDFFQX1 rn_reg_reg_27__2_ ( .D(n397), .SIN(rn_reg[33]), .SMC(test_se), .C(
        net12613), .Q(rn_reg[34]) );
  SDFFQX1 rn_reg_reg_31__5_ ( .D(n2812), .SIN(rn_reg[4]), .SMC(test_se), .C(
        net12633), .Q(rn_reg[5]) );
  SDFFQX1 rn_reg_reg_31__2_ ( .D(n395), .SIN(rn_reg[1]), .SMC(test_se), .C(
        net12633), .Q(rn_reg[2]) );
  SDFFQX1 rn_reg_reg_11__5_ ( .D(n388), .SIN(rn_reg[164]), .SMC(test_se), .C(
        net12533), .Q(rn_reg[165]) );
  SDFFQX1 rn_reg_reg_11__2_ ( .D(n396), .SIN(rn_reg[161]), .SMC(test_se), .C(
        net12533), .Q(rn_reg[162]) );
  SDFFQX1 rn_reg_reg_15__5_ ( .D(n388), .SIN(rn_reg[132]), .SMC(test_se), .C(
        net12553), .Q(rn_reg[133]) );
  SDFFQX1 rn_reg_reg_15__2_ ( .D(n397), .SIN(rn_reg[129]), .SMC(test_se), .C(
        net12553), .Q(rn_reg[130]) );
  SDFFQX1 rn_reg_reg_0__2_ ( .D(n395), .SIN(rn_reg[249]), .SMC(test_se), .C(
        net12478), .Q(rn_reg[250]) );
  SDFFQX1 rn_reg_reg_4__2_ ( .D(n396), .SIN(rn_reg[217]), .SMC(test_se), .C(
        net12498), .Q(rn_reg[218]) );
  SDFFQX1 rn_reg_reg_0__5_ ( .D(n389), .SIN(rn_reg[252]), .SMC(test_se), .C(
        net12478), .Q(rn_reg[253]) );
  SDFFQX1 rn_reg_reg_4__5_ ( .D(n389), .SIN(rn_reg[220]), .SMC(test_se), .C(
        net12498), .Q(rn_reg[221]) );
  SDFFQX1 rn_reg_reg_16__5_ ( .D(n388), .SIN(rn_reg[124]), .SMC(test_se), .C(
        net12558), .Q(rn_reg[125]) );
  SDFFQX1 rn_reg_reg_16__2_ ( .D(n397), .SIN(rn_reg[121]), .SMC(test_se), .C(
        net12558), .Q(rn_reg[122]) );
  SDFFQX1 rn_reg_reg_20__2_ ( .D(n397), .SIN(rn_reg[89]), .SMC(test_se), .C(
        net12578), .Q(rn_reg[90]) );
  SDFFQX1 rn_reg_reg_24__5_ ( .D(n2812), .SIN(rn_reg[60]), .SMC(test_se), .C(
        net12598), .Q(rn_reg[61]) );
  SDFFQX1 rn_reg_reg_24__2_ ( .D(n395), .SIN(rn_reg[57]), .SMC(test_se), .C(
        net12598), .Q(rn_reg[58]) );
  SDFFQX1 rn_reg_reg_8__5_ ( .D(n388), .SIN(rn_reg[188]), .SMC(test_se), .C(
        net12518), .Q(rn_reg[189]) );
  SDFFQX1 rn_reg_reg_8__2_ ( .D(n396), .SIN(rn_reg[185]), .SMC(test_se), .C(
        net12518), .Q(rn_reg[186]) );
  SDFFQX1 rn_reg_reg_1__2_ ( .D(n395), .SIN(rn_reg[241]), .SMC(test_se), .C(
        net12483), .Q(rn_reg[242]) );
  SDFFQX1 rn_reg_reg_5__2_ ( .D(n396), .SIN(rn_reg[209]), .SMC(test_se), .C(
        net12503), .Q(rn_reg[210]) );
  SDFFQX1 rn_reg_reg_1__5_ ( .D(n389), .SIN(rn_reg[244]), .SMC(test_se), .C(
        net12483), .Q(rn_reg[245]) );
  SDFFQX1 rn_reg_reg_17__5_ ( .D(n388), .SIN(rn_reg[116]), .SMC(test_se), .C(
        net12563), .Q(rn_reg[117]) );
  SDFFQX1 rn_reg_reg_17__2_ ( .D(n397), .SIN(rn_reg[113]), .SMC(test_se), .C(
        net12563), .Q(rn_reg[114]) );
  SDFFQX1 rn_reg_reg_21__2_ ( .D(n397), .SIN(rn_reg[81]), .SMC(test_se), .C(
        net12583), .Q(rn_reg[82]) );
  SDFFQX1 rn_reg_reg_25__5_ ( .D(n389), .SIN(rn_reg[52]), .SMC(test_se), .C(
        net12603), .Q(rn_reg[53]) );
  SDFFQX1 rn_reg_reg_25__2_ ( .D(n394), .SIN(rn_reg[49]), .SMC(test_se), .C(
        net12603), .Q(rn_reg[50]) );
  SDFFQX1 rn_reg_reg_29__5_ ( .D(n387), .SIN(rn_reg[20]), .SMC(test_se), .C(
        net12623), .Q(rn_reg[21]) );
  SDFFQX1 rn_reg_reg_29__2_ ( .D(n2813), .SIN(rn_reg[17]), .SMC(test_se), .C(
        net12623), .Q(rn_reg[18]) );
  SDFFQX1 rn_reg_reg_9__5_ ( .D(n388), .SIN(rn_reg[180]), .SMC(test_se), .C(
        net12523), .Q(rn_reg[181]) );
  SDFFQX1 rn_reg_reg_9__2_ ( .D(n396), .SIN(rn_reg[177]), .SMC(test_se), .C(
        net12523), .Q(rn_reg[178]) );
  SDFFQX1 rn_reg_reg_13__5_ ( .D(n388), .SIN(rn_reg[148]), .SMC(test_se), .C(
        net12543), .Q(rn_reg[149]) );
  SDFFQX1 rn_reg_reg_13__2_ ( .D(n397), .SIN(rn_reg[145]), .SMC(test_se), .C(
        net12543), .Q(rn_reg[146]) );
  SDFFQX1 rn_reg_reg_2__2_ ( .D(n395), .SIN(rn_reg[233]), .SMC(test_se), .C(
        net12488), .Q(rn_reg[234]) );
  SDFFQX1 rn_reg_reg_2__5_ ( .D(n389), .SIN(rn_reg[236]), .SMC(test_se), .C(
        net12488), .Q(rn_reg[237]) );
  SDFFQX1 rn_reg_reg_18__5_ ( .D(n387), .SIN(rn_reg[108]), .SMC(test_se), .C(
        net12568), .Q(rn_reg[109]) );
  SDFFQX1 rn_reg_reg_18__2_ ( .D(n397), .SIN(rn_reg[105]), .SMC(test_se), .C(
        net12568), .Q(rn_reg[106]) );
  SDFFQX1 dpl_reg_reg_3__3_ ( .D(N12596), .SIN(dpl_reg[26]), .SMC(test_se), 
        .C(net12408), .Q(dpl_reg[27]) );
  SDFFQX1 dpl_reg_reg_7__3_ ( .D(N12632), .SIN(dpl_reg[58]), .SMC(test_se), 
        .C(net12388), .Q(dpl_reg[59]) );
  SDFFQX1 dpl_reg_reg_2__3_ ( .D(N12587), .SIN(dpl_reg[18]), .SMC(test_se), 
        .C(net12413), .Q(dpl_reg[19]) );
  SDFFQX1 dpl_reg_reg_6__3_ ( .D(N12623), .SIN(dpl_reg[50]), .SMC(test_se), 
        .C(net12393), .Q(dpl_reg[51]) );
  SDFFQX1 rn_reg_reg_3__7_ ( .D(n406), .SIN(rn_reg[230]), .SMC(test_se), .C(
        net12493), .Q(rn_reg[231]) );
  SDFFQX1 rn_reg_reg_7__7_ ( .D(n407), .SIN(rn_reg[198]), .SMC(test_se), .C(
        net12513), .Q(rn_reg[199]) );
  SDFFQX1 rn_reg_reg_19__7_ ( .D(n408), .SIN(rn_reg[102]), .SMC(test_se), .C(
        net12573), .Q(rn_reg[103]) );
  SDFFQX1 rn_reg_reg_23__7_ ( .D(n406), .SIN(rn_reg[70]), .SMC(test_se), .C(
        net12593), .Q(rn_reg[71]) );
  SDFFQX1 rn_reg_reg_27__7_ ( .D(n408), .SIN(rn_reg[38]), .SMC(test_se), .C(
        net12613), .Q(rn_reg[39]) );
  SDFFQX1 rn_reg_reg_31__7_ ( .D(n406), .SIN(rn_reg[6]), .SMC(test_se), .C(
        net12633), .Q(rn_reg[7]) );
  SDFFQX1 rn_reg_reg_11__7_ ( .D(n407), .SIN(rn_reg[166]), .SMC(test_se), .C(
        net12533), .Q(rn_reg[167]) );
  SDFFQX1 rn_reg_reg_15__7_ ( .D(n408), .SIN(rn_reg[134]), .SMC(test_se), .C(
        net12553), .Q(rn_reg[135]) );
  SDFFQX1 rn_reg_reg_0__7_ ( .D(n406), .SIN(rn_reg[254]), .SMC(test_se), .C(
        net12478), .Q(rn_reg[255]) );
  SDFFQX1 rn_reg_reg_4__7_ ( .D(n407), .SIN(rn_reg[222]), .SMC(test_se), .C(
        net12498), .Q(rn_reg[223]) );
  SDFFQX1 rn_reg_reg_16__7_ ( .D(n408), .SIN(rn_reg[126]), .SMC(test_se), .C(
        net12558), .Q(rn_reg[127]) );
  SDFFQX1 rn_reg_reg_20__7_ ( .D(n408), .SIN(rn_reg[94]), .SMC(test_se), .C(
        net12578), .Q(rn_reg[95]) );
  SDFFQX1 rn_reg_reg_24__7_ ( .D(n406), .SIN(rn_reg[62]), .SMC(test_se), .C(
        net12598), .Q(rn_reg[63]) );
  SDFFQX1 rn_reg_reg_8__7_ ( .D(n407), .SIN(rn_reg[190]), .SMC(test_se), .C(
        net12518), .Q(rn_reg[191]) );
  SDFFQX1 rn_reg_reg_1__7_ ( .D(n406), .SIN(rn_reg[246]), .SMC(test_se), .C(
        net12483), .Q(rn_reg[247]) );
  SDFFQX1 rn_reg_reg_5__7_ ( .D(n407), .SIN(rn_reg[214]), .SMC(test_se), .C(
        net12503), .Q(rn_reg[215]) );
  SDFFQX1 rn_reg_reg_17__7_ ( .D(n408), .SIN(rn_reg[118]), .SMC(test_se), .C(
        net12563), .Q(rn_reg[119]) );
  SDFFQX1 rn_reg_reg_21__7_ ( .D(n408), .SIN(rn_reg[86]), .SMC(test_se), .C(
        net12583), .Q(rn_reg[87]) );
  SDFFQX1 rn_reg_reg_25__7_ ( .D(n2831), .SIN(rn_reg[54]), .SMC(test_se), .C(
        net12603), .Q(rn_reg[55]) );
  SDFFQX1 rn_reg_reg_29__7_ ( .D(n2831), .SIN(rn_reg[22]), .SMC(test_se), .C(
        net12623), .Q(rn_reg[23]) );
  SDFFQX1 rn_reg_reg_9__7_ ( .D(n407), .SIN(rn_reg[182]), .SMC(test_se), .C(
        net12523), .Q(rn_reg[183]) );
  SDFFQX1 rn_reg_reg_13__7_ ( .D(n407), .SIN(rn_reg[150]), .SMC(test_se), .C(
        net12543), .Q(rn_reg[151]) );
  SDFFQX1 rn_reg_reg_2__7_ ( .D(n406), .SIN(rn_reg[238]), .SMC(test_se), .C(
        net12488), .Q(rn_reg[239]) );
  SDFFQX1 rn_reg_reg_18__7_ ( .D(n408), .SIN(rn_reg[110]), .SMC(test_se), .C(
        net12568), .Q(rn_reg[111]) );
  SDFFQX1 rn_reg_reg_26__7_ ( .D(n408), .SIN(rn_reg[46]), .SMC(test_se), .C(
        net12608), .Q(rn_reg[47]) );
  SDFFQX1 rn_reg_reg_30__7_ ( .D(n406), .SIN(rn_reg[14]), .SMC(test_se), .C(
        net12628), .Q(rn_reg[15]) );
  SDFFQX1 rn_reg_reg_10__7_ ( .D(n407), .SIN(rn_reg[174]), .SMC(test_se), .C(
        net12528), .Q(rn_reg[175]) );
  SDFFQX1 rn_reg_reg_14__7_ ( .D(n408), .SIN(rn_reg[142]), .SMC(test_se), .C(
        net12548), .Q(rn_reg[143]) );
  SDFFQX1 dpl_reg_reg_5__3_ ( .D(N12614), .SIN(dpl_reg[42]), .SMC(test_se), 
        .C(net12398), .Q(dpl_reg[43]) );
  SDFFQX1 dpl_reg_reg_5__2_ ( .D(N12613), .SIN(dpl_reg[41]), .SMC(test_se), 
        .C(net12398), .Q(dpl_reg[42]) );
  SDFFQX1 sp_reg_reg_6_ ( .D(N12703), .SIN(sp[5]), .SMC(test_se), .C(net12372), 
        .Q(sp[6]) );
  SDFFQX1 sp_reg_reg_7_ ( .D(N12704), .SIN(sp[6]), .SMC(test_se), .C(net12372), 
        .Q(sp[7]) );
  SDFFQX1 dpl_reg_reg_1__3_ ( .D(N12578), .SIN(dpl_reg[10]), .SMC(test_se), 
        .C(net12418), .Q(dpl_reg[11]) );
  SDFFQX1 dpl_reg_reg_1__2_ ( .D(N12577), .SIN(dpl_reg[9]), .SMC(test_se), .C(
        net12418), .Q(dpl_reg[10]) );
  SDFFQX1 dpl_reg_reg_0__3_ ( .D(N12569), .SIN(dpl_reg[2]), .SMC(test_se), .C(
        net12423), .Q(dpl_reg[3]) );
  SDFFQX1 dpl_reg_reg_0__2_ ( .D(N12568), .SIN(dpl_reg[1]), .SMC(test_se), .C(
        net12423), .Q(dpl_reg[2]) );
  SDFFQX1 dpl_reg_reg_4__3_ ( .D(N12605), .SIN(dpl_reg[34]), .SMC(test_se), 
        .C(net12403), .Q(dpl_reg[35]) );
  SDFFQX1 dpl_reg_reg_4__2_ ( .D(N12604), .SIN(dpl_reg[33]), .SMC(test_se), 
        .C(net12403), .Q(dpl_reg[34]) );
  SDFFQX1 waitcnt_reg_1_ ( .D(N12975), .SIN(waitcnt_0_), .SMC(test_se), .C(
        net12473), .Q(waitcnt_1_) );
  SDFFQX1 ckcon_r_reg_5_ ( .D(N12970), .SIN(ckcon[4]), .SMC(test_se), .C(
        net12372), .Q(ckcon[5]) );
  SDFFQX1 memrd_s_reg ( .D(N584), .SIN(n2864), .SMC(test_se), .C(net12372), 
        .Q(memrd) );
  SDFFQX1 dec_cop_reg_1_ ( .D(N10583), .SIN(dec_cop[0]), .SMC(test_se), .C(
        net12372), .Q(dec_cop[1]) );
  SDFFQX1 ckcon_r_reg_4_ ( .D(N12969), .SIN(ckcon[3]), .SMC(test_se), .C(
        net12372), .Q(ckcon[4]) );
  SDFFQX1 ramdatao_r_reg_6_ ( .D(N11504), .SIN(ramdatao[5]), .SMC(test_se), 
        .C(net12372), .Q(ramdatao[6]) );
  SDFFQX1 rn_reg_reg_28__4_ ( .D(n405), .SIN(rn_reg[27]), .SMC(test_se), .C(
        net12618), .Q(rn_reg[28]) );
  SDFFQX1 rn_reg_reg_28__3_ ( .D(n393), .SIN(rn_reg[26]), .SMC(test_se), .C(
        net12618), .Q(rn_reg[27]) );
  SDFFQX1 rn_reg_reg_28__1_ ( .D(n398), .SIN(rn_reg[24]), .SMC(test_se), .C(
        net12618), .Q(rn_reg[25]) );
  SDFFQX1 rn_reg_reg_28__0_ ( .D(n412), .SIN(rn_reg[39]), .SMC(test_se), .C(
        net12618), .Q(rn_reg[24]) );
  SDFFQX1 rn_reg_reg_12__4_ ( .D(n404), .SIN(rn_reg[155]), .SMC(test_se), .C(
        net12538), .Q(rn_reg[156]) );
  SDFFQX1 rn_reg_reg_12__3_ ( .D(n392), .SIN(rn_reg[154]), .SMC(test_se), .C(
        net12538), .Q(rn_reg[155]) );
  SDFFQX1 rn_reg_reg_12__1_ ( .D(n399), .SIN(rn_reg[152]), .SMC(test_se), .C(
        net12538), .Q(rn_reg[153]) );
  SDFFQX1 rn_reg_reg_12__0_ ( .D(n411), .SIN(rn_reg[167]), .SMC(test_se), .C(
        net12538), .Q(rn_reg[152]) );
  SDFFQX1 rn_reg_reg_6__3_ ( .D(n391), .SIN(rn_reg[202]), .SMC(test_se), .C(
        net12508), .Q(rn_reg[203]) );
  SDFFQX1 rn_reg_reg_6__1_ ( .D(n400), .SIN(rn_reg[200]), .SMC(test_se), .C(
        net12508), .Q(rn_reg[201]) );
  SDFFQX1 rn_reg_reg_6__0_ ( .D(n410), .SIN(rn_reg[215]), .SMC(test_se), .C(
        net12508), .Q(rn_reg[200]) );
  SDFFQX1 rn_reg_reg_6__4_ ( .D(n403), .SIN(rn_reg[203]), .SMC(test_se), .C(
        net12508), .Q(rn_reg[204]) );
  SDFFQX1 rn_reg_reg_22__4_ ( .D(n403), .SIN(rn_reg[75]), .SMC(test_se), .C(
        net12588), .Q(rn_reg[76]) );
  SDFFQX1 rn_reg_reg_22__3_ ( .D(n391), .SIN(rn_reg[74]), .SMC(test_se), .C(
        net12588), .Q(rn_reg[75]) );
  SDFFQX1 rn_reg_reg_22__1_ ( .D(n401), .SIN(rn_reg[72]), .SMC(test_se), .C(
        net12588), .Q(rn_reg[73]) );
  SDFFQX1 rn_reg_reg_22__0_ ( .D(n412), .SIN(rn_reg[87]), .SMC(test_se), .C(
        net12588), .Q(rn_reg[72]) );
  SDFFQX1 rn_reg_reg_7__5_ ( .D(n389), .SIN(rn_reg[196]), .SMC(test_se), .C(
        net12513), .Q(rn_reg[197]) );
  SDFFQX1 rn_reg_reg_23__5_ ( .D(n389), .SIN(rn_reg[68]), .SMC(test_se), .C(
        net12593), .Q(rn_reg[69]) );
  SDFFQX1 rn_reg_reg_20__5_ ( .D(n387), .SIN(rn_reg[92]), .SMC(test_se), .C(
        net12578), .Q(rn_reg[93]) );
  SDFFQX1 rn_reg_reg_5__5_ ( .D(n389), .SIN(rn_reg[212]), .SMC(test_se), .C(
        net12503), .Q(rn_reg[213]) );
  SDFFQX1 rn_reg_reg_21__5_ ( .D(n387), .SIN(rn_reg[84]), .SMC(test_se), .C(
        net12583), .Q(rn_reg[85]) );
  SDFFQX1 rn_reg_reg_26__5_ ( .D(n387), .SIN(rn_reg[44]), .SMC(test_se), .C(
        net12608), .Q(rn_reg[45]) );
  SDFFQX1 rn_reg_reg_26__2_ ( .D(n395), .SIN(rn_reg[41]), .SMC(test_se), .C(
        net12608), .Q(rn_reg[42]) );
  SDFFQX1 rn_reg_reg_30__5_ ( .D(n2812), .SIN(rn_reg[12]), .SMC(test_se), .C(
        net12628), .Q(rn_reg[13]) );
  SDFFQX1 rn_reg_reg_30__2_ ( .D(n395), .SIN(rn_reg[9]), .SMC(test_se), .C(
        net12628), .Q(rn_reg[10]) );
  SDFFQX1 rn_reg_reg_10__5_ ( .D(n388), .SIN(rn_reg[172]), .SMC(test_se), .C(
        net12528), .Q(rn_reg[173]) );
  SDFFQX1 rn_reg_reg_10__2_ ( .D(n396), .SIN(rn_reg[169]), .SMC(test_se), .C(
        net12528), .Q(rn_reg[170]) );
  SDFFQX1 rn_reg_reg_14__5_ ( .D(n388), .SIN(rn_reg[140]), .SMC(test_se), .C(
        net12548), .Q(rn_reg[141]) );
  SDFFQX1 rn_reg_reg_14__2_ ( .D(n397), .SIN(rn_reg[137]), .SMC(test_se), .C(
        net12548), .Q(rn_reg[138]) );
  SDFFQX1 dpl_reg_reg_3__2_ ( .D(N12595), .SIN(dpl_reg[25]), .SMC(test_se), 
        .C(net12408), .Q(dpl_reg[26]) );
  SDFFQX1 dpl_reg_reg_3__1_ ( .D(N12594), .SIN(dpl_reg[24]), .SMC(test_se), 
        .C(net12408), .Q(dpl_reg[25]) );
  SDFFQX1 dpl_reg_reg_7__2_ ( .D(N12631), .SIN(dpl_reg[57]), .SMC(test_se), 
        .C(net12388), .Q(dpl_reg[58]) );
  SDFFQX1 dpl_reg_reg_2__2_ ( .D(N12586), .SIN(dpl_reg[17]), .SMC(test_se), 
        .C(net12413), .Q(dpl_reg[18]) );
  SDFFQX1 dpl_reg_reg_2__1_ ( .D(N12585), .SIN(dpl_reg[16]), .SMC(test_se), 
        .C(net12413), .Q(dpl_reg[17]) );
  SDFFQX1 dpl_reg_reg_6__2_ ( .D(N12622), .SIN(dpl_reg[49]), .SMC(test_se), 
        .C(net12393), .Q(dpl_reg[50]) );
  SDFFQX1 rn_reg_reg_3__3_ ( .D(n391), .SIN(rn_reg[226]), .SMC(test_se), .C(
        net12493), .Q(rn_reg[227]) );
  SDFFQX1 rn_reg_reg_3__1_ ( .D(n400), .SIN(rn_reg[224]), .SMC(test_se), .C(
        net12493), .Q(rn_reg[225]) );
  SDFFQX1 rn_reg_reg_3__0_ ( .D(n410), .SIN(rn_reg[239]), .SMC(test_se), .C(
        net12493), .Q(rn_reg[224]) );
  SDFFQX1 rn_reg_reg_7__3_ ( .D(n391), .SIN(rn_reg[194]), .SMC(test_se), .C(
        net12513), .Q(rn_reg[195]) );
  SDFFQX1 rn_reg_reg_7__1_ ( .D(n400), .SIN(rn_reg[192]), .SMC(test_se), .C(
        net12513), .Q(rn_reg[193]) );
  SDFFQX1 rn_reg_reg_7__0_ ( .D(n411), .SIN(rn_reg[207]), .SMC(test_se), .C(
        net12513), .Q(rn_reg[192]) );
  SDFFQX1 rn_reg_reg_7__4_ ( .D(n403), .SIN(rn_reg[195]), .SMC(test_se), .C(
        net12513), .Q(rn_reg[196]) );
  SDFFQX1 rn_reg_reg_3__4_ ( .D(n403), .SIN(rn_reg[227]), .SMC(test_se), .C(
        net12493), .Q(rn_reg[228]) );
  SDFFQX1 rn_reg_reg_19__4_ ( .D(n405), .SIN(rn_reg[99]), .SMC(test_se), .C(
        net12573), .Q(rn_reg[100]) );
  SDFFQX1 rn_reg_reg_19__3_ ( .D(n393), .SIN(rn_reg[98]), .SMC(test_se), .C(
        net12573), .Q(rn_reg[99]) );
  SDFFQX1 rn_reg_reg_19__1_ ( .D(n398), .SIN(rn_reg[96]), .SMC(test_se), .C(
        net12573), .Q(rn_reg[97]) );
  SDFFQX1 rn_reg_reg_19__0_ ( .D(n412), .SIN(rn_reg[111]), .SMC(test_se), .C(
        net12573), .Q(rn_reg[96]) );
  SDFFQX1 rn_reg_reg_23__4_ ( .D(n403), .SIN(rn_reg[67]), .SMC(test_se), .C(
        net12593), .Q(rn_reg[68]) );
  SDFFQX1 rn_reg_reg_23__3_ ( .D(n391), .SIN(rn_reg[66]), .SMC(test_se), .C(
        net12593), .Q(rn_reg[67]) );
  SDFFQX1 rn_reg_reg_23__1_ ( .D(n400), .SIN(rn_reg[64]), .SMC(test_se), .C(
        net12593), .Q(rn_reg[65]) );
  SDFFQX1 rn_reg_reg_23__0_ ( .D(n410), .SIN(rn_reg[79]), .SMC(test_se), .C(
        net12593), .Q(rn_reg[64]) );
  SDFFQX1 rn_reg_reg_27__4_ ( .D(n405), .SIN(rn_reg[35]), .SMC(test_se), .C(
        net12613), .Q(rn_reg[36]) );
  SDFFQX1 rn_reg_reg_27__3_ ( .D(n393), .SIN(rn_reg[34]), .SMC(test_se), .C(
        net12613), .Q(rn_reg[35]) );
  SDFFQX1 rn_reg_reg_27__1_ ( .D(n398), .SIN(rn_reg[32]), .SMC(test_se), .C(
        net12613), .Q(rn_reg[33]) );
  SDFFQX1 rn_reg_reg_27__0_ ( .D(n412), .SIN(rn_reg[47]), .SMC(test_se), .C(
        net12613), .Q(rn_reg[32]) );
  SDFFQX1 rn_reg_reg_31__4_ ( .D(n402), .SIN(rn_reg[3]), .SMC(test_se), .C(
        net12633), .Q(rn_reg[4]) );
  SDFFQX1 rn_reg_reg_31__3_ ( .D(n390), .SIN(rn_reg[2]), .SMC(test_se), .C(
        net12633), .Q(rn_reg[3]) );
  SDFFQX1 rn_reg_reg_31__1_ ( .D(n401), .SIN(rn_reg[0]), .SMC(test_se), .C(
        net12633), .Q(rn_reg[1]) );
  SDFFQX1 rn_reg_reg_31__0_ ( .D(n410), .SIN(rn_reg[15]), .SMC(test_se), .C(
        net12633), .Q(rn_reg[0]) );
  SDFFQX1 rn_reg_reg_11__4_ ( .D(n404), .SIN(rn_reg[163]), .SMC(test_se), .C(
        net12533), .Q(rn_reg[164]) );
  SDFFQX1 rn_reg_reg_11__3_ ( .D(n392), .SIN(rn_reg[162]), .SMC(test_se), .C(
        net12533), .Q(rn_reg[163]) );
  SDFFQX1 rn_reg_reg_11__1_ ( .D(n399), .SIN(rn_reg[160]), .SMC(test_se), .C(
        net12533), .Q(rn_reg[161]) );
  SDFFQX1 rn_reg_reg_11__0_ ( .D(n411), .SIN(rn_reg[175]), .SMC(test_se), .C(
        net12533), .Q(rn_reg[160]) );
  SDFFQX1 rn_reg_reg_15__4_ ( .D(n404), .SIN(rn_reg[131]), .SMC(test_se), .C(
        net12553), .Q(rn_reg[132]) );
  SDFFQX1 rn_reg_reg_15__3_ ( .D(n392), .SIN(rn_reg[130]), .SMC(test_se), .C(
        net12553), .Q(rn_reg[131]) );
  SDFFQX1 rn_reg_reg_15__1_ ( .D(n399), .SIN(rn_reg[128]), .SMC(test_se), .C(
        net12553), .Q(rn_reg[129]) );
  SDFFQX1 rn_reg_reg_15__0_ ( .D(n411), .SIN(rn_reg[143]), .SMC(test_se), .C(
        net12553), .Q(rn_reg[128]) );
  SDFFQX1 rn_reg_reg_0__3_ ( .D(n391), .SIN(rn_reg[250]), .SMC(test_se), .C(
        net12478), .Q(rn_reg[251]) );
  SDFFQX1 rn_reg_reg_0__1_ ( .D(n400), .SIN(rn_reg[248]), .SMC(test_se), .C(
        net12478), .Q(rn_reg[249]) );
  SDFFQX1 rn_reg_reg_0__0_ ( .D(n410), .SIN(rmwinstr), .SMC(test_se), .C(
        net12478), .Q(rn_reg[248]) );
  SDFFQX1 rn_reg_reg_4__3_ ( .D(n391), .SIN(rn_reg[218]), .SMC(test_se), .C(
        net12498), .Q(rn_reg[219]) );
  SDFFQX1 rn_reg_reg_4__1_ ( .D(n400), .SIN(rn_reg[216]), .SMC(test_se), .C(
        net12498), .Q(rn_reg[217]) );
  SDFFQX1 rn_reg_reg_4__0_ ( .D(n410), .SIN(rn_reg[231]), .SMC(test_se), .C(
        net12498), .Q(rn_reg[216]) );
  SDFFQX1 rn_reg_reg_0__4_ ( .D(n403), .SIN(rn_reg[251]), .SMC(test_se), .C(
        net12478), .Q(rn_reg[252]) );
  SDFFQX1 rn_reg_reg_4__4_ ( .D(n403), .SIN(rn_reg[219]), .SMC(test_se), .C(
        net12498), .Q(rn_reg[220]) );
  SDFFQX1 rn_reg_reg_16__4_ ( .D(n404), .SIN(rn_reg[123]), .SMC(test_se), .C(
        net12558), .Q(rn_reg[124]) );
  SDFFQX1 rn_reg_reg_16__3_ ( .D(n392), .SIN(rn_reg[122]), .SMC(test_se), .C(
        net12558), .Q(rn_reg[123]) );
  SDFFQX1 rn_reg_reg_16__1_ ( .D(n399), .SIN(rn_reg[120]), .SMC(test_se), .C(
        net12558), .Q(rn_reg[121]) );
  SDFFQX1 rn_reg_reg_16__0_ ( .D(n411), .SIN(rn_reg[135]), .SMC(test_se), .C(
        net12558), .Q(rn_reg[120]) );
  SDFFQX1 rn_reg_reg_20__4_ ( .D(n405), .SIN(rn_reg[91]), .SMC(test_se), .C(
        net12578), .Q(rn_reg[92]) );
  SDFFQX1 rn_reg_reg_20__3_ ( .D(n393), .SIN(rn_reg[90]), .SMC(test_se), .C(
        net12578), .Q(rn_reg[91]) );
  SDFFQX1 rn_reg_reg_20__1_ ( .D(n398), .SIN(rn_reg[88]), .SMC(test_se), .C(
        net12578), .Q(rn_reg[89]) );
  SDFFQX1 rn_reg_reg_20__0_ ( .D(n412), .SIN(rn_reg[103]), .SMC(test_se), .C(
        net12578), .Q(rn_reg[88]) );
  SDFFQX1 rn_reg_reg_24__4_ ( .D(n402), .SIN(rn_reg[59]), .SMC(test_se), .C(
        net12598), .Q(rn_reg[60]) );
  SDFFQX1 rn_reg_reg_24__3_ ( .D(n390), .SIN(rn_reg[58]), .SMC(test_se), .C(
        net12598), .Q(rn_reg[59]) );
  SDFFQX1 rn_reg_reg_24__1_ ( .D(n401), .SIN(rn_reg[56]), .SMC(test_se), .C(
        net12598), .Q(rn_reg[57]) );
  SDFFQX1 rn_reg_reg_24__0_ ( .D(n410), .SIN(rn_reg[71]), .SMC(test_se), .C(
        net12598), .Q(rn_reg[56]) );
  SDFFQX1 rn_reg_reg_8__4_ ( .D(n404), .SIN(rn_reg[187]), .SMC(test_se), .C(
        net12518), .Q(rn_reg[188]) );
  SDFFQX1 rn_reg_reg_8__3_ ( .D(n392), .SIN(rn_reg[186]), .SMC(test_se), .C(
        net12518), .Q(rn_reg[187]) );
  SDFFQX1 rn_reg_reg_8__1_ ( .D(n399), .SIN(rn_reg[184]), .SMC(test_se), .C(
        net12518), .Q(rn_reg[185]) );
  SDFFQX1 rn_reg_reg_8__0_ ( .D(n411), .SIN(rn_reg[199]), .SMC(test_se), .C(
        net12518), .Q(rn_reg[184]) );
  SDFFQX1 rn_reg_reg_1__3_ ( .D(n391), .SIN(rn_reg[242]), .SMC(test_se), .C(
        net12483), .Q(rn_reg[243]) );
  SDFFQX1 rn_reg_reg_1__1_ ( .D(n400), .SIN(rn_reg[240]), .SMC(test_se), .C(
        net12483), .Q(rn_reg[241]) );
  SDFFQX1 rn_reg_reg_1__0_ ( .D(n410), .SIN(rn_reg[255]), .SMC(test_se), .C(
        net12483), .Q(rn_reg[240]) );
  SDFFQX1 rn_reg_reg_5__3_ ( .D(n391), .SIN(rn_reg[210]), .SMC(test_se), .C(
        net12503), .Q(rn_reg[211]) );
  SDFFQX1 rn_reg_reg_5__1_ ( .D(n400), .SIN(rn_reg[208]), .SMC(test_se), .C(
        net12503), .Q(rn_reg[209]) );
  SDFFQX1 rn_reg_reg_5__0_ ( .D(n410), .SIN(rn_reg[223]), .SMC(test_se), .C(
        net12503), .Q(rn_reg[208]) );
  SDFFQX1 rn_reg_reg_5__4_ ( .D(n403), .SIN(rn_reg[211]), .SMC(test_se), .C(
        net12503), .Q(rn_reg[212]) );
  SDFFQX1 rn_reg_reg_1__4_ ( .D(n403), .SIN(rn_reg[243]), .SMC(test_se), .C(
        net12483), .Q(rn_reg[244]) );
  SDFFQX1 rn_reg_reg_17__4_ ( .D(n404), .SIN(rn_reg[115]), .SMC(test_se), .C(
        net12563), .Q(rn_reg[116]) );
  SDFFQX1 rn_reg_reg_17__3_ ( .D(n392), .SIN(rn_reg[114]), .SMC(test_se), .C(
        net12563), .Q(rn_reg[115]) );
  SDFFQX1 rn_reg_reg_17__1_ ( .D(n399), .SIN(rn_reg[112]), .SMC(test_se), .C(
        net12563), .Q(rn_reg[113]) );
  SDFFQX1 rn_reg_reg_17__0_ ( .D(n412), .SIN(rn_reg[127]), .SMC(test_se), .C(
        net12563), .Q(rn_reg[112]) );
  SDFFQX1 rn_reg_reg_21__4_ ( .D(n405), .SIN(rn_reg[83]), .SMC(test_se), .C(
        net12583), .Q(rn_reg[84]) );
  SDFFQX1 rn_reg_reg_21__3_ ( .D(n393), .SIN(rn_reg[82]), .SMC(test_se), .C(
        net12583), .Q(rn_reg[83]) );
  SDFFQX1 rn_reg_reg_21__1_ ( .D(n398), .SIN(rn_reg[80]), .SMC(test_se), .C(
        net12583), .Q(rn_reg[81]) );
  SDFFQX1 rn_reg_reg_21__0_ ( .D(n412), .SIN(rn_reg[95]), .SMC(test_se), .C(
        net12583), .Q(rn_reg[80]) );
  SDFFQX1 rn_reg_reg_25__4_ ( .D(n405), .SIN(rn_reg[51]), .SMC(test_se), .C(
        net12603), .Q(rn_reg[52]) );
  SDFFQX1 rn_reg_reg_25__3_ ( .D(n393), .SIN(rn_reg[50]), .SMC(test_se), .C(
        net12603), .Q(rn_reg[51]) );
  SDFFQX1 rn_reg_reg_25__1_ ( .D(n398), .SIN(rn_reg[48]), .SMC(test_se), .C(
        net12603), .Q(rn_reg[49]) );
  SDFFQX1 rn_reg_reg_25__0_ ( .D(n409), .SIN(rn_reg[63]), .SMC(test_se), .C(
        net12603), .Q(rn_reg[48]) );
  SDFFQX1 rn_reg_reg_29__4_ ( .D(n405), .SIN(rn_reg[19]), .SMC(test_se), .C(
        net12623), .Q(rn_reg[20]) );
  SDFFQX1 rn_reg_reg_29__3_ ( .D(n393), .SIN(rn_reg[18]), .SMC(test_se), .C(
        net12623), .Q(rn_reg[19]) );
  SDFFQX1 rn_reg_reg_29__1_ ( .D(n398), .SIN(rn_reg[16]), .SMC(test_se), .C(
        net12623), .Q(rn_reg[17]) );
  SDFFQX1 rn_reg_reg_29__0_ ( .D(n412), .SIN(rn_reg[31]), .SMC(test_se), .C(
        net12623), .Q(rn_reg[16]) );
  SDFFQX1 rn_reg_reg_9__4_ ( .D(n404), .SIN(rn_reg[179]), .SMC(test_se), .C(
        net12523), .Q(rn_reg[180]) );
  SDFFQX1 rn_reg_reg_9__3_ ( .D(n392), .SIN(rn_reg[178]), .SMC(test_se), .C(
        net12523), .Q(rn_reg[179]) );
  SDFFQX1 rn_reg_reg_9__1_ ( .D(n399), .SIN(rn_reg[176]), .SMC(test_se), .C(
        net12523), .Q(rn_reg[177]) );
  SDFFQX1 rn_reg_reg_9__0_ ( .D(n411), .SIN(rn_reg[191]), .SMC(test_se), .C(
        net12523), .Q(rn_reg[176]) );
  SDFFQX1 rn_reg_reg_13__4_ ( .D(n404), .SIN(rn_reg[147]), .SMC(test_se), .C(
        net12543), .Q(rn_reg[148]) );
  SDFFQX1 rn_reg_reg_13__3_ ( .D(n392), .SIN(rn_reg[146]), .SMC(test_se), .C(
        net12543), .Q(rn_reg[147]) );
  SDFFQX1 rn_reg_reg_13__1_ ( .D(n399), .SIN(rn_reg[144]), .SMC(test_se), .C(
        net12543), .Q(rn_reg[145]) );
  SDFFQX1 rn_reg_reg_13__0_ ( .D(n411), .SIN(rn_reg[159]), .SMC(test_se), .C(
        net12543), .Q(rn_reg[144]) );
  SDFFQX1 rn_reg_reg_2__3_ ( .D(n391), .SIN(rn_reg[234]), .SMC(test_se), .C(
        net12488), .Q(rn_reg[235]) );
  SDFFQX1 rn_reg_reg_2__1_ ( .D(n400), .SIN(rn_reg[232]), .SMC(test_se), .C(
        net12488), .Q(rn_reg[233]) );
  SDFFQX1 rn_reg_reg_2__0_ ( .D(n410), .SIN(rn_reg[247]), .SMC(test_se), .C(
        net12488), .Q(rn_reg[232]) );
  SDFFQX1 rn_reg_reg_2__4_ ( .D(n403), .SIN(rn_reg[235]), .SMC(test_se), .C(
        net12488), .Q(rn_reg[236]) );
  SDFFQX1 rn_reg_reg_18__4_ ( .D(n405), .SIN(rn_reg[107]), .SMC(test_se), .C(
        net12568), .Q(rn_reg[108]) );
  SDFFQX1 rn_reg_reg_18__3_ ( .D(n393), .SIN(rn_reg[106]), .SMC(test_se), .C(
        net12568), .Q(rn_reg[107]) );
  SDFFQX1 rn_reg_reg_18__1_ ( .D(n398), .SIN(rn_reg[104]), .SMC(test_se), .C(
        net12568), .Q(rn_reg[105]) );
  SDFFQX1 rn_reg_reg_18__0_ ( .D(n412), .SIN(rn_reg[119]), .SMC(test_se), .C(
        net12568), .Q(rn_reg[104]) );
  SDFFQX1 dpl_reg_reg_3__0_ ( .D(N12593), .SIN(dpl_reg[23]), .SMC(test_se), 
        .C(net12408), .Q(dpl_reg[24]) );
  SDFFQX1 dpl_reg_reg_7__1_ ( .D(N12630), .SIN(dpl_reg[56]), .SMC(test_se), 
        .C(net12388), .Q(dpl_reg[57]) );
  SDFFQX1 dpl_reg_reg_7__0_ ( .D(N12629), .SIN(dpl_reg[55]), .SMC(test_se), 
        .C(net12388), .Q(dpl_reg[56]) );
  SDFFQX1 dpl_reg_reg_2__0_ ( .D(N12584), .SIN(dpl_reg[15]), .SMC(test_se), 
        .C(net12413), .Q(dpl_reg[16]) );
  SDFFQX1 dpl_reg_reg_6__1_ ( .D(N12621), .SIN(dpl_reg[48]), .SMC(test_se), 
        .C(net12393), .Q(dpl_reg[49]) );
  SDFFQX1 dpl_reg_reg_6__0_ ( .D(N12620), .SIN(dpl_reg[47]), .SMC(test_se), 
        .C(net12393), .Q(dpl_reg[48]) );
  SDFFQX1 dec_cop_reg_4_ ( .D(N10586), .SIN(dec_cop[3]), .SMC(test_se), .C(
        net12372), .Q(dec_cop[4]) );
  SDFFQX1 sp_reg_reg_5_ ( .D(N12702), .SIN(sp[4]), .SMC(test_se), .C(net12372), 
        .Q(sp[5]) );
  SDFFQX1 dec_cop_reg_3_ ( .D(N10585), .SIN(dec_cop[2]), .SMC(test_se), .C(
        net12372), .Q(dec_cop[3]) );
  SDFFQX1 dpl_reg_reg_5__1_ ( .D(N12612), .SIN(dpl_reg[40]), .SMC(test_se), 
        .C(net12398), .Q(dpl_reg[41]) );
  SDFFQX1 dpl_reg_reg_5__0_ ( .D(N12611), .SIN(dpl_reg[39]), .SMC(test_se), 
        .C(net12398), .Q(dpl_reg[40]) );
  SDFFQX1 dpl_reg_reg_1__1_ ( .D(N12576), .SIN(dpl_reg[8]), .SMC(test_se), .C(
        net12418), .Q(dpl_reg[9]) );
  SDFFQX1 dpl_reg_reg_1__0_ ( .D(N12575), .SIN(dpl_reg[7]), .SMC(test_se), .C(
        net12418), .Q(dpl_reg[8]) );
  SDFFQX1 dpl_reg_reg_0__1_ ( .D(N12567), .SIN(dpl_reg[0]), .SMC(test_se), .C(
        net12423), .Q(dpl_reg[1]) );
  SDFFQX1 dpl_reg_reg_0__0_ ( .D(N12566), .SIN(dph_reg[63]), .SMC(test_se), 
        .C(net12423), .Q(dpl_reg[0]) );
  SDFFQX1 dpl_reg_reg_4__1_ ( .D(N12603), .SIN(dpl_reg[32]), .SMC(test_se), 
        .C(net12403), .Q(dpl_reg[33]) );
  SDFFQX1 dpl_reg_reg_4__0_ ( .D(N12602), .SIN(dpl_reg[31]), .SMC(test_se), 
        .C(net12403), .Q(dpl_reg[32]) );
  SDFFQX1 dec_cop_reg_7_ ( .D(N10589), .SIN(dec_cop[6]), .SMC(test_se), .C(
        net12372), .Q(dec_cop[7]) );
  SDFFQX1 ckcon_r_reg_3_ ( .D(N12968), .SIN(ckcon[2]), .SMC(test_se), .C(
        net12372), .Q(ckcon[3]) );
  SDFFQX1 ckcon_r_reg_7_ ( .D(N12972), .SIN(ckcon[6]), .SMC(test_se), .C(
        net12372), .Q(ckcon[7]) );
  SDFFQX1 pmw_reg_reg ( .D(n2830), .SIN(phase[5]), .SMC(test_se), .C(net12372), 
        .Q(pmw) );
  SDFFQX1 temp2_reg_7_ ( .D(N12730), .SIN(temp2_comb[6]), .SMC(test_se), .C(
        net12372), .Q(temp2_comb[7]) );
  SDFFQX1 waitcnt_reg_0_ ( .D(N12974), .SIN(temp[7]), .SMC(test_se), .C(
        net12473), .Q(waitcnt_0_) );
  SDFFQX1 dec_accop_reg_17_ ( .D(n2824), .SIN(dec_accop[16]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[17]) );
  SDFFQX1 ramdatao_r_reg_5_ ( .D(N11503), .SIN(ramdatao[4]), .SMC(test_se), 
        .C(net12372), .Q(ramdatao[5]) );
  SDFFQX1 ramdatao_r_reg_7_ ( .D(N11505), .SIN(ramdatao[6]), .SMC(test_se), 
        .C(net12372), .Q(ramdatao[7]) );
  SDFFQX1 rn_reg_reg_26__4_ ( .D(n402), .SIN(rn_reg[43]), .SMC(test_se), .C(
        net12608), .Q(rn_reg[44]) );
  SDFFQX1 rn_reg_reg_26__3_ ( .D(n390), .SIN(rn_reg[42]), .SMC(test_se), .C(
        net12608), .Q(rn_reg[43]) );
  SDFFQX1 rn_reg_reg_26__1_ ( .D(n400), .SIN(rn_reg[40]), .SMC(test_se), .C(
        net12608), .Q(rn_reg[41]) );
  SDFFQX1 rn_reg_reg_26__0_ ( .D(n2832), .SIN(rn_reg[55]), .SMC(test_se), .C(
        net12608), .Q(rn_reg[40]) );
  SDFFQX1 rn_reg_reg_30__4_ ( .D(n402), .SIN(rn_reg[11]), .SMC(test_se), .C(
        net12628), .Q(rn_reg[12]) );
  SDFFQX1 rn_reg_reg_30__3_ ( .D(n390), .SIN(rn_reg[10]), .SMC(test_se), .C(
        net12628), .Q(rn_reg[11]) );
  SDFFQX1 rn_reg_reg_30__1_ ( .D(n401), .SIN(rn_reg[8]), .SMC(test_se), .C(
        net12628), .Q(rn_reg[9]) );
  SDFFQX1 rn_reg_reg_30__0_ ( .D(n412), .SIN(rn_reg[23]), .SMC(test_se), .C(
        net12628), .Q(rn_reg[8]) );
  SDFFQX1 rn_reg_reg_10__4_ ( .D(n404), .SIN(rn_reg[171]), .SMC(test_se), .C(
        net12528), .Q(rn_reg[172]) );
  SDFFQX1 rn_reg_reg_10__3_ ( .D(n392), .SIN(rn_reg[170]), .SMC(test_se), .C(
        net12528), .Q(rn_reg[171]) );
  SDFFQX1 rn_reg_reg_10__1_ ( .D(n399), .SIN(rn_reg[168]), .SMC(test_se), .C(
        net12528), .Q(rn_reg[169]) );
  SDFFQX1 rn_reg_reg_10__0_ ( .D(n411), .SIN(rn_reg[183]), .SMC(test_se), .C(
        net12528), .Q(rn_reg[168]) );
  SDFFQX1 rn_reg_reg_14__4_ ( .D(n404), .SIN(rn_reg[139]), .SMC(test_se), .C(
        net12548), .Q(rn_reg[140]) );
  SDFFQX1 rn_reg_reg_14__3_ ( .D(n392), .SIN(rn_reg[138]), .SMC(test_se), .C(
        net12548), .Q(rn_reg[139]) );
  SDFFQX1 rn_reg_reg_14__1_ ( .D(n399), .SIN(rn_reg[136]), .SMC(test_se), .C(
        net12548), .Q(rn_reg[137]) );
  SDFFQX1 rn_reg_reg_14__0_ ( .D(n411), .SIN(rn_reg[151]), .SMC(test_se), .C(
        net12548), .Q(rn_reg[136]) );
  SDFFQX1 dec_accop_reg_12_ ( .D(N10575), .SIN(dec_accop[11]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[12]) );
  SDFFQX1 dec_cop_reg_6_ ( .D(N10588), .SIN(dec_cop[5]), .SMC(test_se), .C(
        net12372), .Q(dec_cop[6]) );
  SDFFQX1 temp2_reg_6_ ( .D(N12729), .SIN(temp2_comb[5]), .SMC(test_se), .C(
        net12372), .Q(temp2_comb[6]) );
  SDFFQX1 sp_reg_reg_4_ ( .D(N12701), .SIN(sp[3]), .SMC(test_se), .C(net12372), 
        .Q(sp[4]) );
  SDFFQX1 dec_accop_reg_15_ ( .D(N10578), .SIN(dec_accop[14]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[15]) );
  SDFFQX1 dec_cop_reg_5_ ( .D(N10587), .SIN(dec_cop[4]), .SMC(test_se), .C(
        net12372), .Q(dec_cop[5]) );
  SDFFQX1 temp_reg_2_ ( .D(N12716), .SIN(temp[1]), .SMC(test_se), .C(net12468), 
        .Q(temp[2]) );
  SDFFQX1 temp_reg_0_ ( .D(N12714), .SIN(temp2_comb[7]), .SMC(test_se), .C(
        net12468), .Q(temp[0]) );
  SDFFQX1 temp_reg_4_ ( .D(N12718), .SIN(temp[3]), .SMC(test_se), .C(net12468), 
        .Q(temp[4]) );
  SDFFQX1 temp_reg_1_ ( .D(N12715), .SIN(temp[0]), .SMC(test_se), .C(net12468), 
        .Q(temp[1]) );
  SDFFQX1 temp_reg_3_ ( .D(N12717), .SIN(temp[2]), .SMC(test_se), .C(net12468), 
        .Q(temp[3]) );
  SDFFQX1 temp_reg_7_ ( .D(N12721), .SIN(temp[6]), .SMC(test_se), .C(net12468), 
        .Q(temp[7]) );
  SDFFQX1 dec_accop_reg_13_ ( .D(N10576), .SIN(dec_accop[12]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[13]) );
  SDFFQX1 temp_reg_5_ ( .D(N12719), .SIN(temp[4]), .SMC(test_se), .C(net12468), 
        .Q(temp[5]) );
  SDFFQX1 temp_reg_6_ ( .D(N12720), .SIN(temp[5]), .SMC(test_se), .C(net12468), 
        .Q(temp[6]) );
  SDFFQX1 bitno_reg_2_ ( .D(n2837), .SIN(N344), .SMC(test_se), .C(net12383), 
        .Q(N345) );
  SDFFQX1 divtempreg_reg_6_ ( .D(N13373), .SIN(divtempreg[5]), .SMC(test_se), 
        .C(net12643), .Q(divtempreg[6]) );
  SDFFQX1 ramwe_r_reg ( .D(N11487), .SIN(ramsfrwe), .SMC(test_se), .C(net12372), .Q(ramwe) );
  SDFFQX1 temp2_reg_5_ ( .D(N12728), .SIN(temp2_comb[4]), .SMC(test_se), .C(
        net12372), .Q(temp2_comb[5]) );
  SDFFQX1 temp2_reg_4_ ( .D(N12727), .SIN(temp2_comb[3]), .SMC(test_se), .C(
        net12372), .Q(temp2_comb[4]) );
  SDFFQX1 sp_reg_reg_3_ ( .D(N12700), .SIN(sp[2]), .SMC(test_se), .C(net12372), 
        .Q(sp[3]) );
  SDFFQX1 dec_accop_reg_11_ ( .D(N10574), .SIN(dec_accop[10]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[11]) );
  SDFFQX1 sp_reg_reg_2_ ( .D(N12699), .SIN(sp[1]), .SMC(test_se), .C(net12372), 
        .Q(sp[2]) );
  SDFFQX1 sp_reg_reg_0_ ( .D(N12697), .SIN(sfrwe_r), .SMC(test_se), .C(
        net12372), .Q(sp[0]) );
  SDFFQX1 dec_accop_reg_3_ ( .D(N10566), .SIN(dec_accop[2]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[3]) );
  SDFFQX1 bitno_reg_0_ ( .D(n2835), .SIN(b[7]), .SMC(test_se), .C(net12383), 
        .Q(N343) );
  SDFFQX1 temp2_reg_3_ ( .D(N12726), .SIN(temp2_comb[2]), .SMC(test_se), .C(
        net12372), .Q(temp2_comb[3]) );
  SDFFQX1 dec_accop_reg_4_ ( .D(N10567), .SIN(dec_accop[3]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[4]) );
  SDFFQX1 sp_reg_reg_1_ ( .D(N12698), .SIN(sp[0]), .SMC(test_se), .C(net12372), 
        .Q(sp[1]) );
  SDFFQX1 dec_accop_reg_1_ ( .D(N10564), .SIN(dec_accop[0]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[1]) );
  SDFFQX1 bitno_reg_1_ ( .D(n2836), .SIN(N343), .SMC(test_se), .C(net12383), 
        .Q(N344) );
  SDFFQX1 phase_reg_2_ ( .D(N681), .SIN(n214), .SMC(test_se), .C(net12372), 
        .Q(phase[2]) );
  SDFFQX1 accactv_reg ( .D(N10562), .SIN(acc[7]), .SMC(test_se), .C(net12372), 
        .Q(accactv) );
  SDFFQX1 dps_reg_reg_0_ ( .D(N12693), .SIN(dpl_reg[63]), .SMC(test_se), .C(
        net12372), .Q(dps[0]) );
  SDFFQX1 acc_reg_reg_5_ ( .D(n2823), .SIN(acc[4]), .SMC(test_se), .C(net12372), .Q(acc[5]) );
  SDFFQX1 acc_reg_reg_4_ ( .D(n2820), .SIN(acc[3]), .SMC(test_se), .C(net12372), .Q(acc[4]) );
  SDFFQX1 interrupt_reg ( .D(n2841), .SIN(instr[7]), .SMC(test_se), .C(
        net12378), .Q(interrupt) );
  SDFFQX1 ramdatao_r_reg_2_ ( .D(N11500), .SIN(ramdatao[1]), .SMC(test_se), 
        .C(net12372), .Q(ramdatao[2]) );
  SDFFQX1 dps_reg_reg_1_ ( .D(N12694), .SIN(dps[0]), .SMC(test_se), .C(
        net12372), .Q(dps[1]) );
  SDFFQX1 b_reg_reg_7_ ( .D(N12484), .SIN(b[6]), .SMC(test_se), .C(net12372), 
        .Q(b[7]) );
  SDFFQX1 pc_reg_2_ ( .D(N482), .SIN(pc_o[1]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[2]) );
  SDFFQX1 temp2_reg_2_ ( .D(N12725), .SIN(temp2_comb[1]), .SMC(test_se), .C(
        net12372), .Q(temp2_comb[2]) );
  SDFFQX1 ramsfraddr_s_reg_5_ ( .D(N11483), .SIN(ramsfraddr[4]), .SMC(test_se), 
        .C(net12372), .Q(ramsfraddr[5]) );
  SDFFQX1 divtempreg_reg_5_ ( .D(N13372), .SIN(divtempreg[4]), .SMC(test_se), 
        .C(net12643), .Q(divtempreg[5]) );
  SDFFQX1 instr_reg_4_ ( .D(N674), .SIN(instr[3]), .SMC(test_se), .C(net12378), 
        .Q(n2869) );
  SDFFQX1 temp2_reg_1_ ( .D(N12724), .SIN(temp2_comb[0]), .SMC(test_se), .C(
        net12372), .Q(temp2_comb[1]) );
  SDFFQX1 divtempreg_reg_3_ ( .D(N13370), .SIN(divtempreg[2]), .SMC(test_se), 
        .C(net12643), .Q(divtempreg[3]) );
  SDFFQX1 divtempreg_reg_4_ ( .D(N13371), .SIN(divtempreg[3]), .SMC(test_se), 
        .C(net12643), .Q(divtempreg[4]) );
  SDFFQX1 ramsfraddr_s_reg_3_ ( .D(N11481), .SIN(ramsfraddr[2]), .SMC(test_se), 
        .C(net12372), .Q(ramsfraddr[3]) );
  SDFFQX1 b_reg_reg_6_ ( .D(N12483), .SIN(b[5]), .SMC(test_se), .C(net12372), 
        .Q(b[6]) );
  SDFFQX1 b_reg_reg_4_ ( .D(N12481), .SIN(b[3]), .SMC(test_se), .C(net12372), 
        .Q(b[4]) );
  SDFFQX1 dec_accop_reg_9_ ( .D(N10572), .SIN(dec_accop[8]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[9]) );
  SDFFQX1 dec_accop_reg_7_ ( .D(N10570), .SIN(dec_accop[6]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[7]) );
  SDFFQX1 ac_reg_reg ( .D(N12706), .SIN(test_si), .SMC(test_se), .C(net12372), 
        .Q(ac) );
  SDFFQX1 b_reg_reg_5_ ( .D(N12482), .SIN(b[4]), .SMC(test_se), .C(net12372), 
        .Q(b[5]) );
  SDFFQX1 acc_reg_reg_3_ ( .D(N12472), .SIN(acc[2]), .SMC(test_se), .C(
        net12372), .Q(acc[3]) );
  SDFFQX1 instr_reg_2_ ( .D(N672), .SIN(instr[1]), .SMC(test_se), .C(net12378), 
        .Q(n2871) );
  SDFFQXL dec_accop_reg_0_ ( .D(N10563), .SIN(d_hold), .SMC(test_se), .C(
        net12372), .Q(dec_accop[0]) );
  SDFFQXL dec_accop_reg_2_ ( .D(N10565), .SIN(dec_accop[1]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[2]) );
  SDFFQXL dec_accop_reg_14_ ( .D(N10577), .SIN(dec_accop[13]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[14]) );
  SDFFQX1 phase_reg_1_ ( .D(N680), .SIN(n2549), .SMC(test_se), .C(net12372), 
        .Q(phase[1]) );
  SDFFQX1 dps_reg_reg_3_ ( .D(n1884), .SIN(n207), .SMC(test_se), .C(net12372), 
        .Q(dps[3]) );
  SDFFQX1 ramdatao_r_reg_0_ ( .D(N11498), .SIN(pmw), .SMC(test_se), .C(
        net12372), .Q(ramdatao[0]) );
  SDFFQX1 rs_reg_reg_0_ ( .D(N12709), .SIN(rn_reg[7]), .SMC(test_se), .C(
        net12372), .Q(rs[0]) );
  SDFFQX1 rs_reg_reg_1_ ( .D(N12710), .SIN(rs[0]), .SMC(test_se), .C(net12372), 
        .Q(rs[1]) );
  SDFFQX1 ramdatao_r_reg_1_ ( .D(N11499), .SIN(ramdatao[0]), .SMC(test_se), 
        .C(net12372), .Q(ramdatao[1]) );
  SDFFQX1 pc_reg_3_ ( .D(N483), .SIN(pc_o[2]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[3]) );
  SDFFQX1 dps_reg_reg_2_ ( .D(N12695), .SIN(dps[1]), .SMC(test_se), .C(
        net12372), .Q(dps[2]) );
  SDFFQX1 dec_accop_reg_6_ ( .D(N10569), .SIN(dec_accop[5]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[6]) );
  SDFFQX1 acc_reg_reg_6_ ( .D(n2822), .SIN(acc[5]), .SMC(test_se), .C(net12372), .Q(acc[6]) );
  SDFFQX1 pc_reg_4_ ( .D(N484), .SIN(pc_o[3]), .SMC(test_se), .C(net12372), 
        .Q(pc_o[4]) );
  SDFFQX1 ramsfraddr_s_reg_1_ ( .D(N11479), .SIN(ramsfraddr[0]), .SMC(test_se), 
        .C(net12372), .Q(ramsfraddr[1]) );
  SDFFQX1 divtempreg_reg_1_ ( .D(N13368), .SIN(divtempreg[0]), .SMC(test_se), 
        .C(net12643), .Q(divtempreg[1]) );
  SDFFQX1 temp2_reg_0_ ( .D(N12723), .SIN(stop), .SMC(test_se), .C(net12372), 
        .Q(temp2_comb[0]) );
  SDFFQX1 divtempreg_reg_0_ ( .D(N13367), .SIN(dec_cop[7]), .SMC(test_se), .C(
        net12643), .Q(divtempreg[0]) );
  SDFFQX1 dec_accop_reg_10_ ( .D(N10573), .SIN(dec_accop[9]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[10]) );
  SDFFQX1 dec_accop_reg_8_ ( .D(N10571), .SIN(dec_accop[7]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[8]) );
  SDFFQX1 dec_accop_reg_16_ ( .D(n2825), .SIN(dec_accop[15]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[16]) );
  SDFFQX1 instr_reg_5_ ( .D(N675), .SIN(n2869), .SMC(test_se), .C(net12378), 
        .Q(n2868) );
  SDFFQX1 instr_reg_1_ ( .D(N671), .SIN(instr[0]), .SMC(test_se), .C(net12378), 
        .Q(n2872) );
  SDFFQX1 ramdatao_r_reg_3_ ( .D(N11501), .SIN(ramdatao[2]), .SMC(test_se), 
        .C(net12372), .Q(ramdatao[3]) );
  SDFFQX1 phase_reg_0_ ( .D(N679), .SIN(phase0_ff), .SMC(test_se), .C(net12372), .Q(phase[0]) );
  SDFFQX1 instr_reg_3_ ( .D(N673), .SIN(instr[2]), .SMC(test_se), .C(net12378), 
        .Q(n2870) );
  SDFFQX1 instr_reg_0_ ( .D(N670), .SIN(idle), .SMC(test_se), .C(net12378), 
        .Q(n2873) );
  SDFFQX1 instr_reg_7_ ( .D(N677), .SIN(instr[6]), .SMC(test_se), .C(net12378), 
        .Q(n2866) );
  SDFFQX1 pc_reg_0_ ( .D(N480), .SIN(p), .SMC(test_se), .C(net12372), .Q(n2865) );
  SDFFQX1 pc_reg_1_ ( .D(N481), .SIN(memaddr[0]), .SMC(test_se), .C(net12372), 
        .Q(memaddr[1]) );
  SDFFQX1 dec_accop_reg_18_ ( .D(N10581), .SIN(dec_accop[17]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[18]) );
  SDFFQX1 ramdatao_r_reg_4_ ( .D(N11502), .SIN(ramdatao[3]), .SMC(test_se), 
        .C(net12372), .Q(ramdatao[4]) );
  SDFFQX1 ramsfraddr_s_reg_6_ ( .D(N11484), .SIN(ramsfraddr[5]), .SMC(test_se), 
        .C(net12372), .Q(ramsfraddr[6]) );
  SDFFQX1 ramsfrwe_reg ( .D(n2829), .SIN(ramsfraddr[7]), .SMC(test_se), .C(
        net12372), .Q(ramsfrwe) );
  SDFFQX1 b_reg_reg_1_ ( .D(N12478), .SIN(b[0]), .SMC(test_se), .C(net12372), 
        .Q(b[1]) );
  SDFFQX1 b_reg_reg_0_ ( .D(N12477), .SIN(accactv), .SMC(test_se), .C(net12372), .Q(b[0]) );
  SDFFQX1 acc_reg_reg_7_ ( .D(n2816), .SIN(acc[6]), .SMC(test_se), .C(net12372), .Q(acc[7]) );
  SDFFQX1 dec_accop_reg_5_ ( .D(N10568), .SIN(dec_accop[4]), .SMC(test_se), 
        .C(net12372), .Q(dec_accop[5]) );
  SDFFQX1 ramsfraddr_s_reg_0_ ( .D(N11478), .SIN(ramoe), .SMC(test_se), .C(
        net12372), .Q(ramsfraddr[0]) );
  SDFFQX1 ramsfraddr_s_reg_4_ ( .D(N11482), .SIN(ramsfraddr[3]), .SMC(test_se), 
        .C(net12372), .Q(ramsfraddr[4]) );
  SDFFQX1 ramsfraddr_s_reg_7_ ( .D(n2834), .SIN(ramsfraddr[6]), .SMC(test_se), 
        .C(net12372), .Q(ramsfraddr[7]) );
  SDFFQX1 divtempreg_reg_2_ ( .D(N13369), .SIN(divtempreg[1]), .SMC(test_se), 
        .C(net12643), .Q(divtempreg[2]) );
  SDFFQX1 ramsfraddr_s_reg_2_ ( .D(N11480), .SIN(ramsfraddr[1]), .SMC(test_se), 
        .C(net12372), .Q(ramsfraddr[2]) );
  SDFFQX1 b_reg_reg_3_ ( .D(N12480), .SIN(b[2]), .SMC(test_se), .C(net12372), 
        .Q(b[3]) );
  SDFFQX1 b_reg_reg_2_ ( .D(N12479), .SIN(b[1]), .SMC(test_se), .C(net12372), 
        .Q(b[2]) );
  SDFFQX1 acc_reg_reg_2_ ( .D(n2821), .SIN(n193), .SMC(test_se), .C(net12372), 
        .Q(acc[2]) );
  SDFFQX1 acc_reg_reg_1_ ( .D(N12470), .SIN(n170), .SMC(test_se), .C(net12372), 
        .Q(acc[1]) );
  SDFFQX1 acc_reg_reg_0_ ( .D(N12469), .SIN(ac), .SMC(test_se), .C(net12372), 
        .Q(acc[0]) );
  SDFFQX1 instr_reg_6_ ( .D(N676), .SIN(instr[5]), .SMC(test_se), .C(net12378), 
        .Q(n2867) );
  SDFFQX1 c_reg_reg ( .D(N12705), .SIN(N345), .SMC(test_se), .C(net12372), .Q(
        c) );
  BUFXL U9 ( .A(n276), .Y(n1) );
  INVX2 U10 ( .A(memdatai[6]), .Y(n2491) );
  INVX2 U11 ( .A(memdatai[1]), .Y(n1297) );
  INVX2 U12 ( .A(memdatai[7]), .Y(n1218) );
  XNOR2X1 U13 ( .A(n783), .B(ramsfraddr[3]), .Y(n318) );
  OAI221X4 U14 ( .A(n156), .B(n655), .C(n970), .D(n654), .E(n220), .Y(n656) );
  OAI222X4 U15 ( .A(n2185), .B(n2228), .C(n1183), .D(n2165), .E(n1173), .F(
        n1181), .Y(n2636) );
  OAI222X1 U16 ( .A(n2185), .B(n1297), .C(n1183), .D(n2180), .E(n1175), .F(
        n1181), .Y(n2637) );
  OAI222X1 U17 ( .A(n1184), .B(n2165), .C(n2491), .D(n1183), .E(n1182), .F(
        n1181), .Y(n2639) );
  INVX2 U18 ( .A(memdatai[0]), .Y(n2228) );
  XOR2X1 U19 ( .A(n1867), .B(n345), .Y(n1440) );
  MUX2X2 U20 ( .D0(memaddr[5]), .D1(n2685), .S(n362), .Y(memaddr_comb[5]) );
  MUX2IX2 U21 ( .D0(n53), .D1(n106), .S(n2690), .Y(memaddr_comb[1]) );
  NOR21X2 U22 ( .B(n291), .A(n1035), .Y(n2662) );
  INVX1 U23 ( .A(sfrdatai[1]), .Y(n1305) );
  INVX2 U24 ( .A(n1760), .Y(n2097) );
  NAND5X2 U25 ( .A(n523), .B(n2554), .C(n522), .D(n521), .E(n520), .Y(n561) );
  NAND21X2 U26 ( .B(dec_accop[9]), .A(n1055), .Y(n1082) );
  INVX2 U27 ( .A(n1080), .Y(n1055) );
  NOR32X2 U28 ( .B(n2679), .C(n422), .A(n2678), .Y(n88) );
  AOI221X1 U29 ( .A(rn_reg[72]), .B(n975), .C(rn_reg[24]), .D(n974), .E(n671), 
        .Y(n687) );
  OAI221X4 U30 ( .A(n156), .B(n670), .C(n970), .D(n669), .E(n968), .Y(n671) );
  OAI221X1 U31 ( .A(n156), .B(n700), .C(n970), .D(n699), .E(n220), .Y(n701) );
  INVX2 U32 ( .A(memdatai[4]), .Y(n2180) );
  MUX2IX4 U33 ( .D0(n67), .D1(n2504), .S(n1179), .Y(n2618) );
  INVX2 U34 ( .A(n1218), .Y(n67) );
  NAND21X2 U35 ( .B(n276), .A(n1980), .Y(n2481) );
  INVX2 U36 ( .A(n2618), .Y(n2644) );
  AND2X2 U37 ( .A(n272), .B(n1747), .Y(n1429) );
  AOI221X1 U38 ( .A(rn_reg[75]), .B(n975), .C(rn_reg[27]), .D(n974), .E(n760), 
        .Y(n776) );
  OAI221XL U39 ( .A(n156), .B(n759), .C(n970), .D(n758), .E(n968), .Y(n760) );
  AOI221X1 U40 ( .A(rn_reg[73]), .B(n975), .C(rn_reg[25]), .D(n974), .E(n805), 
        .Y(n821) );
  INVX2 U41 ( .A(n1083), .Y(n1424) );
  NAND2X1 U42 ( .A(n10), .B(n11), .Y(n102) );
  NOR2X2 U43 ( .A(n1009), .B(n1343), .Y(n220) );
  AOI221X1 U44 ( .A(rn_reg[200]), .B(n975), .C(rn_reg[152]), .D(n974), .E(n656), .Y(n691) );
  AOI21BBX1 U45 ( .B(n85), .C(n333), .A(n216), .Y(n1432) );
  INVX2 U46 ( .A(n2639), .Y(n1185) );
  OAI221X1 U47 ( .A(n293), .B(n1440), .C(n1918), .D(n2329), .E(n1439), .Y(
        n1441) );
  XOR2X2 U48 ( .A(n1868), .B(n2206), .Y(n1867) );
  AOI221X1 U49 ( .A(rn_reg[203]), .B(n975), .C(rn_reg[155]), .D(n974), .E(n745), .Y(n780) );
  AOI221X1 U50 ( .A(rn_reg[201]), .B(n975), .C(rn_reg[153]), .D(n974), .E(n790), .Y(n825) );
  AOI221X1 U51 ( .A(rn_reg[76]), .B(n975), .C(rn_reg[28]), .D(n974), .E(n716), 
        .Y(n732) );
  OAI221XL U52 ( .A(n156), .B(n715), .C(n970), .D(n714), .E(n968), .Y(n716) );
  AOI221X1 U53 ( .A(rn_reg[204]), .B(n975), .C(rn_reg[156]), .D(n974), .E(n701), .Y(n736) );
  MUX2BXL U54 ( .D0(n1904), .D1(n1190), .S(acc[0]), .Y(n1191) );
  NAND21X1 U55 ( .B(n1845), .A(n334), .Y(n1067) );
  INVX1 U56 ( .A(n878), .Y(n1175) );
  OR2X1 U57 ( .A(n508), .B(n507), .Y(n876) );
  NAND21X1 U58 ( .B(n507), .A(n508), .Y(n875) );
  INVX2 U59 ( .A(dec_accop[18]), .Y(n1076) );
  INVX1 U60 ( .A(n2659), .Y(n97) );
  INVX1 U61 ( .A(temp2_comb[1]), .Y(n2459) );
  INVX1 U62 ( .A(n881), .Y(n1182) );
  INVX2 U63 ( .A(n561), .Y(n1009) );
  NOR3XL U64 ( .A(n1865), .B(n1071), .C(n294), .Y(n293) );
  INVX1 U65 ( .A(n1769), .Y(n1071) );
  INVX1 U66 ( .A(n873), .Y(n946) );
  AO21X1 U67 ( .B(n1158), .C(n214), .A(n1046), .Y(n951) );
  AOI21X1 U68 ( .B(n1063), .C(n1850), .A(n1845), .Y(n287) );
  INVX1 U69 ( .A(n1703), .Y(n68) );
  INVX1 U70 ( .A(n1068), .Y(n1075) );
  NAND21X1 U71 ( .B(dec_accop[5]), .A(n1078), .Y(n1068) );
  OA222XL U72 ( .A(n293), .B(n1194), .C(n1193), .D(n2094), .E(n1791), .F(n2383), .Y(n1195) );
  AO21X1 U73 ( .B(ramdatao[2]), .C(n1906), .A(n1745), .Y(n1751) );
  NAND21X1 U74 ( .B(n1096), .A(n503), .Y(n1046) );
  INVX1 U75 ( .A(n1097), .Y(n503) );
  INVX1 U76 ( .A(n345), .Y(n77) );
  INVXL U77 ( .A(n2206), .Y(n75) );
  AO2222X1 U78 ( .A(n2287), .B(n1012), .C(n2351), .D(n1013), .E(temp[5]), .F(
        n1011), .G(ramsfraddr[5]), .H(n1010), .Y(n879) );
  NAND2XL U79 ( .A(n258), .B(n2112), .Y(n10) );
  INVX3 U80 ( .A(ramsfraddr[7]), .Y(n2554) );
  INVX1 U81 ( .A(n1870), .Y(n91) );
  INVX1 U82 ( .A(n1871), .Y(n90) );
  NAND21X1 U83 ( .B(n1067), .A(dec_accop[13]), .Y(n1909) );
  OA222X1 U84 ( .A(n1918), .B(n1965), .C(n1086), .D(n2459), .E(n293), .F(n1085), .Y(n1087) );
  INVX1 U85 ( .A(n1610), .Y(n1622) );
  OAI221X1 U86 ( .A(n875), .B(n2159), .C(n2569), .D(n876), .E(n784), .Y(n881)
         );
  OAI221X1 U87 ( .A(n875), .B(n2233), .C(n234), .D(n1157), .E(n829), .Y(n878)
         );
  INVX1 U88 ( .A(n1179), .Y(n2) );
  OAI221X1 U89 ( .A(n875), .B(n2382), .C(n234), .D(n1254), .E(n739), .Y(n1178)
         );
  INVX1 U90 ( .A(acc[6]), .Y(n2329) );
  NAND21X1 U91 ( .B(n1117), .A(n469), .Y(n1610) );
  NAND43X1 U92 ( .B(n1708), .C(n221), .D(n222), .A(n1707), .Y(n2158) );
  OA222XL U93 ( .A(n1918), .B(n2263), .C(n1706), .D(n2160), .E(n293), .F(n1705), .Y(n1707) );
  MUX2X1 U94 ( .D0(memrd), .D1(n2650), .S(n420), .Y(memrd_comb) );
  OA222X1 U95 ( .A(n27), .B(n2496), .C(n2852), .D(n26), .E(n2337), .F(n2423), 
        .Y(n299) );
  NAND32X1 U96 ( .B(dec_accop[11]), .C(n1068), .A(n1065), .Y(n1051) );
  OA222X1 U97 ( .A(n2259), .B(n2423), .C(n26), .D(n2260), .E(n27), .F(n2261), 
        .Y(n2113) );
  OAI221X1 U98 ( .A(n1347), .B(n2028), .C(n1034), .D(n185), .E(n2106), .Y(
        n2112) );
  INVX1 U99 ( .A(n2667), .Y(n104) );
  INVX1 U100 ( .A(n498), .Y(n928) );
  NAND21X1 U101 ( .B(dec_accop[8]), .A(n1763), .Y(n1080) );
  AOI221XL U102 ( .A(rn_reg[77]), .B(n173), .C(rn_reg[29]), .D(n195), .E(n847), 
        .Y(n863) );
  AOI221XL U103 ( .A(rn_reg[205]), .B(n173), .C(rn_reg[157]), .D(n195), .E(
        n832), .Y(n867) );
  AO21X1 U104 ( .B(ramdatao[1]), .C(n1906), .A(n1056), .Y(n1088) );
  AOI221XL U105 ( .A(rn_reg[78]), .B(n173), .C(rn_reg[30]), .D(n195), .E(n900), 
        .Y(n916) );
  AOI221XL U106 ( .A(rn_reg[206]), .B(n173), .C(rn_reg[158]), .D(n195), .E(
        n885), .Y(n920) );
  OA222X1 U107 ( .A(n2390), .B(n2423), .C(n27), .D(n2391), .E(n2854), .F(n26), 
        .Y(n2309) );
  OA222X1 U108 ( .A(n27), .B(n2304), .C(n2853), .D(n2422), .E(n2303), .F(n2423), .Y(n298) );
  NAND2X1 U109 ( .A(n1910), .B(n2201), .Y(n1902) );
  AOI221XL U110 ( .A(rn_reg[79]), .B(n975), .C(rn_reg[31]), .D(n974), .E(n973), 
        .Y(n1003) );
  AOI221XL U111 ( .A(rn_reg[207]), .B(n975), .C(rn_reg[159]), .D(n974), .E(
        n954), .Y(n1007) );
  MUX2IX1 U112 ( .D0(n1412), .D1(n2278), .S(n1537), .Y(n226) );
  AO2222XL U113 ( .A(n2611), .B(n2767), .C(n2607), .D(n2769), .E(n2610), .F(
        n2768), .G(n2606), .H(n2770), .Y(n1408) );
  MUX2IX1 U114 ( .D0(n1485), .D1(n2277), .S(n1537), .Y(n224) );
  NAND21X1 U115 ( .B(n2871), .A(n151), .Y(n1953) );
  INVX1 U116 ( .A(n951), .Y(n511) );
  INVX1 U117 ( .A(n2112), .Y(n8) );
  AND2X1 U118 ( .A(n99), .B(n1022), .Y(n262) );
  INVX1 U119 ( .A(n2431), .Y(n1041) );
  NAND21X1 U120 ( .B(n2866), .A(n1124), .Y(n2012) );
  INVX1 U121 ( .A(n2042), .Y(n2044) );
  MUX2BXL U122 ( .D0(n2032), .D1(n2031), .S(codefetch_s), .Y(n2045) );
  OA222X1 U123 ( .A(n2306), .B(n2423), .C(n27), .D(n2305), .E(n2855), .F(n2422), .Y(n2308) );
  INVX1 U124 ( .A(n500), .Y(n1098) );
  INVX1 U125 ( .A(n1357), .Y(n501) );
  INVX1 U126 ( .A(ramsfraddr[1]), .Y(n2561) );
  INVX1 U127 ( .A(temp2_comb[0]), .Y(n2094) );
  AO21X1 U128 ( .B(n1258), .C(n1343), .A(n1257), .Y(n1269) );
  MUX2AXL U129 ( .D0(rs[0]), .D1(n2275), .S(n1775), .Y(n783) );
  INVX1 U130 ( .A(n2595), .Y(n1252) );
  INVX1 U131 ( .A(dec_accop[10]), .Y(n1763) );
  AOI221XL U132 ( .A(rn_reg[202]), .B(n173), .C(rn_reg[154]), .D(n195), .E(
        n533), .Y(n649) );
  AOI221XL U133 ( .A(rn_reg[74]), .B(n173), .C(rn_reg[26]), .D(n195), .E(n565), 
        .Y(n645) );
  MUX2AXL U134 ( .D0(sp[0]), .D1(n2278), .S(n947), .Y(n785) );
  MUX2BXL U135 ( .D0(sp[1]), .D1(n2277), .S(n947), .Y(n332) );
  INVX1 U136 ( .A(acc[2]), .Y(n2263) );
  INVX1 U137 ( .A(N13353), .Y(n1197) );
  OA222X1 U138 ( .A(n1918), .B(n1964), .C(n1749), .D(n2257), .E(n293), .F(
        n1748), .Y(n1750) );
  INVX1 U139 ( .A(n1960), .Y(n1132) );
  NAND21X1 U140 ( .B(n2573), .A(n1252), .Y(n1410) );
  NAND21X1 U141 ( .B(b[7]), .A(n2193), .Y(n2194) );
  NAND41X1 U142 ( .D(n2554), .A(n313), .B(ramsfrwe), .C(ramsfraddr[6]), .Y(
        n1816) );
  INVX1 U143 ( .A(ramsfraddr[5]), .Y(n2555) );
  NAND21X1 U144 ( .B(ramsfraddr[3]), .A(ramsfraddr[4]), .Y(n2594) );
  OA222X1 U145 ( .A(n2062), .B(n2285), .C(n2303), .D(n2061), .E(n2060), .F(
        n2313), .Y(n1806) );
  NAND21X1 U146 ( .B(n1041), .A(n2440), .Y(n1224) );
  NAND21X1 U147 ( .B(n1721), .A(n2015), .Y(n2011) );
  INVX1 U148 ( .A(n2439), .Y(n2103) );
  NAND32X1 U149 ( .B(n186), .C(n419), .A(n502), .Y(n2431) );
  INVX1 U150 ( .A(n1287), .Y(n502) );
  OA222X1 U151 ( .A(interrupt), .B(n1166), .C(instr[0]), .D(n483), .E(instr[7]), .F(n1018), .Y(n489) );
  NAND21X1 U152 ( .B(n2045), .A(n2044), .Y(n2455) );
  OR2X1 U153 ( .A(n73), .B(n2041), .Y(n2458) );
  INVX1 U154 ( .A(n2170), .Y(n73) );
  NAND2X1 U155 ( .A(n2045), .B(n2044), .Y(n2460) );
  INVX1 U156 ( .A(n1224), .Y(n1100) );
  MUX2X1 U157 ( .D0(ramsfraddr[1]), .D1(n79), .S(waitstaten), .Y(
        ramsfraddr_comb[1]) );
  OA222X1 U158 ( .A(n2062), .B(n2180), .C(n2390), .D(n2061), .E(n2060), .F(
        n2396), .Y(n1698) );
  INVX1 U159 ( .A(n2867), .Y(n1124) );
  INVX1 U160 ( .A(n1869), .Y(n92) );
  OA222X1 U161 ( .A(n2062), .B(n1297), .C(n2472), .D(n2061), .E(n2060), .F(
        n2459), .Y(n1153) );
  INVX1 U162 ( .A(n1269), .Y(n2084) );
  NOR2X1 U163 ( .A(n1323), .B(n325), .Y(n324) );
  NAND5XL U164 ( .A(n1910), .B(n1909), .C(n1769), .D(n1791), .E(n1768), .Y(
        n1819) );
  MUX2X1 U165 ( .D0(n1489), .D1(n2278), .S(n1256), .Y(n1509) );
  AND2X1 U166 ( .A(n946), .B(n740), .Y(n742) );
  INVX1 U167 ( .A(temp2_comb[4]), .Y(n2396) );
  INVX1 U168 ( .A(ramdatao[4]), .Y(n2628) );
  GEN2XL U169 ( .D(n2845), .E(pc_o[5]), .C(n1531), .B(memaddr[6]), .A(n1524), 
        .Y(n1525) );
  OA222X1 U170 ( .A(n2062), .B(n2165), .C(n2306), .D(n2061), .E(n2060), .F(
        n2160), .Y(n1709) );
  MUX2AXL U171 ( .D0(n925), .D1(n924), .S(n1176), .Y(n225) );
  OAI31XL U172 ( .A(n495), .B(n2535), .C(n2522), .D(mempsrd), .Y(n2517) );
  ENOX1 U173 ( .A(n1183), .B(n2285), .C(n653), .D(n1179), .Y(n2183) );
  INVX1 U174 ( .A(n63), .Y(n2642) );
  AND2X1 U175 ( .A(n378), .B(n1614), .Y(N10574) );
  OAI21BBX1 U176 ( .A(n2185), .B(n1218), .C(n2), .Y(n1184) );
  NOR32X4 U177 ( .B(n422), .C(n2679), .A(n2678), .Y(n84) );
  NAND2X1 U178 ( .A(n3), .B(n8), .Y(n11) );
  INVX1 U179 ( .A(n258), .Y(n3) );
  NOR21X2 U180 ( .B(n1202), .A(n98), .Y(n258) );
  MUX2IXL U181 ( .D0(n57), .D1(n110), .S(n2690), .Y(memaddr_comb[2]) );
  NAND21X1 U182 ( .B(n2662), .A(n2661), .Y(n2663) );
  OA33X1 U183 ( .A(ramsfraddr[7]), .B(n1447), .C(n1149), .D(n1129), .E(n1128), 
        .F(n1146), .Y(n12) );
  AOI21X1 U184 ( .B(n1021), .C(n1047), .A(n1037), .Y(n13) );
  INVX1 U185 ( .A(n2869), .Y(n418) );
  INVX1 U186 ( .A(n418), .Y(instr[4]) );
  INVX1 U187 ( .A(n2205), .Y(n294) );
  INVX1 U188 ( .A(n2132), .Y(n72) );
  NAND2X1 U189 ( .A(n72), .B(stop), .Y(n14) );
  MUX2AXL U190 ( .D0(rs[1]), .D1(n2628), .S(n1775), .Y(n1254) );
  NOR2X1 U191 ( .A(n1033), .B(n1032), .Y(n15) );
  AO21X1 U192 ( .B(n1009), .C(n2277), .A(n826), .Y(n2472) );
  INVX1 U193 ( .A(n2472), .Y(n96) );
  INVX1 U194 ( .A(n2112), .Y(n2428) );
  NOR4XL U195 ( .A(n2449), .B(n2448), .C(n2447), .D(n239), .Y(n17) );
  NOR4XL U196 ( .A(n2349), .B(n2348), .C(n2347), .D(n240), .Y(n18) );
  NAND32X1 U197 ( .B(ramsfraddr[2]), .C(ramsfraddr[0]), .A(n2561), .Y(n2134)
         );
  INVX1 U198 ( .A(n2134), .Y(n313) );
  AOI21X1 U199 ( .B(n179), .C(n48), .A(n383), .Y(n19) );
  AOI21X1 U200 ( .B(n1225), .C(pc_i[9]), .A(n1572), .Y(n20) );
  AOI21X1 U201 ( .B(n1225), .C(pc_i[15]), .A(n1550), .Y(n21) );
  AOI21X1 U202 ( .B(n1225), .C(pc_i[11]), .A(n1568), .Y(n22) );
  AOI21X1 U203 ( .B(n1225), .C(pc_i[13]), .A(n1564), .Y(n23) );
  INVX1 U204 ( .A(n441), .Y(n422) );
  INVXL U205 ( .A(n13), .Y(n24) );
  INVXL U206 ( .A(n2422), .Y(n25) );
  INVXL U207 ( .A(n25), .Y(n26) );
  INVXL U208 ( .A(n15), .Y(n27) );
  INVXL U209 ( .A(n1979), .Y(n28) );
  INVXL U210 ( .A(n1979), .Y(n29) );
  INVXL U211 ( .A(n1978), .Y(n30) );
  INVXL U212 ( .A(n1978), .Y(n31) );
  INVXL U213 ( .A(pc_o[15]), .Y(n32) );
  INVXL U214 ( .A(n32), .Y(memaddr[15]) );
  INVXL U215 ( .A(n1283), .Y(n34) );
  INVXL U216 ( .A(n34), .Y(n35) );
  INVXL U217 ( .A(n48), .Y(n36) );
  INVXL U218 ( .A(pc_o[7]), .Y(n37) );
  INVXL U219 ( .A(n37), .Y(memaddr[7]) );
  INVXL U220 ( .A(pc_o[4]), .Y(n39) );
  INVXL U221 ( .A(n39), .Y(memaddr[4]) );
  INVXL U222 ( .A(pc_o[12]), .Y(n41) );
  INVXL U223 ( .A(n41), .Y(memaddr[12]) );
  INVXL U224 ( .A(pc_o[6]), .Y(n43) );
  INVXL U225 ( .A(n43), .Y(memaddr[6]) );
  INVXL U226 ( .A(pc_o[5]), .Y(n45) );
  INVXL U227 ( .A(n45), .Y(memaddr[5]) );
  INVXL U228 ( .A(n2482), .Y(n47) );
  INVXL U229 ( .A(n47), .Y(n48) );
  INVXL U230 ( .A(pc_o[13]), .Y(n49) );
  INVXL U231 ( .A(n49), .Y(memaddr[13]) );
  INVXL U232 ( .A(pc_o[8]), .Y(n51) );
  INVXL U233 ( .A(n51), .Y(memaddr[8]) );
  INVXL U234 ( .A(memaddr[1]), .Y(n53) );
  INVXL U235 ( .A(n53), .Y(pc_o[1]) );
  INVXL U236 ( .A(n19), .Y(n55) );
  INVXL U237 ( .A(n19), .Y(n56) );
  INVXL U238 ( .A(pc_o[2]), .Y(n57) );
  INVXL U239 ( .A(n57), .Y(memaddr[2]) );
  INVXL U240 ( .A(pc_o[3]), .Y(n59) );
  INVXL U241 ( .A(n59), .Y(memaddr[3]) );
  INVXL U242 ( .A(n2865), .Y(n61) );
  INVXL U243 ( .A(n61), .Y(memaddr[0]) );
  GEN2X1 U244 ( .D(n1955), .E(n1949), .C(n1948), .B(n1947), .A(n1946), .Y(
        n1977) );
  ENOXL U245 ( .A(n1184), .B(n2180), .C(n1178), .D(n1179), .Y(n2640) );
  NAND21XL U246 ( .B(n2237), .A(n2455), .Y(n2484) );
  INVXL U247 ( .A(n2455), .Y(n2238) );
  AOI22CXL U248 ( .C(n923), .D(n1179), .A(n2491), .B(n1184), .Y(n63) );
  OAI21AX1 U249 ( .B(n1435), .C(n2459), .A(n1428), .Y(n274) );
  BUFXL U250 ( .A(n2636), .Y(n64) );
  BUFXL U251 ( .A(memdatai[4]), .Y(n65) );
  EORXL U252 ( .A(sfrdatai[2]), .B(n1037), .C(n24), .D(n2260), .Y(n66) );
  AO2222XL U253 ( .A(alu_out[1]), .B(n2481), .C(memdatai[1]), .D(n2454), .E(
        n2453), .F(ramdatai[1]), .G(n2452), .H(n96), .Y(n2462) );
  AO2222XL U254 ( .A(alu_out[2]), .B(n2481), .C(memdatai[2]), .D(n2454), .E(
        n2452), .F(n2148), .G(n2453), .H(ramdatai[2]), .Y(n2151) );
  AO2222XL U255 ( .A(alu_out[0]), .B(n2481), .C(memdatai[0]), .D(n2454), .E(
        n2453), .F(ramdatai[0]), .G(n2452), .H(n2091), .Y(n2096) );
  ENOX1 U256 ( .A(n86), .B(n2264), .C(n94), .D(n2669), .Y(n271) );
  INVX1 U257 ( .A(n653), .Y(n2505) );
  AOI21AX1 U258 ( .B(n1704), .C(n333), .A(n68), .Y(n216) );
  BUFXL U259 ( .A(n67), .Y(n69) );
  OAI221X1 U260 ( .A(n1965), .B(n1874), .C(n2411), .D(n1873), .E(n1872), .Y(
        n1875) );
  INVXL U261 ( .A(n2285), .Y(n70) );
  NAND8X1 U262 ( .A(n2636), .B(n2638), .C(n1187), .D(n63), .E(n2637), .F(n1186), .G(sfrwe_comb_s), .H(n1185), .Y(n2666) );
  INVX3 U263 ( .A(sfrdatai[0]), .Y(n2230) );
  INVX2 U264 ( .A(n2666), .Y(n2132) );
  NAND32X1 U265 ( .B(n1174), .C(n1172), .A(n1218), .Y(n1183) );
  OA222XL U266 ( .A(n2062), .B(n2491), .C(n2337), .D(n2061), .E(n2060), .F(
        n2344), .Y(n2063) );
  BUFXL U267 ( .A(n2618), .Y(n71) );
  NAND5X1 U268 ( .A(n36), .B(n2040), .C(n2169), .D(n2168), .E(n2039), .Y(n2041) );
  ENOX1 U269 ( .A(n2230), .B(n2314), .C(ramdatai[0]), .D(n13), .Y(n1200) );
  BUFXL U270 ( .A(n66), .Y(n74) );
  AND2XL U271 ( .A(n386), .B(n2639), .Y(N11481) );
  INVXL U272 ( .A(sfrdatai[2]), .Y(n2261) );
  AO22AX1 U273 ( .A(n1867), .B(n77), .C(n75), .D(n1868), .Y(n2207) );
  INVXL U274 ( .A(n2165), .Y(n76) );
  NAND2X1 U275 ( .A(n1037), .B(sfrdatai[1]), .Y(n99) );
  OA21X1 U276 ( .B(n270), .C(n271), .A(n2319), .Y(n269) );
  NOR32X4 U277 ( .B(n2679), .C(n422), .A(n2678), .Y(n2690) );
  OAI221XL U278 ( .A(n1388), .B(n185), .C(n2644), .D(n1387), .E(n2645), .Y(n78) );
  AND2XL U279 ( .A(n386), .B(n2642), .Y(N11484) );
  BUFXL U280 ( .A(n2637), .Y(n79) );
  BUFXL U281 ( .A(n2662), .Y(n80) );
  INVXL U282 ( .A(n2491), .Y(n81) );
  AO2222XL U283 ( .A(alu_out[3]), .B(n2481), .C(n76), .D(n2454), .E(
        ramdatai[3]), .F(n2453), .G(n2452), .H(n2157), .Y(n2156) );
  BUFXL U284 ( .A(n258), .Y(n82) );
  EORX1 U285 ( .A(n95), .B(n1037), .C(n2227), .D(n24), .Y(n83) );
  INVX2 U286 ( .A(n2230), .Y(n95) );
  INVX4 U287 ( .A(n2677), .Y(n2678) );
  OAI22X1 U288 ( .A(n272), .B(n1747), .C(n1429), .D(n326), .Y(n85) );
  EORX1 U289 ( .A(sfrdatai[2]), .B(n1037), .C(n24), .D(n2260), .Y(n86) );
  MUX2X1 U290 ( .D0(memaddr[4]), .D1(n2684), .S(n84), .Y(memaddr_comb[4]) );
  MUX2BX1 U291 ( .D0(pc_o[3]), .D1(n101), .S(n84), .Y(memaddr_comb[3]) );
  AOI21AXL U292 ( .B(n103), .C(n15), .A(n107), .Y(n87) );
  INVX1 U293 ( .A(n1201), .Y(n107) );
  NAND32X2 U294 ( .B(n72), .C(n2676), .A(n2663), .Y(n2679) );
  INVXL U295 ( .A(n2660), .Y(n89) );
  OA222X1 U296 ( .A(n2201), .B(n90), .C(n1831), .D(n91), .E(n92), .F(n93), .Y(
        n1872) );
  XNOR2X1 U297 ( .A(n2207), .B(n1866), .Y(n93) );
  INVX3 U298 ( .A(n1913), .Y(n1435) );
  AOI211X4 U299 ( .C(sfrdatai[0]), .D(n15), .A(n2430), .B(n1203), .Y(n1204) );
  OAI22X1 U300 ( .A(n2230), .B(n2314), .C(n2227), .D(n24), .Y(n94) );
  AO222X1 U301 ( .A(sfrdatai[1]), .B(n15), .C(n25), .D(ramdatai[1]), .E(n96), 
        .F(n1033), .Y(n2110) );
  AND2XL U302 ( .A(n1447), .B(n69), .Y(n1450) );
  INVX1 U303 ( .A(n2682), .Y(n110) );
  INVXL U304 ( .A(n2686), .Y(n105) );
  INVX2 U305 ( .A(n2481), .Y(n2169) );
  NAND32X1 U306 ( .B(n2660), .C(n97), .A(n2658), .Y(n2661) );
  NAND21X2 U307 ( .B(n269), .A(n2673), .Y(n2674) );
  NAND21XL U308 ( .B(n2065), .A(n95), .Y(n1245) );
  NAND2X2 U309 ( .A(n2664), .B(n104), .Y(n100) );
  INVX1 U310 ( .A(n2683), .Y(n101) );
  AOI21AX1 U311 ( .B(sfrdatai[0]), .C(n15), .A(n107), .Y(n98) );
  OA33X1 U312 ( .A(n1037), .B(n2419), .C(n1036), .D(sfrdatai[1]), .E(n2419), 
        .F(n1036), .Y(n1107) );
  NAND6X2 U313 ( .A(n1206), .B(n1208), .C(n2623), .D(n2515), .E(n2132), .F(
        n1222), .Y(n2664) );
  NAND3X4 U314 ( .A(n100), .B(n2674), .C(n14), .Y(n2675) );
  MUX2IX1 U315 ( .D0(n61), .D1(n109), .S(n88), .Y(memaddr_comb[0]) );
  XOR2X1 U316 ( .A(n102), .B(n2110), .Y(n1035) );
  BUFXL U317 ( .A(n95), .Y(n103) );
  INVX1 U318 ( .A(n2681), .Y(n106) );
  MUX2IX1 U319 ( .D0(n43), .D1(n105), .S(n88), .Y(memaddr_comb[6]) );
  NAND21XL U320 ( .B(n71), .A(n373), .Y(n1217) );
  INVX1 U321 ( .A(n2680), .Y(n109) );
  NOR21XL U322 ( .B(n2332), .A(n1200), .Y(n108) );
  AOI31X1 U323 ( .A(n364), .B(n2384), .C(n2119), .D(n83), .Y(n363) );
  INVXL U324 ( .A(n108), .Y(n1227) );
  OA22X1 U325 ( .A(n2474), .B(n1889), .C(n2065), .D(n1305), .Y(n1154) );
  MUX2XL U326 ( .D0(n2412), .D1(n199), .S(n74), .Y(n2269) );
  OAI21X1 U327 ( .B(n2665), .C(n262), .A(n1023), .Y(n270) );
  NAND21X2 U328 ( .B(n2676), .A(n2675), .Y(n2677) );
  AOI21X1 U329 ( .B(n147), .C(n48), .A(n382), .Y(n1608) );
  INVX1 U330 ( .A(n1608), .Y(n111) );
  INVX1 U331 ( .A(n1608), .Y(n112) );
  BUFX3 U332 ( .A(n1602), .Y(n113) );
  AOI21X1 U333 ( .B(n2604), .C(n2482), .A(n383), .Y(n1592) );
  INVX1 U334 ( .A(n1592), .Y(n114) );
  INVX1 U335 ( .A(n1592), .Y(n115) );
  INVX1 U336 ( .A(n1629), .Y(n116) );
  NAND21X1 U337 ( .B(n204), .A(n1617), .Y(n1655) );
  BUFX3 U338 ( .A(n1609), .Y(n117) );
  AOI21X1 U339 ( .B(n2608), .C(n48), .A(n383), .Y(n2087) );
  INVX1 U340 ( .A(n2087), .Y(n118) );
  INVX1 U341 ( .A(n2087), .Y(n119) );
  INVX1 U342 ( .A(n2868), .Y(n120) );
  INVX1 U343 ( .A(n169), .Y(instr[0]) );
  BUFX3 U344 ( .A(n1593), .Y(n122) );
  AOI21X1 U345 ( .B(n2605), .C(n2482), .A(n383), .Y(n1594) );
  INVX1 U346 ( .A(n1594), .Y(n123) );
  INVX1 U347 ( .A(n1594), .Y(n124) );
  INVX1 U348 ( .A(n2849), .Y(pc_o[11]) );
  INVX1 U349 ( .A(n1787), .Y(n126) );
  NAND21X1 U350 ( .B(n2870), .A(n2872), .Y(n1725) );
  BUFX3 U351 ( .A(n2088), .Y(n127) );
  AOI21X1 U352 ( .B(n2609), .C(n2482), .A(n383), .Y(n2280) );
  INVX1 U353 ( .A(n2280), .Y(n128) );
  INVX1 U354 ( .A(n2280), .Y(n129) );
  BUFX3 U355 ( .A(n991), .Y(n130) );
  BUFXL U356 ( .A(n2481), .Y(n131) );
  INVX1 U357 ( .A(n2801), .Y(n132) );
  INVX1 U358 ( .A(n132), .Y(n133) );
  INVX1 U359 ( .A(n132), .Y(n134) );
  INVX1 U360 ( .A(n2275), .Y(n135) );
  INVX1 U361 ( .A(ramdatao[3]), .Y(n2275) );
  AO21XL U362 ( .B(ramdatao[3]), .C(n1906), .A(n1701), .Y(n1708) );
  INVX1 U363 ( .A(n1033), .Y(n136) );
  INVX1 U364 ( .A(n1124), .Y(instr[6]) );
  NAND21X1 U365 ( .B(n2867), .A(instr[7]), .Y(n1166) );
  BUFX3 U366 ( .A(n1595), .Y(n138) );
  AOI21X1 U367 ( .B(n163), .C(n48), .A(n383), .Y(n1596) );
  INVX1 U368 ( .A(n1596), .Y(n139) );
  INVX1 U369 ( .A(n1596), .Y(n140) );
  OR2X1 U370 ( .A(n536), .B(n547), .Y(n141) );
  OAI221XL U371 ( .A(n156), .B(n744), .C(n970), .D(n743), .E(n220), .Y(n745)
         );
  OR2X1 U372 ( .A(n536), .B(n547), .Y(n970) );
  NAND21X1 U373 ( .B(n2873), .A(n2182), .Y(n536) );
  BUFX3 U374 ( .A(n993), .Y(n142) );
  BUFX3 U375 ( .A(n979), .Y(n143) );
  INVX1 U376 ( .A(n1157), .Y(instr[1]) );
  INVX1 U377 ( .A(n2604), .Y(n145) );
  OA2222XL U378 ( .A(dpl_reg[8]), .B(n1584), .C(dpl_reg[0]), .D(n1583), .E(
        dpl_reg[40]), .F(n1582), .G(dpl_reg[32]), .H(n1581), .Y(n1407) );
  OA2222XL U379 ( .A(dpl_reg[9]), .B(n1584), .C(dpl_reg[1]), .D(n1583), .E(
        dpl_reg[41]), .F(n1582), .G(dpl_reg[33]), .H(n1581), .Y(n1483) );
  NAND2X1 U380 ( .A(n1509), .B(n1271), .Y(n1583) );
  INVX1 U381 ( .A(n2489), .Y(pc_o[14]) );
  INVX1 U382 ( .A(n1552), .Y(n147) );
  INVX1 U383 ( .A(n2802), .Y(n148) );
  INVX1 U384 ( .A(n148), .Y(n149) );
  INVX1 U385 ( .A(n1903), .Y(n150) );
  BUFXL U386 ( .A(n2870), .Y(instr[3]) );
  INVX1 U387 ( .A(instr[3]), .Y(n151) );
  INVX1 U388 ( .A(instr[3]), .Y(n152) );
  BUFX3 U389 ( .A(n2282), .Y(n153) );
  AOI21X1 U390 ( .B(n203), .C(n2482), .A(n383), .Y(n1598) );
  INVX1 U391 ( .A(n1598), .Y(n154) );
  INVX1 U392 ( .A(n1598), .Y(n155) );
  NOR2XL U393 ( .A(n554), .B(n536), .Y(n972) );
  INVX1 U394 ( .A(n972), .Y(n156) );
  INVX1 U395 ( .A(n972), .Y(n157) );
  BUFX3 U396 ( .A(n987), .Y(n158) );
  BUFX3 U397 ( .A(n997), .Y(n159) );
  BUFX3 U398 ( .A(n981), .Y(n160) );
  INVX1 U399 ( .A(n2850), .Y(pc_o[9]) );
  INVX1 U400 ( .A(n2605), .Y(n162) );
  INVX1 U401 ( .A(n1551), .Y(n163) );
  INVX1 U402 ( .A(n2798), .Y(n164) );
  INVX1 U403 ( .A(n164), .Y(n165) );
  INVX1 U404 ( .A(n164), .Y(n166) );
  INVX1 U405 ( .A(n213), .Y(n167) );
  NAND21X1 U406 ( .B(n2028), .A(n501), .Y(n2439) );
  INVX1 U407 ( .A(n2195), .Y(n168) );
  BUFX3 U408 ( .A(n1626), .Y(n169) );
  INVX1 U409 ( .A(n1965), .Y(n170) );
  XOR2XL U410 ( .A(n1436), .B(acc[0]), .Y(n1422) );
  BUFX3 U411 ( .A(n1599), .Y(n171) );
  INVX1 U412 ( .A(n1923), .Y(n172) );
  INVX1 U413 ( .A(n524), .Y(n173) );
  NAND21XL U414 ( .B(n547), .A(n538), .Y(n524) );
  BUFX3 U415 ( .A(n989), .Y(n174) );
  BUFX3 U416 ( .A(n995), .Y(n175) );
  BUFX3 U417 ( .A(n977), .Y(n176) );
  NAND21X1 U418 ( .B(n545), .A(n539), .Y(n977) );
  INVX1 U419 ( .A(n1216), .Y(n177) );
  INVX1 U420 ( .A(n2609), .Y(n178) );
  INVX1 U421 ( .A(n1541), .Y(n179) );
  INVX1 U422 ( .A(n2800), .Y(n180) );
  INVX1 U423 ( .A(n180), .Y(n181) );
  INVX1 U424 ( .A(n180), .Y(n182) );
  BUFXL U425 ( .A(n2866), .Y(n183) );
  BUFX1 U426 ( .A(n2866), .Y(instr[7]) );
  BUFX3 U427 ( .A(phase[0]), .Y(n2549) );
  INVX1 U428 ( .A(n2549), .Y(n185) );
  INVX1 U429 ( .A(n2549), .Y(n186) );
  INVX1 U430 ( .A(n2549), .Y(n187) );
  OAI211X1 U431 ( .C(n504), .D(n187), .A(n511), .B(n2645), .Y(n1013) );
  INVX1 U432 ( .A(n2440), .Y(n188) );
  NAND32X1 U433 ( .B(n2022), .C(n2647), .A(n1622), .Y(n2440) );
  INVX1 U434 ( .A(n2864), .Y(n189) );
  INVX1 U435 ( .A(n189), .Y(mempswr) );
  BUFX3 U436 ( .A(n1845), .Y(n191) );
  INVX1 U437 ( .A(n1721), .Y(instr[2]) );
  NAND21X1 U438 ( .B(instr[4]), .A(n2871), .Y(n1117) );
  INVX1 U439 ( .A(n1964), .Y(n193) );
  BUFX3 U440 ( .A(n1597), .Y(n194) );
  INVX1 U441 ( .A(n526), .Y(n195) );
  BUFX3 U442 ( .A(n999), .Y(n196) );
  BUFX3 U443 ( .A(n985), .Y(n197) );
  BUFX3 U444 ( .A(n983), .Y(n198) );
  NAND21X1 U445 ( .B(n1972), .A(n2037), .Y(n199) );
  NAND21XL U446 ( .B(n1953), .A(n1612), .Y(n1972) );
  INVX1 U447 ( .A(n1266), .Y(n200) );
  INVX1 U448 ( .A(n2608), .Y(n201) );
  AO21X1 U449 ( .B(n1258), .C(n2182), .A(n1253), .Y(n1272) );
  INVX1 U450 ( .A(n2255), .Y(pc_o[10]) );
  INVX1 U451 ( .A(n1542), .Y(n203) );
  AO2222XL U452 ( .A(n2606), .B(n2774), .C(n2607), .D(n2773), .E(n2610), .F(
        n2772), .G(n2611), .H(n2771), .Y(n1484) );
  BUFX3 U453 ( .A(n2868), .Y(n204) );
  BUFX3 U454 ( .A(n2868), .Y(instr[5]) );
  INVX1 U455 ( .A(dps[2]), .Y(n206) );
  INVX1 U456 ( .A(n206), .Y(n207) );
  INVX1 U457 ( .A(n206), .Y(n209) );
  INVX1 U458 ( .A(phase[1]), .Y(n212) );
  INVX1 U459 ( .A(n212), .Y(n213) );
  INVX1 U460 ( .A(n212), .Y(n214) );
  GEN2XL U461 ( .D(n2038), .E(n2037), .C(n2538), .B(n214), .A(n2036), .Y(n2170) );
  INVX1 U462 ( .A(n213), .Y(n2028) );
  NAND21XL U463 ( .B(n498), .A(n1028), .Y(n499) );
  NAND21XL U464 ( .B(n1254), .A(n561), .Y(n562) );
  MUX2X1 U465 ( .D0(N13337), .D1(divtempreg[0]), .S(N13343), .Y(n315) );
  AO21X1 U466 ( .B(n946), .C(n872), .A(n870), .Y(n922) );
  NAND21X1 U467 ( .B(n528), .A(n535), .Y(n554) );
  INVXL U468 ( .A(n2871), .Y(n1721) );
  NAND21XL U469 ( .B(n535), .A(n528), .Y(n556) );
  INVX3 U470 ( .A(n695), .Y(n1173) );
  OAI221XL U471 ( .A(n157), .B(n971), .C(n141), .D(n969), .E(n968), .Y(n973)
         );
  AO2222XL U472 ( .A(n2353), .B(n1013), .C(n1012), .D(n2362), .E(temp[7]), .F(
        n1011), .G(n1010), .H(ramsfraddr[7]), .Y(n2504) );
  NAND21XL U473 ( .B(n1248), .A(n2644), .Y(n1180) );
  XOR2X1 U474 ( .A(n1178), .B(n1182), .Y(n877) );
  INVX1 U475 ( .A(n1977), .Y(n277) );
  INVX1 U476 ( .A(n291), .Y(n2430) );
  MUX2IXL U477 ( .D0(n787), .D1(n786), .S(n332), .Y(n227) );
  INVX1 U478 ( .A(n418), .Y(n416) );
  AO21X4 U479 ( .B(n1009), .C(n2275), .A(n781), .Y(n2306) );
  NAND42X1 U480 ( .C(n1751), .D(n231), .A(n285), .B(n1750), .Y(n1939) );
  AO21X1 U481 ( .B(n1009), .C(n2633), .A(n1008), .Y(n2424) );
  AO21X1 U482 ( .B(n1009), .C(n2630), .A(n868), .Y(n2303) );
  INVX1 U483 ( .A(n1166), .Y(n1384) );
  MUX2BXL U484 ( .D0(N13336), .D1(n2411), .S(N13343), .Y(n312) );
  INVX1 U485 ( .A(accactv), .Y(n1845) );
  INVX1 U486 ( .A(n546), .Y(n555) );
  MUX2IXL U487 ( .D0(n329), .D1(n330), .S(n1256), .Y(n1257) );
  NAND21X1 U488 ( .B(n1657), .A(n1989), .Y(n1956) );
  INVXL U489 ( .A(n1657), .Y(n1781) );
  NAND21X1 U490 ( .B(n554), .A(n538), .Y(n979) );
  AO21X1 U491 ( .B(n1615), .C(n1629), .A(n1971), .Y(n2108) );
  INVX1 U492 ( .A(n2623), .Y(n2624) );
  INVX1 U493 ( .A(n2356), .Y(n1256) );
  INVX1 U494 ( .A(n1764), .Y(n1918) );
  AO21X1 U495 ( .B(n1198), .C(n1940), .A(n2624), .Y(n1102) );
  INVX1 U496 ( .A(n505), .Y(n1990) );
  AND2X1 U497 ( .A(n437), .B(n2697), .Y(n438) );
  OA222X1 U498 ( .A(n1984), .B(n2526), .C(n1975), .D(n212), .E(n2528), .F(
        n2000), .Y(n280) );
  INVXL U499 ( .A(n1313), .Y(n693) );
  NAND21X1 U500 ( .B(n553), .A(n555), .Y(n997) );
  NAND21XL U501 ( .B(n545), .A(n544), .Y(n987) );
  NAND21XL U502 ( .B(n556), .A(n555), .Y(n993) );
  NAND21X1 U503 ( .B(n325), .A(n1731), .Y(n1374) );
  INVX1 U504 ( .A(n696), .Y(n286) );
  INVX1 U505 ( .A(n534), .Y(n528) );
  NAND21X1 U506 ( .B(n1370), .A(n473), .Y(n2315) );
  GEN2XL U507 ( .D(n1092), .E(n1091), .C(n2028), .B(n1090), .A(n1089), .Y(
        n2656) );
  INVX1 U508 ( .A(n1973), .Y(n1944) );
  NAND21XL U509 ( .B(n120), .A(n1617), .Y(n1959) );
  NAND21X1 U510 ( .B(n1941), .A(n1896), .Y(n465) );
  INVX1 U511 ( .A(n2517), .Y(codefetch_s) );
  AND2XL U512 ( .A(n944), .B(n943), .Y(n950) );
  AO21X1 U513 ( .B(n1438), .C(n1910), .A(n2438), .Y(n1439) );
  AOI221X1 U514 ( .A(acc[3]), .B(n1907), .C(multemp2[1]), .D(n2192), .E(n1441), 
        .Y(n1442) );
  MUX2IX1 U515 ( .D0(n309), .D1(n310), .S(n422), .Y(ramwe_comb) );
  INVX2 U516 ( .A(dec_accop[6]), .Y(n1078) );
  MUX2XL U517 ( .D0(N13338), .D1(divtempreg[1]), .S(N13343), .Y(n316) );
  INVXL U518 ( .A(n2873), .Y(n1626) );
  OA2222XL U519 ( .A(dpl_reg[10]), .B(n1584), .C(dpl_reg[2]), .D(n1583), .E(
        dpl_reg[42]), .F(n1582), .G(dpl_reg[34]), .H(n1581), .Y(n1480) );
  INVXL U520 ( .A(n444), .Y(n1731) );
  INVX1 U521 ( .A(ramdatao[0]), .Y(n2278) );
  NAND2X1 U522 ( .A(n207), .B(n1255), .Y(n329) );
  INVXL U523 ( .A(instr[5]), .Y(n1941) );
  INVX1 U524 ( .A(dps[3]), .Y(n1255) );
  AO21XL U525 ( .B(n384), .C(n163), .A(n428), .Y(N12547) );
  INVXL U526 ( .A(n1043), .Y(n1983) );
  NAND21XL U527 ( .B(n1657), .A(n928), .Y(n1038) );
  INVXL U528 ( .A(n1044), .Y(n1346) );
  INVXL U529 ( .A(n869), .Y(n1012) );
  NAND2XL U530 ( .A(n509), .B(n930), .Y(n1289) );
  INVXL U531 ( .A(n441), .Y(waitstaten) );
  NAND21XL U532 ( .B(n2624), .A(n420), .Y(n2634) );
  INVXL U533 ( .A(n441), .Y(n423) );
  NAND21XL U534 ( .B(n145), .A(n1543), .Y(n1593) );
  INVXL U535 ( .A(n1583), .Y(n2604) );
  NAND21XL U536 ( .B(n424), .A(n420), .Y(n2545) );
  NAND21XL U537 ( .B(n2228), .A(n373), .Y(n1887) );
  AND2XL U538 ( .A(n386), .B(n79), .Y(N11479) );
  AND3XL U539 ( .A(n386), .B(n1754), .C(n1781), .Y(N10581) );
  AND2XL U540 ( .A(n386), .B(n2641), .Y(N11483) );
  AND2XL U541 ( .A(n2829), .B(n2644), .Y(N11489) );
  AO21XL U542 ( .B(n384), .C(n147), .A(n427), .Y(N12556) );
  AO21XL U543 ( .B(n384), .C(n179), .A(n427), .Y(N12520) );
  AO21XL U544 ( .B(n384), .C(n203), .A(n428), .Y(N12511) );
  AND2XL U545 ( .A(n378), .B(n64), .Y(N11478) );
  AND2XL U546 ( .A(n386), .B(n2640), .Y(N11482) );
  NAND21XL U547 ( .B(n1657), .A(n1613), .Y(n2408) );
  INVX2 U548 ( .A(memdatai[5]), .Y(n2285) );
  INVX2 U549 ( .A(memdatai[3]), .Y(n2165) );
  INVXL U550 ( .A(n1430), .Y(n1689) );
  NAND21XL U551 ( .B(n1509), .A(n1271), .Y(n1584) );
  NAND21XL U552 ( .B(n1), .A(codefetch_s), .Y(n2676) );
  NAND32XL U553 ( .B(n1501), .C(n2084), .A(n1509), .Y(n1551) );
  INVXL U554 ( .A(n1818), .Y(n1865) );
  NAND21XL U555 ( .B(n1016), .A(n1015), .Y(n2292) );
  NAND21XL U556 ( .B(n1959), .A(n928), .Y(n496) );
  NAND21XL U557 ( .B(n1061), .A(n1060), .Y(n1817) );
  INVXL U558 ( .A(n1029), .Y(n1732) );
  INVXL U559 ( .A(n1958), .Y(n1016) );
  INVXL U560 ( .A(n1874), .Y(n1821) );
  NAND21XL U561 ( .B(n1718), .A(n2015), .Y(n2013) );
  INVXL U562 ( .A(n2251), .Y(n1198) );
  INVXL U563 ( .A(n1030), .Y(n1651) );
  NAND21XL U564 ( .B(n2013), .A(n1028), .Y(n2106) );
  INVXL U565 ( .A(n1997), .Y(n1341) );
  INVXL U566 ( .A(n1192), .Y(n1864) );
  OR2XL U567 ( .A(n2090), .B(n2061), .Y(n1244) );
  NAND21XL U568 ( .B(n1781), .A(n505), .Y(n1664) );
  INVXL U569 ( .A(n697), .Y(n740) );
  OAI21BBXL U570 ( .A(n1292), .B(n1896), .C(n930), .Y(n931) );
  INVXL U571 ( .A(n2007), .Y(n2001) );
  NAND21XL U572 ( .B(n472), .A(n2009), .Y(n1165) );
  NAND21XL U573 ( .B(n1615), .A(n1671), .Y(n1616) );
  NAND21XL U574 ( .B(n188), .A(n1042), .Y(n2445) );
  INVXL U575 ( .A(n2022), .Y(n1787) );
  OAI21BBX1 U576 ( .A(n1127), .B(n1126), .C(n1677), .Y(n1150) );
  NAND21XL U577 ( .B(n2022), .A(n1654), .Y(n2000) );
  NAND21XL U578 ( .B(n2022), .A(n2017), .Y(n1112) );
  NAND32XL U579 ( .B(n2005), .C(n2004), .A(n2003), .Y(n2006) );
  AND2XL U580 ( .A(n1207), .B(n1833), .Y(n1155) );
  INVXL U581 ( .A(n2039), .Y(n2453) );
  OAI22XL U582 ( .A(n17), .B(n2451), .C(n2623), .D(n2450), .Y(N11505) );
  OAI22XL U583 ( .A(n18), .B(n2451), .C(n2623), .D(n2350), .Y(N11504) );
  NOR32XL U584 ( .B(n2415), .C(n2384), .A(n215), .Y(n2385) );
  MUX2IX1 U585 ( .D0(n199), .D1(n2412), .S(n305), .Y(n215) );
  OAI22XL U586 ( .A(n2629), .B(n2451), .C(n2623), .D(n2405), .Y(N11502) );
  OAI22XL U587 ( .A(n2632), .B(n2451), .C(n2623), .D(n2327), .Y(N11503) );
  XOR3X1 U588 ( .A(n2100), .B(n2099), .C(n2130), .Y(n2101) );
  AND2XL U589 ( .A(n2521), .B(n76), .Y(N673) );
  AND2XL U590 ( .A(n2521), .B(n81), .Y(N676) );
  AND2XL U591 ( .A(n2521), .B(n65), .Y(N674) );
  OAI22XL U592 ( .A(n241), .B(n2451), .C(n2623), .D(n2274), .Y(N11500) );
  AND2XL U593 ( .A(n377), .B(n1760), .Y(N12470) );
  NAND21XL U594 ( .B(n2623), .A(n420), .Y(n2635) );
  NAND21XL U595 ( .B(n178), .A(n1543), .Y(n2282) );
  NAND21XL U596 ( .B(n201), .A(n1543), .Y(n2088) );
  NAND21XL U597 ( .B(n126), .A(n1759), .Y(n1756) );
  OAI22AXL U598 ( .D(n2183), .C(n2545), .A(n2185), .B(n2184), .Y(N11480) );
  INVXL U599 ( .A(memdatai[2]), .Y(n2247) );
  AO21XL U600 ( .B(n380), .C(n1307), .A(n427), .Y(N12699) );
  AND2XL U601 ( .A(n386), .B(n2352), .Y(N12703) );
  AND2XL U602 ( .A(n377), .B(n2182), .Y(N12709) );
  AND2XL U603 ( .A(n377), .B(n1344), .Y(N12701) );
  AND2XL U604 ( .A(n377), .B(n2351), .Y(N12702) );
  AND2XL U605 ( .A(n378), .B(n1343), .Y(N12710) );
  AND2XL U606 ( .A(n1759), .B(n1629), .Y(N10568) );
  AND2XL U607 ( .A(n1788), .B(n1629), .Y(N10564) );
  AND3XL U608 ( .A(n1347), .B(n1346), .C(n1958), .Y(n1348) );
  INVXL U609 ( .A(n2541), .Y(n2544) );
  XOR2XL U610 ( .A(n2206), .B(n2207), .Y(n2208) );
  INVXL U611 ( .A(n1582), .Y(n2609) );
  INVXL U612 ( .A(n1581), .Y(n2608) );
  INVXL U613 ( .A(n1761), .Y(n1762) );
  NAND31XL U614 ( .C(n2202), .A(n2201), .B(n2200), .Y(n2203) );
  AO21XL U615 ( .B(n1665), .C(n1651), .A(n1650), .Y(n1652) );
  NAND21XL U616 ( .B(n424), .A(n1633), .Y(n941) );
  NAND21XL U617 ( .B(n424), .A(n2189), .Y(n1808) );
  MUX2XL U618 ( .D0(n2864), .D1(n2653), .S(n420), .Y(mempswr_comb) );
  OA21XL U619 ( .B(n1435), .C(n2344), .A(n1434), .Y(n1437) );
  INVXL U620 ( .A(n1427), .Y(n273) );
  NOR8X1 U621 ( .A(n1940), .B(n1939), .C(n1938), .D(n2158), .E(n2372), .F(
        n1937), .G(n1936), .H(n2057), .Y(n1955) );
  OA21XL U622 ( .B(n1435), .C(n2313), .A(n1434), .Y(n1433) );
  INVXL U623 ( .A(n2090), .Y(n2091) );
  OA2222XL U624 ( .A(n2460), .B(n43), .C(n2344), .D(n2458), .E(n36), .F(n2050), 
        .G(n2455), .H(n2346), .Y(n2051) );
  OA2222XL U625 ( .A(n57), .B(n2460), .C(n2257), .D(n2458), .E(n36), .F(n2149), 
        .G(n2455), .H(n2254), .Y(n2150) );
  INVXL U626 ( .A(n2259), .Y(n2148) );
  NAND21X1 U627 ( .B(n2170), .A(n2043), .Y(n2042) );
  INVXL U628 ( .A(n1976), .Y(n278) );
  NAND4XL U629 ( .A(n2505), .B(n225), .C(n2619), .D(n2504), .Y(n281) );
  INVX2 U630 ( .A(n562), .Y(n968) );
  AO21X4 U631 ( .B(n1009), .C(n2628), .A(n737), .Y(n2390) );
  OA2222XL U632 ( .A(n999), .B(n967), .C(n997), .D(n966), .E(n995), .F(n965), 
        .G(n993), .H(n964), .Y(n1004) );
  OA2222XL U633 ( .A(n999), .B(n998), .C(n997), .D(n996), .E(n995), .F(n994), 
        .G(n993), .H(n992), .Y(n1000) );
  NAND43X1 U634 ( .B(n1196), .C(n217), .D(n218), .A(n1195), .Y(n1920) );
  OAI22X1 U635 ( .A(n263), .B(n1964), .C(n1831), .D(n1873), .Y(n217) );
  OAI22XL U636 ( .A(n1192), .B(n2411), .C(n1817), .D(n2263), .Y(n218) );
  OAI21BBXL U637 ( .A(N12808), .B(n951), .C(n219), .Y(n2353) );
  MUX2IX1 U638 ( .D0(n950), .D1(n949), .S(n211), .Y(n219) );
  OAI22XL U639 ( .A(n1964), .B(n168), .C(n263), .D(n2383), .Y(n221) );
  OAI22XL U640 ( .A(n1817), .B(n2294), .C(n1791), .D(n2411), .Y(n222) );
  NAND32XL U641 ( .B(n1509), .C(n2084), .A(n1272), .Y(n1552) );
  MUX2IX1 U642 ( .D0(n1482), .D1(n2625), .S(n1537), .Y(n223) );
  NAND32XL U643 ( .B(n1509), .C(n1269), .A(n1272), .Y(n1541) );
  NAND32XL U644 ( .B(n1816), .C(n2555), .A(n2136), .Y(n1059) );
  NAND21X1 U645 ( .B(n1906), .A(n1057), .Y(n1820) );
  NAND32XL U646 ( .B(n1501), .C(n1269), .A(n1509), .Y(n1542) );
  MUX2X1 U647 ( .D0(n880), .D1(n879), .S(n1175), .Y(n882) );
  AND3X1 U648 ( .A(n1173), .B(n1177), .C(n1178), .Y(n880) );
  INVXL U649 ( .A(n1272), .Y(n1501) );
  INVX1 U650 ( .A(n1270), .Y(n1271) );
  NAND21X1 U651 ( .B(n418), .A(n2171), .Y(n500) );
  NAND21X1 U652 ( .B(n167), .A(n2005), .Y(n2645) );
  OAI211XL U653 ( .C(n1845), .D(n1076), .A(n334), .B(n1860), .Y(n1061) );
  INVX1 U654 ( .A(n510), .Y(n514) );
  INVXL U655 ( .A(n1909), .Y(n1903) );
  NOR2XL U656 ( .A(n1845), .B(n1054), .Y(n288) );
  OAI21BBXL U657 ( .A(N12802), .B(n951), .C(n227), .Y(n1308) );
  OAI21BBXL U658 ( .A(N12801), .B(n951), .C(n228), .Y(n1313) );
  MUX2IXL U659 ( .D0(n946), .D1(n870), .S(n259), .Y(n228) );
  OAI211X1 U660 ( .C(n1983), .D(n167), .A(n1038), .B(n1019), .Y(n1020) );
  OAI21BBXL U661 ( .A(n286), .B(n343), .C(n872), .Y(n698) );
  MUX2IXL U662 ( .D0(n742), .D1(n741), .S(n343), .Y(n282) );
  OAI21BBXL U663 ( .A(N12804), .B(n951), .C(n282), .Y(n1345) );
  INVXL U664 ( .A(n545), .Y(n538) );
  NAND43X1 U665 ( .B(n1088), .C(n229), .D(n230), .A(n1087), .Y(n1940) );
  OAI22XL U666 ( .A(N13343), .B(n1922), .C(n263), .D(n2263), .Y(n229) );
  OAI22XL U667 ( .A(n1817), .B(n2116), .C(n1791), .D(n2294), .Y(n230) );
  OAI22XL U668 ( .A(n1922), .B(n1965), .C(n263), .D(n2116), .Y(n231) );
  MUX2IX1 U669 ( .D0(n1472), .D1(n2275), .S(n1537), .Y(n232) );
  MUX2IX1 U670 ( .D0(n1461), .D1(n2628), .S(n1537), .Y(n233) );
  INVXL U671 ( .A(n465), .Y(n473) );
  AO21XL U672 ( .B(n1903), .C(n2438), .A(n1902), .Y(n1415) );
  INVX1 U673 ( .A(n497), .Y(n1096) );
  INVX1 U674 ( .A(n515), .Y(n870) );
  NAND21XL U675 ( .B(n951), .A(n514), .Y(n515) );
  MUX2AXL U676 ( .D0(n1920), .D1(n2224), .S(n1980), .Y(n1921) );
  NAND32XL U677 ( .B(n1265), .C(n1778), .A(n1949), .Y(n1266) );
  OAI32XL U678 ( .A(n1621), .B(n2022), .C(n167), .D(n283), .E(n186), .Y(n518)
         );
  NAND21X1 U679 ( .B(n1721), .A(n416), .Y(n1718) );
  NAND21XL U680 ( .B(n553), .A(n552), .Y(n999) );
  INVXL U681 ( .A(n1928), .Y(n2050) );
  INVXL U682 ( .A(n1929), .Y(n2288) );
  NOR2XL U683 ( .A(n1356), .B(n235), .Y(n234) );
  AOI21X1 U684 ( .B(n506), .C(n1260), .A(n1375), .Y(n235) );
  NAND32XL U685 ( .B(n1370), .C(n1972), .A(n1941), .Y(n1017) );
  INVXL U686 ( .A(n2522), .Y(n2508) );
  INVXL U687 ( .A(n1922), .Y(n2195) );
  INVXL U688 ( .A(n1688), .Y(n1691) );
  OA21XL U689 ( .B(n926), .C(n1629), .A(n1989), .Y(n927) );
  INVXL U690 ( .A(n1793), .Y(n1796) );
  NAND21XL U691 ( .B(n35), .A(n1896), .Y(n1640) );
  INVXL U692 ( .A(n462), .Y(n1811) );
  INVXL U693 ( .A(ramdatai[0]), .Y(n2227) );
  OR2XL U694 ( .A(n1128), .B(n1030), .Y(n292) );
  XOR3XL U695 ( .A(n1427), .B(n1079), .C(n236), .Y(n1085) );
  OAI22XL U696 ( .A(n1425), .B(n1424), .C(n1084), .D(n1422), .Y(n236) );
  NAND21XL U697 ( .B(n1865), .A(n2205), .Y(n1869) );
  OA21XL U698 ( .B(n1711), .C(n1953), .A(n1109), .Y(n476) );
  AOI211XL U699 ( .C(n324), .D(n1988), .A(n1987), .B(n1986), .Y(n1995) );
  AND4XL U700 ( .A(n295), .B(n1985), .C(n1984), .D(n1983), .Y(n1996) );
  NAND32XL U701 ( .B(n2561), .C(n2562), .A(n2559), .Y(n2558) );
  NAND32XL U702 ( .B(n419), .C(n1640), .A(n1941), .Y(n1264) );
  MUX2IX1 U703 ( .D0(n1538), .D1(n2630), .S(n1537), .Y(n237) );
  MUX2IX1 U704 ( .D0(n1528), .D1(n2811), .S(n1537), .Y(n238) );
  NAND21XL U705 ( .B(n1124), .A(n1789), .Y(n1260) );
  NAND21XL U706 ( .B(n24), .A(ramdatai[1]), .Y(n1022) );
  NAND21XL U707 ( .B(n1711), .A(n2016), .Y(n1333) );
  AOI211XL U708 ( .C(n1382), .D(n152), .A(n2869), .B(n1166), .Y(n481) );
  INVXL U709 ( .A(n1840), .Y(n1847) );
  OAI221XL U710 ( .A(n1115), .B(n186), .C(n1114), .D(n2028), .E(n1113), .Y(
        n1447) );
  INVXL U711 ( .A(n1935), .Y(n2093) );
  OAI31XL U712 ( .A(n1810), .B(n187), .C(n35), .D(n1500), .Y(n2482) );
  NAND32XL U713 ( .B(n35), .C(n1718), .A(n152), .Y(n1671) );
  INVXL U714 ( .A(n1409), .Y(n2580) );
  INVXL U715 ( .A(ramdatai[1]), .Y(n2468) );
  NAND21XL U716 ( .B(n1323), .A(n1324), .Y(n1810) );
  INVXL U717 ( .A(n1370), .Y(n1292) );
  NAND21XL U718 ( .B(n152), .A(n1789), .Y(n1618) );
  NAND21XL U719 ( .B(n12), .A(ramdatai[0]), .Y(n1246) );
  NAND21XL U720 ( .B(n186), .A(n1713), .Y(n2471) );
  INVXL U721 ( .A(n1323), .Y(n1369) );
  NAND21XL U722 ( .B(n1993), .A(n1615), .Y(n1130) );
  NAND21XL U723 ( .B(n1711), .A(n2017), .Y(n1730) );
  NAND21XL U724 ( .B(n1166), .A(n1360), .Y(n1131) );
  NAND21XL U725 ( .B(n35), .A(n2016), .Y(n1656) );
  OR2XL U726 ( .A(n35), .B(n1260), .Y(n1952) );
  OR2XL U727 ( .A(n1265), .B(n1110), .Y(n1278) );
  OR2XL U728 ( .A(n2554), .B(n1031), .Y(n1032) );
  OR2XL U729 ( .A(n2094), .B(n2060), .Y(n1243) );
  AND3XL U730 ( .A(n1716), .B(n1323), .C(n1720), .Y(n484) );
  AND3XL U731 ( .A(n2017), .B(n1899), .C(n152), .Y(n466) );
  AND3XL U732 ( .A(n1974), .B(n1973), .C(n1972), .Y(n1975) );
  AND2XL U733 ( .A(n1167), .B(n1166), .Y(n1168) );
  OAI211XL U734 ( .C(n1973), .D(n1972), .A(n1047), .B(n1039), .Y(n2291) );
  NAND21XL U735 ( .B(n2265), .A(n2668), .Y(n2384) );
  INVXL U736 ( .A(n483), .Y(n1094) );
  NAND21XL U737 ( .B(n2265), .A(n2665), .Y(n2296) );
  NAND21XL U738 ( .B(n1166), .A(n1611), .Y(n2003) );
  NAND21XL U739 ( .B(n152), .A(n1136), .Y(n1137) );
  NAND21XL U740 ( .B(n483), .A(n1654), .Y(n485) );
  INVXL U741 ( .A(n2109), .Y(n1034) );
  NAND21XL U742 ( .B(n35), .A(n1322), .Y(n1945) );
  NAND32XL U743 ( .B(n185), .C(n2548), .A(n2648), .Y(n2550) );
  OAI22XL U744 ( .A(n2314), .B(n2305), .C(n2855), .D(n24), .Y(n2117) );
  NAND32XL U745 ( .B(n269), .C(n1026), .A(n2671), .Y(n2249) );
  AND3XL U746 ( .A(n2319), .B(n2436), .C(n2117), .Y(n1026) );
  NAND21XL U747 ( .B(n2668), .A(n1207), .Y(n1229) );
  AND2XL U748 ( .A(n2509), .B(n2517), .Y(n1396) );
  OAI222XL U749 ( .A(n2445), .B(n32), .C(n2444), .D(n2443), .E(n2442), .F(
        n2441), .Y(n239) );
  OAI222XL U750 ( .A(n2445), .B(n2489), .C(n2444), .D(n2346), .E(n2442), .F(
        n2345), .Y(n240) );
  OAI22XL U751 ( .A(n2314), .B(n2496), .C(n2852), .D(n24), .Y(n2333) );
  OAI221XL U752 ( .A(n2386), .B(n2668), .C(n2317), .D(n2665), .E(n2316), .Y(
        n2318) );
  OAI22XL U753 ( .A(n2314), .B(n2421), .C(n2851), .D(n24), .Y(n2418) );
  XNOR3X1 U754 ( .A(n2428), .B(n2389), .C(n2392), .Y(n2393) );
  OAI22XL U755 ( .A(n2314), .B(n2391), .C(n2854), .D(n24), .Y(n2388) );
  OAI22XL U756 ( .A(n2314), .B(n2304), .C(n2853), .D(n24), .Y(n2302) );
  NOR3XL U757 ( .A(n2273), .B(n2272), .C(n242), .Y(n241) );
  OAI222XL U758 ( .A(n2430), .B(n2271), .C(n2270), .D(n2269), .E(n74), .F(
        n2268), .Y(n242) );
  XNOR3X1 U759 ( .A(n2428), .B(n2258), .C(n243), .Y(n2271) );
  OAI222XL U760 ( .A(n27), .B(n2261), .C(n26), .D(n2260), .E(n2259), .F(n136), 
        .Y(n243) );
  MUX2IX1 U761 ( .D0(n1520), .D1(n2633), .S(n1537), .Y(n244) );
  AOI21XL U762 ( .B(n2544), .C(n2510), .A(n2517), .Y(n300) );
  AND2XL U763 ( .A(n2547), .B(n2541), .Y(n2511) );
  MUX2IX1 U764 ( .D0(n1588), .D1(n2278), .S(n1587), .Y(n245) );
  MUX2IX1 U765 ( .D0(n1575), .D1(n2277), .S(n1587), .Y(n246) );
  MUX2IX1 U766 ( .D0(n1277), .D1(n2625), .S(n1587), .Y(n247) );
  MUX2IX1 U767 ( .D0(n1571), .D1(n2275), .S(n1587), .Y(n248) );
  MUX2IX1 U768 ( .D0(n1394), .D1(n2628), .S(n1587), .Y(n249) );
  MUX2IX1 U769 ( .D0(n1567), .D1(n2630), .S(n1587), .Y(n250) );
  MUX2IX1 U770 ( .D0(n1563), .D1(n2811), .S(n1587), .Y(n251) );
  OAI22XL U771 ( .A(n358), .B(n1597), .C(n2050), .D(n139), .Y(N12626) );
  OAI22XL U772 ( .A(n358), .B(n1599), .C(n2050), .D(n154), .Y(N12590) );
  OAI22XL U773 ( .A(n358), .B(n2282), .C(n2050), .D(n128), .Y(N12617) );
  OAI22XL U774 ( .A(n358), .B(n1595), .C(n2050), .D(n123), .Y(N12581) );
  OAI22XL U775 ( .A(n358), .B(n2088), .C(n2050), .D(n118), .Y(N12608) );
  OAI22XL U776 ( .A(n358), .B(n1593), .C(n2050), .D(n114), .Y(N12572) );
  OAI22XL U777 ( .A(n358), .B(n1609), .C(n2050), .D(n111), .Y(N12635) );
  OAI22XL U778 ( .A(n358), .B(n1602), .C(n2050), .D(n55), .Y(N12599) );
  OAI22XL U779 ( .A(n1544), .B(n1597), .C(n2046), .D(n139), .Y(N12624) );
  OAI22XL U780 ( .A(n1544), .B(n1599), .C(n2046), .D(n154), .Y(N12588) );
  OAI22XL U781 ( .A(n1544), .B(n2282), .C(n2046), .D(n128), .Y(N12615) );
  OAI22XL U782 ( .A(n1544), .B(n1595), .C(n2046), .D(n123), .Y(N12579) );
  OAI22XL U783 ( .A(n1544), .B(n2088), .C(n2046), .D(n118), .Y(N12606) );
  OAI22XL U784 ( .A(n1544), .B(n1593), .C(n2046), .D(n114), .Y(N12570) );
  OAI22XL U785 ( .A(n1544), .B(n1609), .C(n2046), .D(n111), .Y(N12633) );
  OAI22XL U786 ( .A(n1544), .B(n1602), .C(n2046), .D(n56), .Y(N12597) );
  NAND21XL U787 ( .B(n2573), .A(n2572), .Y(n2574) );
  NAND32XL U788 ( .B(n2569), .C(n2568), .A(n2567), .Y(n2570) );
  NAND32XL U789 ( .B(n2569), .C(n2567), .A(n2572), .Y(n2556) );
  NAND21XL U790 ( .B(n2594), .A(n2572), .Y(n2565) );
  NOR21XL U791 ( .B(n2508), .A(n252), .Y(N12912) );
  AOI21X1 U792 ( .B(n380), .C(n2507), .A(n2506), .Y(n252) );
  NOR21XL U793 ( .B(n1752), .A(n253), .Y(n1753) );
  OAI222XL U794 ( .A(n2259), .B(n2471), .C(n2260), .D(n2467), .E(n2252), .F(
        n2473), .Y(n253) );
  NAND21XL U795 ( .B(n2517), .A(n373), .Y(n2614) );
  NAND32XL U796 ( .B(n2535), .C(n382), .A(n2517), .Y(n1221) );
  INVXL U797 ( .A(ramdatai[4]), .Y(n2854) );
  NAND21XL U798 ( .B(n1778), .A(n375), .Y(n1779) );
  AND2XL U799 ( .A(n2824), .B(n2522), .Y(N372) );
  AND2XL U800 ( .A(n2825), .B(n2522), .Y(N371) );
  AND2XL U801 ( .A(n377), .B(n78), .Y(N11486) );
  AND2XL U802 ( .A(n1759), .B(n324), .Y(N10577) );
  AND3XL U803 ( .A(memack), .B(n2697), .C(n2703), .Y(n2699) );
  INVXL U804 ( .A(n2057), .Y(n2494) );
  INVXL U805 ( .A(n1938), .Y(n2394) );
  INVXL U806 ( .A(n1936), .Y(n2300) );
  MUX2IXL U807 ( .D0(n2329), .D1(n2328), .S(n2409), .Y(n304) );
  INVXL U808 ( .A(n2297), .Y(n2298) );
  NAND21XL U809 ( .B(n2265), .A(n2124), .Y(n2414) );
  AO21XL U810 ( .B(n2292), .C(n2671), .A(n2291), .Y(n2330) );
  INVXL U811 ( .A(n2697), .Y(n2585) );
  AO22XL U812 ( .A(n2583), .B(mempsack), .C(n2703), .D(memack), .Y(n2584) );
  NAND21XL U813 ( .B(n2265), .A(n2264), .Y(n2266) );
  MUX2XL U814 ( .D0(n2263), .D1(n2262), .S(n2409), .Y(n2270) );
  AOI211XL U815 ( .C(n1732), .D(n1899), .A(n1660), .B(n1659), .Y(n1667) );
  AO21XL U816 ( .B(n1737), .C(n1736), .A(n185), .Y(n2473) );
  OR4X1 U817 ( .A(n1591), .B(n1712), .C(n1291), .D(n254), .Y(n2373) );
  AOI21XL U818 ( .B(n2002), .C(n1999), .A(n186), .Y(n254) );
  OA21XL U819 ( .B(n1733), .C(n1732), .A(n1731), .Y(n1734) );
  NOR43XL U820 ( .B(n1771), .C(n1770), .D(n2200), .A(n1819), .Y(n1773) );
  NAND32XL U821 ( .B(n1821), .C(n1764), .A(n2209), .Y(n1765) );
  OAI21BBXL U822 ( .A(n1732), .B(n1684), .C(n1661), .Y(n1662) );
  NAND21XL U823 ( .B(n418), .A(n2237), .Y(n2469) );
  NAND32XL U824 ( .B(n325), .C(n1647), .A(n1991), .Y(n1757) );
  INVXL U825 ( .A(n2557), .Y(n2575) );
  NAND32XL U826 ( .B(n2559), .C(n2562), .A(n2561), .Y(n2560) );
  INVXL U827 ( .A(n2668), .Y(n2669) );
  INVXL U828 ( .A(ramwe), .Y(n309) );
  NAND43X1 U829 ( .B(n1445), .C(n1444), .D(n1443), .A(n1442), .Y(n2372) );
  OAI22XL U830 ( .A(n1922), .B(n2294), .C(n1831), .D(n1874), .Y(n1443) );
  XNOR2X1 U831 ( .A(n1436), .B(n311), .Y(n1425) );
  NAND2XL U832 ( .A(c), .B(n1080), .Y(n311) );
  INVX1 U833 ( .A(n1875), .Y(n1942) );
  AND2XL U834 ( .A(n1911), .B(n1910), .Y(n1917) );
  MUX2XL U835 ( .D0(n1909), .D1(n1908), .S(acc[6]), .Y(n1911) );
  OAI211XL U836 ( .C(dec_accop[7]), .D(n1082), .A(n1070), .B(n1767), .Y(n2205)
         );
  OAI221XL U837 ( .A(n157), .B(n789), .C(n141), .D(n788), .E(n220), .Y(n790)
         );
  XNOR2XL U838 ( .A(n1254), .B(ramsfraddr[4]), .Y(n317) );
  AO222X1 U839 ( .A(n1540), .B(temp[4]), .C(dptr_inc[4]), .D(n1590), .E(n1539), 
        .F(n233), .Y(n1930) );
  AO222X1 U840 ( .A(n1540), .B(temp[3]), .C(dptr_inc[3]), .D(n1590), .E(n1539), 
        .F(n232), .Y(n1931) );
  AO222X1 U841 ( .A(n1540), .B(temp[2]), .C(dptr_inc[2]), .D(n1590), .E(n1539), 
        .F(n223), .Y(n1932) );
  NAND43X1 U842 ( .B(n2022), .C(n1610), .D(n2533), .A(n213), .Y(n2035) );
  MUX2XL U843 ( .D0(pc_o[1]), .D1(n1933), .S(n1934), .Y(N12842) );
  AND2XL U844 ( .A(n1792), .B(n1910), .Y(n1798) );
  AND2XL U845 ( .A(n1687), .B(n1910), .Y(n1693) );
  OAI22XL U846 ( .A(n1922), .B(n2116), .C(n263), .D(n2329), .Y(n1801) );
  INVX1 U847 ( .A(n450), .Y(n2135) );
  XOR2XL U848 ( .A(n525), .B(ramsfraddr[1]), .Y(n523) );
  NAND21X1 U849 ( .B(n1256), .A(dps[3]), .Y(n2358) );
  INVXL U850 ( .A(n1908), .Y(n1766) );
  NAND32X1 U851 ( .B(n1864), .C(n1863), .A(n1862), .Y(n1870) );
  AND4XL U852 ( .A(n1861), .B(n1860), .C(n1859), .D(n1858), .Y(n1863) );
  INVX1 U853 ( .A(n2202), .Y(n1862) );
  AOI211XL U854 ( .C(accactv), .D(n1857), .A(n1856), .B(n1855), .Y(n1858) );
  NAND31XL U855 ( .C(n1067), .A(dec_accop[2]), .B(n1062), .Y(n1791) );
  INVXL U856 ( .A(instr[7]), .Y(n325) );
  NAND21XL U857 ( .B(n2870), .A(n1135), .Y(n1331) );
  OA2222XL U858 ( .A(n991), .B(n813), .C(n989), .D(n812), .E(n987), .F(n811), 
        .G(n985), .H(n810), .Y(n819) );
  OA2222XL U859 ( .A(n999), .B(n817), .C(n997), .D(n816), .E(n995), .F(n815), 
        .G(n993), .H(n814), .Y(n818) );
  NAND21XL U860 ( .B(n2871), .A(n416), .Y(n1358) );
  INVX1 U861 ( .A(n512), .Y(n2581) );
  MUX2AXL U862 ( .D0(sp[2]), .D1(n2625), .S(n947), .Y(n516) );
  NAND43X1 U863 ( .B(n1104), .C(n1103), .D(n1102), .A(n1101), .Y(n2657) );
  INVX1 U864 ( .A(n537), .Y(n552) );
  INVXL U865 ( .A(n923), .Y(n1176) );
  AND3XL U866 ( .A(n1282), .B(n1958), .C(n447), .Y(n494) );
  AO22AXL U867 ( .A(phase[0]), .B(n1342), .C(phase[1]), .D(n1349), .Y(n2643)
         );
  INVXL U868 ( .A(ramdatao[2]), .Y(n2625) );
  OR2X1 U869 ( .A(n185), .B(n337), .Y(n2423) );
  NOR2XL U870 ( .A(dec_accop[2]), .B(dec_accop[14]), .Y(n344) );
  NAND21XL U871 ( .B(N343), .A(N344), .Y(n2264) );
  NAND21XL U872 ( .B(n1024), .A(N343), .Y(n2124) );
  OAI31XL U873 ( .A(dec_accop[7]), .B(n1069), .C(n1082), .D(accactv), .Y(n1860) );
  MUX2XL U874 ( .D0(n1940), .D1(temp[1]), .S(n1980), .Y(N12825) );
  NAND2XL U875 ( .A(dec_accop[0]), .B(accactv), .Y(n1057) );
  MUX2XL U876 ( .D0(n1939), .D1(temp[2]), .S(n1980), .Y(N12826) );
  INVXL U877 ( .A(ramdatao[1]), .Y(n2277) );
  NAND43XL U878 ( .B(ramsfraddr[4]), .C(n2558), .D(n2595), .A(ramsfraddr[3]), 
        .Y(n1632) );
  INVXL U879 ( .A(dps[0]), .Y(n1489) );
  NAND21XL U880 ( .B(n1845), .A(dec_accop[17]), .Y(n1826) );
  NAND21X1 U881 ( .B(n185), .A(interrupt), .Y(n2647) );
  OAI31XL U882 ( .A(n1027), .B(n1341), .C(n2108), .D(n214), .Y(n1031) );
  INVXL U883 ( .A(n1351), .Y(n1027) );
  INVXL U884 ( .A(dec_accop[3]), .Y(n1063) );
  NAND21XL U885 ( .B(n1493), .A(dps[2]), .Y(n2801) );
  OAI221XL U886 ( .A(n489), .B(n488), .C(n487), .D(n1029), .E(n486), .Y(n490)
         );
  NAND21XL U887 ( .B(n209), .A(n2600), .Y(n2807) );
  NAND21XL U888 ( .B(n1262), .A(n1324), .Y(n1500) );
  NAND21XL U889 ( .B(n191), .A(dec_cop[2]), .Y(n1859) );
  INVXL U890 ( .A(n1356), .Y(n1379) );
  AO21XL U891 ( .B(n1839), .C(n1838), .A(n1845), .Y(n1854) );
  OR2XL U892 ( .A(dps[0]), .B(dps[1]), .Y(n1493) );
  INVXL U893 ( .A(dec_accop[1]), .Y(n1851) );
  NAND21XL U894 ( .B(n191), .A(dec_cop[1]), .Y(n1832) );
  NAND21XL U895 ( .B(n1490), .A(dps[2]), .Y(n2798) );
  NAND21XL U896 ( .B(n1491), .A(n209), .Y(n2800) );
  NAND21XL U897 ( .B(n1492), .A(n209), .Y(n2802) );
  OAI211XL U898 ( .C(n1899), .D(n2009), .A(n1898), .B(phase[0]), .Y(n1923) );
  NAND21XL U899 ( .B(dps[2]), .A(n2603), .Y(n365) );
  NAND21XL U900 ( .B(dps[2]), .A(n2602), .Y(n367) );
  NAND21XL U901 ( .B(dps[2]), .A(n2603), .Y(n2804) );
  NAND21XL U902 ( .B(n209), .A(n2602), .Y(n368) );
  NAND21XL U903 ( .B(dps[2]), .A(n2602), .Y(n2806) );
  NAND21XL U904 ( .B(n209), .A(n2603), .Y(n366) );
  NAND21XL U905 ( .B(dps[2]), .A(n2601), .Y(n370) );
  NAND21XL U906 ( .B(n209), .A(n2600), .Y(n371) );
  NAND21XL U907 ( .B(n209), .A(n2601), .Y(n369) );
  NAND21XL U908 ( .B(n209), .A(n2601), .Y(n2808) );
  NAND21XL U909 ( .B(dps[2]), .A(n2600), .Y(n372) );
  AO21XL U910 ( .B(N345), .C(n2292), .A(n2291), .Y(n2267) );
  NAND21XL U911 ( .B(dps[0]), .A(dps[1]), .Y(n1491) );
  NAND21XL U912 ( .B(n1489), .A(dps[1]), .Y(n1490) );
  NAND21XL U913 ( .B(dps[1]), .A(dps[0]), .Y(n1492) );
  NOR21XL U914 ( .B(n448), .A(n255), .Y(n449) );
  XNOR2XL U915 ( .A(instr[7]), .B(instr[1]), .Y(n255) );
  INVXL U916 ( .A(temp[0]), .Y(n2224) );
  INVXL U917 ( .A(temp[4]), .Y(n2382) );
  INVXL U918 ( .A(temp[3]), .Y(n2159) );
  INVXL U919 ( .A(temp[1]), .Y(n2233) );
  INVXL U920 ( .A(temp[2]), .Y(n2262) );
  MUX2IX1 U921 ( .D0(state[0]), .D1(n1397), .S(n2809), .Y(n1398) );
  AO222XL U922 ( .A(n1540), .B(temp[7]), .C(dptr_inc[7]), .D(n1590), .E(n1539), 
        .F(n244), .Y(n1927) );
  AO222XL U923 ( .A(n1591), .B(temp[0]), .C(dptr_inc[8]), .D(n200), .E(n1589), 
        .F(n245), .Y(n1926) );
  AO222XL U924 ( .A(n1591), .B(temp[1]), .C(dptr_inc[9]), .D(n200), .E(n1589), 
        .F(n246), .Y(n1925) );
  AO222XL U925 ( .A(n1591), .B(temp[2]), .C(dptr_inc[10]), .D(n200), .E(n1589), 
        .F(n247), .Y(n1924) );
  AO222XL U926 ( .A(n1591), .B(temp[3]), .C(dptr_inc[11]), .D(n200), .E(n1589), 
        .F(n248), .Y(n2172) );
  AO222XL U927 ( .A(n1591), .B(temp[4]), .C(dptr_inc[12]), .D(n200), .E(n1589), 
        .F(n249), .Y(n2178) );
  AO222XL U928 ( .A(n1591), .B(temp[5]), .C(dptr_inc[13]), .D(n200), .E(n1589), 
        .F(n250), .Y(n2283) );
  AO222XL U929 ( .A(n1591), .B(temp[6]), .C(dptr_inc[14]), .D(n200), .E(n1589), 
        .F(n251), .Y(n2483) );
  AOI211XL U930 ( .C(n2518), .D(n2517), .A(n425), .B(n2547), .Y(n2519) );
  AO222XL U931 ( .A(n1591), .B(temp[7]), .C(dptr_inc[15]), .D(n200), .E(n1589), 
        .F(n2139), .Y(n2380) );
  INVXL U932 ( .A(temp[7]), .Y(n2410) );
  NAND2XL U933 ( .A(n2501), .B(n435), .Y(n354) );
  NAND21XL U934 ( .B(n209), .A(n2599), .Y(n2597) );
  AND2XL U935 ( .A(n209), .B(n2599), .Y(n353) );
  AOI22AXL U936 ( .A(pc_o[4]), .B(n1456), .D(n2387), .C(n1216), .Y(n1457) );
  AOI21X1 U937 ( .B(n1225), .C(pc_i[1]), .A(n1488), .Y(n256) );
  NAND21XL U938 ( .B(n1462), .A(memaddr[4]), .Y(n1530) );
  INVXL U939 ( .A(temp[6]), .Y(n2328) );
  MUX2AXL U940 ( .D0(n1414), .D1(n1413), .S(n2865), .Y(n257) );
  INVXL U941 ( .A(temp[5]), .Y(n2293) );
  AND3XL U942 ( .A(n2197), .B(n2196), .C(n2195), .Y(n2198) );
  OAI211XL U943 ( .C(n2033), .D(n1813), .A(n2038), .B(n1812), .Y(n1814) );
  INVX1 U944 ( .A(n381), .Y(n374) );
  INVX1 U945 ( .A(n381), .Y(n373) );
  INVX1 U946 ( .A(n381), .Y(n375) );
  INVX1 U947 ( .A(n381), .Y(n376) );
  INVX1 U948 ( .A(n381), .Y(n378) );
  INVX1 U949 ( .A(n381), .Y(n379) );
  INVX1 U950 ( .A(n2545), .Y(n380) );
  INVX1 U951 ( .A(n2545), .Y(n377) );
  INVX1 U952 ( .A(n385), .Y(n381) );
  INVX1 U953 ( .A(n385), .Y(n382) );
  AND2X1 U954 ( .A(n377), .B(n1950), .Y(N10572) );
  INVX1 U955 ( .A(n384), .Y(n383) );
  INVX1 U956 ( .A(n1288), .Y(n2845) );
  INVX1 U957 ( .A(n1956), .Y(n1971) );
  INVX1 U958 ( .A(n1289), .Y(n1092) );
  INVX1 U959 ( .A(n2004), .Y(n1984) );
  NAND21X1 U960 ( .B(n1673), .A(n260), .Y(n1950) );
  NAND21X1 U961 ( .B(n2175), .A(n375), .Y(n1979) );
  NAND21X1 U962 ( .B(n382), .A(n2175), .Y(n1978) );
  AND2X1 U963 ( .A(n2622), .B(n379), .Y(N11499) );
  INVX1 U964 ( .A(n2327), .Y(n2823) );
  INVX1 U965 ( .A(n2274), .Y(n2821) );
  INVX1 U966 ( .A(n1222), .Y(n1223) );
  INVX1 U967 ( .A(n2146), .Y(n398) );
  INVX1 U968 ( .A(n2190), .Y(n394) );
  INVX1 U969 ( .A(n2186), .Y(n409) );
  INVX1 U970 ( .A(n2146), .Y(n399) );
  INVX1 U971 ( .A(n2357), .Y(n392) );
  INVX1 U972 ( .A(n2143), .Y(n404) );
  INVX1 U973 ( .A(n2186), .Y(n412) );
  INVX1 U974 ( .A(n2137), .Y(n408) );
  INVX1 U975 ( .A(n2143), .Y(n403) );
  INVX1 U976 ( .A(n2186), .Y(n411) );
  INVX1 U977 ( .A(n2137), .Y(n407) );
  INVX1 U978 ( .A(n2186), .Y(n410) );
  INVX1 U979 ( .A(n2146), .Y(n400) );
  INVX1 U980 ( .A(n2357), .Y(n391) );
  INVX1 U981 ( .A(n2842), .Y(n388) );
  INVX1 U982 ( .A(n2190), .Y(n397) );
  INVX1 U983 ( .A(n2842), .Y(n389) );
  INVX1 U984 ( .A(n2190), .Y(n396) );
  INVX1 U985 ( .A(n2146), .Y(n401) );
  INVX1 U986 ( .A(n2140), .Y(n415) );
  INVX1 U987 ( .A(n2140), .Y(n414) );
  INVX1 U988 ( .A(n2190), .Y(n395) );
  INVX1 U989 ( .A(n2357), .Y(n393) );
  INVX1 U990 ( .A(n2143), .Y(n405) );
  INVX1 U991 ( .A(n2184), .Y(n2837) );
  INVX1 U992 ( .A(n1887), .Y(n2835) );
  INVX1 U993 ( .A(n2545), .Y(n385) );
  INVX1 U994 ( .A(n2545), .Y(n386) );
  AO21X1 U995 ( .B(n384), .C(n2604), .A(n428), .Y(N12493) );
  AO21X1 U996 ( .B(n384), .C(n2605), .A(n428), .Y(N12502) );
  AND2X1 U997 ( .A(n1782), .B(n1781), .Y(N10582) );
  INVX1 U998 ( .A(n2478), .Y(n2836) );
  INVX1 U999 ( .A(n2545), .Y(n384) );
  INVX1 U1000 ( .A(n1685), .Y(n2058) );
  NOR2X1 U1001 ( .A(n2839), .B(n2840), .Y(n1288) );
  NAND21X1 U1002 ( .B(n1654), .A(n1638), .Y(n1620) );
  INVX1 U1003 ( .A(n2641), .Y(n1187) );
  INVXL U1004 ( .A(n72), .Y(n2672) );
  NAND21X1 U1005 ( .B(n2229), .A(n1446), .Y(n1242) );
  INVX1 U1006 ( .A(n1937), .Y(n2229) );
  NAND21X1 U1007 ( .B(n1657), .A(n1132), .Y(n509) );
  NAND21XL U1008 ( .B(n2229), .A(n1198), .Y(n1222) );
  INVX1 U1009 ( .A(n1551), .Y(n2610) );
  INVX1 U1010 ( .A(n496), .Y(n2005) );
  INVX1 U1011 ( .A(n556), .Y(n539) );
  INVX1 U1012 ( .A(n1817), .Y(n2192) );
  INVX1 U1013 ( .A(n875), .Y(n1011) );
  INVX1 U1014 ( .A(n876), .Y(n1010) );
  INVX1 U1015 ( .A(n1014), .Y(n1158) );
  NAND43X1 U1016 ( .B(n1971), .C(n1970), .D(n1969), .A(n260), .Y(n2004) );
  INVX1 U1017 ( .A(n1616), .Y(n1638) );
  INVX1 U1018 ( .A(n1181), .Y(n1179) );
  AOI21X1 U1019 ( .B(n1787), .C(n1616), .A(n1713), .Y(n260) );
  INVX1 U1020 ( .A(n2292), .Y(n2265) );
  INVX1 U1021 ( .A(n2419), .Y(n2332) );
  INVX1 U1022 ( .A(n2013), .Y(n1654) );
  INVX1 U1023 ( .A(n1199), .Y(n2412) );
  INVX1 U1024 ( .A(n2108), .Y(n1347) );
  INVX1 U1025 ( .A(n1112), .Y(n1141) );
  NAND2X1 U1026 ( .A(n1150), .B(n2062), .Y(n2061) );
  INVX1 U1027 ( .A(n2000), .Y(n1673) );
  INVX1 U1028 ( .A(n1202), .Y(n1230) );
  INVX1 U1029 ( .A(n1281), .Y(n1134) );
  INVX1 U1030 ( .A(n2486), .Y(n2175) );
  INVX1 U1031 ( .A(n1402), .Y(n2622) );
  NAND21X1 U1032 ( .B(n199), .A(n2121), .Y(n2122) );
  AO21X1 U1033 ( .B(n2837), .C(n1215), .A(n2841), .Y(N672) );
  AO21X1 U1034 ( .B(n2835), .C(n1215), .A(n2841), .Y(N670) );
  NAND21X1 U1035 ( .B(n2626), .A(n375), .Y(n2274) );
  NAND21X1 U1036 ( .B(n2631), .A(n373), .Y(n2327) );
  INVX1 U1037 ( .A(n2350), .Y(n2822) );
  INVX1 U1038 ( .A(n2405), .Y(n2820) );
  INVX1 U1039 ( .A(n2450), .Y(n2816) );
  INVX1 U1040 ( .A(n1584), .Y(n2605) );
  NAND21X1 U1041 ( .B(n162), .A(n1543), .Y(n1595) );
  NAND21X1 U1042 ( .B(n1551), .A(n1543), .Y(n1597) );
  NAND21X1 U1043 ( .B(n2247), .A(n373), .Y(n2184) );
  NAND21X1 U1044 ( .B(n1297), .A(n373), .Y(n2478) );
  INVX1 U1045 ( .A(n1263), .Y(n1543) );
  NAND21X1 U1046 ( .B(n36), .A(n374), .Y(n1263) );
  NAND21X1 U1047 ( .B(n2624), .A(n374), .Y(n2451) );
  NAND21X1 U1048 ( .B(n390), .A(n434), .Y(N12690) );
  NAND21X1 U1049 ( .B(n402), .A(n433), .Y(N12691) );
  INVX1 U1050 ( .A(n2357), .Y(n390) );
  INVX1 U1051 ( .A(n2842), .Y(n387) );
  AND2X1 U1052 ( .A(n377), .B(n2098), .Y(N12469) );
  INVX1 U1053 ( .A(n1380), .Y(n2829) );
  INVX1 U1054 ( .A(n1756), .Y(n2825) );
  INVX1 U1055 ( .A(n2137), .Y(n406) );
  INVX1 U1056 ( .A(n2140), .Y(n413) );
  INVX1 U1057 ( .A(n2143), .Y(n402) );
  NAND21X1 U1058 ( .B(n1775), .A(n375), .Y(n2216) );
  AO21X1 U1059 ( .B(n386), .C(n2608), .A(n428), .Y(N12529) );
  AO21X1 U1060 ( .B(n384), .C(n2609), .A(n427), .Y(N12538) );
  AND3X1 U1061 ( .A(n376), .B(n1990), .C(n1754), .Y(N10565) );
  AND3X1 U1062 ( .A(n376), .B(n1789), .C(n1946), .Y(N10588) );
  AND2X1 U1063 ( .A(n1788), .B(n1728), .Y(N10567) );
  AND2X1 U1064 ( .A(n1782), .B(n1651), .Y(N10563) );
  AND2X1 U1065 ( .A(n1788), .B(n1787), .Y(N10589) );
  AND2X1 U1066 ( .A(n1782), .B(n1990), .Y(N10583) );
  NOR21XL U1067 ( .B(n377), .A(n261), .Y(N10571) );
  AOI21X1 U1068 ( .B(n1728), .C(n1620), .A(n1659), .Y(n261) );
  INVX1 U1069 ( .A(n1631), .Y(n1782) );
  NAND21X1 U1070 ( .B(n382), .A(n1665), .Y(n1631) );
  NAND21XL U1071 ( .B(n423), .A(n434), .Y(N370) );
  NAND21X1 U1072 ( .B(n1446), .A(n2408), .Y(n1685) );
  NAND21X1 U1073 ( .B(n2839), .A(n1239), .Y(n1455) );
  INVX1 U1074 ( .A(n1239), .Y(n2840) );
  INVX1 U1075 ( .A(n1238), .Y(n2839) );
  INVX1 U1076 ( .A(n1216), .Y(n2838) );
  INVX1 U1077 ( .A(n2442), .Y(n2104) );
  INVX1 U1078 ( .A(n1557), .Y(n1545) );
  INVX1 U1079 ( .A(n1225), .Y(n1579) );
  INVX1 U1080 ( .A(n2445), .Y(n2105) );
  INVX1 U1081 ( .A(n2367), .Y(n2463) );
  INVX1 U1082 ( .A(n434), .Y(n424) );
  INVX1 U1083 ( .A(n2477), .Y(n2365) );
  INVX1 U1084 ( .A(n434), .Y(n425) );
  INVX1 U1085 ( .A(n433), .Y(n432) );
  OR2X1 U1086 ( .A(n1732), .B(n1620), .Y(n1683) );
  INVX1 U1087 ( .A(n433), .Y(n427) );
  INVX1 U1088 ( .A(n434), .Y(n431) );
  INVX1 U1089 ( .A(n433), .Y(n430) );
  INVX1 U1090 ( .A(n435), .Y(n429) );
  INVX1 U1091 ( .A(n434), .Y(n428) );
  INVX1 U1092 ( .A(n435), .Y(n426) );
  NAND21X1 U1093 ( .B(n2623), .A(n2097), .Y(n2658) );
  INVX3 U1094 ( .A(n2667), .Y(n2670) );
  INVX1 U1095 ( .A(n1180), .Y(sfrwe_comb_s) );
  INVX1 U1096 ( .A(n2640), .Y(n1186) );
  AO21X1 U1097 ( .B(n2195), .C(n1197), .A(n1920), .Y(n1937) );
  OAI221X1 U1098 ( .A(n1184), .B(n2285), .C(n1177), .D(n1181), .E(n1183), .Y(
        n2641) );
  INVX1 U1099 ( .A(n441), .Y(n420) );
  INVX1 U1100 ( .A(n2041), .Y(n2043) );
  INVX1 U1101 ( .A(n2454), .Y(n2040) );
  INVX1 U1102 ( .A(n2189), .Y(n1775) );
  NAND43X1 U1103 ( .B(n1042), .C(n1098), .D(n2103), .A(n1100), .Y(n1097) );
  AO21XL U1104 ( .B(n946), .C(n697), .A(n870), .Y(n741) );
  NAND21XL U1105 ( .B(n2062), .A(memdatai[0]), .Y(n1241) );
  INVX1 U1106 ( .A(n2011), .Y(n1613) );
  INVX1 U1107 ( .A(n2303), .Y(n2287) );
  NAND21X1 U1108 ( .B(n1374), .A(n416), .Y(n1657) );
  NAND21X1 U1109 ( .B(n525), .A(n528), .Y(n547) );
  NAND32X1 U1110 ( .B(n1013), .C(n518), .A(n234), .Y(n507) );
  NAND21X1 U1111 ( .B(n514), .A(n511), .Y(n873) );
  INVX1 U1112 ( .A(n1542), .Y(n2606) );
  INVX1 U1113 ( .A(n1541), .Y(n2607) );
  INVX1 U1114 ( .A(n1552), .Y(n2611) );
  AO21XL U1115 ( .B(n946), .C(n259), .A(n870), .Y(n786) );
  INVX1 U1116 ( .A(n524), .Y(n975) );
  INVX1 U1117 ( .A(n1059), .Y(n1906) );
  INVX1 U1118 ( .A(n2424), .Y(n2362) );
  INVX1 U1119 ( .A(n499), .Y(n2171) );
  INVX1 U1120 ( .A(n2337), .Y(n2053) );
  INVX1 U1121 ( .A(n525), .Y(n535) );
  INVX1 U1122 ( .A(n1820), .Y(n1770) );
  INVX1 U1123 ( .A(n1067), .Y(n1767) );
  INVX1 U1124 ( .A(n1013), .Y(n828) );
  AO21X1 U1125 ( .B(n1732), .C(n1629), .A(n1125), .Y(n2109) );
  NAND21X1 U1126 ( .B(n1075), .A(n288), .Y(n1769) );
  NAND21X1 U1127 ( .B(n1960), .A(n1990), .Y(n1014) );
  NAND21X1 U1128 ( .B(n1811), .A(n416), .Y(n464) );
  NAND21XL U1129 ( .B(n1046), .A(n2430), .Y(n1089) );
  OAI211X1 U1130 ( .C(n1642), .D(n1972), .A(n1017), .B(n475), .Y(n1044) );
  AND2X1 U1131 ( .A(n1015), .B(n1038), .Y(n475) );
  INVX1 U1132 ( .A(n1718), .Y(n2017) );
  AO21XL U1133 ( .B(n946), .C(n208), .A(n922), .Y(n945) );
  XNOR2XL U1134 ( .A(n1202), .B(n1201), .Y(n1203) );
  AO21XL U1135 ( .B(n946), .C(n210), .A(n945), .Y(n949) );
  AOI21X1 U1136 ( .B(n1416), .C(n1059), .A(n1821), .Y(n263) );
  INVX1 U1137 ( .A(n553), .Y(n544) );
  INVX1 U1138 ( .A(n1672), .Y(n1615) );
  INVX1 U1139 ( .A(n1951), .Y(n1125) );
  INVX1 U1140 ( .A(n1333), .Y(n1989) );
  INVX1 U1141 ( .A(n472), .Y(n2033) );
  INVX1 U1142 ( .A(n2501), .Y(n1815) );
  INVX1 U1143 ( .A(n1045), .Y(n1091) );
  NAND32X1 U1144 ( .B(n1044), .C(n1043), .A(n1958), .Y(n1045) );
  NAND2X1 U1145 ( .A(n518), .B(n234), .Y(n869) );
  NAND21X1 U1146 ( .B(n1972), .A(n2037), .Y(n2419) );
  NAND21X1 U1147 ( .B(n2612), .A(n2185), .Y(n1181) );
  NAND21X1 U1148 ( .B(n2011), .A(n1136), .Y(n930) );
  OAI211XL U1149 ( .C(n2022), .D(n1621), .A(n1014), .B(n1161), .Y(n1043) );
  INVX1 U1150 ( .A(n1962), .Y(n1789) );
  INVX1 U1151 ( .A(n1411), .Y(n1537) );
  NAND21X1 U1152 ( .B(n1410), .A(n2580), .Y(n1411) );
  INVX1 U1153 ( .A(n1940), .Y(n2474) );
  OAI31XL U1154 ( .A(instr[4]), .B(n1960), .C(n1959), .D(n1958), .Y(n1969) );
  INVX1 U1155 ( .A(n942), .Y(n1136) );
  INVX1 U1156 ( .A(n1159), .Y(n1371) );
  NAND21XL U1157 ( .B(n1158), .A(n1314), .Y(n1159) );
  INVX1 U1158 ( .A(n471), .Y(n1642) );
  NAND21X1 U1159 ( .B(n1784), .A(n1777), .Y(n471) );
  AND3X1 U1160 ( .A(n2002), .B(n2001), .C(n2000), .Y(n2029) );
  NAND21XL U1161 ( .B(n1097), .A(n1096), .Y(n2444) );
  NAND21X1 U1162 ( .B(n1033), .A(n1032), .Y(n2422) );
  NAND21XL U1163 ( .B(n1615), .A(n1610), .Y(n1988) );
  NAND21XL U1164 ( .B(n1611), .A(n1610), .Y(n1635) );
  NAND21X1 U1165 ( .B(n1618), .A(n1612), .Y(n1109) );
  OA21X1 U1166 ( .B(n1789), .C(n2011), .A(n1165), .Y(n467) );
  INVX1 U1167 ( .A(n1959), .Y(n1728) );
  INVX1 U1168 ( .A(n1972), .Y(n1322) );
  INVX1 U1169 ( .A(n1405), .Y(n1540) );
  INVX1 U1170 ( .A(n1649), .Y(n1611) );
  INVX1 U1171 ( .A(n1406), .Y(n1539) );
  NAND21X1 U1172 ( .B(n1590), .A(n1405), .Y(n1406) );
  INVX1 U1173 ( .A(n2306), .Y(n2157) );
  INVX1 U1174 ( .A(n2390), .Y(n1982) );
  INVX1 U1175 ( .A(n1618), .Y(n1360) );
  INVX1 U1176 ( .A(n1131), .Y(n1713) );
  INVX1 U1177 ( .A(n1290), .Y(n1999) );
  NAND32X1 U1178 ( .B(n1404), .C(n1289), .A(n1287), .Y(n1290) );
  INVX1 U1179 ( .A(n1963), .Y(n1970) );
  NAND21X1 U1180 ( .B(n1962), .A(n1961), .Y(n1963) );
  NAND21XL U1181 ( .B(n1224), .A(n1098), .Y(n2442) );
  AO21X1 U1182 ( .B(n1148), .C(n1147), .A(n1146), .Y(n1152) );
  NAND21X1 U1183 ( .B(n1944), .A(n2428), .Y(n1202) );
  NAND2X1 U1184 ( .A(n1017), .B(n1897), .Y(n1199) );
  INVXL U1185 ( .A(n2440), .Y(n2591) );
  NAND21X1 U1186 ( .B(n1374), .A(n1148), .Y(n1378) );
  NAND32XL U1187 ( .B(n1990), .C(n1653), .A(n1259), .Y(n1126) );
  INVX1 U1188 ( .A(n1447), .Y(n2062) );
  INVX1 U1189 ( .A(n1671), .Y(n1623) );
  INVX1 U1190 ( .A(n2471), .Y(n2363) );
  INVX1 U1191 ( .A(n1952), .Y(n1991) );
  INVX1 U1192 ( .A(n1889), .Y(n1446) );
  INVX1 U1193 ( .A(n1656), .Y(n1754) );
  INVX1 U1194 ( .A(n2006), .Y(n2527) );
  INVX1 U1195 ( .A(n1130), .Y(n1987) );
  INVX1 U1196 ( .A(n1120), .Y(n1715) );
  NAND21X1 U1197 ( .B(instr[4]), .A(n1369), .Y(n1259) );
  NAND21X1 U1198 ( .B(n1944), .A(n1961), .Y(n1281) );
  MUX2X1 U1199 ( .D0(n2412), .D1(n2419), .S(n1108), .Y(n1040) );
  INVX1 U1200 ( .A(n1228), .Y(n1205) );
  INVX1 U1201 ( .A(n1621), .Y(n2008) );
  INVX1 U1202 ( .A(n1640), .Y(n1946) );
  NAND21X1 U1203 ( .B(n2171), .A(n1981), .Y(n2454) );
  INVX1 U1204 ( .A(n1810), .Y(n2038) );
  INVX1 U1205 ( .A(n1278), .Y(n2538) );
  INVX1 U1206 ( .A(n2315), .Y(n1023) );
  OR2XL U1207 ( .A(n2534), .B(n2676), .Y(n2486) );
  OAI31XL U1208 ( .A(n1155), .B(n89), .C(n80), .D(n2658), .Y(n1402) );
  NAND21X1 U1209 ( .B(n2175), .A(n2460), .Y(n2485) );
  INVX1 U1210 ( .A(n2168), .Y(n2452) );
  INVX1 U1211 ( .A(n2249), .Y(n1207) );
  INVX1 U1212 ( .A(sfrdatai[3]), .Y(n2305) );
  NOR2X1 U1213 ( .A(n2175), .B(n2244), .Y(n264) );
  NOR2X1 U1214 ( .A(n2175), .B(n2241), .Y(n265) );
  AND2X1 U1215 ( .A(n2646), .B(n416), .Y(retiinstr) );
  INVX1 U1216 ( .A(n2645), .Y(n2646) );
  INVX1 U1217 ( .A(n2460), .Y(n2239) );
  XOR3X1 U1218 ( .A(n2428), .B(n299), .C(n2425), .Y(n2339) );
  OAI22XL U1219 ( .A(n82), .B(n2112), .C(n2111), .D(n2110), .Y(n2258) );
  AND2XL U1220 ( .A(n82), .B(n2112), .Y(n2111) );
  GEN2XL U1221 ( .D(n2437), .E(n2343), .C(n2342), .B(n2434), .A(n2341), .Y(
        n2348) );
  MUX2X1 U1222 ( .D0(n2336), .D1(n2335), .S(n2334), .Y(n2342) );
  OAI22XL U1223 ( .A(n2431), .B(n2340), .C(n2430), .D(n2339), .Y(n2341) );
  AND2X1 U1224 ( .A(n2332), .B(n304), .Y(n2335) );
  GEN2XL U1225 ( .D(n2437), .E(n2436), .C(n2435), .B(n2434), .A(n2433), .Y(
        n2448) );
  OAI32X1 U1226 ( .A(n2420), .B(n199), .C(n2418), .D(n2417), .E(n2416), .Y(
        n2435) );
  OAI22XL U1227 ( .A(n2432), .B(n2431), .C(n2430), .D(n2429), .Y(n2433) );
  AND3X1 U1228 ( .A(n2415), .B(n2414), .C(n2413), .Y(n2416) );
  INVX1 U1229 ( .A(sfrdatai[4]), .Y(n2391) );
  OA222X1 U1230 ( .A(n2430), .B(n2311), .C(n2853), .D(n2408), .E(n2431), .F(
        n2310), .Y(n2323) );
  XOR3X1 U1231 ( .A(n2428), .B(n298), .C(n2338), .Y(n2311) );
  INVX1 U1232 ( .A(sfrdatai[5]), .Y(n2304) );
  INVX1 U1233 ( .A(sfrdatai[6]), .Y(n2496) );
  INVX1 U1234 ( .A(n2243), .Y(n2480) );
  INVX1 U1235 ( .A(n2307), .Y(n2115) );
  INVX1 U1236 ( .A(sfrdatai[7]), .Y(n2421) );
  INVX1 U1237 ( .A(n2398), .Y(n2437) );
  INVX1 U1238 ( .A(n2388), .Y(n2386) );
  INVX1 U1239 ( .A(n2302), .Y(n2317) );
  INVX1 U1240 ( .A(n2117), .Y(n2121) );
  INVX1 U1241 ( .A(n2333), .Y(n2334) );
  INVX1 U1242 ( .A(n2418), .Y(n2417) );
  OA22XL U1243 ( .A(n2431), .B(n2387), .C(n2386), .D(n2385), .Y(n2403) );
  OA22X1 U1244 ( .A(n2317), .B(n2301), .C(n2300), .D(n2406), .Y(n2325) );
  AND3X1 U1245 ( .A(n2415), .B(n2296), .C(n2295), .Y(n2301) );
  MUX2X1 U1246 ( .D0(n199), .D1(n2412), .S(n306), .Y(n2295) );
  INVX1 U1247 ( .A(n1214), .Y(n2521) );
  NAND21X1 U1248 ( .B(n2614), .A(n1215), .Y(n1214) );
  NAND6XL U1249 ( .A(n1246), .B(n1245), .C(n1244), .D(n1243), .E(n1242), .F(
        n1241), .Y(n2098) );
  NAND21X1 U1250 ( .B(n2065), .A(sfrdatai[7]), .Y(n1452) );
  AND3X1 U1251 ( .A(n2836), .B(codefetch_s), .C(n1215), .Y(N671) );
  INVX1 U1252 ( .A(n1220), .Y(n1215) );
  OAI31XL U1253 ( .A(n1220), .B(n2285), .C(n2545), .D(n1219), .Y(N675) );
  OAI31XL U1254 ( .A(n1220), .B(n1218), .C(n382), .D(n1219), .Y(N677) );
  INVX1 U1255 ( .A(n1219), .Y(n2841) );
  INVX1 U1256 ( .A(n2099), .Y(n2626) );
  INVX1 U1257 ( .A(n2730), .Y(n2631) );
  NOR21XL U1258 ( .B(n379), .A(n2101), .Y(N12905) );
  XOR3XL U1259 ( .A(n2098), .B(n2097), .C(n957), .Y(n2100) );
  XNOR2XL U1260 ( .A(n266), .B(n267), .Y(n957) );
  XNOR2XL U1261 ( .A(n2728), .B(n2727), .Y(n266) );
  XNOR2XL U1262 ( .A(n2730), .B(n2729), .Y(n267) );
  OAI22X1 U1263 ( .A(codefetch_s), .B(n2613), .C(n2547), .D(n2614), .Y(N679)
         );
  INVX1 U1264 ( .A(n1276), .Y(n1587) );
  NAND21X1 U1265 ( .B(n1410), .A(n2579), .Y(n1276) );
  INVX1 U1266 ( .A(n1267), .Y(n1591) );
  INVX1 U1267 ( .A(n1268), .Y(n1589) );
  NAND21X1 U1268 ( .B(n1590), .A(n1267), .Y(n1268) );
  NAND21X1 U1269 ( .B(n2728), .A(n375), .Y(n2450) );
  NAND21X1 U1270 ( .B(n2729), .A(n374), .Y(n2405) );
  NAND21X1 U1271 ( .B(n2727), .A(n375), .Y(n2350) );
  AND2X1 U1272 ( .A(n377), .B(n2130), .Y(N12472) );
  INVX1 U1273 ( .A(n1025), .Y(n2319) );
  NAND21X1 U1274 ( .B(n1542), .A(n1543), .Y(n1599) );
  NAND21X1 U1275 ( .B(n1552), .A(n1543), .Y(n1609) );
  NAND21X1 U1276 ( .B(n1541), .A(n1543), .Y(n1602) );
  NAND21X1 U1277 ( .B(n1248), .A(n373), .Y(n1380) );
  INVX1 U1278 ( .A(n1624), .Y(n1759) );
  NAND21X1 U1279 ( .B(n1649), .A(n375), .Y(n1624) );
  NAND21X1 U1280 ( .B(n2174), .A(n375), .Y(n2188) );
  AO21X1 U1281 ( .B(n2564), .C(n2575), .A(n432), .Y(N13014) );
  AO21X1 U1282 ( .B(n2564), .C(n2576), .A(n432), .Y(N13023) );
  AO21X1 U1283 ( .B(n2564), .C(n2577), .A(n432), .Y(N13032) );
  AO21X1 U1284 ( .B(n2564), .C(n2579), .A(n432), .Y(N13050) );
  AO21X1 U1285 ( .B(n2564), .C(n2580), .A(n432), .Y(N13059) );
  AO21X1 U1286 ( .B(n2564), .C(n313), .A(n431), .Y(N13077) );
  AO21X1 U1287 ( .B(n2566), .C(n2575), .A(n431), .Y(N13086) );
  AO21X1 U1288 ( .B(n2566), .C(n2576), .A(n431), .Y(N13095) );
  AO21X1 U1289 ( .B(n2566), .C(n2577), .A(n431), .Y(N13104) );
  AO21X1 U1290 ( .B(n2566), .C(n2579), .A(n431), .Y(N13122) );
  AO21X1 U1291 ( .B(n2566), .C(n2580), .A(n431), .Y(N13131) );
  AO21X1 U1292 ( .B(n2566), .C(n313), .A(n431), .Y(N13149) );
  AO21X1 U1293 ( .B(n2571), .C(n2575), .A(n430), .Y(N13158) );
  AO21X1 U1294 ( .B(n2571), .C(n2576), .A(n430), .Y(N13167) );
  AO21X1 U1295 ( .B(n2571), .C(n2577), .A(n430), .Y(N13176) );
  AO21X1 U1296 ( .B(n2571), .C(n2579), .A(n430), .Y(N13194) );
  AO21X1 U1297 ( .B(n2571), .C(n2580), .A(n430), .Y(N13203) );
  AO21X1 U1298 ( .B(n2571), .C(n313), .A(n430), .Y(N13221) );
  AO21X1 U1299 ( .B(n2582), .C(n2575), .A(n430), .Y(N13230) );
  AO21X1 U1300 ( .B(n2582), .C(n2576), .A(n429), .Y(N13239) );
  AO21X1 U1301 ( .B(n2577), .C(n2582), .A(n429), .Y(N13248) );
  AO21X1 U1302 ( .B(n2582), .C(n2579), .A(n429), .Y(N13266) );
  AO21X1 U1303 ( .B(n2582), .C(n2580), .A(n429), .Y(N13275) );
  AO21X1 U1304 ( .B(n2582), .C(n313), .A(n429), .Y(N13293) );
  OAI22X1 U1305 ( .A(n2851), .B(n2408), .C(n2407), .D(n2406), .Y(n2449) );
  INVX1 U1306 ( .A(n2842), .Y(n2812) );
  INVX1 U1307 ( .A(n2190), .Y(n2813) );
  INVX1 U1308 ( .A(n2137), .Y(n2831) );
  INVX1 U1309 ( .A(n2140), .Y(n2833) );
  INVX1 U1310 ( .A(n2146), .Y(n2828) );
  INVX1 U1311 ( .A(n2186), .Y(n2832) );
  INVX1 U1312 ( .A(n1755), .Y(n2824) );
  NAND32X1 U1313 ( .B(n2546), .C(n383), .A(n2544), .Y(n2613) );
  INVX1 U1314 ( .A(n1217), .Y(n2834) );
  AO21X1 U1315 ( .B(n380), .C(n1313), .A(n432), .Y(N12697) );
  AO21X1 U1316 ( .B(n384), .C(n1308), .A(n432), .Y(N12698) );
  AO21X1 U1317 ( .B(n380), .C(n2592), .A(n429), .Y(N12722) );
  NAND43X1 U1318 ( .B(n2591), .C(n2590), .D(n2589), .A(n2588), .Y(n2592) );
  AO21X1 U1319 ( .B(n380), .C(n2612), .A(n427), .Y(N11491) );
  INVX1 U1320 ( .A(n1981), .Y(n2237) );
  AND3X1 U1321 ( .A(n376), .B(n1946), .C(n1949), .Y(N10587) );
  AND3X1 U1322 ( .A(n376), .B(n1728), .C(n1682), .Y(N10570) );
  AND3X1 U1323 ( .A(n376), .B(n2009), .C(n1682), .Y(N10576) );
  AND3X1 U1324 ( .A(n376), .B(n1899), .C(n1683), .Y(N10573) );
  AND3X1 U1325 ( .A(n376), .B(n1684), .C(n1683), .Y(N10575) );
  AND2X1 U1326 ( .A(n378), .B(n1345), .Y(N12700) );
  AND2X1 U1327 ( .A(n1784), .B(n1783), .Y(N10586) );
  AND2X1 U1328 ( .A(n1758), .B(n378), .Y(N10578) );
  INVX1 U1329 ( .A(n1757), .Y(n1758) );
  AND2X1 U1330 ( .A(n1786), .B(n378), .Y(N10585) );
  INVX1 U1331 ( .A(n1785), .Y(n1786) );
  AND2X1 U1332 ( .A(n2650), .B(n378), .Y(N584) );
  AND2X1 U1333 ( .A(n1780), .B(n1783), .Y(N10584) );
  INVX1 U1334 ( .A(n1777), .Y(n1780) );
  AND2X1 U1335 ( .A(n1650), .B(n379), .Y(N10566) );
  AND2X1 U1336 ( .A(n377), .B(n2353), .Y(N12704) );
  INVX1 U1337 ( .A(n1625), .Y(n1788) );
  NAND21X1 U1338 ( .B(n1897), .A(n375), .Y(n1625) );
  NAND31X1 U1339 ( .C(n425), .A(n2613), .B(n2614), .Y(N685) );
  NAND2X1 U1340 ( .A(n435), .B(n2842), .Y(N12692) );
  AOI31XL U1341 ( .A(n1956), .B(n1951), .C(n1661), .D(n2545), .Y(N10569) );
  AOI31X1 U1342 ( .A(n1351), .B(n1349), .C(n1348), .D(n2545), .Y(N690) );
  OAI22X1 U1343 ( .A(n2852), .B(n2408), .C(n2494), .D(n2406), .Y(n2349) );
  OR2X1 U1344 ( .A(n2061), .B(n2424), .Y(n1448) );
  INVX1 U1345 ( .A(n1939), .Y(n2252) );
  INVX1 U1346 ( .A(n2158), .Y(n2166) );
  INVX1 U1347 ( .A(n2656), .Y(n2434) );
  INVX1 U1348 ( .A(n2330), .Y(n2415) );
  INVX1 U1349 ( .A(n2546), .Y(n2542) );
  MUX2X1 U1350 ( .D0(n2412), .D1(n199), .S(n2420), .Y(n2413) );
  OR3XL U1351 ( .A(n2331), .B(n2330), .C(n268), .Y(n2336) );
  MUX2IX1 U1352 ( .D0(n199), .D1(n2412), .S(n304), .Y(n268) );
  MUX2X1 U1353 ( .D0(n2412), .D1(n199), .S(n2123), .Y(n2118) );
  NAND3X1 U1354 ( .A(dpc[1]), .B(n2846), .C(n2827), .Y(n1239) );
  NAND3X1 U1355 ( .A(dpc[1]), .B(dpc[2]), .C(n2827), .Y(n1238) );
  INVX1 U1356 ( .A(n1231), .Y(n2827) );
  AOI221XL U1357 ( .A(n1329), .B(n2839), .C(n1330), .D(n2840), .E(n1231), .Y(
        n1327) );
  INVX1 U1358 ( .A(n1464), .Y(n1465) );
  INVX1 U1359 ( .A(n1514), .Y(n2817) );
  OAI221X1 U1360 ( .A(n1239), .B(n2819), .C(n1238), .D(n2818), .E(n2827), .Y(
        n1514) );
  NAND21X1 U1361 ( .B(n2838), .A(n1285), .Y(n1557) );
  OAI22X1 U1362 ( .A(n1239), .B(n1330), .C(n1238), .D(n1329), .Y(n1336) );
  NOR3XL U1363 ( .A(n2846), .B(dpc[1]), .C(n1231), .Y(n1216) );
  NOR3XL U1364 ( .A(dpc[1]), .B(dpc[2]), .C(n1231), .Y(n1225) );
  NAND21X1 U1365 ( .B(n177), .A(n1337), .Y(n1576) );
  NAND21X1 U1366 ( .B(n2588), .A(n1742), .Y(n2367) );
  OR2X1 U1367 ( .A(n2588), .B(n2590), .Y(n2488) );
  INVX1 U1368 ( .A(n2373), .Y(n2492) );
  INVX1 U1369 ( .A(n1738), .Y(n1742) );
  NAND5XL U1370 ( .A(n2471), .B(n2440), .C(n2467), .D(n2473), .E(n2477), .Y(
        n1738) );
  INVX1 U1371 ( .A(dpc[2]), .Y(n2846) );
  NAND21X1 U1372 ( .B(instr[4]), .A(n2171), .Y(n2477) );
  INVX1 U1373 ( .A(n2368), .Y(n2465) );
  INVX1 U1374 ( .A(n2366), .Y(n2466) );
  INVX1 U1375 ( .A(n1722), .Y(n1723) );
  INVX1 U1376 ( .A(n1619), .Y(n1659) );
  NAND21X1 U1377 ( .B(n1618), .A(n1617), .Y(n1619) );
  INVX1 U1378 ( .A(n2473), .Y(n2364) );
  INVX1 U1379 ( .A(n1630), .Y(n1665) );
  INVX1 U1380 ( .A(rst), .Y(n434) );
  INVX1 U1381 ( .A(n2467), .Y(n1674) );
  INVX1 U1382 ( .A(n1822), .Y(n1829) );
  INVX1 U1383 ( .A(rst), .Y(n435) );
  INVX1 U1384 ( .A(n1808), .Y(n1809) );
  INVX1 U1385 ( .A(rst), .Y(n433) );
  INVX1 U1386 ( .A(n2250), .Y(n1473) );
  INVX1 U1387 ( .A(n2558), .Y(n2576) );
  MUX2X1 U1388 ( .D0(memwr), .D1(n2649), .S(waitstaten), .Y(memwr_comb) );
  AND4XL U1389 ( .A(n2624), .B(n1244), .C(n1243), .D(n2515), .Y(n1209) );
  AND4X1 U1390 ( .A(n1242), .B(n1241), .C(n1246), .D(n1208), .Y(n1210) );
  OAI211X1 U1391 ( .C(n12), .D(n2468), .A(n1154), .B(n1153), .Y(n1760) );
  NAND21X1 U1392 ( .B(n2657), .A(n2656), .Y(n2659) );
  INVX1 U1393 ( .A(n2655), .Y(n2660) );
  OAI221X1 U1394 ( .A(n1108), .B(n1107), .C(n262), .D(n1106), .E(n1105), .Y(
        n2655) );
  AND3X1 U1395 ( .A(n2119), .B(n2296), .C(n1040), .Y(n1106) );
  INVX1 U1396 ( .A(n2657), .Y(n1105) );
  OAI221X1 U1397 ( .A(mempsack), .B(n440), .C(memack), .D(n439), .E(n438), .Y(
        n441) );
  INVX1 U1398 ( .A(n2587), .Y(n437) );
  NAND21X1 U1399 ( .B(n2151), .A(n2150), .Y(n2682) );
  NAND21X1 U1400 ( .B(n2048), .A(n2047), .Y(n2684) );
  AO2222XL U1401 ( .A(alu_out[4]), .B(n2481), .C(n65), .D(n2454), .E(n2453), 
        .F(ramdatai[4]), .G(n2452), .H(n1982), .Y(n2048) );
  OA2222XL U1402 ( .A(n39), .B(n2460), .C(n2396), .D(n2458), .E(n36), .F(n2046), .G(n2455), .H(n2397), .Y(n2047) );
  NAND21X1 U1403 ( .B(n2052), .A(n2051), .Y(n2686) );
  AO2222XL U1404 ( .A(alu_out[6]), .B(n2481), .C(n81), .D(n2454), .E(n2453), 
        .F(ramdatai[6]), .G(n2452), .H(n2053), .Y(n2052) );
  NAND32XL U1405 ( .B(n1082), .C(n1078), .A(n1081), .Y(n1430) );
  OAI22X1 U1406 ( .A(n272), .B(n1747), .C(n1429), .D(n326), .Y(n1704) );
  INVX1 U1407 ( .A(n1945), .Y(n1947) );
  MUX2X1 U1408 ( .D0(n1944), .D1(n1943), .S(n1942), .Y(n1948) );
  AND2X1 U1409 ( .A(n416), .B(n1941), .Y(n1943) );
  MAJ3X1 U1410 ( .A(n275), .B(n274), .C(n273), .Y(n272) );
  OAI21X1 U1411 ( .B(n1425), .C(n1424), .A(n1423), .Y(n275) );
  NAND21X1 U1412 ( .B(n2462), .A(n2461), .Y(n2681) );
  OA2222XL U1413 ( .A(n53), .B(n2460), .C(n2459), .D(n2458), .E(n36), .F(n2457), .G(n2456), .H(n2455), .Y(n2461) );
  NAND21X1 U1414 ( .B(n2096), .A(n2095), .Y(n2680) );
  OA2222XL U1415 ( .A(n2460), .B(n61), .C(n2094), .D(n2458), .E(n36), .F(n2093), .G(n2455), .H(n2092), .Y(n2095) );
  NAND21X1 U1416 ( .B(n2156), .A(n2155), .Y(n2683) );
  OA2222XL U1417 ( .A(n59), .B(n2460), .C(n2160), .D(n2458), .E(n47), .F(n2154), .G(n2455), .H(n2153), .Y(n2155) );
  NAND21X1 U1418 ( .B(n2290), .A(n2289), .Y(n2685) );
  AO2222XL U1419 ( .A(alu_out[5]), .B(n2481), .C(n70), .D(n2454), .E(n2453), 
        .F(ramdatai[5]), .G(n2452), .H(n2287), .Y(n2290) );
  OA2222XL U1420 ( .A(n45), .B(n2460), .C(n2313), .D(n2458), .E(n47), .F(n2288), .G(n2455), .H(n2320), .Y(n2289) );
  OA21XL U1421 ( .B(n1435), .C(n2396), .A(n1430), .Y(n1431) );
  AO21X1 U1422 ( .B(n1424), .C(n1425), .A(n1422), .Y(n1423) );
  INVX1 U1423 ( .A(n1077), .Y(n1420) );
  NAND32XL U1424 ( .B(n1076), .C(n1082), .A(n1081), .Y(n1077) );
  OAI221X1 U1425 ( .A(n1435), .B(n2094), .C(n1082), .D(n1081), .E(n1430), .Y(
        n1083) );
  AOI31X1 U1426 ( .A(n277), .B(n278), .C(n279), .D(n280), .Y(n276) );
  MUX2IX1 U1427 ( .D0(n1969), .D1(n1970), .S(n1968), .Y(n279) );
  NAND32X1 U1428 ( .B(n1816), .C(n2594), .A(n2555), .Y(n2189) );
  AO21X1 U1429 ( .B(n1009), .C(n2278), .A(n692), .Y(n2090) );
  AO44X1 U1430 ( .A(n691), .B(n690), .C(n689), .D(n688), .E(n687), .F(n686), 
        .G(n685), .H(n684), .Y(n692) );
  OA2222XL U1431 ( .A(n983), .B(n660), .C(n981), .D(n659), .E(n979), .F(n658), 
        .G(n977), .H(n657), .Y(n690) );
  OA2222XL U1432 ( .A(n983), .B(n675), .C(n981), .D(n674), .E(n979), .F(n673), 
        .G(n977), .H(n672), .Y(n686) );
  AO44X1 U1433 ( .A(n825), .B(n824), .C(n823), .D(n822), .E(n821), .F(n820), 
        .G(n819), .H(n818), .Y(n826) );
  OA2222XL U1434 ( .A(n198), .B(n794), .C(n160), .D(n793), .E(n143), .F(n792), 
        .G(n176), .H(n791), .Y(n824) );
  OA2222XL U1435 ( .A(n983), .B(n809), .C(n981), .D(n808), .E(n979), .F(n807), 
        .G(n977), .H(n806), .Y(n820) );
  AO44X1 U1436 ( .A(n736), .B(n735), .C(n734), .D(n733), .E(n732), .F(n731), 
        .G(n730), .H(n729), .Y(n737) );
  OA2222XL U1437 ( .A(n983), .B(n705), .C(n981), .D(n704), .E(n979), .F(n703), 
        .G(n977), .H(n702), .Y(n735) );
  OA2222XL U1438 ( .A(n983), .B(n720), .C(n981), .D(n719), .E(n979), .F(n718), 
        .G(n977), .H(n717), .Y(n731) );
  AO44X1 U1439 ( .A(n780), .B(n779), .C(n778), .D(n777), .E(n776), .F(n775), 
        .G(n774), .H(n773), .Y(n781) );
  OA2222XL U1440 ( .A(n983), .B(n749), .C(n981), .D(n748), .E(n979), .F(n747), 
        .G(n977), .H(n746), .Y(n779) );
  OA2222XL U1441 ( .A(n983), .B(n764), .C(n981), .D(n763), .E(n979), .F(n762), 
        .G(n977), .H(n761), .Y(n775) );
  NAND31X1 U1442 ( .C(n2507), .A(n281), .B(irq), .Y(n2541) );
  OA222X1 U1443 ( .A(n2567), .B(n876), .C(n828), .D(n738), .E(n869), .F(n2390), 
        .Y(n739) );
  INVX1 U1444 ( .A(n1344), .Y(n738) );
  OA222X1 U1445 ( .A(n234), .B(n783), .C(n828), .D(n782), .E(n869), .F(n2306), 
        .Y(n784) );
  INVX1 U1446 ( .A(n1345), .Y(n782) );
  OA222X1 U1447 ( .A(n2561), .B(n876), .C(n828), .D(n827), .E(n869), .F(n2472), 
        .Y(n829) );
  INVX1 U1448 ( .A(n1308), .Y(n827) );
  AO21X1 U1449 ( .B(memdatai[2]), .C(n1174), .A(n2183), .Y(n2638) );
  AND2XL U1450 ( .A(n882), .B(n881), .Y(n924) );
  NAND43X1 U1451 ( .B(n1173), .C(n877), .D(n878), .A(n1177), .Y(n925) );
  AOI31XL U1452 ( .A(n1957), .B(n1974), .C(n1956), .D(n1955), .Y(n1976) );
  INVX1 U1453 ( .A(n1950), .Y(n1957) );
  OAI221X1 U1454 ( .A(n875), .B(n2224), .C(n234), .D(n169), .E(n694), .Y(n695)
         );
  OA222X1 U1455 ( .A(n2559), .B(n876), .C(n828), .D(n693), .E(n869), .F(n2090), 
        .Y(n694) );
  AO21XL U1456 ( .B(n1009), .C(n2625), .A(n650), .Y(n2259) );
  AO44X1 U1457 ( .A(n649), .B(n648), .C(n647), .D(n646), .E(n645), .F(n644), 
        .G(n643), .H(n642), .Y(n650) );
  OA2222XL U1458 ( .A(n198), .B(n543), .C(n160), .D(n542), .E(n143), .F(n541), 
        .G(n176), .H(n540), .Y(n648) );
  OA2222XL U1459 ( .A(n198), .B(n573), .C(n160), .D(n572), .E(n143), .F(n571), 
        .G(n176), .H(n570), .Y(n644) );
  AO44X1 U1460 ( .A(n867), .B(n866), .C(n865), .D(n864), .E(n863), .F(n862), 
        .G(n861), .H(n860), .Y(n868) );
  OA2222XL U1461 ( .A(n196), .B(n844), .C(n159), .D(n843), .E(n175), .F(n842), 
        .G(n142), .H(n841), .Y(n864) );
  OA2222XL U1462 ( .A(n196), .B(n859), .C(n159), .D(n858), .E(n175), .F(n857), 
        .G(n142), .H(n856), .Y(n860) );
  NAND21X1 U1463 ( .B(n1157), .A(n283), .Y(n525) );
  INVX1 U1464 ( .A(n1725), .Y(n2015) );
  INVX1 U1465 ( .A(n783), .Y(n2182) );
  OAI31XL U1466 ( .A(N13353), .B(n1980), .C(n1922), .D(n1921), .Y(N12824) );
  INVX1 U1467 ( .A(n2035), .Y(n1042) );
  INVX3 U1468 ( .A(n879), .Y(n1177) );
  AOI21XL U1469 ( .B(n324), .C(n2015), .A(n1613), .Y(n283) );
  OAI221X1 U1470 ( .A(n875), .B(n2262), .C(n234), .D(n1721), .E(n652), .Y(n653) );
  OA222X1 U1471 ( .A(n2562), .B(n876), .C(n828), .D(n651), .E(n869), .F(n2259), 
        .Y(n652) );
  INVX1 U1472 ( .A(n1307), .Y(n651) );
  NAND32XL U1473 ( .B(n2084), .C(n1272), .A(n1509), .Y(n1581) );
  NAND32XL U1474 ( .B(n1509), .C(n1272), .A(n1269), .Y(n1582) );
  NAND21X1 U1475 ( .B(n1941), .A(n1384), .Y(n2022) );
  NAND21XL U1476 ( .B(n547), .A(n555), .Y(n985) );
  NAND21XL U1477 ( .B(n547), .A(n552), .Y(n981) );
  NAND21XL U1478 ( .B(n556), .A(n552), .Y(n989) );
  AO44X1 U1479 ( .A(n1007), .B(n1006), .C(n1005), .D(n1004), .E(n1003), .F(
        n1002), .G(n1001), .H(n1000), .Y(n1008) );
  NAND21XL U1480 ( .B(n536), .A(n544), .Y(n983) );
  NAND21XL U1481 ( .B(n554), .A(n552), .Y(n991) );
  NAND21XL U1482 ( .B(n554), .A(n555), .Y(n995) );
  NAND32X1 U1483 ( .B(n1060), .C(n1061), .A(n1826), .Y(n2201) );
  NAND32XL U1484 ( .B(n1068), .C(n1065), .A(n288), .Y(n1908) );
  AO222X1 U1485 ( .A(n741), .B(n286), .C(n946), .D(n698), .E(N12805), .F(n951), 
        .Y(n1344) );
  NAND21XL U1486 ( .B(n1655), .A(n928), .Y(n1287) );
  OA22X1 U1487 ( .A(n2383), .B(n1817), .C(n1791), .D(n2329), .Y(n285) );
  NAND21X1 U1488 ( .B(n1283), .A(n2034), .Y(n1960) );
  AO21XL U1489 ( .B(n1009), .C(n2811), .A(n921), .Y(n2337) );
  AO44X1 U1490 ( .A(n920), .B(n919), .C(n918), .D(n917), .E(n916), .F(n915), 
        .G(n914), .H(n913), .Y(n921) );
  OA2222XL U1491 ( .A(n196), .B(n897), .C(n159), .D(n896), .E(n175), .F(n895), 
        .G(n142), .H(n894), .Y(n917) );
  OA2222XL U1492 ( .A(n196), .B(n912), .C(n159), .D(n911), .E(n175), .F(n910), 
        .G(n142), .H(n909), .Y(n913) );
  NAND21XL U1493 ( .B(n2526), .A(n2005), .Y(n2039) );
  NAND21X1 U1494 ( .B(n1058), .A(n1770), .Y(n1064) );
  NAND21X1 U1495 ( .B(n519), .A(n2135), .Y(n2595) );
  NAND21X1 U1496 ( .B(n1953), .A(n1321), .Y(n498) );
  NAND32XL U1497 ( .B(n1820), .C(n1819), .A(n1818), .Y(n2202) );
  NAND32X1 U1498 ( .B(n259), .C(n332), .A(n516), .Y(n697) );
  NAND32X1 U1499 ( .B(n343), .C(n697), .A(n696), .Y(n872) );
  AND2XL U1500 ( .A(n946), .B(n785), .Y(n787) );
  NAND21X1 U1501 ( .B(n1331), .A(n1018), .Y(n1357) );
  OR2X1 U1502 ( .A(n1064), .B(n287), .Y(n1054) );
  AND2XL U1503 ( .A(n509), .B(n496), .Y(n504) );
  OAI22XL U1504 ( .A(n333), .B(n85), .C(n1690), .D(n1703), .Y(n1761) );
  AND2XL U1505 ( .A(n333), .B(n85), .Y(n1690) );
  INVX1 U1506 ( .A(n785), .Y(n259) );
  INVX1 U1507 ( .A(n1912), .Y(n1434) );
  NAND21X1 U1508 ( .B(n1408), .A(n1407), .Y(n1412) );
  INVX1 U1509 ( .A(n2012), .Y(n1617) );
  INVX1 U1510 ( .A(n526), .Y(n974) );
  NAND21XL U1511 ( .B(n536), .A(n539), .Y(n526) );
  INVX1 U1512 ( .A(n1382), .Y(n1321) );
  INVX1 U1513 ( .A(n513), .Y(n947) );
  NAND21X1 U1514 ( .B(n1410), .A(n2581), .Y(n513) );
  INVX1 U1515 ( .A(n1711), .Y(n1135) );
  INVX1 U1516 ( .A(n1372), .Y(n1028) );
  INVX1 U1517 ( .A(n516), .Y(n284) );
  INVX1 U1518 ( .A(n1254), .Y(n1343) );
  INVX1 U1519 ( .A(n1358), .Y(n1018) );
  NAND21X1 U1520 ( .B(n1481), .A(n1480), .Y(n1482) );
  AO2222XL U1521 ( .A(n2611), .B(n2777), .C(n2607), .D(n2779), .E(n2610), .F(
        n2778), .G(n2606), .H(n2780), .Y(n1481) );
  NAND21X1 U1522 ( .B(n1484), .A(n1483), .Y(n1485) );
  NAND21X1 U1523 ( .B(n1272), .A(n2084), .Y(n1270) );
  INVX1 U1524 ( .A(n1331), .Y(n469) );
  OAI211X1 U1525 ( .C(n167), .D(n509), .A(n2645), .B(n2039), .Y(n510) );
  AO222XL U1526 ( .A(n786), .B(n284), .C(n946), .D(n517), .E(N12803), .F(n951), 
        .Y(n1307) );
  AO21XL U1527 ( .B(n284), .C(n332), .A(n740), .Y(n517) );
  NAND21X1 U1528 ( .B(n483), .A(n1944), .Y(n505) );
  NAND21X1 U1529 ( .B(n151), .A(n1781), .Y(n1951) );
  NAND32XL U1530 ( .B(n1067), .C(n1076), .A(n1860), .Y(n1818) );
  NAND21XL U1531 ( .B(n535), .A(n534), .Y(n553) );
  NAND21X1 U1532 ( .B(n1331), .A(n2017), .Y(n1672) );
  NAND32XL U1533 ( .B(n151), .C(n2022), .A(n419), .Y(n1997) );
  NAND21XL U1534 ( .B(n1820), .A(n1058), .Y(n1874) );
  NAND21XL U1535 ( .B(n1655), .A(n1622), .Y(n1351) );
  OR2XL U1536 ( .A(n2557), .B(n1410), .Y(n2501) );
  NAND5XL U1537 ( .A(n2430), .B(n1100), .C(n2445), .D(n2439), .E(n1099), .Y(
        n2623) );
  AND4X1 U1538 ( .A(n2656), .B(n2297), .C(n2444), .D(n2442), .Y(n1099) );
  NAND21XL U1539 ( .B(n1157), .A(n416), .Y(n472) );
  NAND21X1 U1540 ( .B(n1864), .A(n1873), .Y(n1764) );
  NAND21XL U1541 ( .B(n151), .A(n416), .Y(n1029) );
  OR3XL U1542 ( .A(n1845), .B(n1063), .C(n1064), .Y(n1192) );
  NAND32XL U1543 ( .B(n2594), .C(n1409), .A(n1252), .Y(n2356) );
  INVX1 U1544 ( .A(n461), .Y(n1324) );
  NAND21X1 U1545 ( .B(n325), .A(n2034), .Y(n461) );
  XNOR3XL U1546 ( .A(n272), .B(n326), .C(n1747), .Y(n1748) );
  XOR3XL U1547 ( .A(n1703), .B(n85), .C(n333), .Y(n1705) );
  OAI211X1 U1548 ( .C(n1091), .D(n167), .A(n1090), .B(n1049), .Y(n2251) );
  AND2X1 U1549 ( .A(n1048), .B(n1047), .Y(n1049) );
  INVX1 U1550 ( .A(n1089), .Y(n1048) );
  OAI22XL U1551 ( .A(n2028), .B(n1997), .C(n1375), .D(n1655), .Y(n1356) );
  OAI22XL U1552 ( .A(n2090), .B(n2423), .C(n2227), .D(n26), .Y(n1201) );
  NAND6XL U1553 ( .A(n1999), .B(n1998), .C(n1997), .D(n1996), .E(n1995), .F(
        n1994), .Y(n2007) );
  OA21X1 U1554 ( .B(n1993), .C(n2013), .A(n1992), .Y(n1994) );
  INVX1 U1555 ( .A(n1953), .Y(n2034) );
  NAND21X1 U1556 ( .B(n2508), .A(cpu_hold), .Y(n1208) );
  OAI21BBXL U1557 ( .A(N12807), .B(n951), .C(n289), .Y(n2352) );
  MUX2IXL U1558 ( .D0(n944), .D1(n945), .S(n210), .Y(n289) );
  OAI21BBXL U1559 ( .A(N12806), .B(n951), .C(n290), .Y(n2351) );
  AOI21XL U1560 ( .B(n922), .C(n208), .A(n944), .Y(n290) );
  INVX1 U1561 ( .A(n948), .Y(n211) );
  NAND4X1 U1562 ( .A(n1031), .B(n2106), .C(n2423), .D(n292), .Y(n291) );
  INVX1 U1563 ( .A(n1778), .Y(n1896) );
  INVX1 U1564 ( .A(n1647), .Y(n2016) );
  INVX1 U1565 ( .A(n1632), .Y(n1633) );
  INVX1 U1566 ( .A(n2665), .Y(n1833) );
  INVX1 U1567 ( .A(n1664), .Y(n506) );
  INVX1 U1568 ( .A(n1655), .Y(n1629) );
  INVX1 U1569 ( .A(n1047), .Y(n508) );
  INVX1 U1570 ( .A(n2124), .Y(n2436) );
  INVX1 U1571 ( .A(n2264), .Y(n2343) );
  NAND21X1 U1572 ( .B(n1471), .A(n1470), .Y(n1472) );
  AO2222XL U1573 ( .A(n2611), .B(n2781), .C(n2607), .D(n2783), .E(n2610), .F(
        n2782), .G(n2606), .H(n2784), .Y(n1471) );
  NAND21X1 U1574 ( .B(n1460), .A(n1459), .Y(n1461) );
  AO2222XL U1575 ( .A(n2611), .B(n2785), .C(n2607), .D(n2787), .E(n2610), .F(
        n2786), .G(n2606), .H(n2788), .Y(n1460) );
  NAND21X1 U1576 ( .B(n1536), .A(n1535), .Y(n1538) );
  AO2222XL U1577 ( .A(n2611), .B(n2789), .C(n2607), .D(n2791), .E(n2610), .F(
        n2790), .G(n2606), .H(n2792), .Y(n1536) );
  NAND21X1 U1578 ( .B(n1527), .A(n1526), .Y(n1528) );
  AO2222XL U1579 ( .A(n2611), .B(n2793), .C(n2607), .D(n2795), .E(n2610), .F(
        n2794), .G(n2606), .H(n2796), .Y(n1527) );
  INVX1 U1580 ( .A(n1791), .Y(n1907) );
  INVX1 U1581 ( .A(n2573), .Y(n2136) );
  INVX1 U1582 ( .A(n874), .Y(n944) );
  NAND32XL U1583 ( .B(n873), .C(n872), .A(n871), .Y(n874) );
  NAND21XL U1584 ( .B(n187), .A(n501), .Y(n497) );
  INVX1 U1585 ( .A(n2358), .Y(n1258) );
  INVX1 U1586 ( .A(n478), .Y(n1985) );
  OAI211X1 U1587 ( .C(n477), .D(n1655), .A(n1346), .B(n476), .Y(n478) );
  INVX1 U1588 ( .A(n1988), .Y(n477) );
  INVX1 U1589 ( .A(n474), .Y(n1015) );
  OAI221XL U1590 ( .A(n1110), .B(n1370), .C(n498), .D(n505), .E(n2315), .Y(
        n474) );
  NAND21XL U1591 ( .B(n1941), .A(n416), .Y(n1962) );
  NAND32XL U1592 ( .B(n419), .C(n1655), .A(n1132), .Y(n1958) );
  NAND32X1 U1593 ( .B(n1941), .C(n1627), .A(n1626), .Y(n1777) );
  NAND21XL U1594 ( .B(n1117), .A(n2015), .Y(n1621) );
  NAND21XL U1595 ( .B(n1716), .A(n1622), .Y(n1161) );
  NAND21XL U1596 ( .B(n2012), .A(n1944), .Y(n1030) );
  NAND21XL U1597 ( .B(n1166), .A(n1944), .Y(n942) );
  XOR3XL U1598 ( .A(n1422), .B(n1425), .C(n1424), .Y(n1194) );
  OA222X1 U1599 ( .A(n1642), .B(n1778), .C(n1641), .D(n1640), .E(n1639), .F(
        n1638), .Y(n1643) );
  AND2X1 U1600 ( .A(n1637), .B(n1962), .Y(n1641) );
  INVX1 U1601 ( .A(n1653), .Y(n1639) );
  AOI21BBXL U1602 ( .B(cpu_resume), .C(irq), .A(n424), .Y(N13379) );
  NAND43X1 U1603 ( .B(n481), .C(n480), .D(n479), .A(n1985), .Y(n491) );
  OAI211X1 U1604 ( .C(n348), .D(n1331), .A(n468), .B(n467), .Y(n479) );
  GEN2XL U1605 ( .D(n1324), .E(n1731), .C(n473), .B(n1157), .A(n466), .Y(n480)
         );
  INVX1 U1606 ( .A(n1932), .Y(n2149) );
  INVX1 U1607 ( .A(n1931), .Y(n2154) );
  INVX1 U1608 ( .A(n1930), .Y(n2046) );
  INVX1 U1609 ( .A(n1720), .Y(n1612) );
  INVX1 U1610 ( .A(n1174), .Y(n2185) );
  INVX1 U1611 ( .A(n871), .Y(n208) );
  INVX1 U1612 ( .A(n943), .Y(n210) );
  INVX1 U1613 ( .A(n1861), .Y(n1060) );
  INVX1 U1614 ( .A(n2523), .Y(n2027) );
  AND2XL U1615 ( .A(n1424), .B(n1425), .Y(n1084) );
  INVX1 U1616 ( .A(n470), .Y(n1784) );
  NAND21XL U1617 ( .B(n1973), .A(n1321), .Y(n470) );
  INVX1 U1618 ( .A(n1646), .Y(n1998) );
  OAI211X1 U1619 ( .C(n1645), .D(n1644), .A(n1785), .B(n1643), .Y(n1646) );
  AND3XL U1620 ( .A(n1993), .B(n1959), .C(n1636), .Y(n1644) );
  INVX1 U1621 ( .A(n1635), .Y(n1645) );
  OA22X1 U1622 ( .A(n1636), .B(n1897), .C(n2419), .D(n1626), .Y(n295) );
  NAND32XL U1623 ( .B(n1626), .C(n1725), .A(n1018), .Y(n1897) );
  NAND32XL U1624 ( .B(n1117), .C(n35), .A(n152), .Y(n1649) );
  NAND21X1 U1625 ( .B(n2526), .A(n1404), .Y(n1405) );
  NAND32XL U1626 ( .B(n1157), .C(n2022), .A(n1156), .Y(n1314) );
  NAND32X1 U1627 ( .B(n1899), .C(n1728), .A(n1636), .Y(n1653) );
  INVX1 U1628 ( .A(n1022), .Y(n1036) );
  OAI32X1 U1629 ( .A(n2701), .B(n439), .C(n2700), .D(n440), .E(n2698), .Y(
        n2587) );
  GEN2XL U1630 ( .D(n929), .E(n1626), .C(n928), .B(n1731), .A(n927), .Y(n937)
         );
  AND2XL U1631 ( .A(n1324), .B(instr[4]), .Y(n929) );
  INVXL U1632 ( .A(n1374), .Y(n926) );
  INVX1 U1633 ( .A(n1266), .Y(n1590) );
  INVX1 U1634 ( .A(n1933), .Y(n2457) );
  INVX1 U1635 ( .A(ramdatai[2]), .Y(n2260) );
  INVX1 U1636 ( .A(n1993), .Y(n2009) );
  INVX1 U1637 ( .A(n1264), .Y(n1404) );
  INVXL U1638 ( .A(n1117), .Y(n1156) );
  INVX1 U1639 ( .A(n1637), .Y(n1949) );
  INVX1 U1640 ( .A(n1627), .Y(n2037) );
  INVX1 U1641 ( .A(n1716), .Y(n1899) );
  INVX1 U1642 ( .A(n2423), .Y(n1033) );
  INVX1 U1643 ( .A(n1133), .Y(n1961) );
  NAND21XL U1644 ( .B(n2012), .A(n1132), .Y(n1133) );
  INVX1 U1645 ( .A(n2314), .Y(n1037) );
  INVX1 U1646 ( .A(n1854), .Y(n1855) );
  INVX1 U1647 ( .A(n1057), .Y(n1416) );
  INVX1 U1648 ( .A(n1172), .Y(n2612) );
  INVX1 U1649 ( .A(n2619), .Y(n1248) );
  INVX1 U1650 ( .A(n1020), .Y(n1021) );
  AND3X1 U1651 ( .A(n2265), .B(n2412), .C(n2419), .Y(n1019) );
  INVX1 U1652 ( .A(n936), .Y(n2698) );
  NAND21X1 U1653 ( .B(n1152), .A(n1151), .Y(n2060) );
  AO21X1 U1654 ( .B(n1279), .C(n1141), .A(n2363), .Y(n2589) );
  OR2X1 U1655 ( .A(n1151), .B(n1152), .Y(n1889) );
  NAND32XL U1656 ( .B(instr[4]), .C(n1810), .A(n1711), .Y(n2548) );
  NAND32X1 U1657 ( .B(n1941), .C(n1972), .A(n1292), .Y(n1785) );
  OR2X1 U1658 ( .A(n1941), .B(n1386), .Y(n1120) );
  AND3X1 U1659 ( .A(n2548), .B(n1130), .C(n1278), .Y(n1114) );
  INVX1 U1660 ( .A(n2589), .Y(n1113) );
  AOI221XL U1661 ( .A(n1623), .B(n1384), .C(n1754), .D(n1714), .E(n1138), .Y(
        n1115) );
  NAND21XL U1662 ( .B(n1265), .A(n2034), .Y(n1630) );
  INVX1 U1663 ( .A(n1137), .Y(n1986) );
  OAI31XL U1664 ( .A(n1993), .B(n1157), .C(n1718), .D(n1109), .Y(n1138) );
  INVX1 U1665 ( .A(n1923), .Y(n1934) );
  OA22X1 U1666 ( .A(n181), .B(n2768), .C(n165), .D(n2767), .Y(n602) );
  OA22X1 U1667 ( .A(n181), .B(n2732), .C(n165), .D(n2731), .Y(n634) );
  OA22X1 U1668 ( .A(n181), .B(n2778), .C(n165), .D(n2777), .Y(n594) );
  INVX1 U1669 ( .A(n1901), .Y(n1980) );
  INVX1 U1670 ( .A(n2267), .Y(n2119) );
  NAND32X1 U1671 ( .B(n1447), .C(n1150), .A(n1149), .Y(n1146) );
  INVX1 U1672 ( .A(pc_i[9]), .Y(n2470) );
  INVX1 U1673 ( .A(n1491), .Y(n2602) );
  INVX1 U1674 ( .A(n1490), .Y(n2603) );
  INVX1 U1675 ( .A(n1492), .Y(n2601) );
  INVX1 U1676 ( .A(n1493), .Y(n2600) );
  NAND4X1 U1677 ( .A(n1361), .B(n1362), .C(n1363), .D(n1364), .Y(dpc[2]) );
  OA22X1 U1678 ( .A(n368), .B(n2718), .C(n2804), .D(n2717), .Y(n1363) );
  OA22X1 U1679 ( .A(n370), .B(n2720), .C(n372), .D(n2719), .Y(n1364) );
  OA22X1 U1680 ( .A(n181), .B(n2716), .C(n165), .D(n2715), .Y(n1361) );
  INVX1 U1681 ( .A(n1128), .Y(n1148) );
  INVX1 U1682 ( .A(n1265), .Y(n1895) );
  INVX1 U1683 ( .A(n1636), .Y(n1684) );
  MUX2IXL U1684 ( .D0(n2528), .D1(n167), .S(n1811), .Y(n296) );
  AND2X1 U1685 ( .A(n1983), .B(n1038), .Y(n1039) );
  NAND4X1 U1686 ( .A(n1352), .B(n1353), .C(n1354), .D(n1355), .Y(dpc[0]) );
  OA22X1 U1687 ( .A(n2806), .B(n2724), .C(n365), .D(n2723), .Y(n1354) );
  OA22X1 U1688 ( .A(n2808), .B(n2726), .C(n2807), .D(n2725), .Y(n1355) );
  OA22X1 U1689 ( .A(n181), .B(n2722), .C(n165), .D(n2721), .Y(n1352) );
  AOI32XL U1690 ( .A(n1991), .B(n2016), .C(n325), .D(n1990), .E(n1989), .Y(
        n1992) );
  AOI31XL U1691 ( .A(n1728), .B(n2034), .C(n169), .D(n446), .Y(n447) );
  INVX1 U1692 ( .A(n2003), .Y(n446) );
  INVX1 U1693 ( .A(n487), .Y(n932) );
  MUX2X1 U1694 ( .D0(n1964), .D1(n2233), .S(n2409), .Y(n1108) );
  MUX2X1 U1695 ( .D0(n1965), .D1(n2224), .S(n2409), .Y(n1228) );
  NAND32X1 U1696 ( .B(n1265), .C(n1972), .A(n1962), .Y(n1349) );
  NAND21XL U1697 ( .B(n1117), .A(n1727), .Y(n1722) );
  NAND21XL U1698 ( .B(n187), .A(n1125), .Y(n1677) );
  OR3XL U1699 ( .A(n2554), .B(n1447), .C(n1149), .Y(n2065) );
  OA22X1 U1700 ( .A(n368), .B(n2744), .C(n2804), .D(n2743), .Y(n628) );
  OA22X1 U1701 ( .A(n181), .B(n2742), .C(n165), .D(n2741), .Y(n626) );
  NAND21X1 U1702 ( .B(n1612), .A(n1116), .Y(n1714) );
  INVX1 U1703 ( .A(n1090), .Y(n2409) );
  INVX1 U1704 ( .A(n1116), .Y(n1727) );
  NAND4X1 U1705 ( .A(n1365), .B(n1366), .C(n1367), .D(n1368), .Y(dpc[1]) );
  OA22X1 U1706 ( .A(n367), .B(n2712), .C(n366), .D(n2711), .Y(n1367) );
  OA22X1 U1707 ( .A(n369), .B(n2714), .C(n371), .D(n2713), .Y(n1368) );
  OA22X1 U1708 ( .A(n181), .B(n2710), .C(n165), .D(n2709), .Y(n1365) );
  NAND4X1 U1709 ( .A(n630), .B(n631), .C(n632), .D(n633), .Y(dph[1]) );
  OA22X1 U1710 ( .A(n367), .B(n2738), .C(n366), .D(n2737), .Y(n632) );
  OA22X1 U1711 ( .A(n370), .B(n2740), .C(n372), .D(n2739), .Y(n633) );
  OA22X1 U1712 ( .A(n181), .B(n2736), .C(n165), .D(n2735), .Y(n630) );
  INVX1 U1713 ( .A(n2583), .Y(n440) );
  NAND4X1 U1714 ( .A(n598), .B(n599), .C(n600), .D(n601), .Y(dpl[1]) );
  OA22X1 U1715 ( .A(n2806), .B(n2774), .C(n365), .D(n2773), .Y(n600) );
  OA22X1 U1716 ( .A(n369), .B(n2776), .C(n371), .D(n2775), .Y(n601) );
  OA22X1 U1717 ( .A(n181), .B(n2772), .C(n165), .D(n2771), .Y(n598) );
  INVX1 U1718 ( .A(n1284), .Y(n2002) );
  OAI211XL U1719 ( .C(n1973), .D(n1640), .A(n1945), .B(n1951), .Y(n1284) );
  OAI221XL U1720 ( .A(n419), .B(n1167), .C(n1789), .D(n1124), .E(n1959), .Y(
        n1147) );
  INVX1 U1721 ( .A(n1375), .Y(n1127) );
  INVX1 U1722 ( .A(n2550), .Y(n2650) );
  INVX1 U1723 ( .A(n2703), .Y(n439) );
  OAI31XL U1724 ( .A(n1110), .B(n1370), .C(n1831), .D(n1038), .Y(n1025) );
  INVX1 U1725 ( .A(pc_i[6]), .Y(n2346) );
  INVX1 U1726 ( .A(pc_i[1]), .Y(n2456) );
  INVX1 U1727 ( .A(n2219), .Y(n2809) );
  NAND32XL U1728 ( .B(n186), .C(n1711), .A(n2034), .Y(n1981) );
  NAND21X1 U1729 ( .B(n1810), .A(n1279), .Y(n2168) );
  INVX1 U1730 ( .A(pc_i[4]), .Y(n2397) );
  INVX1 U1731 ( .A(pc_i[5]), .Y(n2320) );
  INVX1 U1732 ( .A(pc_i[3]), .Y(n2153) );
  INVX1 U1733 ( .A(n2512), .Y(n2534) );
  INVX1 U1734 ( .A(pc_i[2]), .Y(n2254) );
  GEN2XL U1735 ( .D(codefetch_s), .E(n2516), .C(n2509), .B(n2534), .A(n1396), 
        .Y(n1397) );
  NAND21X1 U1736 ( .B(n2361), .A(n2360), .Y(n2687) );
  AO2222XL U1737 ( .A(alu_out[7]), .B(n131), .C(n69), .D(n2454), .E(n2453), 
        .F(ramdatai[7]), .G(n2452), .H(n2362), .Y(n2361) );
  OA2222XL U1738 ( .A(n37), .B(n2460), .C(n2438), .D(n2458), .E(n36), .F(n2359), .G(n2455), .H(n2443), .Y(n2360) );
  INVX1 U1739 ( .A(n2543), .Y(n2810) );
  INVX1 U1740 ( .A(pc_i[0]), .Y(n2092) );
  OAI31XL U1741 ( .A(n2453), .B(n2171), .C(n2170), .D(n2169), .Y(n2243) );
  XNOR3X1 U1742 ( .A(n2428), .B(n297), .C(n2427), .Y(n2429) );
  OAI222XL U1743 ( .A(n2424), .B(n2423), .C(n2851), .D(n2422), .E(n27), .F(
        n2421), .Y(n297) );
  OAI222XL U1744 ( .A(n2728), .B(n2635), .C(n17), .D(n2634), .E(n423), .F(
        n2633), .Y(ramdatao_comb[7]) );
  OAI222XL U1745 ( .A(n2727), .B(n2635), .C(n18), .D(n2634), .E(n2811), .F(
        waitstaten), .Y(ramdatao_comb[6]) );
  OAI22XL U1746 ( .A(n43), .B(n2440), .C(n2439), .D(n2344), .Y(n2347) );
  OAI22XL U1747 ( .A(n37), .B(n2440), .C(n2439), .D(n2438), .Y(n2447) );
  OA222X1 U1748 ( .A(n2394), .B(n2406), .C(n2854), .D(n2408), .E(n2430), .F(
        n2393), .Y(n2401) );
  OAI222XL U1749 ( .A(n2854), .B(n2422), .C(n27), .D(n2391), .E(n2390), .F(
        n136), .Y(n2392) );
  OAI222XL U1750 ( .A(n2629), .B(n2634), .C(n2729), .D(n2635), .E(waitstaten), 
        .F(n2628), .Y(ramdatao_comb[4]) );
  OAI222XL U1751 ( .A(n2632), .B(n2634), .C(n2631), .D(n2635), .E(waitstaten), 
        .F(n2630), .Y(ramdatao_comb[5]) );
  INVX1 U1752 ( .A(n2404), .Y(n2629) );
  NAND5XL U1753 ( .A(n2403), .B(n2402), .C(n2401), .D(n2400), .E(n2399), .Y(
        n2404) );
  OA222X1 U1754 ( .A(n2439), .B(n2396), .C(n2442), .D(n2395), .E(n39), .F(
        n2440), .Y(n2400) );
  NAND32X1 U1755 ( .B(n199), .C(n2388), .A(n305), .Y(n2402) );
  INVX1 U1756 ( .A(n2326), .Y(n2632) );
  NAND5XL U1757 ( .A(n2325), .B(n2324), .C(n2323), .D(n2322), .E(n2321), .Y(
        n2326) );
  OA222X1 U1758 ( .A(n2439), .B(n2313), .C(n2442), .D(n2312), .E(n45), .F(
        n2440), .Y(n2322) );
  NAND32X1 U1759 ( .B(n199), .C(n2302), .A(n306), .Y(n2324) );
  AO21X1 U1760 ( .B(n2319), .C(n2318), .A(n2671), .Y(n2398) );
  AOI221XL U1761 ( .A(n2436), .B(n2418), .C(n2343), .D(n2333), .E(n2315), .Y(
        n2316) );
  OA222X1 U1762 ( .A(n2430), .B(n2126), .C(n2125), .D(n2656), .E(n2166), .F(
        n2251), .Y(n2127) );
  OA222X1 U1763 ( .A(n2124), .B(n2249), .C(n2123), .D(n2122), .E(n2121), .F(
        n2120), .Y(n2125) );
  XOR3X1 U1764 ( .A(n2428), .B(n2115), .C(n2114), .Y(n2126) );
  AND3X1 U1765 ( .A(n2119), .B(n2414), .C(n2118), .Y(n2120) );
  OA222X1 U1766 ( .A(n2668), .B(n2398), .C(n2444), .D(n2397), .E(n41), .F(
        n2445), .Y(n2399) );
  OA222X1 U1767 ( .A(n2665), .B(n2398), .C(n2444), .D(n2320), .E(n49), .F(
        n2445), .Y(n2321) );
  OAI222XL U1768 ( .A(n2626), .B(n2635), .C(n241), .D(n2634), .E(waitstaten), 
        .F(n2625), .Y(ramdatao_comb[2]) );
  INVX1 U1769 ( .A(n1924), .Y(n2242) );
  INVX1 U1770 ( .A(n1927), .Y(n2359) );
  INVX1 U1771 ( .A(n1926), .Y(n2223) );
  AOI211X1 U1772 ( .C(pc_i[0]), .D(n1234), .A(n1233), .B(n1232), .Y(n1235) );
  INVX1 U1773 ( .A(n2444), .Y(n1234) );
  AOI211XL U1774 ( .C(n1230), .D(n87), .A(n2430), .B(n82), .Y(n1232) );
  INVX1 U1775 ( .A(n1229), .Y(n1233) );
  OAI222XL U1776 ( .A(n2855), .B(n26), .C(n27), .D(n2305), .E(n2306), .F(n136), 
        .Y(n2114) );
  OAI222XL U1777 ( .A(n2252), .B(n2251), .C(n2431), .D(n2250), .E(n2264), .F(
        n2249), .Y(n2273) );
  NAND21X1 U1778 ( .B(n1519), .A(n1518), .Y(n1520) );
  AO2222XL U1779 ( .A(n2611), .B(n2797), .C(n2607), .D(n2803), .E(n2610), .F(
        n2799), .G(n2606), .H(n2805), .Y(n1519) );
  NAND21X1 U1780 ( .B(n1586), .A(n1585), .Y(n1588) );
  AO2222XL U1781 ( .A(n2611), .B(n2731), .C(n2606), .D(n2733), .E(n2610), .F(
        n2732), .G(n2607), .H(n2734), .Y(n1586) );
  AND2X1 U1782 ( .A(n385), .B(n2654), .Y(N582) );
  OAI221XL U1783 ( .A(n2439), .B(n2257), .C(n57), .D(n2440), .E(n2256), .Y(
        n2272) );
  NAND32X1 U1784 ( .B(n2219), .C(n383), .A(n2810), .Y(n2503) );
  GEN2XL U1785 ( .D(n2514), .E(n2512), .C(n2511), .B(n2535), .A(codefetch_s), 
        .Y(n2513) );
  OAI211X1 U1786 ( .C(n12), .D(n2855), .A(n1710), .B(n1709), .Y(n2130) );
  OA22X1 U1787 ( .A(n2166), .B(n1889), .C(n2065), .D(n2305), .Y(n1710) );
  INVX1 U1788 ( .A(n1925), .Y(n2236) );
  NAND21X1 U1789 ( .B(n1574), .A(n1573), .Y(n1575) );
  AO2222XL U1790 ( .A(n2611), .B(n2735), .C(n2607), .D(n2737), .E(n2610), .F(
        n2736), .G(n2606), .H(n2738), .Y(n1574) );
  OAI31XL U1791 ( .A(n2810), .B(cs_run), .C(n2219), .D(n72), .Y(n2498) );
  INVX1 U1792 ( .A(n2510), .Y(n2547) );
  OAI22X1 U1793 ( .A(n2503), .B(n2516), .C(n527), .D(n1400), .Y(n1880) );
  OAI22X1 U1794 ( .A(n2503), .B(n2515), .C(n527), .D(n2502), .Y(n1879) );
  AND2X1 U1795 ( .A(n1403), .B(n435), .Y(N515) );
  OAI22XL U1796 ( .A(n72), .B(n1402), .C(n1401), .D(n2498), .Y(n1403) );
  AND2X1 U1797 ( .A(n2516), .B(n1400), .Y(n1401) );
  AND2X1 U1798 ( .A(n2500), .B(n435), .Y(N512) );
  OAI22XL U1799 ( .A(n2499), .B(n72), .C(n2667), .D(n2498), .Y(n2500) );
  INVX1 U1800 ( .A(n2621), .Y(n2499) );
  NAND2X1 U1801 ( .A(n433), .B(n529), .Y(n527) );
  OAI21X1 U1802 ( .B(n2810), .C(n530), .A(n2809), .Y(n529) );
  NOR43XL U1803 ( .B(n1454), .C(n1453), .D(n1452), .A(n1451), .Y(n2728) );
  NAND21XL U1804 ( .B(n2059), .A(ramdatai[7]), .Y(n1454) );
  NAND21X1 U1805 ( .B(n2407), .A(n1685), .Y(n1453) );
  NAND31X1 U1806 ( .C(n1450), .A(n1449), .B(n1448), .Y(n1451) );
  NAND21X1 U1807 ( .B(n2544), .A(n2510), .Y(n1220) );
  OAI211X1 U1808 ( .C(n12), .D(n2260), .A(n1891), .B(n1890), .Y(n2099) );
  OA222X1 U1809 ( .A(n2062), .B(n2247), .C(n2259), .D(n2061), .E(n2060), .F(
        n2257), .Y(n1890) );
  OA22XL U1810 ( .A(n2252), .B(n1889), .C(n2065), .D(n2261), .Y(n1891) );
  OAI211X1 U1811 ( .C(n2065), .D(n2304), .A(n1807), .B(n1806), .Y(n2730) );
  OA22X1 U1812 ( .A(n2059), .B(n2853), .C(n2058), .D(n2300), .Y(n1807) );
  OR2X1 U1813 ( .A(n382), .B(n300), .Y(n1219) );
  INVX1 U1814 ( .A(n1700), .Y(n2729) );
  OAI211X1 U1815 ( .C(n2065), .D(n2391), .A(n1699), .B(n1698), .Y(n1700) );
  OA22X1 U1816 ( .A(n2059), .B(n2854), .C(n2058), .D(n2394), .Y(n1699) );
  NAND21X1 U1817 ( .B(n1274), .A(n1273), .Y(n1277) );
  AO2222XL U1818 ( .A(n147), .B(n2741), .C(n179), .D(n2743), .E(n163), .F(
        n2742), .G(n203), .H(n2744), .Y(n1274) );
  AND2X1 U1819 ( .A(n378), .B(n2543), .Y(N588) );
  INVX1 U1820 ( .A(n2066), .Y(n2727) );
  OAI211X1 U1821 ( .C(n2065), .D(n2496), .A(n2064), .B(n2063), .Y(n2066) );
  OA22X1 U1822 ( .A(n2059), .B(n2852), .C(n2058), .D(n2494), .Y(n2064) );
  NAND21X1 U1823 ( .B(n2173), .A(n2174), .Y(n2244) );
  INVXL U1824 ( .A(ramdatai[3]), .Y(n2855) );
  NAND21X1 U1825 ( .B(n1570), .A(n1569), .Y(n1571) );
  AO2222XL U1826 ( .A(n147), .B(n2747), .C(n179), .D(n2749), .E(n163), .F(
        n2748), .G(n203), .H(n2750), .Y(n1570) );
  AND2X1 U1827 ( .A(n385), .B(n2627), .Y(N11501) );
  NAND21XL U1828 ( .B(n167), .A(n1404), .Y(n1267) );
  OR2X1 U1829 ( .A(n2174), .B(n2173), .Y(n2241) );
  OA22X1 U1830 ( .A(n2806), .B(n2750), .C(n365), .D(n2749), .Y(n624) );
  OA22X1 U1831 ( .A(n182), .B(n2748), .C(n166), .D(n2747), .Y(n622) );
  OA22X1 U1832 ( .A(n182), .B(n2782), .C(n166), .D(n2781), .Y(n590) );
  NAND21X1 U1833 ( .B(n1393), .A(n1392), .Y(n1394) );
  AO2222XL U1834 ( .A(n147), .B(n2751), .C(n179), .D(n2753), .E(n163), .F(
        n2752), .G(n203), .H(n2754), .Y(n1393) );
  NAND21X1 U1835 ( .B(n1566), .A(n1565), .Y(n1567) );
  AO2222XL U1836 ( .A(n147), .B(n2755), .C(n179), .D(n2757), .E(n163), .F(
        n2756), .G(n203), .H(n2758), .Y(n1566) );
  INVX1 U1837 ( .A(n2593), .Y(n2579) );
  AND2X1 U1838 ( .A(n385), .B(n2621), .Y(N11498) );
  INVX1 U1839 ( .A(n1900), .Y(n2826) );
  NAND21X1 U1840 ( .B(n2410), .A(n1980), .Y(n1900) );
  NAND21X1 U1841 ( .B(n1562), .A(n1561), .Y(n1563) );
  AO2222XL U1842 ( .A(n147), .B(n2759), .C(n179), .D(n2761), .E(n163), .F(
        n2760), .G(n203), .H(n2762), .Y(n1562) );
  OA2222XL U1843 ( .A(n2766), .B(n178), .C(n2765), .D(n201), .E(n2763), .F(
        n1552), .G(n2764), .H(n1551), .Y(n1553) );
  INVX1 U1844 ( .A(pc_i[7]), .Y(n2443) );
  NAND21X1 U1845 ( .B(n2379), .A(n2378), .Y(N12721) );
  NAND21X1 U1846 ( .B(n424), .A(n2377), .Y(n2378) );
  NOR21XL U1847 ( .B(sfrdatai[7]), .A(n2495), .Y(n2379) );
  NAND31X1 U1848 ( .C(n2376), .A(n2375), .B(n2374), .Y(n2377) );
  OAI22X1 U1849 ( .A(n424), .B(n2286), .C(n2304), .D(n2495), .Y(N12719) );
  OA2222XL U1850 ( .A(n2300), .B(n2493), .C(n2492), .D(n2285), .E(n2853), .F(
        n2490), .G(n49), .H(n2488), .Y(n2286) );
  OAI22X1 U1851 ( .A(n425), .B(n2497), .C(n2496), .D(n2495), .Y(N12720) );
  OA2222XL U1852 ( .A(n2494), .B(n2493), .C(n2492), .D(n2491), .E(n2490), .F(
        n2852), .G(n2489), .H(n2488), .Y(n2497) );
  OAI22X1 U1853 ( .A(n424), .B(n2167), .C(n2305), .D(n2495), .Y(N12717) );
  OA2222XL U1854 ( .A(n2166), .B(n2493), .C(n2492), .D(n2165), .E(n2855), .F(
        n2490), .G(n2849), .H(n2488), .Y(n2167) );
  OAI22X1 U1855 ( .A(n425), .B(n2181), .C(n2391), .D(n2495), .Y(N12718) );
  OA2222XL U1856 ( .A(n2394), .B(n2493), .C(n2492), .D(n2180), .E(n2854), .F(
        n2490), .G(n41), .H(n2488), .Y(n2181) );
  OA2222XL U1857 ( .A(n2229), .B(n2493), .C(n2492), .D(n2228), .E(n2490), .F(
        n2227), .G(n51), .H(n2488), .Y(n2231) );
  NAND21X1 U1858 ( .B(n2630), .A(n373), .Y(n2842) );
  NAND21X1 U1859 ( .B(n2625), .A(n374), .Y(n2190) );
  NAND21X1 U1860 ( .B(n2275), .A(n374), .Y(n2357) );
  NAND21X1 U1861 ( .B(n2633), .A(n374), .Y(n2137) );
  NAND21X1 U1862 ( .B(n2811), .A(n373), .Y(n2140) );
  NAND21X1 U1863 ( .B(n1716), .A(n1759), .Y(n1755) );
  NAND21X1 U1864 ( .B(n2277), .A(n373), .Y(n2146) );
  NAND21X1 U1865 ( .B(n2278), .A(n374), .Y(n2186) );
  NAND21X1 U1866 ( .B(n2628), .A(n374), .Y(n2143) );
  INVX1 U1867 ( .A(n2565), .Y(n2566) );
  NAND2X1 U1868 ( .A(n1500), .B(n374), .Y(n2083) );
  AO21X1 U1869 ( .B(n2564), .C(n2578), .A(n432), .Y(N13041) );
  AO21X1 U1870 ( .B(n2564), .C(n2581), .A(n431), .Y(N13068) );
  AO21X1 U1871 ( .B(n2566), .C(n2578), .A(n431), .Y(N13113) );
  AO21X1 U1872 ( .B(n2566), .C(n2581), .A(n431), .Y(N13140) );
  AO21X1 U1873 ( .B(n2571), .C(n2578), .A(n430), .Y(N13185) );
  AO21X1 U1874 ( .B(n2571), .C(n2581), .A(n430), .Y(N13212) );
  AO21X1 U1875 ( .B(n2578), .C(n2582), .A(n429), .Y(N13257) );
  AO21X1 U1876 ( .B(n2582), .C(n2581), .A(n430), .Y(N13284) );
  AO21X1 U1877 ( .B(n2598), .C(n2600), .A(n429), .Y(N12637) );
  AO21X1 U1878 ( .B(n2598), .C(n2601), .A(n428), .Y(N12644) );
  AO21X1 U1879 ( .B(n2598), .C(n2602), .A(n429), .Y(N12651) );
  AO21X1 U1880 ( .B(n2598), .C(n2603), .A(n428), .Y(N12658) );
  AO21X1 U1881 ( .B(n353), .C(n2600), .A(n429), .Y(N12665) );
  AO21X1 U1882 ( .B(n353), .C(n2601), .A(n428), .Y(N12672) );
  AO21X1 U1883 ( .B(n353), .C(n2602), .A(n428), .Y(N12679) );
  AO21X1 U1884 ( .B(n353), .C(n2603), .A(n428), .Y(N12686) );
  NAND21X1 U1885 ( .B(n2218), .A(n2217), .Y(N12711) );
  NAND21X1 U1886 ( .B(n2216), .A(n2215), .Y(n2217) );
  NOR2XL U1887 ( .A(n2190), .B(n2189), .Y(n2218) );
  NAND21X1 U1888 ( .B(n2214), .A(n2213), .Y(n2215) );
  INVX1 U1889 ( .A(n2596), .Y(n2599) );
  NAND43X1 U1890 ( .B(n2595), .C(n2594), .D(n2593), .A(n376), .Y(n2596) );
  INVX1 U1891 ( .A(n2568), .Y(n2572) );
  NOR3XL U1892 ( .A(n1829), .B(n1817), .C(n2552), .Y(n301) );
  INVX1 U1893 ( .A(n2372), .Y(n2407) );
  NOR3XL U1894 ( .A(n1829), .B(n1922), .C(n2551), .Y(n302) );
  INVX1 U1895 ( .A(n2570), .Y(n2571) );
  INVX1 U1896 ( .A(n2556), .Y(n2564) );
  INVX1 U1897 ( .A(n2574), .Y(n2582) );
  OAI221X1 U1898 ( .A(n2232), .B(n2188), .C(n2187), .D(n2146), .E(n435), .Y(
        N12486) );
  OAI221X1 U1899 ( .A(n2222), .B(n2188), .C(n2187), .D(n2186), .E(n435), .Y(
        N12485) );
  OAI221X1 U1900 ( .A(n2240), .B(n2188), .C(n2187), .D(n2190), .E(n433), .Y(
        N12487) );
  OAI22XL U1901 ( .A(n1510), .B(n2085), .C(n1509), .D(n2083), .Y(N12693) );
  INVX1 U1902 ( .A(dpc[3]), .Y(n1510) );
  OAI22XL U1903 ( .A(n1942), .B(n2216), .C(n2189), .D(n2137), .Y(N12705) );
  OAI22X1 U1904 ( .A(n1681), .B(n1680), .C(n1679), .D(n382), .Y(N10562) );
  AND3X1 U1905 ( .A(n1678), .B(n1677), .C(n1676), .Y(n1679) );
  AND2X1 U1906 ( .A(n1755), .B(n1756), .Y(n1680) );
  AOI211X1 U1907 ( .C(n1787), .D(n1675), .A(n2363), .B(n1674), .Y(n1676) );
  OAI22X1 U1908 ( .A(n1753), .B(n381), .C(n2477), .D(n2184), .Y(N12725) );
  OA2222XL U1909 ( .A(n2257), .B(n2368), .C(n2253), .D(n2469), .E(n57), .F(
        n2367), .G(n2262), .H(n2366), .Y(n1752) );
  OAI22X1 U1910 ( .A(n256), .B(n1597), .C(n2457), .D(n139), .Y(N12621) );
  OAI22X1 U1911 ( .A(n2147), .B(n1597), .C(n2149), .D(n139), .Y(N12622) );
  OAI22X1 U1912 ( .A(n2152), .B(n1597), .C(n2154), .D(n139), .Y(N12623) );
  OAI22X1 U1913 ( .A(n2147), .B(n1599), .C(n2149), .D(n154), .Y(N12586) );
  OAI22X1 U1914 ( .A(n2152), .B(n1599), .C(n2154), .D(n154), .Y(N12587) );
  OAI22X1 U1915 ( .A(n2147), .B(n2282), .C(n2149), .D(n128), .Y(N12613) );
  OAI22X1 U1916 ( .A(n2152), .B(n2282), .C(n2154), .D(n128), .Y(N12614) );
  OAI22X1 U1917 ( .A(n2147), .B(n1595), .C(n2149), .D(n123), .Y(N12577) );
  OAI22X1 U1918 ( .A(n2152), .B(n1595), .C(n2154), .D(n123), .Y(N12578) );
  OAI22X1 U1919 ( .A(n2147), .B(n2088), .C(n2149), .D(n118), .Y(N12604) );
  OAI22X1 U1920 ( .A(n2152), .B(n2088), .C(n2154), .D(n118), .Y(N12605) );
  OAI22X1 U1921 ( .A(n2147), .B(n1593), .C(n2149), .D(n114), .Y(N12568) );
  OAI22X1 U1922 ( .A(n2152), .B(n1593), .C(n2154), .D(n114), .Y(N12569) );
  OAI22X1 U1923 ( .A(n2147), .B(n1609), .C(n2149), .D(n111), .Y(N12631) );
  OAI22X1 U1924 ( .A(n2152), .B(n1609), .C(n2154), .D(n111), .Y(N12632) );
  OAI22X1 U1925 ( .A(n2147), .B(n1602), .C(n2149), .D(n55), .Y(N12595) );
  OAI22X1 U1926 ( .A(n2152), .B(n1602), .C(n2154), .D(n56), .Y(N12596) );
  OAI22X1 U1927 ( .A(n1600), .B(n1597), .C(n2223), .D(n139), .Y(N12548) );
  OAI22X1 U1928 ( .A(n2049), .B(n1597), .C(n2288), .D(n140), .Y(N12625) );
  OAI22X1 U1929 ( .A(n20), .B(n1597), .C(n2236), .D(n140), .Y(N12549) );
  OAI22X1 U1930 ( .A(n1607), .B(n194), .C(n2242), .D(n140), .Y(N12550) );
  OAI22X1 U1931 ( .A(n2049), .B(n1599), .C(n2288), .D(n154), .Y(N12589) );
  OAI22X1 U1932 ( .A(n20), .B(n1599), .C(n2236), .D(n154), .Y(N12513) );
  OAI22X1 U1933 ( .A(n1607), .B(n1599), .C(n2242), .D(n155), .Y(N12514) );
  OAI22X1 U1934 ( .A(n1600), .B(n1595), .C(n2223), .D(n123), .Y(N12503) );
  OAI22X1 U1935 ( .A(n1600), .B(n2282), .C(n2223), .D(n128), .Y(N12539) );
  OAI22X1 U1936 ( .A(n2049), .B(n2282), .C(n2288), .D(n128), .Y(N12616) );
  OAI22X1 U1937 ( .A(n20), .B(n2282), .C(n2236), .D(n129), .Y(N12540) );
  OAI22X1 U1938 ( .A(n1607), .B(n153), .C(n2242), .D(n129), .Y(N12541) );
  OAI22X1 U1939 ( .A(n2049), .B(n1595), .C(n2288), .D(n123), .Y(N12580) );
  OAI22X1 U1940 ( .A(n20), .B(n1595), .C(n2236), .D(n124), .Y(N12504) );
  OAI22X1 U1941 ( .A(n1607), .B(n138), .C(n2242), .D(n124), .Y(N12505) );
  OAI22X1 U1942 ( .A(n1600), .B(n1593), .C(n2223), .D(n114), .Y(N12494) );
  OAI22X1 U1943 ( .A(n1600), .B(n2088), .C(n2223), .D(n118), .Y(N12530) );
  OAI22X1 U1944 ( .A(n2049), .B(n2088), .C(n2288), .D(n118), .Y(N12607) );
  OAI22X1 U1945 ( .A(n20), .B(n2088), .C(n2236), .D(n119), .Y(N12531) );
  OAI22X1 U1946 ( .A(n1607), .B(n127), .C(n2242), .D(n119), .Y(N12532) );
  OAI22X1 U1947 ( .A(n2049), .B(n1593), .C(n2288), .D(n114), .Y(N12571) );
  OAI22X1 U1948 ( .A(n20), .B(n1593), .C(n2236), .D(n115), .Y(N12495) );
  OAI22X1 U1949 ( .A(n1607), .B(n122), .C(n2242), .D(n115), .Y(N12496) );
  OAI22X1 U1950 ( .A(n1600), .B(n1602), .C(n2223), .D(n55), .Y(N12521) );
  OAI22X1 U1951 ( .A(n1600), .B(n1609), .C(n2223), .D(n111), .Y(N12557) );
  OAI22X1 U1952 ( .A(n2049), .B(n1609), .C(n2288), .D(n111), .Y(N12634) );
  OAI22X1 U1953 ( .A(n20), .B(n1609), .C(n2236), .D(n112), .Y(N12558) );
  OAI22X1 U1954 ( .A(n1607), .B(n117), .C(n2242), .D(n112), .Y(N12559) );
  OAI22X1 U1955 ( .A(n2049), .B(n1602), .C(n2288), .D(n56), .Y(N12598) );
  OAI22X1 U1956 ( .A(n20), .B(n1602), .C(n2236), .D(n55), .Y(N12522) );
  OAI22X1 U1957 ( .A(n1607), .B(n113), .C(n2242), .D(n56), .Y(N12523) );
  OAI22X1 U1958 ( .A(n1600), .B(n171), .C(n2223), .D(n155), .Y(N12512) );
  OAI22X1 U1959 ( .A(n2089), .B(n194), .C(n2359), .D(n140), .Y(N12627) );
  OAI22X1 U1960 ( .A(n2089), .B(n171), .C(n2359), .D(n155), .Y(N12591) );
  OAI22X1 U1961 ( .A(n2089), .B(n153), .C(n2359), .D(n129), .Y(N12618) );
  OAI22X1 U1962 ( .A(n2089), .B(n138), .C(n2359), .D(n124), .Y(N12582) );
  OAI22X1 U1963 ( .A(n2089), .B(n127), .C(n2359), .D(n119), .Y(N12609) );
  OAI22X1 U1964 ( .A(n2089), .B(n122), .C(n2359), .D(n115), .Y(N12573) );
  OAI22X1 U1965 ( .A(n2089), .B(n117), .C(n2359), .D(n112), .Y(N12636) );
  OAI22X1 U1966 ( .A(n2089), .B(n113), .C(n2359), .D(n55), .Y(N12600) );
  OAI22X1 U1967 ( .A(n22), .B(n194), .C(n2177), .D(n140), .Y(N12551) );
  OAI22X1 U1968 ( .A(n22), .B(n171), .C(n2177), .D(n155), .Y(N12515) );
  OAI22X1 U1969 ( .A(n22), .B(n153), .C(n2177), .D(n129), .Y(N12542) );
  OAI22X1 U1970 ( .A(n22), .B(n138), .C(n2177), .D(n124), .Y(N12506) );
  OAI22X1 U1971 ( .A(n22), .B(n127), .C(n2177), .D(n119), .Y(N12533) );
  OAI22X1 U1972 ( .A(n22), .B(n122), .C(n2177), .D(n115), .Y(N12497) );
  OAI22X1 U1973 ( .A(n22), .B(n117), .C(n2177), .D(n112), .Y(N12560) );
  OAI22X1 U1974 ( .A(n22), .B(n113), .C(n2177), .D(n56), .Y(N12524) );
  OAI22X1 U1975 ( .A(n1606), .B(n194), .C(n1605), .D(n140), .Y(N12552) );
  OAI22X1 U1976 ( .A(n23), .B(n194), .C(n2281), .D(n140), .Y(N12553) );
  OAI22X1 U1977 ( .A(n1606), .B(n171), .C(n1605), .D(n155), .Y(N12516) );
  OAI22X1 U1978 ( .A(n23), .B(n171), .C(n2281), .D(n155), .Y(N12517) );
  OAI22X1 U1979 ( .A(n1606), .B(n153), .C(n1605), .D(n129), .Y(N12543) );
  OAI22X1 U1980 ( .A(n23), .B(n153), .C(n2281), .D(n129), .Y(N12544) );
  OAI22X1 U1981 ( .A(n1606), .B(n138), .C(n1605), .D(n124), .Y(N12507) );
  OAI22X1 U1982 ( .A(n23), .B(n138), .C(n2281), .D(n124), .Y(N12508) );
  OAI22X1 U1983 ( .A(n1606), .B(n127), .C(n1605), .D(n119), .Y(N12534) );
  OAI22X1 U1984 ( .A(n23), .B(n127), .C(n2281), .D(n119), .Y(N12535) );
  OAI22X1 U1985 ( .A(n1606), .B(n122), .C(n1605), .D(n115), .Y(N12498) );
  OAI22X1 U1986 ( .A(n23), .B(n122), .C(n2281), .D(n115), .Y(N12499) );
  OAI22X1 U1987 ( .A(n1606), .B(n117), .C(n1605), .D(n112), .Y(N12561) );
  OAI22X1 U1988 ( .A(n23), .B(n117), .C(n2281), .D(n112), .Y(N12562) );
  OAI22X1 U1989 ( .A(n1606), .B(n113), .C(n1605), .D(n55), .Y(N12525) );
  OAI22X1 U1990 ( .A(n23), .B(n113), .C(n2281), .D(n56), .Y(N12526) );
  OAI22X1 U1991 ( .A(n1604), .B(n194), .C(n1603), .D(n140), .Y(N12554) );
  OAI22X1 U1992 ( .A(n21), .B(n194), .C(n1601), .D(n140), .Y(N12555) );
  OAI22X1 U1993 ( .A(n1604), .B(n171), .C(n1603), .D(n155), .Y(N12518) );
  OAI22X1 U1994 ( .A(n21), .B(n171), .C(n1601), .D(n155), .Y(N12519) );
  OAI22X1 U1995 ( .A(n1604), .B(n153), .C(n1603), .D(n129), .Y(N12545) );
  OAI22X1 U1996 ( .A(n21), .B(n153), .C(n1601), .D(n129), .Y(N12546) );
  OAI22X1 U1997 ( .A(n1604), .B(n138), .C(n1603), .D(n124), .Y(N12509) );
  OAI22X1 U1998 ( .A(n21), .B(n138), .C(n1601), .D(n124), .Y(N12510) );
  OAI22X1 U1999 ( .A(n1604), .B(n127), .C(n1603), .D(n119), .Y(N12536) );
  OAI22X1 U2000 ( .A(n21), .B(n127), .C(n1601), .D(n119), .Y(N12537) );
  OAI22X1 U2001 ( .A(n1604), .B(n122), .C(n1603), .D(n115), .Y(N12500) );
  OAI22X1 U2002 ( .A(n21), .B(n122), .C(n1601), .D(n115), .Y(N12501) );
  OAI22X1 U2003 ( .A(n1604), .B(n117), .C(n1603), .D(n112), .Y(N12563) );
  OAI22X1 U2004 ( .A(n21), .B(n117), .C(n1601), .D(n112), .Y(N12564) );
  OAI22X1 U2005 ( .A(n1604), .B(n113), .C(n1603), .D(n55), .Y(N12527) );
  OAI22X1 U2006 ( .A(n21), .B(n113), .C(n1601), .D(n56), .Y(N12528) );
  OAI22XL U2007 ( .A(n425), .B(n2358), .C(n2357), .D(n2356), .Y(n1884) );
  OAI22XL U2008 ( .A(n1502), .B(n2085), .C(n1501), .D(n2083), .Y(N12694) );
  INVX1 U2009 ( .A(dpc[4]), .Y(n1502) );
  OAI22XL U2010 ( .A(n2086), .B(n2085), .C(n2084), .D(n2083), .Y(N12695) );
  INVX1 U2011 ( .A(dpc[5]), .Y(n2086) );
  OAI22X1 U2012 ( .A(n2093), .B(n140), .C(n257), .D(n1597), .Y(N12620) );
  OAI22X1 U2013 ( .A(n2093), .B(n155), .C(n257), .D(n1599), .Y(N12584) );
  OAI22X1 U2014 ( .A(n2093), .B(n129), .C(n257), .D(n2282), .Y(N12611) );
  OAI22X1 U2015 ( .A(n2457), .B(n129), .C(n256), .D(n2282), .Y(N12612) );
  OAI22X1 U2016 ( .A(n2093), .B(n124), .C(n257), .D(n1595), .Y(N12575) );
  OAI22X1 U2017 ( .A(n2457), .B(n124), .C(n256), .D(n1595), .Y(N12576) );
  OAI22X1 U2018 ( .A(n2093), .B(n119), .C(n257), .D(n2088), .Y(N12602) );
  OAI22X1 U2019 ( .A(n2457), .B(n119), .C(n256), .D(n2088), .Y(N12603) );
  OAI22X1 U2020 ( .A(n2093), .B(n115), .C(n257), .D(n1593), .Y(N12566) );
  OAI22X1 U2021 ( .A(n2457), .B(n115), .C(n256), .D(n1593), .Y(N12567) );
  OAI22X1 U2022 ( .A(n2093), .B(n112), .C(n257), .D(n1609), .Y(N12629) );
  OAI22X1 U2023 ( .A(n2457), .B(n112), .C(n256), .D(n1609), .Y(N12630) );
  OAI22X1 U2024 ( .A(n2093), .B(n55), .C(n257), .D(n1602), .Y(N12593) );
  OAI22X1 U2025 ( .A(n2457), .B(n155), .C(n256), .D(n1599), .Y(N12585) );
  OAI22X1 U2026 ( .A(n2457), .B(n56), .C(n256), .D(n1602), .Y(N12594) );
  OAI22XL U2027 ( .A(n424), .B(n1306), .C(n2495), .D(n1305), .Y(N12715) );
  OA2222XL U2028 ( .A(n2474), .B(n2493), .C(n2492), .D(n1297), .E(n2490), .F(
        n2468), .G(n2850), .H(n2488), .Y(n1306) );
  OAI22XL U2029 ( .A(n425), .B(n2248), .C(n2261), .D(n2495), .Y(N12716) );
  OA2222XL U2030 ( .A(n2252), .B(n2493), .C(n2492), .D(n2247), .E(n2490), .F(
        n2260), .G(n2255), .H(n2488), .Y(n2248) );
  OAI22XL U2031 ( .A(n1381), .B(n2545), .C(n2644), .D(n1380), .Y(N11487) );
  INVX1 U2032 ( .A(n2617), .Y(n1381) );
  AND4XL U2033 ( .A(n2829), .B(n2505), .C(n225), .D(n2504), .Y(n2506) );
  INVX1 U2034 ( .A(n1221), .Y(n2355) );
  NAND21X1 U2035 ( .B(n1500), .A(n375), .Y(n2085) );
  INVXL U2036 ( .A(ramdatai[5]), .Y(n2853) );
  NAND32X1 U2037 ( .B(n425), .C(n356), .A(n2551), .Y(N13366) );
  NAND32X1 U2038 ( .B(n425), .C(n355), .A(n2552), .Y(N13324) );
  INVXL U2039 ( .A(ramdatai[6]), .Y(n2852) );
  INVX1 U2040 ( .A(n2187), .Y(n2174) );
  AND3X1 U2041 ( .A(n376), .B(n2652), .C(n2648), .Y(N585) );
  AND2X1 U2042 ( .A(n355), .B(multemp2[3]), .Y(N13326) );
  AND2X1 U2043 ( .A(n355), .B(multemp2[7]), .Y(N13330) );
  AND2X1 U2044 ( .A(n355), .B(multemp2[8]), .Y(N13331) );
  AND2X1 U2045 ( .A(n355), .B(multemp2[4]), .Y(N13327) );
  AND2X1 U2046 ( .A(n355), .B(multemp2[2]), .Y(N13325) );
  AND2X1 U2047 ( .A(n355), .B(multemp2[5]), .Y(N13328) );
  AND2X1 U2048 ( .A(n355), .B(multemp2[6]), .Y(N13329) );
  AND2X1 U2049 ( .A(n355), .B(multemp2[9]), .Y(N13332) );
  AND2X1 U2050 ( .A(n2834), .B(n2643), .Y(N11488) );
  AND2X1 U2051 ( .A(n2830), .B(n2652), .Y(N583) );
  OAI21BBX1 U2052 ( .A(n1684), .B(n1635), .C(n1648), .Y(n1614) );
  AND2X1 U2053 ( .A(n356), .B(n1827), .Y(N13369) );
  AND2X1 U2054 ( .A(n356), .B(n2068), .Y(N13370) );
  AND2X1 U2055 ( .A(n356), .B(n2075), .Y(N13371) );
  AND2X1 U2056 ( .A(n356), .B(n2074), .Y(N13372) );
  AND2X1 U2057 ( .A(n356), .B(n2067), .Y(N13368) );
  AND2X1 U2058 ( .A(n356), .B(n357), .Y(N13367) );
  AND2X1 U2059 ( .A(n356), .B(n2076), .Y(N13373) );
  INVX1 U2060 ( .A(n1779), .Y(n1783) );
  INVX1 U2061 ( .A(n2354), .Y(n2830) );
  NAND21X1 U2062 ( .B(n2648), .A(n374), .Y(n2354) );
  OAI211X1 U2063 ( .C(n936), .D(n2703), .A(n2702), .B(n435), .Y(n934) );
  OAI22X1 U2064 ( .A(n2701), .B(n2700), .C(n2699), .D(n2698), .Y(n2702) );
  OA22X1 U2065 ( .A(n367), .B(n2792), .C(n366), .D(n2791), .Y(n584) );
  OA22X1 U2066 ( .A(n2806), .B(n2788), .C(n365), .D(n2787), .Y(n588) );
  OA22X1 U2067 ( .A(n182), .B(n2790), .C(n166), .D(n2789), .Y(n582) );
  OA22X1 U2068 ( .A(n182), .B(n2756), .C(n166), .D(n2755), .Y(n614) );
  OA22X1 U2069 ( .A(n182), .B(n2786), .C(n166), .D(n2785), .Y(n586) );
  OA22X1 U2070 ( .A(n182), .B(n2752), .C(n166), .D(n2751), .Y(n618) );
  INVXL U2071 ( .A(ramdatai[7]), .Y(n2851) );
  AOI211X1 U2072 ( .C(n2706), .D(n2707), .A(n934), .B(n2705), .Y(N12975) );
  INVX1 U2073 ( .A(n933), .Y(n2705) );
  AND2X1 U2074 ( .A(n2704), .B(n2706), .Y(N12974) );
  INVX1 U2075 ( .A(n934), .Y(n2704) );
  OA22X1 U2076 ( .A(n2802), .B(n2766), .C(n134), .D(n2765), .Y(n607) );
  OA22X1 U2077 ( .A(n182), .B(n2760), .C(n166), .D(n2759), .Y(n610) );
  OA22X1 U2078 ( .A(n182), .B(n2794), .C(n166), .D(n2793), .Y(n578) );
  NAND32X1 U2079 ( .B(n425), .C(n2587), .A(n2586), .Y(N12977) );
  NAND21X1 U2080 ( .B(n2585), .A(n2584), .Y(n2586) );
  INVX1 U2081 ( .A(n2483), .Y(n1603) );
  INVX1 U2082 ( .A(n2380), .Y(n1601) );
  NAND21X1 U2083 ( .B(n2514), .A(n2535), .Y(n2546) );
  OA21X1 U2084 ( .B(n2490), .C(n2851), .A(n303), .Y(n2374) );
  NAND2XL U2085 ( .A(n2373), .B(n69), .Y(n303) );
  OA22X1 U2086 ( .A(n2806), .B(n2762), .C(n365), .D(n2761), .Y(n612) );
  OA22X1 U2087 ( .A(n182), .B(n2764), .C(n166), .D(n2763), .Y(n606) );
  OA22X1 U2088 ( .A(n182), .B(n2799), .C(n166), .D(n2797), .Y(n566) );
  NAND21X1 U2089 ( .B(n2299), .A(n2298), .Y(n2406) );
  INVX1 U2090 ( .A(n2408), .Y(n2299) );
  INVX1 U2091 ( .A(n2172), .Y(n2177) );
  INVX1 U2092 ( .A(n2178), .Y(n1605) );
  INVX1 U2093 ( .A(n2283), .Y(n2281) );
  INVX1 U2094 ( .A(n2509), .Y(n2514) );
  MUX2X1 U2095 ( .D0(n2411), .D1(n2410), .S(n2409), .Y(n2420) );
  MUX2X1 U2096 ( .D0(n2116), .D1(n2159), .S(n2409), .Y(n2123) );
  OA222X1 U2097 ( .A(n2445), .B(n2255), .C(n2444), .D(n2254), .E(n2442), .F(
        n2253), .Y(n2256) );
  MUX2XL U2098 ( .D0(N13347), .D1(n315), .S(N13353), .Y(n1827) );
  MUX2XL U2099 ( .D0(N13348), .D1(n316), .S(N13353), .Y(n2068) );
  MUX2XL U2100 ( .D0(N13349), .D1(n314), .S(N13353), .Y(n2075) );
  MUX2XL U2101 ( .D0(N13350), .D1(n323), .S(N13353), .Y(n2074) );
  MUX2XL U2102 ( .D0(N13346), .D1(n312), .S(N13353), .Y(n2067) );
  MUX2XL U2103 ( .D0(N13351), .D1(n322), .S(N13353), .Y(n2076) );
  NAND21X1 U2104 ( .B(n12), .A(n2408), .Y(n2059) );
  NAND21X1 U2105 ( .B(n2493), .A(n2372), .Y(n2375) );
  INVX1 U2106 ( .A(pc_i[10]), .Y(n2253) );
  INVX1 U2107 ( .A(pc_i[12]), .Y(n2395) );
  INVX1 U2108 ( .A(pc_i[14]), .Y(n2345) );
  INVX1 U2109 ( .A(pc_i[13]), .Y(n2312) );
  INVX1 U2110 ( .A(pc_i[15]), .Y(n2441) );
  AOI211X1 U2111 ( .C(n2332), .D(n2270), .A(n2331), .B(n2267), .Y(n2268) );
  INVX1 U2112 ( .A(n2266), .Y(n2331) );
  NAND21X1 U2113 ( .B(n1500), .A(dpc[0]), .Y(n1231) );
  AO21X1 U2114 ( .B(n1455), .C(n1463), .A(n1486), .Y(n1464) );
  AO21X1 U2115 ( .B(n1426), .C(n37), .A(n1337), .Y(n2432) );
  INVX1 U2116 ( .A(pc_i[8]), .Y(n1877) );
  INVX1 U2117 ( .A(n1529), .Y(n1466) );
  NOR2X1 U2118 ( .A(n37), .B(n1426), .Y(n1337) );
  MUX2IX1 U2119 ( .D0(n2383), .D1(n2382), .S(n2409), .Y(n305) );
  MUX2IX1 U2120 ( .D0(n2294), .D1(n2293), .S(n2409), .Y(n306) );
  INVX1 U2121 ( .A(n2648), .Y(n2651) );
  AOI22X1 U2122 ( .A(n2840), .B(n1302), .C(n2839), .D(n1301), .Y(n1293) );
  OAI221X1 U2123 ( .A(n1288), .B(n2850), .C(n1320), .D(n2838), .E(n1327), .Y(
        n1326) );
  OAI221X1 U2124 ( .A(n1288), .B(n37), .C(n1337), .D(n2838), .E(n2817), .Y(
        n1350) );
  OAI221X1 U2125 ( .A(n1288), .B(n2849), .C(n1303), .D(n2838), .E(n2844), .Y(
        n1309) );
  OAI21BBX1 U2126 ( .A(n1216), .B(n1310), .C(n2844), .Y(n1316) );
  OAI21BBX1 U2127 ( .A(n1216), .B(n1294), .C(n2843), .Y(n1298) );
  OAI21BBX1 U2128 ( .A(n1216), .B(n1328), .C(n1327), .Y(n1334) );
  INVX1 U2129 ( .A(n1546), .Y(n1556) );
  OAI221X1 U2130 ( .A(n1285), .B(n2838), .C(n1288), .D(n49), .E(n2843), .Y(
        n1546) );
  INVX1 U2131 ( .A(n1319), .Y(n2844) );
  OAI221X1 U2132 ( .A(n1311), .B(n1238), .C(n1312), .D(n1239), .E(n2827), .Y(
        n1319) );
  INVX1 U2133 ( .A(n1300), .Y(n2843) );
  OAI221X1 U2134 ( .A(n1301), .B(n1238), .C(n1302), .D(n1239), .E(n2827), .Y(
        n1300) );
  INVX1 U2135 ( .A(n530), .Y(cs_run) );
  NOR21XL U2136 ( .B(n2192), .A(n2191), .Y(n2214) );
  NOR8XL U2137 ( .A(multemp2[9]), .B(multemp2[8]), .C(multemp2[7]), .D(
        multemp2[6]), .E(multemp2[5]), .F(multemp2[4]), .G(multemp2[3]), .H(
        multemp2[2]), .Y(n2191) );
  AOI21X1 U2138 ( .B(n2840), .C(n61), .A(n2839), .Y(n307) );
  OAI221X1 U2139 ( .A(n1238), .B(n1523), .C(n1239), .D(n1522), .E(n2827), .Y(
        n1531) );
  INVX1 U2140 ( .A(n1521), .Y(n1522) );
  OAI22X1 U2141 ( .A(n1238), .B(n1513), .C(n1239), .D(n1512), .Y(n1524) );
  OA22XL U2142 ( .A(n2508), .B(n1670), .C(n2028), .D(n1956), .Y(n1678) );
  AND4X1 U2143 ( .A(n1669), .B(n1668), .C(n1667), .D(n1666), .Y(n1670) );
  AOI221XL U2144 ( .A(n1728), .B(n1663), .C(n1654), .D(n1653), .E(n1652), .Y(
        n1668) );
  AO21X1 U2145 ( .B(n1530), .C(n45), .A(n1466), .Y(n2310) );
  OAI21BBX1 U2146 ( .A(n1529), .B(n43), .C(n1426), .Y(n2340) );
  AOI22X1 U2147 ( .A(n2840), .B(n1312), .C(n2839), .D(n1311), .Y(n1318) );
  OA22X1 U2148 ( .A(n1239), .B(n1521), .C(n1238), .D(n1511), .Y(n308) );
  OAI21BBX1 U2149 ( .A(n1462), .B(n39), .C(n1530), .Y(n2387) );
  INVX1 U2150 ( .A(n1860), .Y(n1771) );
  NOR2X1 U2151 ( .A(n1310), .B(n2849), .Y(n1303) );
  NOR2X1 U2152 ( .A(n1328), .B(n2850), .Y(n1320) );
  INVX1 U2153 ( .A(n1511), .Y(n1523) );
  OAI21BBX1 U2154 ( .A(n1474), .B(n59), .C(n1462), .Y(n2102) );
  NOR2X1 U2155 ( .A(n1294), .B(n49), .Y(n1285) );
  INVX1 U2156 ( .A(n1512), .Y(n2819) );
  NAND3X1 U2157 ( .A(n37), .B(n51), .C(n2819), .Y(n1330) );
  NAND2X1 U2158 ( .A(n1743), .B(n1744), .Y(n2366) );
  NAND32X1 U2159 ( .B(n1741), .C(n1743), .A(n1744), .Y(n2368) );
  INVX1 U2160 ( .A(n2469), .Y(n1741) );
  AOI211X1 U2161 ( .C(n1961), .D(n2869), .A(n1735), .B(n1734), .Y(n1736) );
  AOI211X1 U2162 ( .C(n1726), .D(n1725), .A(n1724), .B(n1723), .Y(n1737) );
  MUX2X1 U2163 ( .D0(n1729), .D1(n1728), .S(n34), .Y(n1735) );
  AOI31XL U2164 ( .A(n1282), .B(n1281), .C(n1349), .D(n2028), .Y(n1291) );
  NAND21X1 U2165 ( .B(n1475), .A(n1474), .Y(n2250) );
  OAI2B11XL U2166 ( .D(n1304), .C(n167), .A(n2492), .B(n2645), .Y(n2590) );
  OA222X1 U2167 ( .A(n2160), .B(n2368), .C(n59), .D(n2367), .E(n2159), .F(
        n2366), .Y(n2161) );
  INVX1 U2168 ( .A(n1730), .Y(n1733) );
  INVX1 U2169 ( .A(n1740), .Y(n1744) );
  NAND21X1 U2170 ( .B(n1739), .A(n1742), .Y(n1740) );
  INVX1 U2171 ( .A(n1463), .Y(n1475) );
  INVX1 U2172 ( .A(n1513), .Y(n2818) );
  NAND3X1 U2173 ( .A(n37), .B(n51), .C(n2818), .Y(n1329) );
  NAND21XL U2174 ( .B(n212), .A(n1673), .Y(n2467) );
  NAND32X1 U2175 ( .B(n1739), .C(n2373), .A(n2589), .Y(n2493) );
  AND4X1 U2176 ( .A(n1998), .B(n1649), .C(n1648), .D(n1757), .Y(n1669) );
  INVX1 U2177 ( .A(n1739), .Y(n2588) );
  INVX1 U2178 ( .A(n1765), .Y(n2200) );
  INVX1 U2179 ( .A(n1280), .Y(n1712) );
  NAND21X1 U2180 ( .B(n2526), .A(n1673), .Y(n1280) );
  NAND21X1 U2181 ( .B(n1655), .A(n1623), .Y(n1661) );
  INVX1 U2182 ( .A(n2647), .Y(intcall) );
  INVX1 U2183 ( .A(n1628), .Y(n1650) );
  NAND43X1 U2184 ( .B(n1959), .C(n1627), .D(n169), .A(n2034), .Y(n1628) );
  OAI22XL U2185 ( .A(n1658), .B(n1897), .C(n1657), .D(n1656), .Y(n1660) );
  AND3XL U2186 ( .A(n1959), .B(n126), .C(n116), .Y(n1658) );
  AOI221XL U2187 ( .A(n1665), .B(n1664), .C(n2009), .D(n1663), .E(n1662), .Y(
        n1666) );
  NAND32XL U2188 ( .B(n1622), .C(n1663), .A(n1649), .Y(n1682) );
  OAI21BBX1 U2189 ( .A(n1475), .B(n61), .C(n1474), .Y(n1476) );
  OAI22XL U2190 ( .A(n212), .B(n1672), .C(n187), .D(n1671), .Y(n1675) );
  OR3XL U2191 ( .A(n2594), .B(n2555), .C(n1816), .Y(n1822) );
  NAND21X1 U2192 ( .B(n424), .A(n1632), .Y(n940) );
  OAI22X1 U2193 ( .A(n2815), .B(n940), .C(n941), .D(n2277), .Y(N12966) );
  OAI22X1 U2194 ( .A(n2814), .B(n940), .C(n941), .D(n2625), .Y(N12967) );
  OAI22X1 U2195 ( .A(n2848), .B(n940), .C(n2811), .D(n941), .Y(N12971) );
  INVX1 U2196 ( .A(n2560), .Y(n2577) );
  AND2X1 U2197 ( .A(n2652), .B(n2648), .Y(n2649) );
  AND2X1 U2198 ( .A(n2652), .B(n2651), .Y(n2653) );
  AND2XL U2199 ( .A(n2644), .B(n2643), .Y(sfroe_comb_s) );
  NAND4X1 U2200 ( .A(n594), .B(n595), .C(n596), .D(n597), .Y(dpl[2]) );
  OA22X1 U2201 ( .A(n367), .B(n2780), .C(n366), .D(n2779), .Y(n596) );
  NAND4X1 U2202 ( .A(n602), .B(n603), .C(n604), .D(n605), .Y(dpl[0]) );
  OA22X1 U2203 ( .A(n368), .B(n2770), .C(n2804), .D(n2769), .Y(n604) );
  NAND4X1 U2204 ( .A(n634), .B(n635), .C(n636), .D(n637), .Y(dph[0]) );
  OA22X1 U2205 ( .A(n365), .B(n2734), .C(n367), .D(n2733), .Y(n636) );
  INVX1 U2206 ( .A(N345), .Y(n2671) );
  NAND4X1 U2207 ( .A(n626), .B(n627), .C(n628), .D(n629), .Y(dph[2]) );
  OA22X1 U2208 ( .A(n2808), .B(n2746), .C(n2807), .D(n2745), .Y(n629) );
  AOI21XL U2209 ( .B(n2619), .C(n71), .A(n2617), .Y(n310) );
  MUX2X1 U2210 ( .D0(ramoe), .D1(n2620), .S(n422), .Y(ramoe_comb) );
  MUX2XL U2211 ( .D0(n1417), .D1(ramdatao[7]), .S(n1906), .Y(n1444) );
  MUX2XL U2212 ( .D0(n1904), .D1(n1415), .S(acc[7]), .Y(n1445) );
  NAND5X2 U2213 ( .A(n1075), .B(n1074), .C(n1073), .D(n1076), .E(n1072), .Y(
        n1436) );
  INVXL U2214 ( .A(dec_accop[8]), .Y(n1074) );
  INVX1 U2215 ( .A(dec_accop[7]), .Y(n1073) );
  INVX1 U2216 ( .A(dec_accop[16]), .Y(n1072) );
  INVXL U2217 ( .A(dec_accop[5]), .Y(n1081) );
  AO21XL U2218 ( .B(temp2_comb[2]), .C(n1913), .A(n1428), .Y(n1747) );
  XOR2XL U2219 ( .A(n1436), .B(acc[1]), .Y(n1427) );
  NAND21X1 U2220 ( .B(n2030), .A(mempsrd), .Y(n2032) );
  AND2X1 U2221 ( .A(n2541), .B(n2516), .Y(n2031) );
  OA2222XL U2222 ( .A(n2029), .B(n187), .C(n2527), .D(n2528), .E(n2525), .F(
        n2028), .G(n2027), .H(n2526), .Y(n2030) );
  MUX2XL U2223 ( .D0(N13339), .D1(divtempreg[2]), .S(N13343), .Y(n314) );
  XOR2XL U2224 ( .A(n1626), .B(ramsfraddr[0]), .Y(n522) );
  XOR2XL U2225 ( .A(n534), .B(ramsfraddr[2]), .Y(n521) );
  NAND21X1 U2226 ( .B(acc[1]), .A(n2263), .Y(n1418) );
  NOR41XL U2227 ( .D(ramwe), .A(n317), .B(n318), .C(n519), .Y(n520) );
  OAI221X1 U2228 ( .A(n1388), .B(n185), .C(n2644), .D(n1387), .E(n2645), .Y(
        n2620) );
  OA2222XL U2229 ( .A(n1725), .B(n1386), .C(instr[5]), .D(n2011), .E(instr[3]), 
        .F(n1385), .G(n1384), .H(n1621), .Y(n1388) );
  INVX1 U2230 ( .A(n2643), .Y(n1387) );
  OA22XL U2231 ( .A(n1657), .B(n1383), .C(n1959), .D(n1382), .Y(n1385) );
  INVX1 U2232 ( .A(rn_reg[44]), .Y(n715) );
  INVX1 U2233 ( .A(rn_reg[12]), .Y(n714) );
  INVX1 U2234 ( .A(rn_reg[43]), .Y(n759) );
  INVX1 U2235 ( .A(rn_reg[11]), .Y(n758) );
  INVX1 U2236 ( .A(rn_reg[169]), .Y(n789) );
  INVX1 U2237 ( .A(rn_reg[137]), .Y(n788) );
  INVX1 U2238 ( .A(rn_reg[168]), .Y(n655) );
  INVX1 U2239 ( .A(rn_reg[136]), .Y(n654) );
  INVX1 U2240 ( .A(rn_reg[172]), .Y(n700) );
  INVX1 U2241 ( .A(rn_reg[140]), .Y(n699) );
  INVX1 U2242 ( .A(rn_reg[171]), .Y(n744) );
  INVX1 U2243 ( .A(rn_reg[139]), .Y(n743) );
  NAND4X1 U2244 ( .A(n319), .B(n320), .C(n321), .D(n1919), .Y(n2057) );
  AOI21XL U2245 ( .B(n1906), .C(ramdatao[6]), .A(n1905), .Y(n319) );
  OA22X1 U2246 ( .A(n2383), .B(n1922), .C(n263), .D(n2411), .Y(n320) );
  AOI22XL U2247 ( .A(multemp1_0_), .B(n2192), .C(acc[2]), .D(n1907), .Y(n321)
         );
  NAND21X1 U2248 ( .B(n1124), .A(instr[5]), .Y(n1323) );
  OAI21AX1 U2249 ( .B(sfroe_r), .C(sfrwe_r), .A(sfrack), .Y(n2697) );
  OA222X1 U2250 ( .A(n1918), .B(n2294), .C(n1917), .D(n2344), .E(n293), .F(
        n1916), .Y(n1919) );
  XOR3XL U2251 ( .A(n1915), .B(n346), .C(n1914), .Y(n1916) );
  MUX2XL U2252 ( .D0(N13341), .D1(divtempreg[4]), .S(N13343), .Y(n322) );
  MUX2XL U2253 ( .D0(N13340), .D1(divtempreg[3]), .S(N13343), .Y(n323) );
  OAI221XL U2254 ( .A(n157), .B(n846), .C(n141), .D(n845), .E(n968), .Y(n847)
         );
  INVX1 U2255 ( .A(rn_reg[45]), .Y(n846) );
  INVX1 U2256 ( .A(rn_reg[13]), .Y(n845) );
  XNOR2XL U2257 ( .A(n1436), .B(acc[2]), .Y(n326) );
  OAI221XL U2258 ( .A(n157), .B(n804), .C(n141), .D(n803), .E(n968), .Y(n805)
         );
  INVX1 U2259 ( .A(rn_reg[41]), .Y(n804) );
  INVX1 U2260 ( .A(rn_reg[9]), .Y(n803) );
  INVX1 U2261 ( .A(rn_reg[40]), .Y(n670) );
  INVX1 U2262 ( .A(rn_reg[8]), .Y(n669) );
  OAI221XL U2263 ( .A(n157), .B(n831), .C(n141), .D(n830), .E(n220), .Y(n832)
         );
  INVX1 U2264 ( .A(rn_reg[173]), .Y(n831) );
  INVX1 U2265 ( .A(rn_reg[141]), .Y(n830) );
  OAI221XL U2266 ( .A(n157), .B(n532), .C(n141), .D(n531), .E(n220), .Y(n533)
         );
  INVX1 U2267 ( .A(rn_reg[170]), .Y(n532) );
  INVX1 U2268 ( .A(rn_reg[138]), .Y(n531) );
  GEN2XL U2269 ( .D(acc[7]), .E(n1421), .C(c), .B(n1420), .A(n1689), .Y(n1912)
         );
  NAND32X1 U2270 ( .B(acc[5]), .C(n1419), .A(n2329), .Y(n1421) );
  AND3XL U2271 ( .A(acc[3]), .B(acc[4]), .C(n1418), .Y(n1419) );
  NAND21XL U2272 ( .B(n2872), .A(n1626), .Y(n1283) );
  MUX2IX1 U2273 ( .D0(n327), .D1(n328), .S(n1256), .Y(n1253) );
  NAND2X1 U2274 ( .A(dps[1]), .B(n1255), .Y(n327) );
  MUX2IXL U2275 ( .D0(ramdatao[1]), .D1(rs[0]), .S(ramdatao[3]), .Y(n328) );
  NAND21X1 U2276 ( .B(n2872), .A(n2873), .Y(n1711) );
  INVX1 U2277 ( .A(dec_accop[13]), .Y(n1062) );
  AO222X1 U2278 ( .A(n1540), .B(temp[5]), .C(dptr_inc[5]), .D(n1590), .E(n1539), .F(n237), .Y(n1929) );
  AO222X1 U2279 ( .A(n1540), .B(temp[6]), .C(dptr_inc[6]), .D(n1590), .E(n1539), .F(n238), .Y(n1928) );
  AO222XL U2280 ( .A(n1540), .B(temp[1]), .C(dptr_inc[1]), .D(n1590), .E(n1539), .F(n224), .Y(n1933) );
  MUX2IXL U2281 ( .D0(ramdatao[2]), .D1(rs[1]), .S(n135), .Y(n330) );
  NAND21XL U2282 ( .B(n2015), .A(n2871), .Y(n534) );
  NAND43X1 U2283 ( .B(n1802), .C(n1801), .D(n1800), .A(n1799), .Y(n1936) );
  OAI22XL U2284 ( .A(n1817), .B(n2411), .C(n1791), .D(n1964), .Y(n1800) );
  AO21XL U2285 ( .B(ramdatao[5]), .C(n1906), .A(n1790), .Y(n1802) );
  NAND43X1 U2286 ( .B(n1697), .C(n1696), .D(n1695), .A(n1694), .Y(n1938) );
  OAI22XL U2287 ( .A(n1817), .B(n2329), .C(n1791), .D(n1965), .Y(n1695) );
  OAI22XL U2288 ( .A(n2263), .B(n1922), .C(n263), .D(n2294), .Y(n1696) );
  AO21XL U2289 ( .B(ramdatao[4]), .C(n1906), .A(n1686), .Y(n1697) );
  NAND21XL U2290 ( .B(n2873), .A(n2872), .Y(n1382) );
  NAND21XL U2291 ( .B(n2873), .A(n783), .Y(n545) );
  XOR2XL U2292 ( .A(n1436), .B(acc[3]), .Y(n1703) );
  NAND21XL U2293 ( .B(ramsfraddr[4]), .A(n2569), .Y(n2573) );
  INVX1 U2294 ( .A(n1053), .Y(n1904) );
  NAND43X1 U2295 ( .B(n1067), .C(n1052), .D(dec_accop[13]), .A(n344), .Y(n1053) );
  INVX1 U2296 ( .A(dec_accop[15]), .Y(n1052) );
  NAND21X1 U2297 ( .B(n1655), .A(n213), .Y(n1372) );
  NAND21XL U2298 ( .B(ramsfraddr[6]), .A(n2555), .Y(n519) );
  INVX1 U2299 ( .A(rn_reg[49]), .Y(n817) );
  INVX1 U2300 ( .A(rn_reg[113]), .Y(n816) );
  INVX1 U2301 ( .A(rn_reg[97]), .Y(n815) );
  OA2222XL U2302 ( .A(n999), .B(n683), .C(n997), .D(n682), .E(n995), .F(n681), 
        .G(n993), .H(n680), .Y(n684) );
  INVX1 U2303 ( .A(rn_reg[48]), .Y(n683) );
  INVX1 U2304 ( .A(rn_reg[96]), .Y(n681) );
  INVX1 U2305 ( .A(rn_reg[112]), .Y(n682) );
  OA2222XL U2306 ( .A(n999), .B(n728), .C(n997), .D(n727), .E(n995), .F(n726), 
        .G(n993), .H(n725), .Y(n729) );
  INVX1 U2307 ( .A(rn_reg[52]), .Y(n728) );
  INVX1 U2308 ( .A(rn_reg[116]), .Y(n727) );
  INVX1 U2309 ( .A(rn_reg[100]), .Y(n726) );
  OA2222XL U2310 ( .A(n999), .B(n772), .C(n997), .D(n771), .E(n995), .F(n770), 
        .G(n993), .H(n769), .Y(n773) );
  INVX1 U2311 ( .A(rn_reg[51]), .Y(n772) );
  INVX1 U2312 ( .A(rn_reg[99]), .Y(n770) );
  INVX1 U2313 ( .A(rn_reg[115]), .Y(n771) );
  INVX1 U2314 ( .A(rn_reg[33]), .Y(n813) );
  INVX1 U2315 ( .A(rn_reg[17]), .Y(n812) );
  INVX1 U2316 ( .A(rn_reg[121]), .Y(n811) );
  OA2222XL U2317 ( .A(n991), .B(n679), .C(n989), .D(n678), .E(n987), .F(n677), 
        .G(n985), .H(n676), .Y(n685) );
  INVX1 U2318 ( .A(rn_reg[32]), .Y(n679) );
  INVX1 U2319 ( .A(rn_reg[120]), .Y(n677) );
  INVX1 U2320 ( .A(rn_reg[16]), .Y(n678) );
  OA2222XL U2321 ( .A(n991), .B(n724), .C(n989), .D(n723), .E(n987), .F(n722), 
        .G(n985), .H(n721), .Y(n730) );
  INVX1 U2322 ( .A(rn_reg[36]), .Y(n724) );
  INVX1 U2323 ( .A(rn_reg[20]), .Y(n723) );
  INVX1 U2324 ( .A(rn_reg[124]), .Y(n722) );
  OA2222XL U2325 ( .A(n991), .B(n768), .C(n989), .D(n767), .E(n987), .F(n766), 
        .G(n985), .H(n765), .Y(n774) );
  INVX1 U2326 ( .A(rn_reg[35]), .Y(n768) );
  INVX1 U2327 ( .A(rn_reg[123]), .Y(n766) );
  INVX1 U2328 ( .A(rn_reg[19]), .Y(n767) );
  OA2222XL U2329 ( .A(n196), .B(n802), .C(n159), .D(n801), .E(n175), .F(n800), 
        .G(n142), .H(n799), .Y(n822) );
  INVX1 U2330 ( .A(rn_reg[177]), .Y(n802) );
  INVX1 U2331 ( .A(rn_reg[241]), .Y(n801) );
  INVX1 U2332 ( .A(rn_reg[225]), .Y(n800) );
  OA2222XL U2333 ( .A(n999), .B(n668), .C(n997), .D(n667), .E(n995), .F(n666), 
        .G(n993), .H(n665), .Y(n688) );
  INVX1 U2334 ( .A(rn_reg[176]), .Y(n668) );
  INVX1 U2335 ( .A(rn_reg[224]), .Y(n666) );
  INVX1 U2336 ( .A(rn_reg[240]), .Y(n667) );
  OA2222XL U2337 ( .A(n999), .B(n713), .C(n997), .D(n712), .E(n995), .F(n711), 
        .G(n993), .H(n710), .Y(n733) );
  INVX1 U2338 ( .A(rn_reg[180]), .Y(n713) );
  INVX1 U2339 ( .A(rn_reg[244]), .Y(n712) );
  INVX1 U2340 ( .A(rn_reg[228]), .Y(n711) );
  OA2222XL U2341 ( .A(n999), .B(n757), .C(n997), .D(n756), .E(n995), .F(n755), 
        .G(n993), .H(n754), .Y(n777) );
  INVX1 U2342 ( .A(rn_reg[179]), .Y(n757) );
  INVX1 U2343 ( .A(rn_reg[227]), .Y(n755) );
  INVX1 U2344 ( .A(rn_reg[243]), .Y(n756) );
  OA2222XL U2345 ( .A(n130), .B(n798), .C(n174), .D(n797), .E(n158), .F(n796), 
        .G(n197), .H(n795), .Y(n823) );
  INVX1 U2346 ( .A(rn_reg[161]), .Y(n798) );
  INVX1 U2347 ( .A(rn_reg[145]), .Y(n797) );
  INVX1 U2348 ( .A(rn_reg[249]), .Y(n796) );
  OA2222XL U2349 ( .A(n991), .B(n664), .C(n989), .D(n663), .E(n987), .F(n662), 
        .G(n985), .H(n661), .Y(n689) );
  INVX1 U2350 ( .A(rn_reg[160]), .Y(n664) );
  INVX1 U2351 ( .A(rn_reg[248]), .Y(n662) );
  INVX1 U2352 ( .A(rn_reg[144]), .Y(n663) );
  OA2222XL U2353 ( .A(n991), .B(n709), .C(n989), .D(n708), .E(n987), .F(n707), 
        .G(n985), .H(n706), .Y(n734) );
  INVX1 U2354 ( .A(rn_reg[164]), .Y(n709) );
  INVX1 U2355 ( .A(rn_reg[148]), .Y(n708) );
  INVX1 U2356 ( .A(rn_reg[252]), .Y(n707) );
  OA2222XL U2357 ( .A(n991), .B(n753), .C(n989), .D(n752), .E(n987), .F(n751), 
        .G(n985), .H(n750), .Y(n778) );
  INVX1 U2358 ( .A(rn_reg[163]), .Y(n753) );
  INVX1 U2359 ( .A(rn_reg[251]), .Y(n751) );
  INVX1 U2360 ( .A(rn_reg[147]), .Y(n752) );
  OA222X1 U2361 ( .A(n1918), .B(n2383), .C(n1798), .D(n2313), .E(n293), .F(
        n1797), .Y(n1799) );
  XOR3XL U2362 ( .A(n1796), .B(n1795), .C(n1794), .Y(n1797) );
  MUX2XL U2363 ( .D0(n1909), .D1(n1908), .S(acc[5]), .Y(n1792) );
  OA222X1 U2364 ( .A(n1918), .B(n2116), .C(n1693), .D(n2396), .E(n293), .F(
        n1692), .Y(n1694) );
  XOR3X1 U2365 ( .A(n1691), .B(n349), .C(n1761), .Y(n1692) );
  MUX2XL U2366 ( .D0(n150), .D1(n1908), .S(acc[4]), .Y(n1687) );
  NAND21XL U2367 ( .B(n783), .A(n2873), .Y(n537) );
  MUX2X1 U2368 ( .D0(pc_o[3]), .D1(n1931), .S(n1934), .Y(N12844) );
  MUX2X1 U2369 ( .D0(memaddr[4]), .D1(n1930), .S(n1934), .Y(N12845) );
  MUX2X1 U2370 ( .D0(pc_o[2]), .D1(n1932), .S(n1934), .Y(N12843) );
  MUX2X1 U2371 ( .D0(memaddr[5]), .D1(n1929), .S(n1934), .Y(N12846) );
  MUX2X1 U2372 ( .D0(memaddr[6]), .D1(n1928), .S(n1934), .Y(N12847) );
  AOI211X1 U2373 ( .C(dec_accop[14]), .D(n1767), .A(n1904), .B(n1766), .Y(
        n1768) );
  MUX2XL U2374 ( .D0(n1909), .D1(n1908), .S(temp2_comb[0]), .Y(n1188) );
  NAND21XL U2375 ( .B(n2182), .A(n2873), .Y(n546) );
  MUX2BXL U2376 ( .D0(n1904), .D1(n331), .S(acc[2]), .Y(n1745) );
  AOI21XL U2377 ( .B(n1903), .C(n2257), .A(n1902), .Y(n331) );
  AO21XL U2378 ( .B(ramdatao[0]), .C(n1906), .A(n1191), .Y(n1196) );
  AND2X1 U2379 ( .A(n1189), .B(n1188), .Y(n1190) );
  INVX1 U2380 ( .A(n1902), .Y(n1189) );
  NAND21XL U2381 ( .B(n2868), .A(n2867), .Y(n444) );
  AOI21XL U2382 ( .B(temp2_comb[3]), .C(n1913), .A(n1689), .Y(n333) );
  AOI21X1 U2383 ( .B(accactv), .C(n1051), .A(n1054), .Y(n334) );
  AO2222XL U2384 ( .A(n1010), .B(ramsfraddr[6]), .C(temp[6]), .D(n1011), .E(
        n2053), .F(n1012), .G(n2352), .H(n1013), .Y(n923) );
  INVX1 U2385 ( .A(rn_reg[47]), .Y(n971) );
  INVX1 U2386 ( .A(rn_reg[15]), .Y(n969) );
  MUX2XL U2387 ( .D0(N13342), .D1(divtempreg[5]), .S(N13343), .Y(n335) );
  INVXL U2388 ( .A(ramsfraddr[3]), .Y(n2569) );
  OAI221XL U2389 ( .A(n157), .B(n564), .C(n141), .D(n563), .E(n968), .Y(n565)
         );
  INVX1 U2390 ( .A(rn_reg[42]), .Y(n564) );
  INVX1 U2391 ( .A(rn_reg[10]), .Y(n563) );
  OAI221XL U2392 ( .A(n157), .B(n899), .C(n141), .D(n898), .E(n968), .Y(n900)
         );
  INVX1 U2393 ( .A(rn_reg[46]), .Y(n899) );
  INVX1 U2394 ( .A(rn_reg[14]), .Y(n898) );
  OAI221XL U2395 ( .A(n157), .B(n953), .C(n141), .D(n952), .E(n220), .Y(n954)
         );
  INVX1 U2396 ( .A(rn_reg[175]), .Y(n953) );
  INVX1 U2397 ( .A(rn_reg[143]), .Y(n952) );
  OAI221XL U2398 ( .A(n157), .B(n884), .C(n141), .D(n883), .E(n220), .Y(n885)
         );
  INVX1 U2399 ( .A(rn_reg[174]), .Y(n884) );
  INVX1 U2400 ( .A(rn_reg[142]), .Y(n883) );
  NAND21XL U2401 ( .B(n2554), .A(ramsfrwe), .Y(n450) );
  NAND21X1 U2402 ( .B(N344), .A(N343), .Y(n2665) );
  NAND21X1 U2403 ( .B(N343), .A(n1024), .Y(n2668) );
  MUX4XL U2404 ( .D0(ckcon[7]), .D1(ramdatao[7]), .D2(ckcon[3]), .D3(
        ramdatao[3]), .S0(n1633), .S1(n336), .Y(n462) );
  MUX2IXL U2405 ( .D0(pmw), .D1(ramdatao[4]), .S(n1815), .Y(n336) );
  INVX1 U2406 ( .A(n1069), .Y(n1070) );
  AOI21XL U2407 ( .B(n1651), .C(n2870), .A(n2109), .Y(n337) );
  NAND31XL U2408 ( .C(n1068), .A(dec_accop[11]), .B(n288), .Y(n1910) );
  AO222XL U2409 ( .A(n1540), .B(temp[0]), .C(dptr_inc[0]), .D(n1590), .E(n1539), .F(n226), .Y(n1935) );
  MUX2AXL U2410 ( .D0(sp[4]), .D1(n2628), .S(n947), .Y(n696) );
  NAND21XL U2411 ( .B(n204), .A(n419), .Y(n1973) );
  OA2222XL U2412 ( .A(dpl_reg[11]), .B(n1584), .C(dpl_reg[3]), .D(n1583), .E(
        dpl_reg[43]), .F(n1582), .G(dpl_reg[35]), .H(n1581), .Y(n1470) );
  OA2222XL U2413 ( .A(dpl_reg[12]), .B(n1584), .C(dpl_reg[4]), .D(n1583), .E(
        dpl_reg[44]), .F(n1582), .G(dpl_reg[36]), .H(n1581), .Y(n1459) );
  OA2222XL U2414 ( .A(dpl_reg[13]), .B(n1584), .C(dpl_reg[5]), .D(n1583), .E(
        dpl_reg[45]), .F(n1582), .G(dpl_reg[37]), .H(n1581), .Y(n1535) );
  OA2222XL U2415 ( .A(dpl_reg[14]), .B(n1584), .C(dpl_reg[6]), .D(n1583), .E(
        dpl_reg[46]), .F(n1582), .G(dpl_reg[38]), .H(n1581), .Y(n1526) );
  NAND21XL U2416 ( .B(n2873), .A(n2033), .Y(n1370) );
  NOR42XL U2417 ( .C(n1681), .D(n2528), .A(phase[4]), .B(phase[5]), .Y(n495)
         );
  NAND21XL U2418 ( .B(n2867), .A(n1324), .Y(n1778) );
  MUX2X1 U2419 ( .D0(n1835), .D1(n1834), .S(N345), .Y(n1840) );
  AO2222XL U2420 ( .A(n2343), .B(temp[2]), .C(n1833), .D(temp[1]), .E(n2436), 
        .F(temp[3]), .G(n2669), .H(temp[0]), .Y(n1835) );
  AO2222XL U2421 ( .A(n2343), .B(temp[6]), .C(n1833), .D(temp[5]), .E(n2436), 
        .F(temp[7]), .G(n2669), .H(temp[4]), .Y(n1834) );
  NAND21XL U2422 ( .B(n1092), .A(phase[1]), .Y(n1047) );
  NAND21XL U2423 ( .B(n1124), .A(n183), .Y(n483) );
  NAND21XL U2424 ( .B(n2870), .A(n2871), .Y(n1647) );
  MUX2XL U2425 ( .D0(n1041), .D1(n2591), .S(pc_o[1]), .Y(n1104) );
  OAI22XL U2426 ( .A(n2459), .B(n2439), .C(n2850), .D(n2445), .Y(n1103) );
  OA22X1 U2427 ( .A(n2444), .B(n2456), .C(n2442), .D(n2470), .Y(n1101) );
  NAND5XL U2428 ( .A(dec_accop[17]), .B(n1767), .C(n1861), .D(n1860), .E(n1076), .Y(n1922) );
  NAND21XL U2429 ( .B(instr[5]), .A(n1896), .Y(n1110) );
  XOR2XL U2430 ( .A(n1436), .B(acc[4]), .Y(n1688) );
  XOR2XL U2431 ( .A(n1436), .B(acc[5]), .Y(n1793) );
  AO21X1 U2432 ( .B(n1095), .C(n1378), .A(n2251), .Y(n2297) );
  AOI32XL U2433 ( .A(n1360), .B(phase[0]), .C(n1094), .D(n1990), .E(n1093), 
        .Y(n1095) );
  OAI31XL U2434 ( .A(n1647), .B(n1626), .C(n167), .D(n1375), .Y(n1093) );
  NAND21XL U2435 ( .B(n1275), .A(ramsfraddr[2]), .Y(n2557) );
  NAND21XL U2436 ( .B(n2561), .A(ramsfraddr[0]), .Y(n1275) );
  NAND32XL U2437 ( .B(ramsfraddr[2]), .C(n2561), .A(n2559), .Y(n1409) );
  NAND32X1 U2438 ( .B(dec_accop[15]), .C(dec_accop[13]), .A(n344), .Y(n1069)
         );
  OAI211X1 U2439 ( .C(n494), .D(n2528), .A(n493), .B(n492), .Y(n2522) );
  AOI222XL U2440 ( .A(phase[4]), .B(n2524), .C(phase[1]), .D(n491), .E(
        phase[0]), .F(n490), .Y(n492) );
  AOI22X1 U2441 ( .A(n1127), .B(n460), .C(phase[2]), .D(n459), .Y(n493) );
  OA2222XL U2442 ( .A(n196), .B(n641), .C(n159), .D(n640), .E(n175), .F(n639), 
        .G(n142), .H(n638), .Y(n642) );
  INVX1 U2443 ( .A(rn_reg[50]), .Y(n641) );
  INVX1 U2444 ( .A(rn_reg[114]), .Y(n640) );
  INVX1 U2445 ( .A(rn_reg[98]), .Y(n639) );
  OA2222XL U2446 ( .A(n130), .B(n855), .C(n174), .D(n854), .E(n158), .F(n853), 
        .G(n197), .H(n852), .Y(n861) );
  INVX1 U2447 ( .A(rn_reg[37]), .Y(n855) );
  INVX1 U2448 ( .A(rn_reg[125]), .Y(n853) );
  INVX1 U2449 ( .A(rn_reg[21]), .Y(n854) );
  OA2222XL U2450 ( .A(n130), .B(n577), .C(n174), .D(n576), .E(n158), .F(n575), 
        .G(n197), .H(n574), .Y(n643) );
  INVX1 U2451 ( .A(rn_reg[34]), .Y(n577) );
  INVX1 U2452 ( .A(rn_reg[18]), .Y(n576) );
  INVX1 U2453 ( .A(rn_reg[122]), .Y(n575) );
  OA2222XL U2454 ( .A(n991), .B(n990), .C(n989), .D(n988), .E(n987), .F(n986), 
        .G(n985), .H(n984), .Y(n1001) );
  INVX1 U2455 ( .A(rn_reg[39]), .Y(n990) );
  INVX1 U2456 ( .A(rn_reg[127]), .Y(n986) );
  INVX1 U2457 ( .A(rn_reg[23]), .Y(n988) );
  OA2222XL U2458 ( .A(n130), .B(n908), .C(n174), .D(n907), .E(n158), .F(n906), 
        .G(n197), .H(n905), .Y(n914) );
  INVX1 U2459 ( .A(rn_reg[38]), .Y(n908) );
  INVX1 U2460 ( .A(rn_reg[126]), .Y(n906) );
  INVX1 U2461 ( .A(rn_reg[22]), .Y(n907) );
  OA2222XL U2462 ( .A(n196), .B(n560), .C(n159), .D(n559), .E(n175), .F(n558), 
        .G(n142), .H(n557), .Y(n646) );
  INVX1 U2463 ( .A(rn_reg[178]), .Y(n560) );
  INVX1 U2464 ( .A(rn_reg[242]), .Y(n559) );
  INVX1 U2465 ( .A(rn_reg[226]), .Y(n558) );
  OA2222XL U2466 ( .A(n130), .B(n840), .C(n174), .D(n839), .E(n158), .F(n838), 
        .G(n197), .H(n837), .Y(n865) );
  INVX1 U2467 ( .A(rn_reg[165]), .Y(n840) );
  INVX1 U2468 ( .A(rn_reg[253]), .Y(n838) );
  INVX1 U2469 ( .A(rn_reg[149]), .Y(n839) );
  OA2222XL U2470 ( .A(n130), .B(n551), .C(n174), .D(n550), .E(n158), .F(n549), 
        .G(n197), .H(n548), .Y(n647) );
  INVX1 U2471 ( .A(rn_reg[162]), .Y(n551) );
  INVX1 U2472 ( .A(rn_reg[146]), .Y(n550) );
  INVX1 U2473 ( .A(rn_reg[250]), .Y(n549) );
  OA2222XL U2474 ( .A(n991), .B(n963), .C(n989), .D(n962), .E(n987), .F(n961), 
        .G(n985), .H(n960), .Y(n1005) );
  INVX1 U2475 ( .A(rn_reg[167]), .Y(n963) );
  INVX1 U2476 ( .A(rn_reg[255]), .Y(n961) );
  INVX1 U2477 ( .A(rn_reg[151]), .Y(n962) );
  OA2222XL U2478 ( .A(n130), .B(n893), .C(n174), .D(n892), .E(n158), .F(n891), 
        .G(n197), .H(n890), .Y(n918) );
  INVX1 U2479 ( .A(rn_reg[166]), .Y(n893) );
  INVX1 U2480 ( .A(rn_reg[254]), .Y(n891) );
  INVX1 U2481 ( .A(rn_reg[150]), .Y(n892) );
  OA2222XL U2482 ( .A(n198), .B(n836), .C(n160), .D(n835), .E(n143), .F(n834), 
        .G(n176), .H(n833), .Y(n866) );
  INVX1 U2483 ( .A(rn_reg[189]), .Y(n836) );
  INVX1 U2484 ( .A(rn_reg[237]), .Y(n834) );
  INVX1 U2485 ( .A(rn_reg[133]), .Y(n835) );
  OA2222XL U2486 ( .A(n983), .B(n959), .C(n981), .D(n958), .E(n979), .F(n956), 
        .G(n977), .H(n955), .Y(n1006) );
  INVX1 U2487 ( .A(rn_reg[191]), .Y(n959) );
  INVX1 U2488 ( .A(rn_reg[239]), .Y(n956) );
  INVX1 U2489 ( .A(rn_reg[135]), .Y(n958) );
  OA2222XL U2490 ( .A(n198), .B(n889), .C(n160), .D(n888), .E(n143), .F(n887), 
        .G(n176), .H(n886), .Y(n919) );
  INVX1 U2491 ( .A(rn_reg[190]), .Y(n889) );
  INVX1 U2492 ( .A(rn_reg[238]), .Y(n887) );
  INVX1 U2493 ( .A(rn_reg[134]), .Y(n888) );
  OA2222XL U2494 ( .A(n198), .B(n851), .C(n160), .D(n850), .E(n143), .F(n849), 
        .G(n176), .H(n848), .Y(n862) );
  INVX1 U2495 ( .A(rn_reg[61]), .Y(n851) );
  INVX1 U2496 ( .A(rn_reg[109]), .Y(n849) );
  INVX1 U2497 ( .A(rn_reg[5]), .Y(n850) );
  OA2222XL U2498 ( .A(n983), .B(n982), .C(n981), .D(n980), .E(n979), .F(n978), 
        .G(n977), .H(n976), .Y(n1002) );
  INVX1 U2499 ( .A(rn_reg[63]), .Y(n982) );
  INVX1 U2500 ( .A(rn_reg[111]), .Y(n978) );
  INVX1 U2501 ( .A(rn_reg[7]), .Y(n980) );
  OA2222XL U2502 ( .A(n198), .B(n904), .C(n160), .D(n903), .E(n143), .F(n902), 
        .G(n176), .H(n901), .Y(n915) );
  INVX1 U2503 ( .A(rn_reg[62]), .Y(n904) );
  INVX1 U2504 ( .A(rn_reg[110]), .Y(n902) );
  INVX1 U2505 ( .A(rn_reg[6]), .Y(n903) );
  NAND43X1 U2506 ( .B(dec_accop[3]), .C(n1064), .D(n191), .A(dec_accop[4]), 
        .Y(n1873) );
  MUX2XL U2507 ( .D0(memaddr[0]), .D1(n1935), .S(n1934), .Y(N12841) );
  MUX2XL U2508 ( .D0(n1938), .D1(temp[4]), .S(n1980), .Y(N12828) );
  MUX2XL U2509 ( .D0(n2158), .D1(temp[3]), .S(n1980), .Y(N12827) );
  MUX2XL U2510 ( .D0(n1936), .D1(temp[5]), .S(n1980), .Y(N12829) );
  MUX2XL U2511 ( .D0(n2057), .D1(temp[6]), .S(n1980), .Y(N12830) );
  INVX1 U2512 ( .A(n2014), .Y(n2525) );
  OAI221XL U2513 ( .A(n204), .B(n2013), .C(n2012), .D(n2011), .E(n2010), .Y(
        n2014) );
  AOI211XL U2514 ( .C(n2015), .D(n2009), .A(n2008), .B(n2007), .Y(n2010) );
  GEN2XL U2515 ( .D(n1787), .E(n469), .C(n2023), .B(n458), .A(n2024), .Y(n459)
         );
  MUX2XL U2516 ( .D0(n453), .D1(n2020), .S(instr[6]), .Y(n458) );
  AND2XL U2517 ( .A(interrupt), .B(n1156), .Y(n453) );
  AND2XL U2518 ( .A(sfrwe_r), .B(n422), .Y(sfrwe) );
  XOR2XL U2519 ( .A(n1436), .B(acc[6]), .Y(n1914) );
  XOR2XL U2520 ( .A(n1436), .B(acc[7]), .Y(n1868) );
  MUX2BXL U2521 ( .D0(n1904), .D1(n338), .S(acc[5]), .Y(n1790) );
  AOI21XL U2522 ( .B(n1903), .C(n2313), .A(n1902), .Y(n338) );
  MUX2BXL U2523 ( .D0(n1904), .D1(n339), .S(acc[6]), .Y(n1905) );
  AOI21XL U2524 ( .B(n1903), .C(n2344), .A(n1902), .Y(n339) );
  MUX2BXL U2525 ( .D0(n1904), .D1(n340), .S(acc[4]), .Y(n1686) );
  AOI21XL U2526 ( .B(n1903), .C(n2396), .A(n1902), .Y(n340) );
  MUX2XL U2527 ( .D0(n1909), .D1(n1908), .S(acc[7]), .Y(n1438) );
  MUX2BXL U2528 ( .D0(n1904), .D1(n341), .S(acc[3]), .Y(n1701) );
  AOI21XL U2529 ( .B(n1903), .C(n2160), .A(n1902), .Y(n341) );
  MUX2BXL U2530 ( .D0(n1904), .D1(n342), .S(acc[1]), .Y(n1056) );
  AOI21XL U2531 ( .B(n1903), .C(n2459), .A(n1902), .Y(n342) );
  INVXL U2532 ( .A(n2872), .Y(n1157) );
  OA21XL U2533 ( .B(acc[0]), .C(n1909), .A(n1910), .Y(n1193) );
  GEN3XL U2534 ( .F(dec_cop[6]), .G(c), .E(dec_cop[5]), .D(n1847), .C(n1842), 
        .B(n1854), .A(n1841), .Y(n1844) );
  MUX2XL U2535 ( .D0(n1837), .D1(dec_cop[5]), .S(c), .Y(n1842) );
  OA21XL U2536 ( .B(c), .C(n1840), .A(dec_cop[3]), .Y(n1841) );
  AND3X1 U2537 ( .A(dec_cop[7]), .B(n1852), .C(n1836), .Y(n1837) );
  MUX2BXL U2538 ( .D0(sp[3]), .D1(n2275), .S(n947), .Y(n343) );
  INVX1 U2539 ( .A(phase[2]), .Y(n2526) );
  INVXL U2540 ( .A(ramsfraddr[0]), .Y(n2559) );
  NAND32XL U2541 ( .B(ramsfraddr[2]), .C(n2559), .A(n2561), .Y(n512) );
  OAI221XL U2542 ( .A(n2871), .B(n452), .C(n183), .D(n1383), .E(n1730), .Y(
        n2020) );
  OA21XL U2543 ( .B(n451), .C(n325), .A(n1627), .Y(n452) );
  INVX1 U2544 ( .A(n464), .Y(n451) );
  OAI32X1 U2545 ( .A(n1848), .B(n1856), .C(n1847), .D(n1846), .E(n191), .Y(
        n1871) );
  OA21X1 U2546 ( .B(n1831), .C(n1839), .A(n1859), .Y(n1848) );
  AOI31X1 U2547 ( .A(n1844), .B(n1859), .C(n1843), .D(dec_cop[0]), .Y(n1846)
         );
  INVX1 U2548 ( .A(dec_cop[1]), .Y(n1843) );
  INVXL U2549 ( .A(acc[7]), .Y(n2411) );
  AND2XL U2550 ( .A(n1746), .B(n1910), .Y(n1749) );
  MUX2XL U2551 ( .D0(n1909), .D1(n1908), .S(acc[2]), .Y(n1746) );
  AND2XL U2552 ( .A(n1702), .B(n1910), .Y(n1706) );
  MUX2XL U2553 ( .D0(n1909), .D1(n1908), .S(acc[3]), .Y(n1702) );
  AND2XL U2554 ( .A(n1066), .B(n1910), .Y(n1086) );
  MUX2XL U2555 ( .D0(n1909), .D1(n1908), .S(acc[1]), .Y(n1066) );
  INVX1 U2556 ( .A(n1050), .Y(n1058) );
  NAND21X1 U2557 ( .B(n1845), .A(dec_accop[1]), .Y(n1050) );
  INVXL U2558 ( .A(ramsfraddr[2]), .Y(n2562) );
  INVX1 U2559 ( .A(temp2_comb[5]), .Y(n2313) );
  INVXL U2560 ( .A(n2869), .Y(n419) );
  INVX1 U2561 ( .A(N344), .Y(n1024) );
  INVX1 U2562 ( .A(interrupt), .Y(n2533) );
  INVX1 U2563 ( .A(dec_accop[4]), .Y(n1850) );
  NAND21XL U2564 ( .B(n185), .A(n2870), .Y(n1375) );
  MUX2AXL U2565 ( .D0(sp[5]), .D1(n2630), .S(n947), .Y(n871) );
  NAND21XL U2566 ( .B(n204), .A(n1384), .Y(n1716) );
  MUX2AXL U2567 ( .D0(sp[6]), .D1(n2811), .S(n947), .Y(n943) );
  NAND21XL U2568 ( .B(n1845), .A(dec_accop[16]), .Y(n1861) );
  NAND21XL U2569 ( .B(instr[7]), .A(n2867), .Y(n1720) );
  NAND21XL U2570 ( .B(instr[4]), .A(n2872), .Y(n1627) );
  NAND21XL U2571 ( .B(n2011), .A(n213), .Y(n1128) );
  NAND21X1 U2572 ( .B(n295), .A(phase[2]), .Y(n1090) );
  AO21X1 U2573 ( .B(n2026), .C(n2025), .A(n2024), .Y(n2523) );
  NAND21XL U2574 ( .B(n2023), .A(n2022), .Y(n2025) );
  MUX2XL U2575 ( .D0(n2021), .D1(n2020), .S(instr[6]), .Y(n2026) );
  AND2X1 U2576 ( .A(n2019), .B(n2018), .Y(n2021) );
  AO21XL U2577 ( .B(temp2_comb[1]), .C(n1913), .A(n1428), .Y(n1079) );
  OAI32XL U2578 ( .A(n464), .B(n35), .C(n1810), .D(n463), .E(n1725), .Y(n2524)
         );
  AOI32XL U2579 ( .A(n324), .B(n1018), .C(n462), .D(n183), .E(n1715), .Y(n463)
         );
  AO21XL U2580 ( .B(temp2_comb[5]), .C(n1913), .A(n1912), .Y(n1794) );
  AO21XL U2581 ( .B(n1164), .C(phase[1]), .A(n1163), .Y(n1174) );
  INVX1 U2582 ( .A(n1161), .Y(n1164) );
  OAI32XL U2583 ( .A(instr[4]), .B(n1375), .C(n1166), .D(n1162), .E(n185), .Y(
        n1163) );
  AND4X1 U2584 ( .A(n1371), .B(n1672), .C(n1161), .D(n1160), .Y(n1162) );
  AOI21XL U2585 ( .B(temp2_comb[7]), .C(n1913), .A(n1689), .Y(n345) );
  AOI21XL U2586 ( .B(temp2_comb[6]), .C(n1913), .A(n1912), .Y(n346) );
  INVX1 U2587 ( .A(temp2_comb[6]), .Y(n2344) );
  INVX1 U2588 ( .A(dec_accop[12]), .Y(n1065) );
  INVX1 U2589 ( .A(dec_cop[6]), .Y(n1852) );
  INVX1 U2590 ( .A(dec_cop[5]), .Y(n1836) );
  NAND21XL U2591 ( .B(n1021), .A(ramsfraddr[7]), .Y(n2314) );
  NAND21XL U2592 ( .B(instr[7]), .A(n1731), .Y(n1636) );
  NAND21XL U2593 ( .B(n1626), .A(n2872), .Y(n1265) );
  NAND21XL U2594 ( .B(n183), .A(n1369), .Y(n1993) );
  MUX2AXL U2595 ( .D0(sp[7]), .D1(n2633), .S(n947), .Y(n948) );
  INVX1 U2596 ( .A(dec_cop[3]), .Y(n1838) );
  NAND21XL U2597 ( .B(instr[4]), .A(instr[5]), .Y(n1637) );
  GEN2XL U2598 ( .D(n1684), .E(n2034), .C(n1125), .B(n457), .A(n456), .Y(n2024) );
  NAND32XL U2599 ( .B(n2870), .C(n1895), .A(n35), .Y(n457) );
  AOI21X1 U2600 ( .B(n1383), .C(n455), .A(n454), .Y(n456) );
  AOI32XL U2601 ( .A(n2034), .B(n2872), .C(n932), .D(n1899), .E(n152), .Y(n454) );
  AND2XL U2602 ( .A(b[1]), .B(acc[0]), .Y(N14337) );
  OAI221X1 U2603 ( .A(n1375), .B(n942), .C(n2526), .D(n1349), .E(n939), .Y(
        n2619) );
  AOI32XL U2604 ( .A(n324), .B(phase[0]), .C(n1615), .D(n214), .E(n938), .Y(
        n939) );
  NAND43X1 U2605 ( .B(n1016), .C(n1987), .D(n937), .A(n935), .Y(n938) );
  AOI221XL U2606 ( .A(n2332), .B(n169), .C(n1622), .D(n932), .E(n931), .Y(n935) );
  OAI22XL U2607 ( .A(n2867), .B(n1941), .C(n419), .D(n2012), .Y(n1325) );
  GEN2XL U2608 ( .D(n2873), .E(n204), .C(n1720), .B(n1959), .A(n1647), .Y(n468) );
  OAI211XL U2609 ( .C(n1171), .D(n1170), .A(n169), .B(n1169), .Y(n1172) );
  AND2XL U2610 ( .A(n2034), .B(phase[0]), .Y(n1169) );
  INVX1 U2611 ( .A(n1165), .Y(n1171) );
  MUX2BXL U2612 ( .D0(n1325), .D1(n1168), .S(n2872), .Y(n1170) );
  AOI22AXL U2613 ( .A(n2848), .B(n2069), .D(n2070), .C(test_so), .Y(n936) );
  NOR2X1 U2614 ( .A(n2069), .B(n2848), .Y(n2070) );
  OAI21X1 U2615 ( .B(ckcon[5]), .C(n2071), .A(n2072), .Y(n2069) );
  OAI21BBX1 U2616 ( .A(n2071), .B(ckcon[5]), .C(waitcnt_1_), .Y(n2072) );
  AND2XL U2617 ( .A(b[0]), .B(acc[0]), .Y(N14336) );
  AOI22BXL U2618 ( .B(n149), .A(dpl_reg[40]), .D(n133), .C(dpl_reg[32]), .Y(
        n603) );
  MUX2BXL U2619 ( .D0(n2873), .D1(n347), .S(n183), .Y(n455) );
  OAI22XL U2620 ( .A(n2871), .B(n1265), .C(n1711), .D(n1117), .Y(n347) );
  MUX2X1 U2621 ( .D0(n485), .D1(n1630), .S(n484), .Y(n486) );
  OA21XL U2622 ( .B(n35), .C(n1655), .A(n482), .Y(n488) );
  NAND5XL U2623 ( .A(n1853), .B(n1852), .C(n1851), .D(n1850), .E(n1849), .Y(
        n1857) );
  INVX1 U2624 ( .A(dec_accop[17]), .Y(n1853) );
  INVX1 U2625 ( .A(dec_cop[7]), .Y(n1849) );
  INVX1 U2626 ( .A(ramdatao[5]), .Y(n2630) );
  AOI21XL U2627 ( .B(n2867), .C(n419), .A(n324), .Y(n348) );
  AOI33XL U2628 ( .A(n1094), .B(n2016), .C(n1157), .D(instr[7]), .E(instr[5]), 
        .F(n1622), .Y(n482) );
  AOI32XL U2629 ( .A(n1322), .B(n2872), .C(n1962), .D(n1989), .E(n1166), .Y(
        n1160) );
  AOI21XL U2630 ( .B(temp2_comb[4]), .C(n1913), .A(n1689), .Y(n349) );
  INVX1 U2631 ( .A(n2708), .Y(n2071) );
  NAND21X1 U2632 ( .B(waitcnt_0_), .A(ckcon[4]), .Y(n2708) );
  INVX1 U2633 ( .A(n1832), .Y(n1856) );
  INVX1 U2634 ( .A(dpl_reg[17]), .Y(n2774) );
  INVX1 U2635 ( .A(dpl_reg[56]), .Y(n2767) );
  INVX1 U2636 ( .A(dpl_reg[58]), .Y(n2777) );
  INVX1 U2637 ( .A(dpl_reg[48]), .Y(n2768) );
  INVX1 U2638 ( .A(dpl_reg[50]), .Y(n2778) );
  INVX1 U2639 ( .A(dpl_reg[49]), .Y(n2772) );
  INVX1 U2640 ( .A(dpl_reg[16]), .Y(n2770) );
  INVX1 U2641 ( .A(dpl_reg[18]), .Y(n2780) );
  INVX1 U2642 ( .A(dpl_reg[57]), .Y(n2771) );
  INVX1 U2643 ( .A(dpl_reg[25]), .Y(n2773) );
  INVX1 U2644 ( .A(dpl_reg[24]), .Y(n2769) );
  INVX1 U2645 ( .A(dpl_reg[26]), .Y(n2779) );
  INVX1 U2646 ( .A(dec_cop[4]), .Y(n1839) );
  INVX1 U2647 ( .A(rn_reg[83]), .Y(n769) );
  INVX1 U2648 ( .A(rn_reg[211]), .Y(n754) );
  INVX1 U2649 ( .A(rn_reg[67]), .Y(n765) );
  INVX1 U2650 ( .A(rn_reg[195]), .Y(n750) );
  INVX1 U2651 ( .A(rn_reg[91]), .Y(n761) );
  INVX1 U2652 ( .A(rn_reg[219]), .Y(n746) );
  INVX1 U2653 ( .A(rn_reg[69]), .Y(n852) );
  INVX1 U2654 ( .A(rn_reg[93]), .Y(n848) );
  INVX1 U2655 ( .A(rn_reg[197]), .Y(n837) );
  INVX1 U2656 ( .A(rn_reg[85]), .Y(n856) );
  INVX1 U2657 ( .A(rn_reg[213]), .Y(n841) );
  INVX1 U2658 ( .A(rn_reg[84]), .Y(n725) );
  INVX1 U2659 ( .A(rn_reg[212]), .Y(n710) );
  INVX1 U2660 ( .A(rn_reg[68]), .Y(n721) );
  INVX1 U2661 ( .A(rn_reg[196]), .Y(n706) );
  INVX1 U2662 ( .A(rn_reg[92]), .Y(n717) );
  INVX1 U2663 ( .A(rn_reg[220]), .Y(n702) );
  INVX1 U2664 ( .A(rn_reg[80]), .Y(n680) );
  INVX1 U2665 ( .A(rn_reg[208]), .Y(n665) );
  INVX1 U2666 ( .A(rn_reg[64]), .Y(n676) );
  INVX1 U2667 ( .A(rn_reg[192]), .Y(n661) );
  INVX1 U2668 ( .A(rn_reg[88]), .Y(n672) );
  INVX1 U2669 ( .A(rn_reg[216]), .Y(n657) );
  INVX1 U2670 ( .A(rn_reg[81]), .Y(n814) );
  INVX1 U2671 ( .A(rn_reg[209]), .Y(n799) );
  INVX1 U2672 ( .A(rn_reg[65]), .Y(n810) );
  INVX1 U2673 ( .A(rn_reg[193]), .Y(n795) );
  INVX1 U2674 ( .A(rn_reg[89]), .Y(n806) );
  INVX1 U2675 ( .A(rn_reg[217]), .Y(n791) );
  INVX1 U2676 ( .A(rn_reg[107]), .Y(n762) );
  INVX1 U2677 ( .A(rn_reg[235]), .Y(n747) );
  INVX1 U2678 ( .A(rn_reg[108]), .Y(n718) );
  INVX1 U2679 ( .A(rn_reg[236]), .Y(n703) );
  INVX1 U2680 ( .A(rn_reg[104]), .Y(n673) );
  INVX1 U2681 ( .A(rn_reg[232]), .Y(n658) );
  INVX1 U2682 ( .A(rn_reg[105]), .Y(n807) );
  INVX1 U2683 ( .A(rn_reg[233]), .Y(n792) );
  INVX1 U2684 ( .A(rn_reg[59]), .Y(n764) );
  INVX1 U2685 ( .A(rn_reg[187]), .Y(n749) );
  INVX1 U2686 ( .A(rn_reg[60]), .Y(n720) );
  INVX1 U2687 ( .A(rn_reg[188]), .Y(n705) );
  INVX1 U2688 ( .A(rn_reg[56]), .Y(n675) );
  INVX1 U2689 ( .A(rn_reg[184]), .Y(n660) );
  INVX1 U2690 ( .A(rn_reg[57]), .Y(n809) );
  INVX1 U2691 ( .A(rn_reg[185]), .Y(n794) );
  INVX1 U2692 ( .A(rn_reg[3]), .Y(n763) );
  INVX1 U2693 ( .A(rn_reg[131]), .Y(n748) );
  INVX1 U2694 ( .A(rn_reg[4]), .Y(n719) );
  INVX1 U2695 ( .A(rn_reg[132]), .Y(n704) );
  INVX1 U2696 ( .A(rn_reg[0]), .Y(n674) );
  INVX1 U2697 ( .A(rn_reg[128]), .Y(n659) );
  INVX1 U2698 ( .A(rn_reg[1]), .Y(n808) );
  INVX1 U2699 ( .A(rn_reg[129]), .Y(n793) );
  OA2222XL U2700 ( .A(instr[5]), .B(n1333), .C(n1384), .D(n1610), .E(n1332), 
        .F(n1960), .G(n1331), .H(n1386), .Y(n1338) );
  INVX1 U2701 ( .A(n1325), .Y(n1332) );
  AOI32XL U2702 ( .A(n214), .B(n34), .C(n1261), .D(n1991), .E(n296), .Y(n1262)
         );
  INVX1 U2703 ( .A(n1259), .Y(n1261) );
  NAND21XL U2704 ( .B(instr[5]), .A(instr[7]), .Y(n1167) );
  NAND21XL U2705 ( .B(n2867), .A(n2017), .Y(n1386) );
  NAND21XL U2706 ( .B(n204), .A(n1124), .Y(n487) );
  NAND43X1 U2707 ( .B(n1341), .C(n1340), .D(n1339), .A(n1338), .Y(n1342) );
  INVX1 U2708 ( .A(n1314), .Y(n1340) );
  NAND21XL U2709 ( .B(dec_accop[9]), .A(n1763), .Y(n1866) );
  NAND2X1 U2710 ( .A(n350), .B(n1923), .Y(n1901) );
  NAND4XL U2711 ( .A(n1896), .B(phase[0]), .C(n1944), .D(n1895), .Y(n350) );
  GEN2XL U2712 ( .D(n1324), .E(n1323), .C(n1322), .B(n1321), .A(n1315), .Y(
        n1339) );
  AND4XL U2713 ( .A(n1324), .B(n2867), .C(n1944), .D(n1626), .Y(n1315) );
  NAND6XL U2714 ( .A(n1379), .B(n2440), .C(n2439), .D(n1378), .E(n2035), .F(
        n1377), .Y(n2617) );
  OA2222XL U2715 ( .A(n1376), .B(n186), .C(n1375), .D(n1374), .E(n1373), .F(
        n1372), .G(n1371), .H(n167), .Y(n1377) );
  OA21XL U2716 ( .B(n2870), .C(n1370), .A(n2011), .Y(n1373) );
  AOI22BXL U2717 ( .B(n2808), .A(dpl_reg[8]), .D(n2807), .C(dpl_reg[0]), .Y(
        n605) );
  AOI22BXL U2718 ( .B(n370), .A(dpl_reg[10]), .D(n372), .C(dpl_reg[2]), .Y(
        n597) );
  AOI22BXL U2719 ( .B(n149), .A(dph_reg[40]), .D(n133), .C(dph_reg[32]), .Y(
        n635) );
  AOI22BXL U2720 ( .B(n149), .A(dpl_reg[42]), .D(n133), .C(dpl_reg[34]), .Y(
        n595) );
  AOI22BXL U2721 ( .B(n149), .A(dpc_tab[30]), .D(n133), .C(dpc_tab[24]), .Y(
        n1353) );
  AOI22BXL U2722 ( .B(n149), .A(dpc_tab[32]), .D(n133), .C(dpc_tab[26]), .Y(
        n1362) );
  NAND21XL U2723 ( .B(n2871), .A(n34), .Y(n1383) );
  INVX1 U2724 ( .A(n1145), .Y(n1151) );
  GEN2XL U2725 ( .D(n1144), .E(n1143), .C(n2526), .B(n1142), .A(n1906), .Y(
        n1145) );
  AND3XL U2726 ( .A(n1131), .B(n1951), .C(n1130), .Y(n1144) );
  AOI31XL U2727 ( .A(n1135), .B(instr[2]), .C(n1781), .D(n1134), .Y(n1143) );
  NAND2XL U2728 ( .A(n351), .B(n2035), .Y(n2036) );
  NAND4XL U2729 ( .A(n324), .B(n2034), .C(n2033), .D(n296), .Y(n351) );
  INVXL U2730 ( .A(acc[1]), .Y(n1964) );
  INVX1 U2731 ( .A(ramdatao[7]), .Y(n2633) );
  INVX1 U2732 ( .A(ramdatao[6]), .Y(n2811) );
  INVX1 U2733 ( .A(n1897), .Y(n1898) );
  INVXL U2734 ( .A(ramsfraddr[4]), .Y(n2567) );
  AOI221XL U2735 ( .A(n1654), .B(n1369), .C(n1360), .D(instr[6]), .E(n1359), 
        .Y(n1376) );
  OAI31XL U2736 ( .A(n1358), .B(n1655), .C(n1382), .D(n1357), .Y(n1359) );
  AOI32XL U2737 ( .A(phase[3]), .B(n1141), .C(n152), .D(n214), .E(n1140), .Y(
        n1142) );
  NAND21X1 U2738 ( .B(n1986), .A(n1139), .Y(n1140) );
  INVX1 U2739 ( .A(n1138), .Y(n1139) );
  INVXL U2740 ( .A(temp2_comb[2]), .Y(n2257) );
  OAI211XL U2741 ( .C(n204), .D(n183), .A(n348), .B(n2012), .Y(n460) );
  INVX1 U2742 ( .A(n1147), .Y(n1129) );
  INVXL U2743 ( .A(temp2_comb[3]), .Y(n2160) );
  INVX1 U2744 ( .A(n445), .Y(n1282) );
  OAI211XL U2745 ( .C(instr[1]), .D(n1112), .A(n1131), .B(n1956), .Y(n445) );
  INVX1 U2746 ( .A(waitcnt_1_), .Y(n2707) );
  INVX1 U2747 ( .A(n2073), .Y(n2700) );
  OAI221X1 U2748 ( .A(waitcnt_1_), .B(n2815), .C(test_so), .D(n2814), .E(n2847), .Y(n2073) );
  OAI211X1 U2749 ( .C(ckcon[1]), .D(n2707), .A(ckcon[0]), .B(n2706), .Y(n2847)
         );
  INVX1 U2750 ( .A(dpl_reg[59]), .Y(n2781) );
  INVX1 U2751 ( .A(dpl_reg[51]), .Y(n2782) );
  INVX1 U2752 ( .A(dpl_reg[20]), .Y(n2788) );
  INVX1 U2753 ( .A(dpl_reg[19]), .Y(n2784) );
  INVX1 U2754 ( .A(dpl_reg[27]), .Y(n2783) );
  INVX1 U2755 ( .A(rn_reg[221]), .Y(n833) );
  INVX1 U2756 ( .A(rn_reg[71]), .Y(n984) );
  INVX1 U2757 ( .A(rn_reg[95]), .Y(n976) );
  INVX1 U2758 ( .A(rn_reg[199]), .Y(n960) );
  INVX1 U2759 ( .A(rn_reg[223]), .Y(n955) );
  INVX1 U2760 ( .A(rn_reg[87]), .Y(n992) );
  INVX1 U2761 ( .A(rn_reg[215]), .Y(n964) );
  INVX1 U2762 ( .A(rn_reg[82]), .Y(n638) );
  INVX1 U2763 ( .A(rn_reg[210]), .Y(n557) );
  INVX1 U2764 ( .A(rn_reg[66]), .Y(n574) );
  INVX1 U2765 ( .A(rn_reg[194]), .Y(n548) );
  INVX1 U2766 ( .A(rn_reg[90]), .Y(n570) );
  INVX1 U2767 ( .A(rn_reg[218]), .Y(n540) );
  INVX1 U2768 ( .A(rn_reg[101]), .Y(n857) );
  INVX1 U2769 ( .A(rn_reg[229]), .Y(n842) );
  INVX1 U2770 ( .A(rn_reg[103]), .Y(n994) );
  INVX1 U2771 ( .A(rn_reg[231]), .Y(n965) );
  INVX1 U2772 ( .A(rn_reg[106]), .Y(n571) );
  INVX1 U2773 ( .A(rn_reg[234]), .Y(n541) );
  INVX1 U2774 ( .A(rn_reg[53]), .Y(n859) );
  INVX1 U2775 ( .A(rn_reg[181]), .Y(n844) );
  INVX1 U2776 ( .A(rn_reg[55]), .Y(n998) );
  INVX1 U2777 ( .A(rn_reg[183]), .Y(n967) );
  INVX1 U2778 ( .A(rn_reg[58]), .Y(n573) );
  INVX1 U2779 ( .A(rn_reg[186]), .Y(n543) );
  INVX1 U2780 ( .A(rn_reg[117]), .Y(n858) );
  INVX1 U2781 ( .A(rn_reg[245]), .Y(n843) );
  INVX1 U2782 ( .A(rn_reg[119]), .Y(n996) );
  INVX1 U2783 ( .A(rn_reg[247]), .Y(n966) );
  INVX1 U2784 ( .A(rn_reg[2]), .Y(n572) );
  INVX1 U2785 ( .A(rn_reg[130]), .Y(n542) );
  NAND21XL U2786 ( .B(n183), .A(n204), .Y(n1116) );
  OR2X1 U2787 ( .A(n2864), .B(mempsrd), .Y(n2583) );
  NAND43X1 U2788 ( .B(instr[3]), .C(n2028), .D(instr[1]), .A(n1123), .Y(n1149)
         );
  MUX2BXL U2789 ( .D0(n1122), .D1(n1121), .S(instr[0]), .Y(n1123) );
  AND3XL U2790 ( .A(n1617), .B(n1721), .C(n1973), .Y(n1122) );
  AND3X1 U2791 ( .A(n1722), .B(n1120), .C(n1119), .Y(n1121) );
  INVX1 U2792 ( .A(n1954), .Y(n1974) );
  OAI31XL U2793 ( .A(instr[7]), .B(n1953), .C(n1952), .D(n1951), .Y(n1954) );
  AOI22BXL U2794 ( .B(n369), .A(dph_reg[8]), .D(n371), .C(dph_reg[0]), .Y(n637) );
  AND2XL U2795 ( .A(b[0]), .B(acc[1]), .Y(N14344) );
  AOI22BXL U2796 ( .B(n149), .A(dpl_reg[41]), .D(n133), .C(dpl_reg[33]), .Y(
        n599) );
  AOI22BXL U2797 ( .B(n149), .A(dph_reg[41]), .D(n133), .C(dph_reg[33]), .Y(
        n631) );
  AOI22BXL U2798 ( .B(n149), .A(dph_reg[42]), .D(n133), .C(dph_reg[34]), .Y(
        n627) );
  AOI22BXL U2799 ( .B(n149), .A(dpc_tab[31]), .D(n133), .C(dpc_tab[25]), .Y(
        n1366) );
  MUX2AXL U2800 ( .D0(n352), .D1(n2017), .S(instr[1]), .Y(n2018) );
  NAND2XL U2801 ( .A(interrupt), .B(n418), .Y(n352) );
  AO21XL U2802 ( .B(n2016), .C(instr[0]), .A(n2015), .Y(n2019) );
  NOR32XL U2803 ( .B(n152), .C(n1369), .A(n449), .Y(n2023) );
  XNOR2XL U2804 ( .A(instr[0]), .B(n183), .Y(n448) );
  INVXL U2805 ( .A(acc[0]), .Y(n1965) );
  INVX1 U2806 ( .A(n1111), .Y(n1279) );
  NAND21XL U2807 ( .B(n187), .A(instr[1]), .Y(n1111) );
  INVXL U2808 ( .A(acc[4]), .Y(n2383) );
  AOI32XL U2809 ( .A(n2871), .B(n2867), .C(n1962), .D(n1118), .E(n2017), .Y(
        n1119) );
  INVX1 U2810 ( .A(n1167), .Y(n1118) );
  INVXL U2811 ( .A(acc[3]), .Y(n2116) );
  INVXL U2812 ( .A(acc[5]), .Y(n2294) );
  AND2XL U2813 ( .A(acc[0]), .B(n1416), .Y(n1417) );
  INVXL U2814 ( .A(c), .Y(n1831) );
  INVX1 U2815 ( .A(temp2_comb[7]), .Y(n2438) );
  INVX1 U2816 ( .A(waitcnt_0_), .Y(n2706) );
  INVX1 U2817 ( .A(ckcon[6]), .Y(n2848) );
  INVX1 U2818 ( .A(ckcon[1]), .Y(n2815) );
  INVX1 U2819 ( .A(ckcon[2]), .Y(n2814) );
  INVX1 U2820 ( .A(dpl_reg[60]), .Y(n2785) );
  INVX1 U2821 ( .A(dpl_reg[61]), .Y(n2789) );
  INVX1 U2822 ( .A(dpl_reg[62]), .Y(n2793) );
  INVX1 U2823 ( .A(dph_reg[56]), .Y(n2731) );
  INVX1 U2824 ( .A(dpl_reg[52]), .Y(n2786) );
  INVX1 U2825 ( .A(dpl_reg[53]), .Y(n2790) );
  INVX1 U2826 ( .A(dpl_reg[54]), .Y(n2794) );
  INVX1 U2827 ( .A(dpl_reg[21]), .Y(n2792) );
  INVX1 U2828 ( .A(dph_reg[24]), .Y(n2734) );
  INVX1 U2829 ( .A(dpl_reg[22]), .Y(n2796) );
  INVX1 U2830 ( .A(dpl_reg[28]), .Y(n2787) );
  INVX1 U2831 ( .A(dpl_reg[29]), .Y(n2791) );
  INVX1 U2832 ( .A(dph_reg[16]), .Y(n2733) );
  INVX1 U2833 ( .A(dpl_reg[30]), .Y(n2795) );
  INVX1 U2834 ( .A(rn_reg[70]), .Y(n905) );
  INVX1 U2835 ( .A(rn_reg[94]), .Y(n901) );
  INVX1 U2836 ( .A(rn_reg[198]), .Y(n890) );
  INVX1 U2837 ( .A(rn_reg[222]), .Y(n886) );
  INVX1 U2838 ( .A(rn_reg[86]), .Y(n909) );
  INVX1 U2839 ( .A(rn_reg[214]), .Y(n894) );
  INVX1 U2840 ( .A(dpc_tab[36]), .Y(n2722) );
  INVX1 U2841 ( .A(dpc_tab[6]), .Y(n2726) );
  INVX1 U2842 ( .A(dpc_tab[12]), .Y(n2724) );
  INVX1 U2843 ( .A(dpc_tab[38]), .Y(n2716) );
  INVX1 U2844 ( .A(dpc_tab[8]), .Y(n2720) );
  INVX1 U2845 ( .A(dpc_tab[14]), .Y(n2718) );
  INVX1 U2846 ( .A(dpc_tab[42]), .Y(n2721) );
  INVX1 U2847 ( .A(dpc_tab[0]), .Y(n2725) );
  INVX1 U2848 ( .A(dpc_tab[18]), .Y(n2723) );
  INVX1 U2849 ( .A(dpc_tab[44]), .Y(n2715) );
  INVX1 U2850 ( .A(dpc_tab[2]), .Y(n2719) );
  INVX1 U2851 ( .A(dpc_tab[20]), .Y(n2717) );
  INVX1 U2852 ( .A(rn_reg[102]), .Y(n910) );
  INVX1 U2853 ( .A(rn_reg[230]), .Y(n895) );
  INVX1 U2854 ( .A(rn_reg[54]), .Y(n912) );
  INVX1 U2855 ( .A(rn_reg[182]), .Y(n897) );
  INVX1 U2856 ( .A(rn_reg[118]), .Y(n911) );
  INVX1 U2857 ( .A(rn_reg[246]), .Y(n896) );
  MUX2AXL U2858 ( .D0(pmw), .D1(n2628), .S(n1815), .Y(n2648) );
  OR2X1 U2859 ( .A(memwr), .B(memrd), .Y(n2703) );
  MUX2X1 U2860 ( .D0(n1967), .D1(n1966), .S(N345), .Y(n1968) );
  OA2222XL U2861 ( .A(n2668), .B(n1965), .C(n2124), .D(n2116), .E(n1964), .F(
        n2665), .G(n2263), .H(n2264), .Y(n1967) );
  OA2222XL U2862 ( .A(n2383), .B(n2668), .C(n2411), .D(n2124), .E(n2665), .F(
        n2294), .G(n2264), .H(n2329), .Y(n1966) );
  AO21XL U2863 ( .B(n2005), .C(n2869), .A(israccess), .Y(n2507) );
  INVX1 U2864 ( .A(n436), .Y(n2701) );
  NAND21X1 U2865 ( .B(ckcon[2]), .A(test_so), .Y(n436) );
  INVX1 U2866 ( .A(dph_reg[57]), .Y(n2735) );
  INVX1 U2867 ( .A(dph_reg[58]), .Y(n2741) );
  INVX1 U2868 ( .A(dph_reg[48]), .Y(n2732) );
  INVX1 U2869 ( .A(dph_reg[49]), .Y(n2736) );
  INVX1 U2870 ( .A(dph_reg[50]), .Y(n2742) );
  INVX1 U2871 ( .A(dph_reg[17]), .Y(n2738) );
  INVX1 U2872 ( .A(dph_reg[18]), .Y(n2744) );
  INVX1 U2873 ( .A(dph_reg[25]), .Y(n2737) );
  INVX1 U2874 ( .A(dph_reg[26]), .Y(n2743) );
  INVX1 U2875 ( .A(dpl_reg[1]), .Y(n2775) );
  INVX1 U2876 ( .A(dph_reg[1]), .Y(n2739) );
  INVX1 U2877 ( .A(dph_reg[2]), .Y(n2745) );
  INVX1 U2878 ( .A(dpl_reg[9]), .Y(n2776) );
  INVX1 U2879 ( .A(dph_reg[9]), .Y(n2740) );
  INVX1 U2880 ( .A(dph_reg[10]), .Y(n2746) );
  INVX1 U2881 ( .A(dpc_tab[37]), .Y(n2710) );
  INVX1 U2882 ( .A(dpc_tab[7]), .Y(n2714) );
  INVX1 U2883 ( .A(dpc_tab[13]), .Y(n2712) );
  INVX1 U2884 ( .A(dpc_tab[43]), .Y(n2709) );
  INVX1 U2885 ( .A(dpc_tab[1]), .Y(n2713) );
  INVX1 U2886 ( .A(dpc_tab[19]), .Y(n2711) );
  INVX1 U2887 ( .A(memaddr[9]), .Y(n2850) );
  OR2X1 U2888 ( .A(state[2]), .B(state[1]), .Y(n2219) );
  INVX1 U2889 ( .A(n442), .Y(n1681) );
  NAND32XL U2890 ( .B(phase[1]), .C(phase[0]), .A(n2526), .Y(n442) );
  INVX1 U2891 ( .A(n443), .Y(n2535) );
  NAND21X1 U2892 ( .B(state[0]), .A(n2809), .Y(n443) );
  INVX1 U2893 ( .A(phase[3]), .Y(n2528) );
  MUX2XL U2894 ( .D0(pc_o[11]), .D1(n2692), .S(n420), .Y(memaddr_comb[11]) );
  NAND21X1 U2895 ( .B(n1213), .A(n1212), .Y(n2512) );
  AO21XL U2896 ( .B(n1211), .C(n1229), .A(n2667), .Y(n1212) );
  MUX2XL U2897 ( .D0(stop), .D1(n2622), .S(n2132), .Y(n1213) );
  AO2222XL U2898 ( .A(n264), .B(ramdatao[3]), .C(n2176), .D(n2486), .E(p2[3]), 
        .F(n265), .G(n2485), .H(pc_o[11]), .Y(n2692) );
  AO2222XL U2899 ( .A(n2172), .B(n48), .C(pc_i[11]), .D(n2484), .E(alu_out[11]), .F(n131), .G(n2480), .H(temp[3]), .Y(n2176) );
  MUX2XL U2900 ( .D0(pc_o[12]), .D1(n2693), .S(n420), .Y(memaddr_comb[12]) );
  AO2222XL U2901 ( .A(n264), .B(ramdatao[4]), .C(n2179), .D(n2486), .E(p2[4]), 
        .F(n265), .G(n2485), .H(pc_o[12]), .Y(n2693) );
  AO2222XL U2902 ( .A(pc_i[12]), .B(n2484), .C(n2178), .D(n48), .E(alu_out[12]), .F(n131), .G(n2480), .H(temp[4]), .Y(n2179) );
  INVX1 U2903 ( .A(idle_r), .Y(n2515) );
  INVX1 U2904 ( .A(stop_r), .Y(n2516) );
  INVX1 U2905 ( .A(idle), .Y(n2502) );
  MUX2XL U2906 ( .D0(ramsfraddr[2]), .D1(n2638), .S(n423), .Y(
        ramsfraddr_comb[2]) );
  MUX2XL U2907 ( .D0(pc_o[13]), .D1(n2694), .S(n420), .Y(memaddr_comb[13]) );
  MUX2XL U2908 ( .D0(pc_o[14]), .D1(n2695), .S(n420), .Y(memaddr_comb[14]) );
  NAND21X1 U2909 ( .B(n1399), .A(n1398), .Y(n2543) );
  MUX2X1 U2910 ( .D0(cs_run), .D1(n2535), .S(codefetch_s), .Y(n1399) );
  AO21XL U2911 ( .B(n2542), .C(n2541), .A(n2540), .Y(n2654) );
  GEN3XL U2912 ( .F(n2539), .G(n2651), .E(n2538), .D(n2549), .C(n2537), .B(
        cs_run), .A(n2536), .Y(n2540) );
  INVX1 U2913 ( .A(n2548), .Y(n2539) );
  AND4XL U2914 ( .A(n2535), .B(n2534), .C(n2533), .D(n2532), .Y(n2536) );
  NAND4X1 U2915 ( .A(n590), .B(n591), .C(n592), .D(n593), .Y(dpl[3]) );
  NAND4X1 U2916 ( .A(n622), .B(n623), .C(n624), .D(n625), .Y(dph[3]) );
  OA22X1 U2917 ( .A(n368), .B(n2784), .C(n2804), .D(n2783), .Y(n592) );
  AO2222XL U2918 ( .A(n264), .B(ramdatao[6]), .C(n2487), .D(n2486), .E(p2[6]), 
        .F(n265), .G(pc_o[14]), .H(n2485), .Y(n2695) );
  AO2222XL U2919 ( .A(pc_i[14]), .B(n2484), .C(n2483), .D(n48), .E(alu_out[14]), .F(n131), .G(n2480), .H(temp[6]), .Y(n2487) );
  AO2222XL U2920 ( .A(n264), .B(ramdatao[5]), .C(n2284), .D(n2486), .E(p2[5]), 
        .F(n265), .G(n2485), .H(pc_o[13]), .Y(n2694) );
  AO2222XL U2921 ( .A(pc_i[13]), .B(n2484), .C(n2283), .D(n48), .E(alu_out[13]), .F(n131), .G(n2480), .H(temp[5]), .Y(n2284) );
  MUX2XL U2922 ( .D0(mempsrd), .D1(n2654), .S(n420), .Y(mempsrd_comb) );
  AOI21X1 U2923 ( .B(n2531), .C(n2530), .A(n2810), .Y(n2537) );
  OA222X1 U2924 ( .A(n2529), .B(n2528), .C(n2527), .D(n2526), .E(n2525), .F(
        n186), .Y(n2530) );
  AOI211XL U2925 ( .C(n214), .D(n2523), .A(codefetch_s), .B(n2522), .Y(n2531)
         );
  INVX1 U2926 ( .A(n2524), .Y(n2529) );
  MUX2X1 U2927 ( .D0(pc_o[15]), .D1(n2696), .S(n422), .Y(memaddr_comb[15]) );
  AO2222XL U2928 ( .A(n264), .B(ramdatao[7]), .C(n2381), .D(n2486), .E(p2[7]), 
        .F(n265), .G(pc_o[15]), .H(n2485), .Y(n2696) );
  AO2222XL U2929 ( .A(pc_i[15]), .B(n2484), .C(n2380), .D(n2482), .E(
        alu_out[15]), .F(n131), .G(n2480), .H(temp[7]), .Y(n2381) );
  NAND21X1 U2930 ( .B(n2235), .A(n2234), .Y(n2689) );
  OA2222XL U2931 ( .A(n2277), .B(n2244), .C(n2233), .D(n2243), .E(n36), .F(
        n2236), .G(n2241), .H(n2232), .Y(n2234) );
  AO2222XL U2932 ( .A(n2239), .B(pc_o[9]), .C(n2238), .D(pc_i[9]), .E(
        alu_out[9]), .F(n131), .G(n2237), .H(instr[6]), .Y(n2235) );
  NAND21X1 U2933 ( .B(n2226), .A(n2225), .Y(n2688) );
  OA2222XL U2934 ( .A(n2224), .B(n2243), .C(n47), .D(n2223), .E(n2241), .F(
        n2222), .G(n2278), .H(n2244), .Y(n2225) );
  AO2222XL U2935 ( .A(n2239), .B(pc_o[8]), .C(pc_i[8]), .D(n2238), .E(
        alu_out[8]), .F(n131), .G(n2237), .H(instr[5]), .Y(n2226) );
  MUX2X1 U2936 ( .D0(memaddr[7]), .D1(n1927), .S(n1934), .Y(N12848) );
  AO21XL U2937 ( .B(n1901), .C(n2372), .A(n2826), .Y(N12831) );
  MUX2X1 U2938 ( .D0(pc_o[8]), .D1(n1926), .S(n1934), .Y(N12849) );
  MUX2X1 U2939 ( .D0(pc_o[9]), .D1(n1925), .S(n1934), .Y(N12850) );
  MUX2X1 U2940 ( .D0(memaddr[11]), .D1(n2172), .S(n172), .Y(N12852) );
  MUX2X1 U2941 ( .D0(pc_o[13]), .D1(n2283), .S(n172), .Y(N12854) );
  MUX2X1 U2942 ( .D0(memaddr[10]), .D1(n1924), .S(n172), .Y(N12851) );
  MUX2X1 U2943 ( .D0(pc_o[12]), .D1(n2178), .S(n172), .Y(N12853) );
  MUX2X1 U2944 ( .D0(memaddr[14]), .D1(n2483), .S(n172), .Y(N12855) );
  MUX2XL U2945 ( .D0(ramsfraddr[0]), .D1(n64), .S(n423), .Y(ramsfraddr_comb[0]) );
  NAND21X1 U2946 ( .B(n2246), .A(n2245), .Y(n2691) );
  OA2222XL U2947 ( .A(n2625), .B(n2244), .C(n2262), .D(n2243), .E(n47), .F(
        n2242), .G(n2241), .H(n2240), .Y(n2245) );
  AO2222XL U2948 ( .A(pc_o[10]), .B(n2239), .C(pc_i[10]), .D(n2238), .E(
        alu_out[10]), .F(n131), .G(n2237), .H(n183), .Y(n2246) );
  NAND4X1 U2949 ( .A(n618), .B(n619), .C(n620), .D(n621), .Y(dph[4]) );
  NAND4X1 U2950 ( .A(n586), .B(n587), .C(n588), .D(n589), .Y(dpl[4]) );
  OA22X1 U2951 ( .A(n367), .B(n2754), .C(n366), .D(n2753), .Y(n620) );
  MUX2XL U2952 ( .D0(ramdatao[3]), .D1(n2627), .S(waitstaten), .Y(
        ramdatao_comb[3]) );
  MUX2XL U2953 ( .D0(n2131), .D1(n2130), .S(n2624), .Y(n2627) );
  NAND32X1 U2954 ( .B(n2129), .C(n2128), .A(n2127), .Y(n2131) );
  OAI22XL U2955 ( .A(n2444), .B(n2153), .C(n2431), .D(n2102), .Y(n2129) );
  AO2222XL U2956 ( .A(n2105), .B(pc_o[11]), .C(pc_i[11]), .D(n2104), .E(n2591), 
        .F(pc_o[3]), .G(temp2_comb[3]), .H(n2103), .Y(n2128) );
  OA2222XL U2957 ( .A(dpl_reg[15]), .B(n1584), .C(dpl_reg[7]), .D(n1583), .E(
        dpl_reg[47]), .F(n1582), .G(dpl_reg[39]), .H(n1581), .Y(n1518) );
  OA2222XL U2958 ( .A(dph_reg[8]), .B(n1584), .C(dph_reg[0]), .D(n1583), .E(
        dph_reg[40]), .F(n1582), .G(dph_reg[32]), .H(n1581), .Y(n1585) );
  MUX2XL U2959 ( .D0(n1247), .D1(n2098), .S(n2624), .Y(n2621) );
  NAND43X1 U2960 ( .B(n1240), .C(n1237), .D(n1236), .A(n1235), .Y(n1247) );
  OAI22X1 U2961 ( .A(n51), .B(n2445), .C(n2442), .D(n1877), .Y(n1236) );
  AO21XL U2962 ( .B(n2865), .C(n1224), .A(n1223), .Y(n1240) );
  NAND4X1 U2963 ( .A(n614), .B(n615), .C(n616), .D(n617), .Y(dph[5]) );
  NAND4X1 U2964 ( .A(n582), .B(n583), .C(n584), .D(n585), .Y(dpl[5]) );
  OA22X1 U2965 ( .A(n368), .B(n2758), .C(n2804), .D(n2757), .Y(n616) );
  MUX2XL U2966 ( .D0(ramdatao[0]), .D1(n2621), .S(n423), .Y(ramdatao_comb[0])
         );
  NAND4X1 U2967 ( .A(n578), .B(n579), .C(n580), .D(n581), .Y(dpl[6]) );
  NAND4X1 U2968 ( .A(n610), .B(n611), .C(n612), .D(n613), .Y(dph[6]) );
  OA22X1 U2969 ( .A(n368), .B(n2796), .C(n2804), .D(n2795), .Y(n580) );
  MUX2X1 U2970 ( .D0(n1555), .D1(ramdatao[7]), .S(n1587), .Y(n2139) );
  NAND21X1 U2971 ( .B(n1554), .A(n1553), .Y(n1555) );
  OA2222XL U2972 ( .A(dph_reg[9]), .B(n162), .C(dph_reg[1]), .D(n145), .E(
        dph_reg[41]), .F(n178), .G(dph_reg[33]), .H(n201), .Y(n1573) );
  NAND21X1 U2973 ( .B(pdmode), .A(n2512), .Y(n2510) );
  MUX2XL U2974 ( .D0(ramdatao[1]), .D1(n2622), .S(n423), .Y(ramdatao_comb[1])
         );
  AO222XL U2975 ( .A(n30), .B(pc_o[2]), .C(n28), .D(n2682), .E(pc_ini[2]), .F(
        n426), .Y(N482) );
  AO222XL U2976 ( .A(n30), .B(n2865), .C(n28), .D(n2680), .E(pc_ini[0]), .F(
        n426), .Y(N480) );
  AO222XL U2977 ( .A(n31), .B(memaddr[3]), .C(n29), .D(n2683), .E(pc_ini[3]), 
        .F(n426), .Y(N483) );
  AO222XL U2978 ( .A(n31), .B(pc_o[1]), .C(n29), .D(n2681), .E(pc_ini[1]), .F(
        n426), .Y(N481) );
  AO222X1 U2979 ( .A(n31), .B(pc_o[10]), .C(n29), .D(n2691), .E(pc_ini[10]), 
        .F(n426), .Y(N490) );
  AO222X1 U2980 ( .A(n30), .B(pc_o[9]), .C(n28), .D(n2689), .E(pc_ini[9]), .F(
        n426), .Y(N489) );
  AO222X1 U2981 ( .A(n31), .B(pc_o[8]), .C(n29), .D(n2688), .E(pc_ini[8]), .F(
        n426), .Y(N488) );
  AO222X1 U2982 ( .A(n30), .B(pc_o[7]), .C(n28), .D(n2687), .E(pc_ini[7]), .F(
        n426), .Y(N487) );
  AO222XL U2983 ( .A(n30), .B(pc_o[6]), .C(n28), .D(n2686), .E(pc_ini[6]), .F(
        n425), .Y(N486) );
  AO222XL U2984 ( .A(n31), .B(pc_o[5]), .C(n29), .D(n2685), .E(pc_ini[5]), .F(
        n426), .Y(N485) );
  AO222XL U2985 ( .A(n30), .B(memaddr[4]), .C(n28), .D(n2684), .E(pc_ini[4]), 
        .F(n426), .Y(N484) );
  NAND4X1 U2986 ( .A(n566), .B(n567), .C(n568), .D(n569), .Y(dpl[7]) );
  NAND4X1 U2987 ( .A(n606), .B(n607), .C(n608), .D(n609), .Y(dph[7]) );
  OA22X1 U2988 ( .A(n2806), .B(n2805), .C(n365), .D(n2803), .Y(n568) );
  MUX2X1 U2989 ( .D0(pc_o[15]), .D1(n2380), .S(n172), .Y(N12856) );
  MUX2X1 U2990 ( .D0(n2520), .D1(pdmode), .S(n2519), .Y(n2446) );
  AND2X1 U2991 ( .A(n2513), .B(n434), .Y(n2520) );
  AO21X1 U2992 ( .B(n2516), .C(n2515), .A(n2542), .Y(n2518) );
  AO21X1 U2993 ( .B(n2221), .C(n2512), .A(n2220), .Y(n1878) );
  INVX1 U2994 ( .A(n2503), .Y(n2221) );
  GEN2XL U2995 ( .D(n2810), .E(n2534), .C(n2219), .B(newinstrlock), .A(n432), 
        .Y(n2220) );
  AO22X1 U2996 ( .A(n379), .B(n2696), .C(pc_ini[15]), .D(n427), .Y(N495) );
  AO22X1 U2997 ( .A(n379), .B(n2695), .C(pc_ini[14]), .D(n427), .Y(N494) );
  AO22X1 U2998 ( .A(n379), .B(n2694), .C(pc_ini[13]), .D(n427), .Y(N493) );
  AO22X1 U2999 ( .A(n379), .B(n2693), .C(pc_ini[12]), .D(n427), .Y(N492) );
  AO22X1 U3000 ( .A(n379), .B(n2692), .C(pc_ini[11]), .D(n427), .Y(N491) );
  OA2222XL U3001 ( .A(dph_reg[10]), .B(n162), .C(dph_reg[2]), .D(n145), .E(
        dph_reg[42]), .F(n178), .G(dph_reg[34]), .H(n201), .Y(n1273) );
  AO21X1 U3002 ( .B(n423), .C(n2133), .A(n432), .Y(N520) );
  MUX2XL U3003 ( .D0(p2sel), .D1(n2627), .S(n2132), .Y(n2133) );
  AND2XL U3004 ( .A(sfroe_r), .B(n422), .Y(sfroe) );
  OA2222XL U3005 ( .A(dph_reg[11]), .B(n162), .C(dph_reg[3]), .D(n145), .E(
        dph_reg[43]), .F(n178), .G(dph_reg[35]), .H(n201), .Y(n1569) );
  OR3XL U3006 ( .A(n2170), .B(n2168), .C(p2sel), .Y(n2173) );
  OA2222XL U3007 ( .A(dph_reg[12]), .B(n162), .C(dph_reg[4]), .D(n145), .E(
        dph_reg[44]), .F(n178), .G(dph_reg[36]), .H(n201), .Y(n1392) );
  OA2222XL U3008 ( .A(dph_reg[13]), .B(n162), .C(dph_reg[5]), .D(n145), .E(
        dph_reg[45]), .F(n178), .G(dph_reg[37]), .H(n201), .Y(n1565) );
  NAND21X1 U3009 ( .B(n1508), .A(n1507), .Y(dpc[3]) );
  OA2222XL U3010 ( .A(n2804), .B(n1506), .C(n2806), .D(n1505), .E(n370), .F(
        n1504), .G(n2807), .H(n1503), .Y(n1507) );
  AO2222XL U3011 ( .A(dpc_tab[27]), .B(n132), .C(dpc_tab[33]), .D(n148), .E(
        dpc_tab[39]), .F(n180), .G(dpc_tab[45]), .H(n164), .Y(n1508) );
  INVX1 U3012 ( .A(dpc_tab[21]), .Y(n1506) );
  AOI22BXL U3013 ( .B(n369), .A(dph_reg[11]), .D(n371), .C(dph_reg[3]), .Y(
        n625) );
  AOI22BXL U3014 ( .B(n2808), .A(dpl_reg[11]), .D(n2807), .C(dpl_reg[3]), .Y(
        n593) );
  AOI22BXL U3015 ( .B(n149), .A(dph_reg[43]), .D(n133), .C(dph_reg[35]), .Y(
        n623) );
  AOI22BXL U3016 ( .B(n2802), .A(dpl_reg[43]), .D(n134), .C(dpl_reg[35]), .Y(
        n591) );
  OR2XL U3017 ( .A(ramsfraddr[2]), .B(n1275), .Y(n2593) );
  INVX1 U3018 ( .A(dpl_reg[63]), .Y(n2797) );
  INVX1 U3019 ( .A(dpl_reg[55]), .Y(n2799) );
  INVX1 U3020 ( .A(dpl_reg[23]), .Y(n2805) );
  INVX1 U3021 ( .A(dpl_reg[31]), .Y(n2803) );
  OA2222XL U3022 ( .A(dph_reg[14]), .B(n162), .C(dph_reg[6]), .D(n145), .E(
        dph_reg[46]), .F(n178), .G(dph_reg[38]), .H(n201), .Y(n1561) );
  MUX2XL U3023 ( .D0(ramsfraddr[5]), .D1(n2641), .S(n423), .Y(
        ramsfraddr_comb[5]) );
  MUX2XL U3024 ( .D0(ramsfraddr[3]), .D1(n2639), .S(waitstaten), .Y(
        ramsfraddr_comb[3]) );
  INVX1 U3025 ( .A(dph_reg[59]), .Y(n2747) );
  INVX1 U3026 ( .A(dph_reg[51]), .Y(n2748) );
  INVX1 U3027 ( .A(dph_reg[19]), .Y(n2750) );
  INVX1 U3028 ( .A(dph_reg[27]), .Y(n2749) );
  MUX2XL U3029 ( .D0(ramsfraddr[4]), .D1(n2640), .S(n423), .Y(
        ramsfraddr_comb[4]) );
  MUX2XL U3030 ( .D0(ramsfraddr[7]), .D1(n2644), .S(n423), .Y(
        ramsfraddr_comb[7]) );
  AO2222XL U3031 ( .A(n203), .B(dph_reg[23]), .C(n179), .D(dph_reg[31]), .E(
        n2604), .F(dph_reg[7]), .G(n2605), .H(dph_reg[15]), .Y(n1554) );
  INVX1 U3032 ( .A(dpc_tab[3]), .Y(n1503) );
  INVX1 U3033 ( .A(dpc_tab[9]), .Y(n1504) );
  INVX1 U3034 ( .A(dpc_tab[15]), .Y(n1505) );
  AND2XL U3035 ( .A(phase0_ff), .B(waitstaten), .Y(newinstr) );
  MUX2XL U3036 ( .D0(ramsfraddr[6]), .D1(n2642), .S(waitstaten), .Y(
        ramsfraddr_comb[6]) );
  NAND21X1 U3037 ( .B(n382), .A(finishdiv), .Y(n2551) );
  NAND21X1 U3038 ( .B(n382), .A(finishmul), .Y(n2552) );
  NAND5XL U3039 ( .A(n378), .B(ramwe), .C(n2555), .D(n2554), .E(n2553), .Y(
        n2568) );
  AO2222XL U3040 ( .A(multemp2[4]), .B(n301), .C(n302), .D(n1827), .E(n1829), 
        .F(n394), .G(b[2]), .H(n1828), .Y(N12479) );
  AO2222XL U3041 ( .A(multemp2[5]), .B(n301), .C(n302), .D(n2068), .E(n1829), 
        .F(n390), .G(b[3]), .H(n1828), .Y(N12480) );
  AO2222XL U3042 ( .A(multemp2[6]), .B(n301), .C(n302), .D(n2075), .E(n1829), 
        .F(n402), .G(b[4]), .H(n1828), .Y(N12481) );
  AO2222XL U3043 ( .A(multemp2[8]), .B(n301), .C(n302), .D(n2076), .E(n1829), 
        .F(n413), .G(b[6]), .H(n1828), .Y(N12483) );
  AO2222XL U3044 ( .A(multemp2[7]), .B(n301), .C(n302), .D(n2074), .E(n1829), 
        .F(n387), .G(b[5]), .H(n1828), .Y(N12482) );
  AO2222XL U3045 ( .A(multemp2[9]), .B(n301), .C(n302), .D(n1830), .E(n1829), 
        .F(n406), .G(b[7]), .H(n1828), .Y(N12484) );
  MUX2XL U3046 ( .D0(N13352), .D1(n335), .S(N13353), .Y(n1830) );
  AO2222XL U3047 ( .A(multemp2[2]), .B(n301), .C(n302), .D(n357), .E(n1829), 
        .F(n409), .G(b[0]), .H(n1828), .Y(N12477) );
  AO2222XL U3048 ( .A(multemp2[3]), .B(n301), .C(n302), .D(n2067), .E(n1829), 
        .F(n398), .G(b[1]), .H(n1828), .Y(N12478) );
  MUX2X1 U3049 ( .D0(n398), .D1(f1), .S(n1809), .Y(n1883) );
  MUX2X1 U3050 ( .D0(gf0), .D1(n394), .S(n354), .Y(n1881) );
  MUX2X1 U3051 ( .D0(n387), .D1(f0), .S(n1809), .Y(n1882) );
  OAI221X1 U3052 ( .A(n2144), .B(n2188), .C(n2187), .D(n2143), .E(n433), .Y(
        N12489) );
  INVX1 U3053 ( .A(p2[4]), .Y(n2144) );
  OAI221X1 U3054 ( .A(n2145), .B(n2188), .C(n2187), .D(n2357), .E(n433), .Y(
        N12488) );
  INVX1 U3055 ( .A(p2[3]), .Y(n2145) );
  OAI221X1 U3056 ( .A(n2141), .B(n2188), .C(n2187), .D(n2140), .E(n433), .Y(
        N12491) );
  INVX1 U3057 ( .A(p2[6]), .Y(n2141) );
  OAI221X1 U3058 ( .A(n2138), .B(n2188), .C(n2187), .D(n2137), .E(n434), .Y(
        N12492) );
  INVX1 U3059 ( .A(p2[7]), .Y(n2138) );
  OAI221X1 U3060 ( .A(n2142), .B(n2188), .C(n2842), .D(n2187), .E(n433), .Y(
        N12490) );
  INVX1 U3061 ( .A(p2[5]), .Y(n2142) );
  INVX1 U3062 ( .A(n1825), .Y(n1828) );
  OAI211X1 U3063 ( .C(n1824), .D(n1823), .A(n379), .B(n1822), .Y(n1825) );
  OAI221XL U3064 ( .A(finishmul), .B(n1817), .C(finishdiv), .D(n1922), .E(
        n2201), .Y(n1824) );
  NAND43X1 U3065 ( .B(n294), .C(n1821), .D(n2202), .A(n1918), .Y(n1823) );
  OAI22XL U3066 ( .A(n1776), .B(n2216), .C(n2189), .D(n2140), .Y(N12706) );
  OA22XL U3067 ( .A(n1774), .B(n2205), .C(n1773), .D(n1772), .Y(n1776) );
  INVXL U3068 ( .A(ac), .Y(n1772) );
  MUX2XL U3069 ( .D0(n1866), .D1(n1763), .S(n1762), .Y(n1774) );
  OAI22X1 U3070 ( .A(n1888), .B(n381), .C(n2477), .D(n1887), .Y(N12723) );
  AND2X1 U3071 ( .A(n1886), .B(n1885), .Y(n1888) );
  AOI221XL U3072 ( .A(n2466), .B(temp[0]), .C(n2465), .D(temp2_comb[0]), .E(
        n1876), .Y(n1886) );
  OA2222XL U3073 ( .A(n2229), .B(n2473), .C(n2090), .D(n2471), .E(n1877), .F(
        n2469), .G(n2227), .H(n2467), .Y(n1885) );
  OAI22X1 U3074 ( .A(n2479), .B(n381), .C(n2478), .D(n2477), .Y(N12724) );
  AND2X1 U3075 ( .A(n2476), .B(n2475), .Y(n2479) );
  AOI221XL U3076 ( .A(n2466), .B(temp[1]), .C(n2465), .D(temp2_comb[1]), .E(
        n2464), .Y(n2476) );
  OA2222XL U3077 ( .A(n2474), .B(n2473), .C(n2472), .D(n2471), .E(n2470), .F(
        n2469), .G(n2468), .H(n2467), .Y(n2475) );
  INVX1 U3078 ( .A(n2597), .Y(n2598) );
  NAND5XL U3079 ( .A(n313), .B(n2136), .C(n2553), .D(ramsfraddr[5]), .E(n2135), 
        .Y(n2187) );
  NOR3XL U3080 ( .A(n1861), .B(n382), .C(finishmul), .Y(n355) );
  OA21X1 U3081 ( .B(n2164), .C(n2163), .A(n380), .Y(N12726) );
  OAI221X1 U3082 ( .A(n2162), .B(n2469), .C(n2855), .D(n2467), .E(n2161), .Y(
        n2163) );
  AO2222XL U3083 ( .A(n2365), .B(n76), .C(n2364), .D(n2158), .E(intvect[0]), 
        .F(n2591), .G(n2363), .H(n2157), .Y(n2164) );
  INVX1 U3084 ( .A(pc_i[11]), .Y(n2162) );
  OA21X1 U3085 ( .B(n1894), .C(n1893), .A(n380), .Y(N12727) );
  OAI221X1 U3086 ( .A(n2395), .B(n2469), .C(n2854), .D(n2467), .E(n1892), .Y(
        n1893) );
  AO2222XL U3087 ( .A(n2365), .B(n65), .C(n2364), .D(n1938), .E(intvect[1]), 
        .F(n2591), .G(n2363), .H(n1982), .Y(n1894) );
  OA222X1 U3088 ( .A(n2396), .B(n2368), .C(n39), .D(n2367), .E(n2382), .F(
        n2366), .Y(n1892) );
  OA21X1 U3089 ( .B(n1805), .C(n1804), .A(n380), .Y(N12728) );
  OAI221X1 U3090 ( .A(n2312), .B(n2469), .C(n2853), .D(n2467), .E(n1803), .Y(
        n1804) );
  AO2222XL U3091 ( .A(n2365), .B(n70), .C(n2364), .D(n1936), .E(intvect[2]), 
        .F(n2591), .G(n2363), .H(n2287), .Y(n1805) );
  OA222X1 U3092 ( .A(n2313), .B(n2368), .C(n45), .D(n2367), .E(n2293), .F(
        n2366), .Y(n1803) );
  OA21X1 U3093 ( .B(n2056), .C(n2055), .A(n380), .Y(N12729) );
  OAI221X1 U3094 ( .A(n2345), .B(n2469), .C(n2852), .D(n2467), .E(n2054), .Y(
        n2055) );
  AO2222XL U3095 ( .A(n2365), .B(n81), .C(n2364), .D(n2057), .E(intvect[3]), 
        .F(n2591), .G(n2363), .H(n2053), .Y(n2056) );
  OA222X1 U3096 ( .A(n2344), .B(n2368), .C(n43), .D(n2367), .E(n2328), .F(
        n2366), .Y(n2054) );
  OA21X1 U3097 ( .B(n2371), .C(n2370), .A(n380), .Y(N12730) );
  OAI221X1 U3098 ( .A(n2441), .B(n2469), .C(n2851), .D(n2467), .E(n2369), .Y(
        n2370) );
  AO2222XL U3099 ( .A(n2365), .B(n69), .C(n2364), .D(n2372), .E(intvect[4]), 
        .F(n2591), .G(n2363), .H(n2362), .Y(n2371) );
  OA222X1 U3100 ( .A(n2438), .B(n2368), .C(n37), .D(n2367), .E(n2410), .F(
        n2366), .Y(n2369) );
  NOR3XL U3101 ( .A(n383), .B(n1826), .C(finishdiv), .Y(n356) );
  NOR32XL U3102 ( .B(n376), .C(n2549), .A(newinstrlock), .Y(N689) );
  AND2XL U3103 ( .A(n2355), .B(phase[1]), .Y(N681) );
  AND2XL U3104 ( .A(n2355), .B(n2549), .Y(N680) );
  AND2X1 U3105 ( .A(n2355), .B(phase[2]), .Y(N682) );
  AND2X1 U3106 ( .A(n2355), .B(phase[3]), .Y(N683) );
  AND2X1 U3107 ( .A(n2355), .B(phase[4]), .Y(N684) );
  AND2X1 U3108 ( .A(state[1]), .B(n378), .Y(N589) );
  AND2X1 U3109 ( .A(state[2]), .B(n379), .Y(N590) );
  INVX1 U3110 ( .A(dph_reg[60]), .Y(n2751) );
  INVX1 U3111 ( .A(dph_reg[52]), .Y(n2752) );
  INVX1 U3112 ( .A(dph_reg[21]), .Y(n2758) );
  INVX1 U3113 ( .A(dph_reg[20]), .Y(n2754) );
  INVX1 U3114 ( .A(dph_reg[28]), .Y(n2753) );
  AO21X1 U3115 ( .B(d_hold), .C(n1395), .A(cpu_resume_fff), .Y(n2509) );
  INVX1 U3116 ( .A(cpu_hold), .Y(n1395) );
  NAND21X1 U3117 ( .B(n1499), .A(n1498), .Y(dpc[4]) );
  OA2222XL U3118 ( .A(n366), .B(n1497), .C(n368), .D(n1496), .E(n370), .F(
        n1495), .G(n372), .H(n1494), .Y(n1498) );
  AO2222XL U3119 ( .A(dpc_tab[28]), .B(n132), .C(dpc_tab[34]), .D(n148), .E(
        dpc_tab[40]), .F(n180), .G(dpc_tab[46]), .H(n164), .Y(n1499) );
  INVX1 U3120 ( .A(dpc_tab[22]), .Y(n1497) );
  AOI22BXL U3121 ( .B(n370), .A(dpl_reg[13]), .D(n372), .C(dpl_reg[5]), .Y(
        n585) );
  AOI22BXL U3122 ( .B(n369), .A(dpl_reg[12]), .D(n371), .C(dpl_reg[4]), .Y(
        n589) );
  AOI22BXL U3123 ( .B(n370), .A(dph_reg[12]), .D(n372), .C(dph_reg[4]), .Y(
        n621) );
  AOI22BXL U3124 ( .B(n2802), .A(dpl_reg[45]), .D(n134), .C(dpl_reg[37]), .Y(
        n583) );
  AOI22BXL U3125 ( .B(n2802), .A(dph_reg[45]), .D(n134), .C(dph_reg[37]), .Y(
        n615) );
  AOI22BXL U3126 ( .B(n2802), .A(dpl_reg[44]), .D(n134), .C(dpl_reg[36]), .Y(
        n587) );
  AOI22BXL U3127 ( .B(n2802), .A(dph_reg[44]), .D(n134), .C(dph_reg[36]), .Y(
        n619) );
  AOI221XL U3128 ( .A(phase[0]), .B(n2109), .C(phase[1]), .D(n2108), .E(n2107), 
        .Y(n2426) );
  INVX1 U3129 ( .A(n2106), .Y(n2107) );
  AOI21BX1 U3130 ( .C(test_so), .B(n933), .A(n934), .Y(N12976) );
  INVXL U3131 ( .A(ramsfraddr[6]), .Y(n2553) );
  INVX1 U3132 ( .A(dph_reg[61]), .Y(n2755) );
  INVX1 U3133 ( .A(dph_reg[62]), .Y(n2759) );
  INVX1 U3134 ( .A(dph_reg[53]), .Y(n2756) );
  INVX1 U3135 ( .A(dph_reg[54]), .Y(n2760) );
  INVX1 U3136 ( .A(dph_reg[22]), .Y(n2762) );
  INVX1 U3137 ( .A(dph_reg[30]), .Y(n2761) );
  INVX1 U3138 ( .A(dph_reg[29]), .Y(n2757) );
  NAND21X1 U3139 ( .B(n2082), .A(n2081), .Y(dpc[5]) );
  OA2222XL U3140 ( .A(n365), .B(n2080), .C(n367), .D(n2079), .E(n2808), .F(
        n2078), .G(n371), .H(n2077), .Y(n2081) );
  AO2222XL U3141 ( .A(dpc_tab[29]), .B(n132), .C(dpc_tab[35]), .D(n148), .E(
        dpc_tab[41]), .F(n180), .G(dpc_tab[47]), .H(n164), .Y(n2082) );
  INVX1 U3142 ( .A(dpc_tab[23]), .Y(n2080) );
  AOI22BXL U3143 ( .B(n2808), .A(dph_reg[13]), .D(n2807), .C(dph_reg[5]), .Y(
        n617) );
  AOI22BXL U3144 ( .B(n2802), .A(dph_reg[46]), .D(n134), .C(dph_reg[38]), .Y(
        n611) );
  AOI22BXL U3145 ( .B(n2802), .A(dpl_reg[46]), .D(n134), .C(dpl_reg[38]), .Y(
        n579) );
  INVX1 U3146 ( .A(p2[1]), .Y(n2232) );
  INVX1 U3147 ( .A(p2[0]), .Y(n2222) );
  INVX1 U3148 ( .A(dph_reg[55]), .Y(n2764) );
  INVX1 U3149 ( .A(dph_reg[39]), .Y(n2765) );
  INVX1 U3150 ( .A(dph_reg[47]), .Y(n2766) );
  INVX1 U3151 ( .A(dph_reg[63]), .Y(n2763) );
  INVX1 U3152 ( .A(dpc_tab[4]), .Y(n1494) );
  AOI22BXL U3153 ( .B(n369), .A(dph_reg[14]), .D(n371), .C(dph_reg[6]), .Y(
        n613) );
  AOI22BXL U3154 ( .B(n2808), .A(dpl_reg[14]), .D(n2807), .C(dpl_reg[6]), .Y(
        n581) );
  AOI22BXL U3155 ( .B(n370), .A(dph_reg[15]), .D(n372), .C(dph_reg[7]), .Y(
        n609) );
  AOI22BXL U3156 ( .B(n369), .A(dpl_reg[15]), .D(n371), .C(dpl_reg[7]), .Y(
        n569) );
  AOI22BXL U3157 ( .B(n367), .A(dph_reg[23]), .D(n366), .C(dph_reg[31]), .Y(
        n608) );
  AOI22BXL U3158 ( .B(n2802), .A(dpl_reg[47]), .D(n134), .C(dpl_reg[39]), .Y(
        n567) );
  INVX1 U3159 ( .A(p2[2]), .Y(n2240) );
  INVX1 U3160 ( .A(dpc_tab[5]), .Y(n2077) );
  INVX1 U3161 ( .A(dpc_tab[11]), .Y(n2078) );
  INVX1 U3162 ( .A(dpc_tab[10]), .Y(n1495) );
  INVX1 U3163 ( .A(dpc_tab[17]), .Y(n2079) );
  INVX1 U3164 ( .A(dpc_tab[16]), .Y(n1496) );
  MUX2BXL U3165 ( .D0(N13345), .D1(n2329), .S(N13353), .Y(n357) );
  NAND21X1 U3166 ( .B(n1530), .A(memaddr[5]), .Y(n1529) );
  NAND21XL U3167 ( .B(n1474), .A(pc_o[3]), .Y(n1462) );
  NAND21XL U3168 ( .B(n53), .A(pc_o[2]), .Y(n1474) );
  NOR32XL U3169 ( .B(n2212), .C(n2211), .A(n2210), .Y(n2213) );
  NAND42XL U3170 ( .C(b[4]), .D(b[6]), .A(n2199), .B(n2198), .Y(n2212) );
  NAND21X1 U3171 ( .B(n2204), .A(n2203), .Y(n2211) );
  NOR32XL U3172 ( .B(n294), .C(n2209), .A(n2208), .Y(n2210) );
  INVX1 U3173 ( .A(n1469), .Y(n2152) );
  OAI221X1 U3174 ( .A(n177), .B(n2102), .C(n2153), .D(n1579), .E(n1468), .Y(
        n1469) );
  MUX2XL U3175 ( .D0(n1467), .D1(n1465), .S(memaddr[3]), .Y(n1468) );
  NAND21X1 U3176 ( .B(n307), .A(n1475), .Y(n1467) );
  AO21XL U3177 ( .B(n2865), .C(n2840), .A(n1231), .Y(n1486) );
  MUX2X1 U3178 ( .D0(n1335), .D1(n1334), .S(pc_o[9]), .Y(n1572) );
  OAI21AX1 U3179 ( .B(n1328), .C(n2838), .A(n1336), .Y(n1335) );
  INVX1 U3180 ( .A(n1580), .Y(n1600) );
  OAI211X1 U3181 ( .C(n1877), .D(n1579), .A(n1578), .B(n1577), .Y(n1580) );
  INVX1 U3182 ( .A(n1336), .Y(n1577) );
  MUX2BXL U3183 ( .D0(n1576), .D1(n1350), .S(pc_o[8]), .Y(n1578) );
  NAND21X1 U3184 ( .B(n2060), .A(temp2_comb[7]), .Y(n1449) );
  AO21XL U3185 ( .B(pc_o[3]), .C(n1455), .A(n1464), .Y(n1456) );
  NOR3XL U3186 ( .A(pc_o[13]), .B(pc_o[14]), .C(n1293), .Y(n1286) );
  MUX2X1 U3187 ( .D0(n1317), .D1(n1316), .S(pc_o[11]), .Y(n1568) );
  OAI21X1 U3188 ( .B(n1310), .C(n2838), .A(n1318), .Y(n1317) );
  MUX2X1 U3189 ( .D0(n1299), .D1(n1298), .S(pc_o[13]), .Y(n1564) );
  OAI21X1 U3190 ( .B(n1294), .C(n2838), .A(n1293), .Y(n1299) );
  MUX2BXL U3191 ( .D0(n1549), .D1(n1548), .S(pc_o[15]), .Y(n1550) );
  AO21X1 U3192 ( .B(n1545), .C(pc_o[14]), .A(n1286), .Y(n1549) );
  NAND2X1 U3193 ( .A(pc_o[6]), .B(n1466), .Y(n1426) );
  NAND2X1 U3194 ( .A(state[0]), .B(n2809), .Y(n530) );
  INVX1 U3195 ( .A(n1251), .Y(n1607) );
  OAI211X1 U3196 ( .C(n2253), .D(n1579), .A(n1318), .B(n1250), .Y(n1251) );
  MUX2BXL U3197 ( .D0(n1249), .D1(n1326), .S(pc_o[10]), .Y(n1250) );
  NAND21X1 U3198 ( .B(n177), .A(n1320), .Y(n1249) );
  INVX1 U3199 ( .A(n1391), .Y(n1606) );
  OAI211X1 U3200 ( .C(n2395), .D(n1579), .A(n1293), .B(n1390), .Y(n1391) );
  MUX2BXL U3201 ( .D0(n1389), .D1(n1309), .S(pc_o[12]), .Y(n1390) );
  NAND21X1 U3202 ( .B(n2838), .A(n1303), .Y(n1389) );
  INVX1 U3203 ( .A(n1560), .Y(n1604) );
  OAI211X1 U3204 ( .C(n2345), .D(n1579), .A(n1559), .B(n1558), .Y(n1560) );
  INVX1 U3205 ( .A(n1286), .Y(n1559) );
  MUX2X1 U3206 ( .D0(n1557), .D1(n1556), .S(pc_o[14]), .Y(n1558) );
  INVX1 U3207 ( .A(n1458), .Y(n1544) );
  OAI211X1 U3208 ( .C(n2397), .D(n1579), .A(n308), .B(n1457), .Y(n1458) );
  AND2X1 U3209 ( .A(n1556), .B(n1547), .Y(n1548) );
  MUX2X1 U3210 ( .D0(n2838), .D1(n1288), .S(pc_o[14]), .Y(n1547) );
  AND2XL U3211 ( .A(b[7]), .B(n193), .Y(N14351) );
  AND2XL U3212 ( .A(b[2]), .B(n193), .Y(N14346) );
  AND2XL U3213 ( .A(b[4]), .B(n170), .Y(N14340) );
  AND2XL U3214 ( .A(b[3]), .B(n193), .Y(N14347) );
  AND2XL U3215 ( .A(b[5]), .B(n170), .Y(N14341) );
  AND2XL U3216 ( .A(b[4]), .B(n193), .Y(N14348) );
  AND2XL U3217 ( .A(b[6]), .B(n170), .Y(N14342) );
  AND2XL U3218 ( .A(b[5]), .B(n193), .Y(N14349) );
  AND2XL U3219 ( .A(b[6]), .B(n193), .Y(N14350) );
  AND2XL U3220 ( .A(b[1]), .B(acc[1]), .Y(N14345) );
  AND2XL U3221 ( .A(b[2]), .B(acc[0]), .Y(N14338) );
  AND2XL U3222 ( .A(b[3]), .B(acc[0]), .Y(N14339) );
  AND2XL U3223 ( .A(b[7]), .B(n170), .Y(N14343) );
  NOR2X1 U3224 ( .A(n1525), .B(n359), .Y(n358) );
  OAI22X1 U3225 ( .A(n177), .B(n2340), .C(n2346), .D(n1579), .Y(n359) );
  INVX1 U3226 ( .A(n1517), .Y(n2089) );
  OAI221X1 U3227 ( .A(n2443), .B(n1579), .C(n177), .D(n2432), .E(n1516), .Y(
        n1517) );
  MUX2X1 U3228 ( .D0(n1515), .D1(n2817), .S(memaddr[7]), .Y(n1516) );
  INVX1 U3229 ( .A(n1524), .Y(n1515) );
  INVX1 U3230 ( .A(n1534), .Y(n2049) );
  OAI221X1 U3231 ( .A(n177), .B(n2310), .C(n2320), .D(n1579), .E(n1533), .Y(
        n1534) );
  MUX2X1 U3232 ( .D0(n308), .D1(n1532), .S(memaddr[5]), .Y(n1533) );
  INVX1 U3233 ( .A(n1531), .Y(n1532) );
  MUX2XL U3234 ( .D0(n1487), .D1(n1486), .S(pc_o[1]), .Y(n1488) );
  NAND21X1 U3235 ( .B(n1216), .A(n307), .Y(n1487) );
  INVX1 U3236 ( .A(n1479), .Y(n2147) );
  OAI211X1 U3237 ( .C(n2254), .D(n1579), .A(n1478), .B(n1477), .Y(n1479) );
  MUX2X1 U3238 ( .D0(n1238), .D1(n177), .S(n1473), .Y(n1478) );
  AOI22XL U3239 ( .A(n1476), .B(n2840), .C(pc_o[2]), .D(n1486), .Y(n1477) );
  NOR32XL U3240 ( .B(n41), .C(n1312), .A(pc_o[11]), .Y(n1302) );
  NAND32X1 U3241 ( .B(memaddr[6]), .C(n1521), .A(n45), .Y(n1512) );
  NAND32XL U3242 ( .B(pc_o[3]), .C(n1463), .A(n39), .Y(n1511) );
  NAND21XL U3243 ( .B(memaddr[0]), .A(n1523), .Y(n1521) );
  NAND21XL U3244 ( .B(pc_o[2]), .A(n53), .Y(n1463) );
  NAND21X1 U3245 ( .B(n1225), .A(n1239), .Y(n1414) );
  AND3X1 U3246 ( .A(n1238), .B(n177), .C(n2827), .Y(n1413) );
  NOR3XL U3247 ( .A(pc_o[10]), .B(pc_o[9]), .C(n1330), .Y(n1312) );
  NAND2X1 U3248 ( .A(n1303), .B(pc_o[12]), .Y(n1294) );
  NAND2X1 U3249 ( .A(n1337), .B(pc_o[8]), .Y(n1328) );
  NAND2X1 U3250 ( .A(n1320), .B(pc_o[10]), .Y(n1310) );
  INVX1 U3251 ( .A(pdmode), .Y(n2532) );
  NOR32XL U3252 ( .B(n41), .C(n1311), .A(pc_o[11]), .Y(n1301) );
  NAND32X1 U3253 ( .B(pc_o[6]), .C(n1511), .A(n45), .Y(n1513) );
  INVX1 U3254 ( .A(memaddr[10]), .Y(n2255) );
  MUX2XL U3255 ( .D0(n1715), .D1(n1714), .S(instr[3]), .Y(n1726) );
  AO21XL U3256 ( .B(n2463), .C(memaddr[0]), .A(n2591), .Y(n1876) );
  AO21XL U3257 ( .B(n2463), .C(pc_o[1]), .A(n2591), .Y(n2464) );
  NOR3XL U3258 ( .A(pc_o[10]), .B(pc_o[9]), .C(n1329), .Y(n1311) );
  OAI31XL U3259 ( .A(n204), .B(n1721), .C(n1720), .D(n1719), .Y(n1724) );
  AO21XL U3260 ( .B(n1718), .C(n152), .A(n1716), .Y(n1719) );
  NOR21XL U3261 ( .B(n2645), .A(n1296), .Y(n2490) );
  NOR43XL U3262 ( .B(n2492), .C(phase[1]), .D(n1304), .A(ramsfraddr[7]), .Y(
        n1296) );
  AO21XL U3263 ( .B(n2538), .C(n2549), .A(n2452), .Y(n1739) );
  AO21XL U3264 ( .B(n1713), .C(n214), .A(n1712), .Y(n1743) );
  INVX1 U3265 ( .A(memaddr[14]), .Y(n2489) );
  NOR21XL U3266 ( .B(pc_o[15]), .A(n2488), .Y(n2376) );
  NAND5XL U3267 ( .A(phase[1]), .B(ramsfraddr[7]), .C(n435), .D(n2492), .E(
        n1304), .Y(n2495) );
  INVXL U3268 ( .A(b[3]), .Y(n2197) );
  INVXL U3269 ( .A(b[2]), .Y(n2196) );
  AND2XL U3270 ( .A(n1727), .B(instr[2]), .Y(n1729) );
  INVX1 U3271 ( .A(memaddr[11]), .Y(n2849) );
  AO21XL U3272 ( .B(instr[3]), .C(n418), .A(n2008), .Y(n1663) );
  INVX1 U3273 ( .A(n1814), .Y(n2652) );
  AND2XL U3274 ( .A(n416), .B(n34), .Y(n1813) );
  MUX2XL U3275 ( .D0(n214), .D1(n2549), .S(n1811), .Y(n1812) );
  AO21XL U3276 ( .B(n1946), .C(n204), .A(n1295), .Y(n1304) );
  OAI31XL U3277 ( .A(instr[4]), .B(n1778), .C(n1382), .D(n1785), .Y(n1295) );
  OAI211XL U3278 ( .C(instr[3]), .D(n1613), .A(n1612), .B(n1944), .Y(n1648) );
  NAND21XL U3279 ( .B(dec_accop[10]), .A(dec_accop[9]), .Y(n2209) );
  OAI22X1 U3280 ( .A(n940), .B(n1634), .C(n941), .D(n2633), .Y(N12972) );
  INVX1 U3281 ( .A(ckcon[7]), .Y(n1634) );
  OAI22X1 U3282 ( .A(n940), .B(n2616), .C(n941), .D(n2630), .Y(N12970) );
  INVX1 U3283 ( .A(ckcon[5]), .Y(n2616) );
  OAI22XL U3284 ( .A(n940), .B(n2279), .C(n941), .D(n2278), .Y(N12965) );
  INVX1 U3285 ( .A(ckcon[0]), .Y(n2279) );
  OAI22XL U3286 ( .A(n940), .B(n2615), .C(n941), .D(n2628), .Y(N12969) );
  INVX1 U3287 ( .A(ckcon[4]), .Y(n2615) );
  OAI22XL U3288 ( .A(n940), .B(n2276), .C(n941), .D(n2275), .Y(N12968) );
  INVX1 U3289 ( .A(ckcon[3]), .Y(n2276) );
  NOR3XL U3290 ( .A(b[0]), .B(b[1]), .C(n2194), .Y(n2199) );
  INVXL U3291 ( .A(b[5]), .Y(n2193) );
  AND2X1 U3292 ( .A(cpu_resume_ff1), .B(n434), .Y(N13380) );
  INVX1 U3293 ( .A(stop), .Y(n1400) );
  INVX1 U3294 ( .A(ov), .Y(n2204) );
  NAND21X1 U3295 ( .B(n2707), .A(waitcnt_0_), .Y(n933) );
  INVX1 U3296 ( .A(n2563), .Y(n2578) );
  NAND32XL U3297 ( .B(ramsfraddr[0]), .C(n2562), .A(n2561), .Y(n2563) );
  BUFXL U3298 ( .A(n2865), .Y(pc_o[0]) );
  INVXL U3299 ( .A(n363), .Y(n1226) );
  INVXL U3300 ( .A(n84), .Y(n361) );
  INVX2 U3301 ( .A(n361), .Y(n362) );
  MUX2IX1 U3302 ( .D0(n2332), .D1(n1199), .S(n1205), .Y(n364) );
  INVXL U3303 ( .A(n2664), .Y(n1211) );
  OAI221XL U3304 ( .A(n2094), .B(n2439), .C(n1228), .D(n1227), .E(n1226), .Y(
        n1237) );
  OAI22XL U3305 ( .A(n424), .B(n2231), .C(n2495), .D(n2230), .Y(N12714) );
  AOI211X1 U3306 ( .C(n108), .D(n1205), .A(n363), .B(n1204), .Y(n1206) );
  MUX2XL U3307 ( .D0(pc_o[10]), .D1(n2691), .S(n362), .Y(memaddr_comb[10]) );
  MUX2XL U3308 ( .D0(pc_o[8]), .D1(n2688), .S(n362), .Y(memaddr_comb[8]) );
  MUX2XL U3309 ( .D0(pc_o[9]), .D1(n2689), .S(n362), .Y(memaddr_comb[9]) );
  MUX2XL U3310 ( .D0(pc_o[7]), .D1(n2687), .S(n362), .Y(memaddr_comb[7]) );
  AO21X4 U3311 ( .B(n1081), .C(n1076), .A(n1082), .Y(n1913) );
  GEN2X1 U3312 ( .D(acc[3]), .E(n1418), .C(ac), .B(n1420), .A(n1689), .Y(n1428) );
  AO44X4 U3313 ( .A(n2132), .B(n1245), .C(n1210), .D(n1209), .E(n1208), .F(
        n2666), .G(n2515), .H(n2502), .Y(n2667) );
  MAJ3X1 U3314 ( .A(n1432), .B(n1431), .C(n1688), .Y(n1795) );
  MAJ3X1 U3315 ( .A(n1433), .B(n1795), .C(n1793), .Y(n1915) );
  MAJ3X1 U3316 ( .A(n1915), .B(n1437), .C(n1914), .Y(n2206) );
  MAJ3X1 U3317 ( .A(n2113), .B(n2426), .C(n2258), .Y(n2307) );
  MAJ3X1 U3318 ( .A(n2308), .B(n2426), .C(n2307), .Y(n2389) );
  MAJ3X1 U3319 ( .A(n2426), .B(n2309), .C(n2389), .Y(n2338) );
  MAJ3X1 U3320 ( .A(n2426), .B(n2338), .C(n298), .Y(n2425) );
  MAJ3X1 U3321 ( .A(n2426), .B(n2425), .C(n299), .Y(n2427) );
  AO33X4 U3322 ( .A(n1833), .B(n2672), .C(n2671), .D(n2670), .E(n2669), .F(
        n2671), .Y(n2673) );
endmodule


module mcu51_cpu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n25, n26, n27, n28, n29, n33, n34, n35, n36,
         n38, n40, n41, n42, n43, n45, n48, n54, n103, n104, n105, n106;

  XOR2X1 U2 ( .A(A[8]), .B(B[15]), .Y(n2) );
  FAD1X1 U3 ( .A(B[14]), .B(A[8]), .CI(n11), .CO(n10), .SO(SUM[14]) );
  FAD1X1 U4 ( .A(B[13]), .B(A[8]), .CI(n12), .CO(n11), .SO(SUM[13]) );
  FAD1X1 U5 ( .A(B[12]), .B(A[8]), .CI(n13), .CO(n12), .SO(SUM[12]) );
  FAD1X1 U6 ( .A(B[11]), .B(A[8]), .CI(n14), .CO(n13), .SO(SUM[11]) );
  FAD1X1 U7 ( .A(B[10]), .B(A[8]), .CI(n15), .CO(n14), .SO(SUM[10]) );
  FAD1X1 U8 ( .A(B[9]), .B(A[8]), .CI(n16), .CO(n15), .SO(SUM[9]) );
  FAD1X1 U9 ( .A(B[8]), .B(A[8]), .CI(n17), .CO(n16), .SO(SUM[8]) );
  FAD1X1 U10 ( .A(A[7]), .B(B[7]), .CI(n18), .CO(n17), .SO(SUM[7]) );
  XOR2X1 U11 ( .A(n21), .B(n3), .Y(SUM[6]) );
  OAI21X1 U12 ( .B(n21), .C(n19), .A(n20), .Y(n18) );
  NOR2X1 U15 ( .A(B[6]), .B(A[6]), .Y(n19) );
  XOR2X1 U25 ( .A(n29), .B(n5), .Y(SUM[4]) );
  OAI21X1 U26 ( .B(n29), .C(n27), .A(n28), .Y(n26) );
  NOR2X1 U29 ( .A(B[4]), .B(A[4]), .Y(n27) );
  OAI21X1 U40 ( .B(n1), .C(n35), .A(n36), .Y(n34) );
  AOI21X1 U42 ( .B(n45), .C(n104), .A(n38), .Y(n36) );
  OAI21X1 U50 ( .B(n1), .C(n42), .A(n43), .Y(n41) );
  NOR2X1 U57 ( .A(A[1]), .B(B[1]), .Y(n42) );
  NOR2X1 U62 ( .A(A[0]), .B(B[0]), .Y(n48) );
  NAND2XL U67 ( .A(n104), .B(n40), .Y(n7) );
  NAND2XL U68 ( .A(B[2]), .B(A[2]), .Y(n40) );
  XNOR2XL U69 ( .A(n7), .B(n41), .Y(SUM[2]) );
  OR2X1 U70 ( .A(B[2]), .B(A[2]), .Y(n104) );
  OR2X1 U71 ( .A(B[3]), .B(A[3]), .Y(n105) );
  INVXL U72 ( .A(n43), .Y(n45) );
  INVXL U73 ( .A(n42), .Y(n54) );
  NAND2XL U74 ( .A(n105), .B(n33), .Y(n6) );
  NAND2XL U75 ( .A(n106), .B(n25), .Y(n4) );
  NAND2XL U76 ( .A(B[4]), .B(A[4]), .Y(n28) );
  NAND2XL U77 ( .A(B[6]), .B(A[6]), .Y(n20) );
  NAND2XL U78 ( .A(B[5]), .B(A[5]), .Y(n25) );
  NAND21XL U79 ( .B(n48), .A(n1), .Y(n9) );
  AOI21AX1 U80 ( .B(n34), .C(n105), .A(n33), .Y(n29) );
  AOI21AX1 U81 ( .B(n26), .C(n106), .A(n25), .Y(n21) );
  NAND2X1 U82 ( .A(n54), .B(n104), .Y(n35) );
  NAND21X1 U83 ( .B(n19), .A(n20), .Y(n3) );
  INVX1 U84 ( .A(n40), .Y(n38) );
  XNOR2XL U85 ( .A(n1), .B(n103), .Y(SUM[1]) );
  AND2XL U86 ( .A(n54), .B(n43), .Y(n103) );
  NAND21XL U87 ( .B(n27), .A(n28), .Y(n5) );
  XNOR2XL U88 ( .A(n6), .B(n34), .Y(SUM[3]) );
  XNOR2XL U89 ( .A(n4), .B(n26), .Y(SUM[5]) );
  NAND2X1 U90 ( .A(A[0]), .B(B[0]), .Y(n1) );
  NAND2X1 U91 ( .A(A[1]), .B(B[1]), .Y(n43) );
  OR2X1 U92 ( .A(B[5]), .B(A[5]), .Y(n106) );
  NAND2X1 U93 ( .A(B[3]), .B(A[3]), .Y(n33) );
  INVX1 U94 ( .A(n9), .Y(SUM[0]) );
  XOR2X1 U95 ( .A(n10), .B(n2), .Y(SUM[15]) );
endmodule


module mcu51_cpu_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n15, n16, n17, n18, n19,
         n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n79, n80;

  FAD1X1 U2 ( .A(A[7]), .B(n38), .CI(n8), .CO(n7), .SO(DIFF[7]) );
  XOR2X1 U3 ( .A(n11), .B(n1), .Y(DIFF[6]) );
  OAI21X1 U4 ( .B(n11), .C(n9), .A(n10), .Y(n8) );
  NOR2X1 U7 ( .A(A[6]), .B(n39), .Y(n9) );
  XOR2X1 U17 ( .A(n19), .B(n3), .Y(DIFF[4]) );
  OAI21X1 U18 ( .B(n19), .C(n17), .A(n18), .Y(n16) );
  NOR2X1 U21 ( .A(A[4]), .B(n41), .Y(n17) );
  NOR2X1 U25 ( .A(n22), .B(n25), .Y(n20) );
  NOR2X1 U29 ( .A(A[3]), .B(n42), .Y(n22) );
  XOR2X1 U31 ( .A(n27), .B(n5), .Y(DIFF[2]) );
  OAI21X1 U32 ( .B(n27), .C(n25), .A(n26), .Y(n24) );
  NOR2X1 U35 ( .A(A[2]), .B(n43), .Y(n25) );
  XOR2X1 U37 ( .A(n6), .B(n31), .Y(DIFF[1]) );
  OAI21X1 U39 ( .B(n29), .C(n31), .A(n30), .Y(n28) );
  NOR2X1 U42 ( .A(A[1]), .B(n44), .Y(n29) );
  NOR2X1 U45 ( .A(n45), .B(A[0]), .Y(n31) );
  OR2X1 U57 ( .A(A[5]), .B(n40), .Y(n80) );
  XNOR2XL U58 ( .A(A[0]), .B(n45), .Y(DIFF[0]) );
  OAI21X1 U59 ( .B(n22), .C(n26), .A(n23), .Y(n79) );
  AOI21X1 U60 ( .B(n28), .C(n20), .A(n79), .Y(n19) );
  NAND2XL U61 ( .A(A[4]), .B(n41), .Y(n18) );
  NAND2XL U62 ( .A(A[6]), .B(n39), .Y(n10) );
  INVXL U63 ( .A(n17), .Y(n34) );
  NAND2XL U64 ( .A(n34), .B(n18), .Y(n3) );
  INVXL U65 ( .A(n9), .Y(n32) );
  NAND2XL U66 ( .A(n32), .B(n10), .Y(n1) );
  AOI21AX1 U67 ( .B(n16), .C(n80), .A(n15), .Y(n11) );
  INVXL U68 ( .A(n28), .Y(n27) );
  INVXL U69 ( .A(n22), .Y(n35) );
  INVX2 U70 ( .A(n7), .Y(DIFF[8]) );
  NAND2X1 U71 ( .A(A[2]), .B(n43), .Y(n26) );
  NAND2X1 U72 ( .A(A[1]), .B(n44), .Y(n30) );
  NAND2X1 U73 ( .A(A[3]), .B(n42), .Y(n23) );
  NAND2X1 U74 ( .A(A[5]), .B(n40), .Y(n15) );
  NAND2XL U75 ( .A(n36), .B(n26), .Y(n5) );
  INVXL U76 ( .A(n25), .Y(n36) );
  XNOR2XL U77 ( .A(n4), .B(n24), .Y(DIFF[3]) );
  NAND2X1 U78 ( .A(n35), .B(n23), .Y(n4) );
  XNOR2XL U79 ( .A(n2), .B(n16), .Y(DIFF[5]) );
  NAND2XL U80 ( .A(n80), .B(n15), .Y(n2) );
  NAND2X1 U81 ( .A(n37), .B(n30), .Y(n6) );
  INVX1 U82 ( .A(n29), .Y(n37) );
  INVX1 U83 ( .A(B[7]), .Y(n38) );
  INVXL U84 ( .A(B[1]), .Y(n44) );
  INVXL U85 ( .A(B[2]), .Y(n43) );
  INVXL U86 ( .A(B[3]), .Y(n42) );
  INVXL U87 ( .A(B[0]), .Y(n45) );
  INVXL U88 ( .A(B[4]), .Y(n41) );
  INVXL U89 ( .A(B[5]), .Y(n40) );
  INVXL U90 ( .A(B[6]), .Y(n39) );
endmodule


module mcu51_cpu_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n15, n16, n17, n18, n19,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n38, n39, n40,
         n41, n42, n43, n44, n45, n78, n79;

  XOR2X1 U3 ( .A(n11), .B(n1), .Y(DIFF[6]) );
  OAI21X1 U4 ( .B(n11), .C(n9), .A(n10), .Y(n8) );
  NOR2X1 U7 ( .A(n39), .B(A[6]), .Y(n9) );
  XOR2X1 U17 ( .A(n19), .B(n3), .Y(DIFF[4]) );
  OAI21X1 U18 ( .B(n19), .C(n17), .A(n18), .Y(n16) );
  NOR2X1 U21 ( .A(n41), .B(A[4]), .Y(n17) );
  OAI21X1 U26 ( .B(n22), .C(n26), .A(n23), .Y(n21) );
  NOR2X1 U29 ( .A(n42), .B(A[3]), .Y(n22) );
  XOR2X1 U31 ( .A(n27), .B(n5), .Y(DIFF[2]) );
  OAI21X1 U32 ( .B(n27), .C(n25), .A(n26), .Y(n24) );
  NOR2X1 U35 ( .A(n43), .B(A[2]), .Y(n25) );
  XOR2X1 U37 ( .A(n6), .B(n31), .Y(DIFF[1]) );
  OAI21X1 U39 ( .B(n29), .C(n31), .A(n30), .Y(n28) );
  NOR2X1 U42 ( .A(n44), .B(A[1]), .Y(n29) );
  NOR2X1 U45 ( .A(n45), .B(A[0]), .Y(n31) );
  INVX1 U57 ( .A(B[3]), .Y(n42) );
  INVX1 U58 ( .A(B[5]), .Y(n40) );
  INVX1 U59 ( .A(B[4]), .Y(n41) );
  INVX1 U60 ( .A(B[1]), .Y(n44) );
  INVX1 U61 ( .A(B[6]), .Y(n39) );
  XNOR2XL U62 ( .A(n4), .B(n24), .Y(DIFF[3]) );
  XNOR2XL U63 ( .A(n2), .B(n16), .Y(DIFF[5]) );
  XNOR2XL U64 ( .A(A[0]), .B(n45), .Y(DIFF[0]) );
  OR2X1 U65 ( .A(n40), .B(A[5]), .Y(n78) );
  NAND2X1 U66 ( .A(n44), .B(A[1]), .Y(n30) );
  NOR2XL U67 ( .A(n25), .B(n22), .Y(n79) );
  INVX1 U68 ( .A(B[7]), .Y(n38) );
  INVX3 U69 ( .A(B[2]), .Y(n43) );
  AOI21X1 U70 ( .B(n79), .C(n28), .A(n21), .Y(n19) );
  INVX2 U71 ( .A(n7), .Y(DIFF[8]) );
  NAND2XL U72 ( .A(n40), .B(A[5]), .Y(n15) );
  INVX1 U73 ( .A(n28), .Y(n27) );
  AOI21AX1 U74 ( .B(n16), .C(n78), .A(n15), .Y(n11) );
  NAND21XL U75 ( .B(n29), .A(n30), .Y(n6) );
  NAND21XL U76 ( .B(n25), .A(n26), .Y(n5) );
  NAND21XL U77 ( .B(n17), .A(n18), .Y(n3) );
  NAND21XL U78 ( .B(n22), .A(n23), .Y(n4) );
  NAND2X1 U79 ( .A(n78), .B(n15), .Y(n2) );
  NAND21XL U80 ( .B(n9), .A(n10), .Y(n1) );
  MAJ3X1 U81 ( .A(n38), .B(A[7]), .C(n8), .Y(n7) );
  NAND2XL U82 ( .A(n43), .B(A[2]), .Y(n26) );
  NAND2XL U83 ( .A(n42), .B(A[3]), .Y(n23) );
  INVX3 U84 ( .A(B[0]), .Y(n45) );
  NAND2XL U85 ( .A(n41), .B(A[4]), .Y(n18) );
  NAND2XL U86 ( .A(n39), .B(A[6]), .Y(n10) );
endmodule


module mcu51_cpu_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1XL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  INVXL U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
endmodule


module mcu51_cpu_a0_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVXL U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
endmodule


module mcu51_cpu_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mpb_a0 ( i_rd, i_wr, wdat0, wdat1, addr0, addr1, r_i2c_attr, esfrm_oe, 
        esfrm_we, sfrack, esfrm_wdat, esfrm_adr, mcu_esfr_rdat, delay_rdat, 
        delay_rrdy, esfrm_rrdy, esfrm_rdat, channel_sel, r_pg0_sel, dma_w, 
        dma_r, dma_addr, dma_wdat, dma_ack, memaddr, memaddr_c, memwr, memrd, 
        memrd_c, cpurst, memdatao, memack, hit_xd, hit_xr, hit_ps, hit_ps_c, 
        idat_r, idat_w, idat_adr, idat_wdat, iram_ce, xram_ce, regx_re, 
        iram_we, xram_we, regx_we, iram_a, xram_a, iram_d, xram_d, iram_rdat, 
        xram_rdat, regx_rdat, bist_en, bist_wr, bist_adr, bist_wdat, bist_xram, 
        mclk, srstz, test_si, test_so, test_se );
  input [1:0] i_rd;
  input [1:0] i_wr;
  input [7:0] wdat0;
  input [7:0] wdat1;
  input [7:0] addr0;
  input [7:0] addr1;
  output [7:0] esfrm_wdat;
  output [6:0] esfrm_adr;
  input [7:0] mcu_esfr_rdat;
  input [7:0] delay_rdat;
  output [7:0] esfrm_rdat;
  input [3:0] r_pg0_sel;
  input [10:0] dma_addr;
  input [7:0] dma_wdat;
  input [15:0] memaddr;
  input [15:0] memaddr_c;
  input [7:0] memdatao;
  input [7:0] idat_adr;
  input [7:0] idat_wdat;
  output [10:0] iram_a;
  output [10:0] xram_a;
  output [7:0] iram_d;
  output [7:0] xram_d;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  input [7:0] regx_rdat;
  input [10:0] bist_adr;
  input [7:0] bist_wdat;
  input r_i2c_attr, delay_rrdy, channel_sel, dma_w, dma_r, memwr, memrd,
         memrd_c, cpurst, idat_r, idat_w, bist_en, bist_wr, bist_xram, mclk,
         srstz, test_si, test_se;
  output esfrm_oe, esfrm_we, sfrack, esfrm_rrdy, dma_ack, memack, hit_xd,
         hit_xr, hit_ps, hit_ps_c, iram_ce, xram_ce, regx_re, iram_we, xram_we,
         regx_we, test_so;
  wire   n184, pg0_rdwait, pg0_wrwait, N44, N45, r_pg0_rdrdy, N46,
         xram_rdsel_0_, n62, n65, n66, n67, n80, n107, n109, n111, n126, n127,
         n128, n132, n133, n134, n135, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, net63459, net63462, net63471, net86083, net86087,
         net86095, net86096, net86097, net86098, net86099, net86109, net86112,
         net86116, net86117, net86118, net86120, net86121, net86123, net86124,
         net86125, net86130, net86133, net86136, net86145, net86154, net86157,
         net86159, net86161, net86162, net86164, net86165, net86166, net86167,
         net86170, net86171, net86172, net86173, net86174, net86175, net86176,
         net86178, net86179, net86205, net86208, net86230, net86231, net86246,
         net86247, net86248, net86249, net86257, net86258, net86264, net89000,
         net90956, net91000, net95702, net96925, net97099, net97103, net100914,
         net100995, net101623, net101622, net101621, net86188, net86163, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63,
         n64, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n110, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n129, n130, n131, n136, n137, n138, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183;

  SDFFRQX1 r_pg0_rdrdy_reg ( .D(N46), .SIN(pg0_wrwait), .SMC(test_se), .C(mclk), .XR(srstz), .Q(r_pg0_rdrdy) );
  SDFFRQX1 xram_rdsel_reg_1_ ( .D(n181), .SIN(xram_rdsel_0_), .SMC(test_se), 
        .C(mclk), .XR(srstz), .Q(test_so) );
  SDFFRQX1 xram_rdsel_reg_0_ ( .D(n49), .SIN(n39), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(xram_rdsel_0_) );
  SDFFRQX1 pg0_rdwait_reg ( .D(N45), .SIN(test_si), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(pg0_rdwait) );
  SDFFRQX1 pg0_wrwait_reg ( .D(N44), .SIN(pg0_rdwait), .SMC(test_se), .C(mclk), 
        .XR(srstz), .Q(pg0_wrwait) );
  INVX2 U3 ( .A(n106), .Y(esfrm_adr[0]) );
  BUFXL U4 ( .A(net101621), .Y(n1) );
  INVX3 U5 ( .A(n159), .Y(esfrm_adr[6]) );
  NOR3X1 U6 ( .A(n59), .B(net86097), .C(net95702), .Y(n49) );
  NAND21X2 U7 ( .B(n87), .A(n11), .Y(net86097) );
  BUFX4 U8 ( .A(net86188), .Y(net89000) );
  MUX2X2 U9 ( .D0(addr1[1]), .D1(addr0[1]), .S(net89000), .Y(esfrm_adr[1]) );
  AND2X2 U10 ( .A(net86095), .B(net101621), .Y(esfrm_oe) );
  INVX3 U11 ( .A(net86163), .Y(net86171) );
  BUFX6 U12 ( .A(n184), .Y(xram_a[0]) );
  NAND43X2 U13 ( .B(n116), .C(n115), .D(n51), .A(n113), .Y(xram_a[5]) );
  AND3X2 U14 ( .A(n43), .B(n44), .C(n45), .Y(n117) );
  AO21X1 U15 ( .B(n68), .C(net86098), .A(n49), .Y(net86208) );
  NAND21X1 U16 ( .B(n30), .A(n31), .Y(n35) );
  INVX1 U17 ( .A(r_i2c_attr), .Y(n30) );
  NAND32X1 U18 ( .B(n15), .C(net86205), .A(net90956), .Y(net86163) );
  INVX2 U19 ( .A(net86208), .Y(n15) );
  INVX1 U20 ( .A(net86246), .Y(net86231) );
  INVX1 U21 ( .A(addr1[7]), .Y(net101623) );
  INVX1 U22 ( .A(addr0[7]), .Y(net101622) );
  NAND31X1 U23 ( .C(n27), .A(r_pg0_sel[3]), .B(n28), .Y(n26) );
  INVX1 U24 ( .A(r_pg0_sel[2]), .Y(n27) );
  NAND21X1 U25 ( .B(r_pg0_sel[0]), .A(net86172), .Y(n28) );
  NAND21X1 U26 ( .B(n29), .A(n26), .Y(net86161) );
  INVX1 U27 ( .A(r_pg0_sel[3]), .Y(n29) );
  NAND21X1 U28 ( .B(n21), .A(n22), .Y(net86124) );
  AND2X1 U29 ( .A(net86264), .B(r_pg0_sel[1]), .Y(n21) );
  INVX1 U30 ( .A(i_wr[0]), .Y(n33) );
  INVX1 U31 ( .A(i_rd[0]), .Y(n20) );
  INVX1 U32 ( .A(n37), .Y(net63471) );
  INVX1 U33 ( .A(n26), .Y(n31) );
  OA222X1 U34 ( .A(net63462), .B(n13), .C(net86161), .D(net86162), .E(n12), 
        .F(net86164), .Y(net86159) );
  OAI21BX1 U35 ( .C(n179), .B(n107), .A(n172), .Y(regx_we) );
  NOR2X1 U36 ( .A(n53), .B(n55), .Y(memack) );
  NAND21X1 U37 ( .B(net86157), .A(dma_addr[5]), .Y(n114) );
  NAND21X1 U38 ( .B(pg0_wrwait), .A(n23), .Y(net86116) );
  NAND31X1 U39 ( .C(r_i2c_attr), .A(n34), .B(net100914), .Y(n23) );
  MUX2IX1 U40 ( .D0(net86098), .D1(net86121), .S(n60), .Y(n64) );
  NAND21X1 U41 ( .B(dma_r), .A(n61), .Y(n63) );
  NOR21XL U42 ( .B(n24), .A(n25), .Y(net86166) );
  NOR32XL U43 ( .B(r_pg0_sel[2]), .C(net86170), .A(n31), .Y(n25) );
  NAND2X1 U44 ( .A(net86171), .B(memaddr_c[9]), .Y(n24) );
  INVX1 U45 ( .A(r_pg0_sel[1]), .Y(net86172) );
  OA222X1 U46 ( .A(net86157), .B(net86174), .C(net86175), .D(n12), .E(net86176), .F(n13), .Y(net86173) );
  OAI2B11X1 U47 ( .D(dma_addr[4]), .C(net86157), .A(n152), .B(n112), .Y(
        xram_a[4]) );
  AND3X1 U48 ( .A(n42), .B(n41), .C(n40), .Y(n112) );
  AND3X1 U49 ( .A(n48), .B(n47), .C(n46), .Y(n110) );
  OAI211X1 U50 ( .C(n86), .D(n85), .A(n103), .B(n84), .Y(xram_d[7]) );
  INVX1 U51 ( .A(n114), .Y(n51) );
  INVX1 U52 ( .A(n154), .Y(n115) );
  OAI2B11X1 U53 ( .D(dma_addr[6]), .C(net86157), .A(n157), .B(n117), .Y(
        xram_a[6]) );
  INVX1 U54 ( .A(r_pg0_sel[0]), .Y(net86136) );
  NAND2XL U55 ( .A(memaddr[2]), .B(net86179), .Y(n2) );
  NAND2XL U56 ( .A(net86170), .B(esfrm_adr[2]), .Y(n3) );
  NAND2XL U57 ( .A(memaddr_c[2]), .B(net86171), .Y(n4) );
  AND3X1 U58 ( .A(n2), .B(n3), .C(n4), .Y(n108) );
  INVX4 U59 ( .A(n13), .Y(net86179) );
  NAND2X1 U60 ( .A(net86264), .B(r_pg0_sel[2]), .Y(n22) );
  INVX1 U61 ( .A(n22), .Y(net97103) );
  OAI2B11X1 U62 ( .D(dma_addr[3]), .C(net86157), .A(n149), .B(n110), .Y(
        xram_a[3]) );
  OAI2B11X1 U63 ( .D(dma_addr[2]), .C(net86157), .A(n138), .B(n108), .Y(
        xram_a[2]) );
  OA33X1 U64 ( .A(net86123), .B(net86124), .C(net86125), .D(n167), .E(bist_en), 
        .F(n166), .Y(n5) );
  INVXL U65 ( .A(n22), .Y(n6) );
  INVXL U66 ( .A(net63459), .Y(n7) );
  INVXL U67 ( .A(n7), .Y(n8) );
  INVXL U68 ( .A(n7), .Y(n9) );
  BUFXL U69 ( .A(esfrm_adr[1]), .Y(n10) );
  AO21X1 U70 ( .B(net86130), .C(net86123), .A(n58), .Y(n11) );
  INVXL U71 ( .A(n68), .Y(n181) );
  AOI222XL U72 ( .A(memaddr[1]), .B(net86179), .C(net86170), .D(n10), .E(
        memaddr_c[1]), .F(net86171), .Y(n14) );
  OAI2B11X4 U73 ( .D(dma_addr[1]), .C(net86157), .A(net86154), .B(n14), .Y(
        xram_a[1]) );
  INVX1 U74 ( .A(net86162), .Y(net86170) );
  AOI22XL U75 ( .A(idat_adr[1]), .B(net86117), .C(net86118), .D(n10), .Y(
        net91000) );
  INVXL U76 ( .A(net100995), .Y(net86188) );
  MUX2IXL U77 ( .D0(addr1[4]), .D1(addr0[4]), .S(net86188), .Y(net86145) );
  BUFXL U78 ( .A(net86163), .Y(n12) );
  NAND21XL U79 ( .B(net86205), .A(n15), .Y(net86157) );
  OR3X4 U80 ( .A(n15), .B(net90956), .C(net86205), .Y(n13) );
  NAND21XL U81 ( .B(bist_en), .A(net86096), .Y(net86162) );
  OAI211XL U82 ( .C(net86165), .D(n13), .A(net86166), .B(net86167), .Y(
        xram_a[9]) );
  MUX2IX2 U83 ( .D0(net101622), .D1(net101623), .S(net100995), .Y(net101621)
         );
  NAND32XL U84 ( .B(bist_en), .C(net86208), .A(net86249), .Y(net86248) );
  NAND32XL U85 ( .B(bist_en), .C(net86247), .A(net86208), .Y(net86246) );
  AOI32XL U86 ( .A(net86130), .B(net86096), .C(net86258), .D(net86247), .E(
        test_so), .Y(net86257) );
  OAI32XL U87 ( .A(net86096), .B(net86097), .C(net86098), .D(xram_rdsel_0_), 
        .E(net86099), .Y(dma_ack) );
  INVX1 U88 ( .A(net86096), .Y(net86121) );
  AND3X2 U89 ( .A(net101621), .B(n34), .C(n35), .Y(esfrm_we) );
  MUX2X2 U90 ( .D0(addr1[5]), .D1(addr0[5]), .S(net89000), .Y(esfrm_adr[5]) );
  MUX2X2 U91 ( .D0(addr1[2]), .D1(addr0[2]), .S(net89000), .Y(esfrm_adr[2]) );
  INVX1 U92 ( .A(esfrm_adr[5]), .Y(n156) );
  BUFXL U93 ( .A(esfrm_oe), .Y(n16) );
  INVXL U94 ( .A(n16), .Y(net86087) );
  BUFXL U95 ( .A(esfrm_we), .Y(n17) );
  MUX2IX1 U96 ( .D0(addr1[3]), .D1(addr0[3]), .S(net89000), .Y(n151) );
  NOR21XL U97 ( .B(net86087), .A(n17), .Y(sfrack) );
  INVX2 U98 ( .A(i_rd[1]), .Y(n32) );
  INVXL U99 ( .A(n32), .Y(n36) );
  NAND21X2 U100 ( .B(i_wr[1]), .A(n32), .Y(net100995) );
  INVXL U101 ( .A(n1), .Y(net100914) );
  NAND21XL U102 ( .B(i_wr[1]), .A(n33), .Y(n34) );
  BUFXL U103 ( .A(i_wr[1]), .Y(n37) );
  NAND21X1 U104 ( .B(n36), .A(n20), .Y(net86095) );
  INVXL U105 ( .A(n87), .Y(n88) );
  OAI211X1 U106 ( .C(n106), .D(net86162), .A(n136), .B(n105), .Y(n184) );
  OAI211X1 U107 ( .C(n78), .D(n85), .A(n97), .B(n77), .Y(xram_d[4]) );
  NAND2X1 U108 ( .A(memaddr[6]), .B(net86179), .Y(n43) );
  AND4XL U109 ( .A(memaddr_c[9]), .B(memaddr_c[8]), .C(n49), .D(n181), .Y(n171) );
  NAND2X1 U110 ( .A(memaddr_c[4]), .B(net86171), .Y(n42) );
  MUX2IX1 U111 ( .D0(addr1[0]), .D1(addr0[0]), .S(net89000), .Y(n106) );
  MUX2IX2 U112 ( .D0(addr1[6]), .D1(addr0[6]), .S(net89000), .Y(n159) );
  NAND2X2 U113 ( .A(memaddr_c[6]), .B(net86171), .Y(n45) );
  OA21X1 U114 ( .B(n156), .C(net86162), .A(n50), .Y(n113) );
  NAND2X1 U115 ( .A(memaddr_c[5]), .B(net86171), .Y(n50) );
  MUX2XL U116 ( .D0(net86097), .D1(n178), .S(bist_en), .Y(iram_ce) );
  BUFX3 U117 ( .A(r_pg0_rdrdy), .Y(n39) );
  INVX1 U118 ( .A(net86133), .Y(net97099) );
  NAND21XL U119 ( .B(bist_en), .A(n87), .Y(net86133) );
  INVX1 U120 ( .A(net86125), .Y(net96925) );
  AO22XL U121 ( .A(idat_adr[0]), .B(net86117), .C(net96925), .D(esfrm_adr[0]), 
        .Y(n137) );
  NAND2XL U122 ( .A(net86170), .B(esfrm_adr[4]), .Y(n41) );
  NAND2X1 U123 ( .A(memaddr[4]), .B(net86179), .Y(n40) );
  INVXL U124 ( .A(net86249), .Y(net86247) );
  AOI22X1 U125 ( .A(dma_wdat[4]), .B(net86230), .C(memdatao[4]), .D(net86231), 
        .Y(n77) );
  NAND2XL U126 ( .A(net86170), .B(esfrm_adr[6]), .Y(n44) );
  INVX1 U127 ( .A(net86109), .Y(net86130) );
  INVX1 U128 ( .A(net86257), .Y(net95702) );
  NAND21XL U129 ( .B(dma_w), .A(memrd_c), .Y(n61) );
  NAND2XL U130 ( .A(memaddr[3]), .B(net86179), .Y(n46) );
  NAND2XL U131 ( .A(net86170), .B(esfrm_adr[3]), .Y(n47) );
  NAND2X1 U132 ( .A(memaddr_c[3]), .B(net86171), .Y(n48) );
  NAND21XL U133 ( .B(bist_en), .A(net86247), .Y(n85) );
  INVXL U134 ( .A(net86145), .Y(esfrm_adr[4]) );
  OR2X2 U135 ( .A(idat_r), .B(idat_w), .Y(n87) );
  AND2XL U136 ( .A(memaddr[5]), .B(net86179), .Y(n116) );
  AOI21XL U137 ( .B(xram_rdsel_0_), .C(test_so), .A(n179), .Y(n53) );
  NAND5X1 U138 ( .A(memwr), .B(net86130), .C(net86123), .D(n165), .E(net86098), 
        .Y(n167) );
  NAND32X1 U139 ( .B(n64), .C(net86097), .A(n63), .Y(n68) );
  NAND21XL U140 ( .B(n9), .A(bist_adr[1]), .Y(net86154) );
  NAND21XL U141 ( .B(n9), .A(bist_adr[0]), .Y(n136) );
  OAI221XL U142 ( .A(net86172), .B(net86162), .C(n8), .D(n162), .E(net86173), 
        .Y(xram_a[8]) );
  OAI211XL U143 ( .C(net86136), .D(net86162), .A(n160), .B(n125), .Y(xram_a[7]) );
  INVX1 U144 ( .A(net86157), .Y(net86178) );
  INVX1 U145 ( .A(n56), .Y(n55) );
  INVX1 U146 ( .A(net86133), .Y(net86117) );
  INVX1 U147 ( .A(net86125), .Y(net86118) );
  NAND21XL U148 ( .B(n7), .A(net86121), .Y(net86205) );
  INVX1 U149 ( .A(cpurst), .Y(n56) );
  INVX1 U150 ( .A(n58), .Y(n180) );
  INVX1 U151 ( .A(bist_en), .Y(net63459) );
  NAND21X1 U152 ( .B(n9), .A(bist_wdat[0]), .Y(n89) );
  OAI21X1 U153 ( .B(n66), .C(net86164), .A(n67), .Y(n65) );
  NAND21X1 U154 ( .B(n9), .A(bist_wdat[4]), .Y(n97) );
  INVX1 U155 ( .A(net86164), .Y(net86112) );
  NAND21X1 U156 ( .B(bist_en), .A(n88), .Y(net86125) );
  NAND21X1 U157 ( .B(n9), .A(bist_wdat[1]), .Y(n91) );
  NAND21X1 U158 ( .B(n8), .A(bist_wdat[3]), .Y(n95) );
  NAND21X1 U159 ( .B(n9), .A(bist_wdat[2]), .Y(n93) );
  NAND21X1 U160 ( .B(n8), .A(bist_wdat[6]), .Y(n101) );
  NAND21X1 U161 ( .B(net86083), .A(n58), .Y(n57) );
  INVX1 U162 ( .A(net86248), .Y(net86230) );
  INVX1 U163 ( .A(n66), .Y(n121) );
  INVXL U164 ( .A(n151), .Y(esfrm_adr[3]) );
  INVXL U165 ( .A(net86116), .Y(net86123) );
  INVX1 U166 ( .A(n167), .Y(n179) );
  NAND21XL U167 ( .B(n180), .A(net86116), .Y(net86249) );
  AO21XL U168 ( .B(net86109), .C(n58), .A(net86247), .Y(net86096) );
  NAND21XL U169 ( .B(net86123), .A(net97103), .Y(n172) );
  INVX1 U170 ( .A(n107), .Y(hit_xr) );
  INVX1 U171 ( .A(n78), .Y(esfrm_wdat[4]) );
  INVX1 U172 ( .A(n70), .Y(esfrm_wdat[0]) );
  NAND21X1 U173 ( .B(n6), .A(net86124), .Y(n58) );
  INVX1 U174 ( .A(net86161), .Y(net86264) );
  NOR3XL U175 ( .A(memaddr_c[12]), .B(memaddr_c[13]), .C(memaddr_c[11]), .Y(
        n67) );
  OAI221XL U176 ( .A(n151), .B(net86125), .C(net86133), .D(n150), .E(n149), 
        .Y(iram_a[3]) );
  INVX1 U177 ( .A(idat_adr[3]), .Y(n150) );
  NOR2X1 U178 ( .A(memaddr_c[8]), .B(memaddr_c[9]), .Y(n66) );
  INVX1 U179 ( .A(idat_adr[6]), .Y(n158) );
  OAI221XL U180 ( .A(n156), .B(net86125), .C(net86133), .D(n155), .E(n154), 
        .Y(iram_a[5]) );
  INVX1 U181 ( .A(idat_adr[5]), .Y(n155) );
  OAI221XL U182 ( .A(net86145), .B(net86125), .C(net86133), .D(n153), .E(n152), 
        .Y(iram_a[4]) );
  INVX1 U183 ( .A(idat_adr[4]), .Y(n153) );
  NAND21X1 U184 ( .B(n104), .A(n103), .Y(iram_d[7]) );
  AO22X1 U185 ( .A(idat_wdat[7]), .B(net97099), .C(esfrm_wdat[7]), .D(net86118), .Y(n104) );
  NAND21X1 U186 ( .B(n102), .A(n101), .Y(iram_d[6]) );
  AO22X1 U187 ( .A(idat_wdat[6]), .B(net86117), .C(esfrm_wdat[6]), .D(net86118), .Y(n102) );
  INVX1 U188 ( .A(memaddr_c[10]), .Y(net86164) );
  INVX1 U189 ( .A(memaddr_c[7]), .Y(n120) );
  NAND21X1 U190 ( .B(n98), .A(n97), .Y(iram_d[4]) );
  AO22X1 U191 ( .A(idat_wdat[4]), .B(net86117), .C(net86118), .D(esfrm_wdat[4]), .Y(n98) );
  NAND21X1 U192 ( .B(n100), .A(n99), .Y(iram_d[5]) );
  AO22X1 U193 ( .A(idat_wdat[5]), .B(net86117), .C(esfrm_wdat[5]), .D(net86118), .Y(n100) );
  NAND21X1 U194 ( .B(n96), .A(n95), .Y(iram_d[3]) );
  AO22X1 U195 ( .A(idat_wdat[3]), .B(net86117), .C(esfrm_wdat[3]), .D(net86118), .Y(n96) );
  NAND4X1 U196 ( .A(memaddr_c[14]), .B(memaddr_c[13]), .C(memaddr_c[15]), .D(
        n111), .Y(n109) );
  AND3X1 U197 ( .A(memaddr_c[12]), .B(memaddr_c[7]), .C(memaddr_c[11]), .Y(
        n111) );
  AO21XL U198 ( .B(n6), .C(net86109), .A(n173), .Y(regx_re) );
  NOR43XL U199 ( .B(n172), .C(net86112), .D(n171), .A(n109), .Y(n173) );
  NAND21X1 U200 ( .B(n90), .A(n89), .Y(iram_d[0]) );
  AO22X1 U201 ( .A(idat_wdat[0]), .B(net86117), .C(net86118), .D(esfrm_wdat[0]), .Y(n90) );
  NAND21X1 U202 ( .B(n94), .A(n93), .Y(iram_d[2]) );
  AO22X1 U203 ( .A(idat_wdat[2]), .B(net86117), .C(esfrm_wdat[2]), .D(net86118), .Y(n94) );
  NAND21X1 U204 ( .B(n92), .A(n91), .Y(iram_d[1]) );
  AO22X1 U205 ( .A(idat_wdat[1]), .B(net97099), .C(esfrm_wdat[1]), .D(net96925), .Y(n92) );
  INVX1 U206 ( .A(hit_xd), .Y(n166) );
  NAND21XL U207 ( .B(n16), .A(n54), .Y(esfrm_rrdy) );
  OAI211X1 U208 ( .C(n168), .D(n178), .A(n5), .B(n177), .Y(xram_we) );
  NAND21X1 U209 ( .B(n8), .A(bist_wdat[5]), .Y(n99) );
  INVX1 U210 ( .A(idat_adr[7]), .Y(n161) );
  AND3XL U211 ( .A(net86116), .B(n87), .C(n57), .Y(N44) );
  OA21XL U212 ( .B(net97103), .C(n88), .A(net86109), .Y(N46) );
  AND3XL U213 ( .A(net86109), .B(n87), .C(n57), .Y(N45) );
  NAND21X1 U214 ( .B(n8), .A(bist_wr), .Y(n168) );
  INVX1 U215 ( .A(iram_a[9]), .Y(n129) );
  INVX1 U216 ( .A(net86124), .Y(net86083) );
  OA21X1 U217 ( .B(idat_adr[4]), .C(idat_adr[3]), .A(idat_adr[5]), .Y(n127) );
  AOI31X1 U218 ( .A(idat_adr[4]), .B(idat_adr[6]), .C(idat_adr[5]), .D(
        idat_adr[7]), .Y(n128) );
  INVX1 U219 ( .A(n80), .Y(n119) );
  AOI32XL U220 ( .A(memrd_c), .B(n165), .C(net86098), .D(n60), .E(net86109), 
        .Y(n59) );
  OAI211X1 U221 ( .C(n70), .D(n85), .A(n89), .B(n69), .Y(xram_d[0]) );
  AOI22X1 U222 ( .A(dma_wdat[0]), .B(net86230), .C(memdatao[0]), .D(net86231), 
        .Y(n69) );
  INVX1 U223 ( .A(memaddr[10]), .Y(net63462) );
  INVX1 U224 ( .A(memaddr[11]), .Y(n183) );
  NAND6XL U225 ( .A(memaddr[14]), .B(memaddr[15]), .C(memaddr[13]), .D(
        memaddr[11]), .E(memaddr[12]), .F(n164), .Y(n107) );
  AND4X1 U226 ( .A(memaddr[9]), .B(memaddr[10]), .C(memaddr[8]), .D(memaddr[7]), .Y(n164) );
  AOI211X1 U227 ( .C(memaddr[14]), .D(n134), .A(memaddr[15]), .B(n55), .Y(
        hit_ps) );
  NAND4X1 U228 ( .A(n183), .B(net63462), .C(n80), .D(n135), .Y(n134) );
  NOR3XL U229 ( .A(memaddr[12]), .B(memaddr[7]), .C(memaddr[13]), .Y(n135) );
  NOR2X1 U230 ( .A(memaddr[8]), .B(memaddr[9]), .Y(n80) );
  NOR4XL U231 ( .A(memaddr[14]), .B(memaddr[15]), .C(memaddr[13]), .D(n132), 
        .Y(hit_xd) );
  OAI211X1 U232 ( .C(net63462), .D(n80), .A(n182), .B(n183), .Y(n132) );
  INVX1 U233 ( .A(memaddr[12]), .Y(n182) );
  NAND21X1 U234 ( .B(n8), .A(bist_adr[5]), .Y(n154) );
  INVX1 U235 ( .A(esfrm_wdat[7]), .Y(n86) );
  AOI22XL U236 ( .A(dma_wdat[7]), .B(net86230), .C(memdatao[7]), .D(net86231), 
        .Y(n84) );
  NAND21X1 U237 ( .B(test_so), .A(xram_rdsel_0_), .Y(n60) );
  NAND21X1 U238 ( .B(n8), .A(bist_adr[2]), .Y(n138) );
  NAND21X1 U239 ( .B(n8), .A(bist_adr[3]), .Y(n149) );
  NAND21X1 U240 ( .B(n9), .A(bist_adr[4]), .Y(n152) );
  NAND21X1 U241 ( .B(n9), .A(bist_adr[6]), .Y(n157) );
  OAI211X1 U242 ( .C(n72), .D(n85), .A(n91), .B(n71), .Y(xram_d[1]) );
  INVX1 U243 ( .A(esfrm_wdat[1]), .Y(n72) );
  AOI22XL U244 ( .A(dma_wdat[1]), .B(net86230), .C(memdatao[1]), .D(net86231), 
        .Y(n71) );
  NAND21X1 U245 ( .B(n148), .A(n138), .Y(iram_a[2]) );
  AO22XL U246 ( .A(idat_adr[2]), .B(net86117), .C(net86118), .D(esfrm_adr[2]), 
        .Y(n148) );
  NAND2X1 U247 ( .A(net91000), .B(net86154), .Y(iram_a[1]) );
  OAI211X1 U248 ( .C(n74), .D(n85), .A(n93), .B(n73), .Y(xram_d[2]) );
  INVX1 U249 ( .A(esfrm_wdat[2]), .Y(n74) );
  AOI22XL U250 ( .A(dma_wdat[2]), .B(net86230), .C(memdatao[2]), .D(net86231), 
        .Y(n73) );
  OAI211X1 U251 ( .C(n83), .D(n85), .A(n101), .B(n82), .Y(xram_d[6]) );
  INVX1 U252 ( .A(esfrm_wdat[6]), .Y(n83) );
  AOI22XL U253 ( .A(dma_wdat[6]), .B(net86230), .C(memdatao[6]), .D(net86231), 
        .Y(n82) );
  OAI211X1 U254 ( .C(n81), .D(n85), .A(n99), .B(n79), .Y(xram_d[5]) );
  INVX1 U255 ( .A(esfrm_wdat[5]), .Y(n81) );
  AOI22XL U256 ( .A(dma_wdat[5]), .B(net86230), .C(memdatao[5]), .D(net86231), 
        .Y(n79) );
  OAI211X1 U257 ( .C(n76), .D(n85), .A(n95), .B(n75), .Y(xram_d[3]) );
  INVX1 U258 ( .A(esfrm_wdat[3]), .Y(n76) );
  AOI22XL U259 ( .A(dma_wdat[3]), .B(net86230), .C(memdatao[3]), .D(net86231), 
        .Y(n75) );
  OAI211X1 U260 ( .C(n181), .D(n5), .A(n177), .B(n176), .Y(xram_ce) );
  MUX3IX1 U261 ( .D0(n175), .D1(n174), .D2(bist_xram), .S0(n49), .S1(bist_en), 
        .Y(n176) );
  AND2X1 U262 ( .A(n181), .B(n62), .Y(n175) );
  OAI31XL U263 ( .A(n65), .B(memaddr_c[15]), .C(memaddr_c[14]), .D(n181), .Y(
        n174) );
  AOI211X1 U264 ( .C(memaddr_c[14]), .D(n133), .A(memaddr_c[15]), .B(n55), .Y(
        hit_ps_c) );
  NAND42X1 U265 ( .C(memaddr_c[7]), .D(memaddr_c[10]), .A(n66), .B(n67), .Y(
        n133) );
  INVX1 U266 ( .A(xram_rdsel_0_), .Y(net86258) );
  OAI2B11X1 U267 ( .D(n126), .C(net86133), .A(net86125), .B(n163), .Y(
        iram_a[10]) );
  OAI211X1 U268 ( .C(net86157), .D(n131), .A(n163), .B(net86159), .Y(
        xram_a[10]) );
  OAI211X1 U269 ( .C(n127), .D(idat_adr[6]), .A(n128), .B(channel_sel), .Y(
        n126) );
  NOR2X1 U270 ( .A(memrd), .B(memwr), .Y(net90956) );
  NAND21X1 U271 ( .B(n137), .A(n136), .Y(iram_a[0]) );
  OAI221X1 U272 ( .A(net86125), .B(net86136), .C(net86133), .D(n161), .E(n160), 
        .Y(iram_a[7]) );
  INVX1 U273 ( .A(memaddr[9]), .Y(net86165) );
  OA21X1 U274 ( .B(net86157), .C(n130), .A(n129), .Y(net86167) );
  NAND32X1 U275 ( .B(net96925), .C(net97099), .A(n162), .Y(iram_a[8]) );
  INVX1 U276 ( .A(bist_adr[8]), .Y(n162) );
  INVX1 U277 ( .A(dma_addr[8]), .Y(net86174) );
  INVX1 U278 ( .A(memaddr[8]), .Y(net86176) );
  INVX1 U279 ( .A(memaddr_c[8]), .Y(net86175) );
  AOI222XL U280 ( .A(dma_addr[7]), .B(net86178), .C(net86179), .D(n124), .E(
        net86171), .F(n123), .Y(n125) );
  OAI31XL U281 ( .A(memaddr[10]), .B(n119), .C(n122), .D(n118), .Y(n124) );
  OAI31XL U282 ( .A(net86112), .B(n122), .C(n121), .D(n120), .Y(n123) );
  INVX1 U283 ( .A(channel_sel), .Y(n122) );
  NOR21XL U284 ( .B(delay_rrdy), .A(r_pg0_rdrdy), .Y(n140) );
  AO222X1 U285 ( .A(mcu_esfr_rdat[7]), .B(n54), .C(r_pg0_rdrdy), .D(n139), .E(
        delay_rdat[7]), .F(n140), .Y(esfrm_rdat[7]) );
  AO222XL U286 ( .A(xram_rdat[7]), .B(net86083), .C(iram_rdat[7]), .D(n180), 
        .E(regx_rdat[7]), .F(n6), .Y(n139) );
  NOR2X1 U287 ( .A(r_pg0_rdrdy), .B(delay_rrdy), .Y(n54) );
  AO222XL U288 ( .A(xram_rdat[0]), .B(net86083), .C(iram_rdat[0]), .D(n180), 
        .E(regx_rdat[0]), .F(net97103), .Y(n147) );
  AO222XL U289 ( .A(n178), .B(n170), .C(n169), .D(net86116), .E(idat_w), .F(
        net86117), .Y(iram_we) );
  INVX1 U290 ( .A(n168), .Y(n170) );
  AND2X1 U291 ( .A(net86118), .B(n180), .Y(n169) );
  AO222X1 U292 ( .A(mcu_esfr_rdat[6]), .B(n54), .C(r_pg0_rdrdy), .D(n141), .E(
        delay_rdat[6]), .F(n140), .Y(esfrm_rdat[6]) );
  AO222XL U293 ( .A(xram_rdat[6]), .B(net86083), .C(iram_rdat[6]), .D(n180), 
        .E(regx_rdat[6]), .F(n6), .Y(n141) );
  AO222XL U294 ( .A(mcu_esfr_rdat[1]), .B(n54), .C(r_pg0_rdrdy), .D(n146), .E(
        delay_rdat[1]), .F(n140), .Y(esfrm_rdat[1]) );
  AO222XL U295 ( .A(xram_rdat[1]), .B(net86083), .C(iram_rdat[1]), .D(n180), 
        .E(regx_rdat[1]), .F(n6), .Y(n146) );
  AO222XL U296 ( .A(mcu_esfr_rdat[2]), .B(n54), .C(r_pg0_rdrdy), .D(n145), .E(
        delay_rdat[2]), .F(n140), .Y(esfrm_rdat[2]) );
  AO222XL U297 ( .A(xram_rdat[2]), .B(net86083), .C(iram_rdat[2]), .D(n180), 
        .E(regx_rdat[2]), .F(net97103), .Y(n145) );
  AO222X1 U298 ( .A(mcu_esfr_rdat[5]), .B(n54), .C(r_pg0_rdrdy), .D(n142), .E(
        delay_rdat[5]), .F(n140), .Y(esfrm_rdat[5]) );
  AO222XL U299 ( .A(xram_rdat[5]), .B(net86083), .C(iram_rdat[5]), .D(n180), 
        .E(regx_rdat[5]), .F(net97103), .Y(n142) );
  AO222X1 U300 ( .A(mcu_esfr_rdat[3]), .B(n54), .C(r_pg0_rdrdy), .D(n144), .E(
        delay_rdat[3]), .F(n140), .Y(esfrm_rdat[3]) );
  AO222XL U301 ( .A(xram_rdat[3]), .B(net86083), .C(iram_rdat[3]), .D(n180), 
        .E(regx_rdat[3]), .F(net97103), .Y(n144) );
  AO222X1 U302 ( .A(mcu_esfr_rdat[4]), .B(n54), .C(n39), .D(n143), .E(
        delay_rdat[4]), .F(n140), .Y(esfrm_rdat[4]) );
  AO222XL U303 ( .A(xram_rdat[4]), .B(net86083), .C(iram_rdat[4]), .D(n180), 
        .E(regx_rdat[4]), .F(n6), .Y(n143) );
  NAND21X1 U304 ( .B(n8), .A(bist_wdat[7]), .Y(n103) );
  NOR21XL U305 ( .B(bist_adr[9]), .A(n8), .Y(iram_a[9]) );
  NAND21X1 U306 ( .B(net63459), .A(bist_adr[10]), .Y(n163) );
  NAND21X1 U307 ( .B(n9), .A(bist_adr[7]), .Y(n160) );
  INVX1 U308 ( .A(memaddr[7]), .Y(n118) );
  NAND5XL U309 ( .A(n62), .B(dma_w), .C(n9), .D(net86120), .E(net86121), .Y(
        n177) );
  INVXL U310 ( .A(net86097), .Y(net86120) );
  INVX1 U311 ( .A(test_so), .Y(net86099) );
  INVX1 U312 ( .A(dma_w), .Y(net86098) );
  OAI21X1 U313 ( .B(dma_addr[9]), .C(dma_addr[8]), .A(dma_addr[10]), .Y(n62)
         );
  INVX1 U314 ( .A(dma_r), .Y(n165) );
  INVX1 U315 ( .A(bist_xram), .Y(n178) );
  INVX1 U316 ( .A(dma_addr[10]), .Y(n131) );
  INVX1 U317 ( .A(dma_addr[9]), .Y(n130) );
  AOI222XL U318 ( .A(dma_addr[0]), .B(net86178), .C(memaddr_c[0]), .D(net86171), .E(memaddr[0]), .F(net86179), .Y(n105) );
  AO21XL U319 ( .B(net100914), .C(net86095), .A(pg0_rdwait), .Y(net86109) );
  AO22XL U320 ( .A(wdat1[7]), .B(n37), .C(wdat0[7]), .D(net63471), .Y(
        esfrm_wdat[7]) );
  AO22XL U321 ( .A(wdat1[6]), .B(n37), .C(wdat0[6]), .D(net63471), .Y(
        esfrm_wdat[6]) );
  AO22XL U322 ( .A(wdat1[5]), .B(n37), .C(wdat0[5]), .D(net63471), .Y(
        esfrm_wdat[5]) );
  AO22XL U323 ( .A(wdat1[3]), .B(n37), .C(wdat0[3]), .D(net63471), .Y(
        esfrm_wdat[3]) );
  AO22XL U324 ( .A(wdat1[2]), .B(n37), .C(wdat0[2]), .D(net63471), .Y(
        esfrm_wdat[2]) );
  AO22XL U325 ( .A(wdat1[1]), .B(n37), .C(wdat0[1]), .D(net63471), .Y(
        esfrm_wdat[1]) );
  MUX2IXL U326 ( .D0(wdat0[4]), .D1(wdat1[4]), .S(n37), .Y(n78) );
  MUX2IXL U327 ( .D0(wdat0[0]), .D1(wdat1[0]), .S(n37), .Y(n70) );
  OAI221XL U328 ( .A(n159), .B(net86125), .C(net86133), .D(n158), .E(n157), 
        .Y(iram_a[6]) );
  AO222XL U329 ( .A(mcu_esfr_rdat[0]), .B(n54), .C(r_pg0_rdrdy), .D(n147), .E(
        delay_rdat[0]), .F(n140), .Y(esfrm_rdat[0]) );
endmodule

